VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 8bitdac_layout
  CLASS BLOCK ;
  FOREIGN 8bitdac_layout ;
  ORIGIN 29.390 25.310 ;
  SIZE 528.610 BY 301.560 ;
  PIN x1_vref5
    ANTENNADIFFAREA 1.081500 ;
    PORT
      LAYER nwell ;
        RECT 116.330 14.860 118.250 17.120 ;
        RECT 117.300 14.770 118.150 14.860 ;
      LAYER li1 ;
        RECT 113.550 15.300 113.850 16.300 ;
        RECT 117.600 15.300 117.860 16.850 ;
        RECT 113.500 15.290 118.750 15.300 ;
        RECT 103.380 15.210 103.630 15.220 ;
        RECT 103.380 14.750 104.360 15.210 ;
        RECT 113.500 15.000 118.770 15.290 ;
        RECT 103.380 14.450 103.630 14.750 ;
        RECT 111.350 14.660 113.190 14.670 ;
        RECT 118.600 14.660 118.770 15.000 ;
        RECT 105.090 14.650 105.330 14.660 ;
        RECT 106.170 14.650 118.770 14.660 ;
        RECT 105.090 14.490 118.770 14.650 ;
        RECT 105.090 14.480 116.600 14.490 ;
        RECT 105.080 14.470 111.400 14.480 ;
        RECT 112.950 14.470 116.600 14.480 ;
        RECT 105.080 14.460 106.950 14.470 ;
        RECT 105.080 14.450 105.330 14.460 ;
        RECT 103.380 14.280 105.330 14.450 ;
        RECT 103.380 13.980 103.650 14.280 ;
        RECT 103.390 13.720 103.650 13.980 ;
        RECT 103.370 13.330 103.670 13.720 ;
        RECT 103.360 12.930 103.670 13.330 ;
        RECT 103.360 12.670 103.650 12.930 ;
        RECT 103.340 12.500 103.650 12.670 ;
        RECT 103.340 12.140 103.630 12.500 ;
        RECT 103.330 12.090 103.630 12.140 ;
        RECT 103.330 11.790 103.600 12.090 ;
        RECT 103.000 11.640 103.600 11.790 ;
        RECT 103.000 10.920 103.510 11.640 ;
        RECT 103.050 10.090 103.500 10.920 ;
    END
  END x1_vref5
  PIN x2_vref1
    ANTENNADIFFAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 105.950 256.390 108.730 256.400 ;
        RECT 105.950 256.370 187.300 256.390 ;
        RECT 101.850 256.360 187.300 256.370 ;
        RECT 101.850 256.170 240.770 256.360 ;
        RECT 101.850 256.150 106.950 256.170 ;
        RECT 101.860 256.050 102.260 256.150 ;
        RECT 240.490 253.310 240.770 256.170 ;
        RECT 240.460 252.970 240.790 253.310 ;
        RECT 240.490 252.950 240.770 252.970 ;
        RECT 101.910 247.800 102.280 252.160 ;
        RECT 240.510 251.450 240.800 252.250 ;
        RECT 240.520 251.320 240.800 251.450 ;
        RECT 240.520 251.140 240.810 251.320 ;
        RECT 240.530 250.870 240.810 251.140 ;
        RECT 240.530 250.640 240.830 250.870 ;
        RECT 240.540 250.470 240.830 250.640 ;
        RECT 240.550 249.670 240.810 250.470 ;
        RECT 240.550 249.070 240.800 249.670 ;
        RECT 239.760 248.620 240.800 249.070 ;
        RECT 101.900 130.960 102.300 247.800 ;
        RECT 101.900 130.810 102.330 130.960 ;
        RECT 101.930 14.050 102.330 130.810 ;
        RECT 101.930 11.560 102.360 14.050 ;
        RECT 101.910 11.440 102.360 11.560 ;
        RECT 101.910 9.400 102.340 11.440 ;
        RECT 103.910 9.870 104.370 10.740 ;
        RECT 103.880 9.400 104.390 9.870 ;
        RECT 101.910 8.950 104.420 9.400 ;
        RECT 101.930 8.940 104.420 8.950 ;
      LAYER mcon ;
        RECT 101.995 256.105 102.165 256.275 ;
        RECT 240.555 253.045 240.725 253.215 ;
        RECT 101.995 251.885 102.165 252.055 ;
        RECT 240.595 252.035 240.765 252.205 ;
      LAYER met1 ;
        RECT 101.880 251.790 102.250 256.380 ;
        RECT 240.460 253.290 240.790 253.310 ;
        RECT 240.460 252.970 240.840 253.290 ;
        RECT 240.500 252.280 240.840 252.970 ;
        RECT 240.490 252.060 240.840 252.280 ;
        RECT 240.490 251.940 240.820 252.060 ;
    END
  END x2_vref1
  PIN inp1
    ANTENNADIFFAREA 0.060900 ;
    PORT
      LAYER li1 ;
        RECT 3.980 252.930 4.270 253.360 ;
        RECT 3.980 251.510 4.270 252.310 ;
        RECT 3.990 251.380 4.270 251.510 ;
        RECT 3.990 251.200 4.280 251.380 ;
        RECT 4.000 250.930 4.280 251.200 ;
        RECT 4.000 250.700 4.300 250.930 ;
        RECT 4.010 250.530 4.300 250.700 ;
        RECT 4.020 249.730 4.280 250.530 ;
        RECT 4.020 249.130 4.270 249.730 ;
        RECT 3.230 248.680 4.270 249.130 ;
      LAYER mcon ;
        RECT 4.055 252.955 4.225 253.125 ;
        RECT 4.045 252.085 4.215 252.255 ;
      LAYER met1 ;
        RECT 3.125 253.925 5.265 254.900 ;
        RECT 3.980 252.020 4.270 253.925 ;
      LAYER via ;
        RECT 3.170 254.790 4.015 254.795 ;
        RECT 3.170 253.960 5.155 254.790 ;
        RECT 4.030 253.955 5.155 253.960 ;
      LAYER met2 ;
        RECT 3.795 272.355 4.685 276.250 ;
        RECT 3.125 253.925 5.265 272.355 ;
    END
  END inp1
  PIN inp2
    ANTENNADIFFAREA 1.020600 ;
    PORT
      LAYER nwell ;
        RECT 352.860 14.800 354.780 17.060 ;
        RECT 353.830 14.710 354.680 14.800 ;
      LAYER li1 ;
        RECT 350.080 15.240 350.380 16.240 ;
        RECT 354.130 15.240 354.390 16.790 ;
        RECT 350.030 15.230 355.280 15.240 ;
        RECT 339.910 15.150 340.160 15.160 ;
        RECT 339.910 14.690 340.890 15.150 ;
        RECT 350.030 14.940 355.300 15.230 ;
        RECT 339.910 14.390 340.160 14.690 ;
        RECT 347.880 14.600 349.720 14.610 ;
        RECT 355.130 14.600 355.300 14.940 ;
        RECT 341.620 14.590 341.860 14.600 ;
        RECT 342.700 14.590 355.300 14.600 ;
        RECT 341.620 14.430 355.300 14.590 ;
        RECT 341.620 14.420 353.130 14.430 ;
        RECT 341.610 14.410 347.930 14.420 ;
        RECT 349.480 14.410 353.130 14.420 ;
        RECT 341.610 14.400 343.480 14.410 ;
        RECT 341.610 14.390 341.860 14.400 ;
        RECT 339.910 14.220 341.860 14.390 ;
        RECT 339.910 13.920 340.180 14.220 ;
        RECT 339.920 13.660 340.180 13.920 ;
        RECT 339.900 13.270 340.200 13.660 ;
        RECT 339.890 12.870 340.200 13.270 ;
        RECT 339.890 12.610 340.180 12.870 ;
        RECT 339.870 12.440 340.180 12.610 ;
        RECT 339.870 12.080 340.160 12.440 ;
        RECT 339.860 12.030 340.160 12.080 ;
        RECT 339.860 11.770 340.130 12.030 ;
        RECT 339.045 11.105 341.490 11.770 ;
      LAYER mcon ;
        RECT 339.150 11.400 341.425 11.695 ;
        RECT 339.150 11.230 341.430 11.400 ;
      LAYER met1 ;
        RECT 339.040 -15.045 341.500 12.055 ;
      LAYER via ;
        RECT 339.115 -14.245 339.375 -14.240 ;
        RECT 339.115 -14.250 339.660 -14.245 ;
        RECT 340.265 -14.250 340.525 -14.245 ;
        RECT 339.115 -15.030 340.195 -14.250 ;
        RECT 339.400 -15.035 340.195 -15.030 ;
        RECT 340.265 -15.035 341.345 -14.250 ;
      LAYER met2 ;
        RECT 339.040 -19.450 341.500 -14.220 ;
        RECT 339.785 -25.310 340.365 -19.450 ;
    END
  END inp2
  PIN d7
    ANTENNAGATEAREA 0.271500 ;
    PORT
      LAYER li1 ;
        RECT 469.650 134.150 470.550 134.610 ;
        RECT 469.770 134.140 470.550 134.150 ;
      LAYER mcon ;
        RECT 469.835 134.300 470.005 134.470 ;
      LAYER met1 ;
        RECT 468.515 134.135 470.100 134.610 ;
      LAYER via ;
        RECT 468.550 134.250 469.065 134.510 ;
      LAYER met2 ;
        RECT 467.920 134.135 469.100 134.610 ;
      LAYER via2 ;
        RECT 467.970 134.230 468.250 134.510 ;
        RECT 468.290 134.235 468.570 134.515 ;
        RECT 468.595 134.235 468.875 134.515 ;
      LAYER met3 ;
        RECT 467.920 125.975 469.085 134.610 ;
        RECT 467.920 124.760 497.080 125.975 ;
        RECT 467.920 123.960 499.220 124.760 ;
        RECT 467.920 123.105 497.080 123.960 ;
        RECT 467.920 123.100 469.085 123.105 ;
    END
  END d7
  PIN out_v
    ANTENNADIFFAREA 1.516100 ;
    PORT
      LAYER li1 ;
        RECT 476.620 134.660 476.880 136.270 ;
        RECT 479.170 135.200 479.470 136.250 ;
        RECT 476.610 134.600 476.880 134.660 ;
        RECT 478.160 134.940 479.470 135.200 ;
        RECT 481.600 134.940 482.600 135.260 ;
        RECT 478.160 134.600 478.470 134.940 ;
        RECT 476.610 134.310 478.470 134.600 ;
        RECT 476.610 134.300 476.920 134.310 ;
        RECT 478.160 134.300 478.470 134.310 ;
        RECT 476.620 133.250 476.920 134.300 ;
        RECT 479.220 133.200 479.470 134.940 ;
      LAYER mcon ;
        RECT 479.230 135.010 479.400 135.180 ;
        RECT 481.655 135.010 481.825 135.180 ;
      LAYER met1 ;
        RECT 481.600 135.250 483.290 135.265 ;
        RECT 479.170 134.950 483.290 135.250 ;
        RECT 481.600 134.935 483.290 134.950 ;
        RECT 481.600 134.930 481.930 134.935 ;
      LAYER via ;
        RECT 481.950 134.975 482.860 135.235 ;
        RECT 482.865 134.975 483.125 135.235 ;
      LAYER met2 ;
        RECT 481.600 134.935 485.000 135.265 ;
      LAYER via2 ;
        RECT 483.095 134.960 483.375 135.240 ;
        RECT 483.410 134.955 483.690 135.235 ;
        RECT 483.705 134.955 484.260 135.235 ;
        RECT 484.270 134.955 484.830 135.235 ;
      LAYER met3 ;
        RECT 482.575 135.595 497.005 141.245 ;
        RECT 482.575 134.795 499.220 135.595 ;
        RECT 482.575 129.945 497.005 134.795 ;
    END
  END out_v
  PIN x1_out_v
    ANTENNADIFFAREA 2.463700 ;
    PORT
      LAYER nwell ;
        RECT 475.620 137.050 476.470 137.160 ;
        RECT 475.400 134.820 477.310 137.050 ;
      LAYER li1 ;
        RECT 228.850 257.770 453.900 257.810 ;
        RECT 476.800 257.770 480.920 257.790 ;
        RECT 228.850 257.600 480.920 257.770 ;
        RECT 228.850 256.630 229.120 257.600 ;
        RECT 476.820 257.580 480.920 257.600 ;
        RECT 480.740 257.330 480.920 257.580 ;
        RECT 228.840 249.080 229.090 255.980 ;
        RECT 222.790 137.070 223.050 138.680 ;
        RECT 225.340 137.610 225.640 138.660 ;
        RECT 228.840 137.710 229.080 249.080 ;
        RECT 480.740 246.010 480.950 257.330 ;
        RECT 480.730 138.110 480.950 246.010 ;
        RECT 480.730 137.900 480.980 138.110 ;
        RECT 222.780 137.010 223.050 137.070 ;
        RECT 224.330 137.350 225.640 137.610 ;
        RECT 227.840 137.370 229.080 137.710 ;
        RECT 224.330 137.010 224.640 137.350 ;
        RECT 222.780 136.720 224.640 137.010 ;
        RECT 222.780 136.710 223.090 136.720 ;
        RECT 224.330 136.710 224.640 136.720 ;
        RECT 222.790 135.660 223.090 136.710 ;
        RECT 225.390 135.610 225.640 137.350 ;
        RECT 480.750 136.900 480.980 137.900 ;
        RECT 475.720 136.610 480.980 136.900 ;
        RECT 475.720 136.600 480.970 136.610 ;
        RECT 475.920 135.050 476.170 136.600 ;
        RECT 479.920 135.650 480.220 136.600 ;
      LAYER mcon ;
        RECT 228.885 256.680 229.055 256.850 ;
        RECT 228.885 255.780 229.055 255.950 ;
        RECT 225.400 137.420 225.570 137.590 ;
        RECT 227.960 137.435 228.130 137.605 ;
      LAYER met1 ;
        RECT 228.830 256.860 229.120 256.920 ;
        RECT 228.820 256.630 229.120 256.860 ;
        RECT 228.840 255.960 229.110 256.630 ;
        RECT 228.830 255.700 229.110 255.960 ;
        RECT 227.840 137.660 228.220 137.700 ;
        RECT 225.340 137.370 228.220 137.660 ;
        RECT 225.340 137.360 228.040 137.370 ;
    END
  END x1_out_v
  PIN x2_out_v
    ANTENNADIFFAREA 2.471600 ;
    PORT
      LAYER nwell ;
        RECT 478.650 132.410 480.570 134.670 ;
        RECT 479.620 132.320 480.470 132.410 ;
      LAYER li1 ;
        RECT 459.320 137.010 459.580 138.620 ;
        RECT 461.870 137.550 462.170 138.600 ;
        RECT 465.160 137.650 465.560 137.670 ;
        RECT 459.310 136.950 459.580 137.010 ;
        RECT 460.860 137.290 462.170 137.550 ;
        RECT 464.370 137.310 465.600 137.650 ;
        RECT 460.860 136.950 461.170 137.290 ;
        RECT 459.310 136.660 461.170 136.950 ;
        RECT 459.310 136.650 459.620 136.660 ;
        RECT 460.860 136.650 461.170 136.660 ;
        RECT 459.320 135.600 459.620 136.650 ;
        RECT 461.920 135.550 462.170 137.290 ;
        RECT 465.160 130.480 465.560 137.310 ;
        RECT 475.870 132.850 476.170 133.850 ;
        RECT 479.920 132.850 480.180 134.400 ;
        RECT 475.820 132.550 481.070 132.850 ;
        RECT 480.860 131.820 481.070 132.550 ;
        RECT 480.860 130.600 481.090 131.820 ;
        RECT 480.860 130.500 481.060 130.600 ;
        RECT 467.700 130.480 481.060 130.500 ;
        RECT 465.160 130.150 481.060 130.480 ;
        RECT 465.160 130.130 467.810 130.150 ;
      LAYER mcon ;
        RECT 461.930 137.360 462.100 137.530 ;
        RECT 464.490 137.375 464.660 137.545 ;
      LAYER met1 ;
        RECT 464.370 137.600 464.750 137.640 ;
        RECT 461.870 137.310 464.750 137.600 ;
        RECT 461.870 137.300 464.570 137.310 ;
    END
  END x2_out_v
  PIN d6
    ANTENNAGATEAREA 0.543000 ;
    PORT
      LAYER li1 ;
        RECT 215.680 137.020 216.100 137.040 ;
        RECT 215.610 136.550 216.720 137.020 ;
        RECT 452.210 136.960 452.630 136.980 ;
        RECT 215.610 136.520 216.100 136.550 ;
        RECT 215.610 133.410 215.810 136.520 ;
        RECT 451.880 136.490 453.250 136.960 ;
        RECT 451.880 136.460 452.630 136.490 ;
        RECT 451.880 133.290 452.340 136.460 ;
        RECT 215.550 132.360 215.820 132.630 ;
        RECT 215.580 127.030 215.820 132.360 ;
        RECT 215.550 121.930 215.820 127.030 ;
        RECT 215.510 119.640 215.820 121.930 ;
        RECT 215.510 6.460 215.770 119.640 ;
        RECT 215.460 -0.540 215.790 6.460 ;
        RECT 441.460 -0.510 448.210 -0.490 ;
        RECT 451.880 -0.510 452.170 132.300 ;
        RECT 441.460 -0.540 452.170 -0.510 ;
        RECT 215.450 -0.840 452.170 -0.540 ;
        RECT 215.450 -0.860 425.550 -0.840 ;
        RECT 426.130 -0.860 452.170 -0.840 ;
        RECT 215.450 -0.930 216.180 -0.860 ;
        RECT 441.460 -0.920 452.170 -0.860 ;
      LAYER mcon ;
        RECT 215.620 133.485 215.790 133.655 ;
        RECT 452.005 133.605 452.175 133.775 ;
        RECT 215.600 132.415 215.770 132.585 ;
        RECT 451.945 131.835 452.115 132.005 ;
        RECT 220.835 -0.770 221.005 -0.600 ;
        RECT 221.095 -0.770 221.265 -0.600 ;
        RECT 221.345 -0.770 221.515 -0.600 ;
        RECT 221.605 -0.770 221.775 -0.600 ;
      LAYER met1 ;
        RECT 215.580 133.710 215.810 133.790 ;
        RECT 215.580 133.430 215.820 133.710 ;
        RECT 215.580 132.630 215.810 133.430 ;
        RECT 215.550 132.360 215.810 132.630 ;
        RECT 215.580 132.350 215.810 132.360 ;
        RECT 451.810 131.700 452.340 133.960 ;
        RECT 220.760 -15.035 221.880 -0.495 ;
      LAYER via ;
        RECT 220.895 -14.965 221.740 -14.130 ;
      LAYER met2 ;
        RECT 220.765 -19.465 221.870 -13.990 ;
        RECT 220.960 -25.310 221.540 -19.465 ;
    END
  END d6
  PIN d5
    ANTENNAGATEAREA 1.086000 ;
    PORT
      LAYER li1 ;
        RECT 88.020 134.880 88.430 134.890 ;
        RECT 88.020 134.860 89.130 134.880 ;
        RECT 87.560 134.430 89.130 134.860 ;
        RECT 324.550 134.820 324.960 134.830 ;
        RECT 324.550 134.800 325.660 134.820 ;
        RECT 87.560 79.180 88.160 134.430 ;
        RECT 88.350 134.410 89.130 134.430 ;
        RECT 189.240 134.690 189.740 134.700 ;
        RECT 189.240 134.240 190.440 134.690 ;
        RECT 189.240 78.750 189.450 134.240 ;
        RECT 189.660 134.220 190.440 134.240 ;
        RECT 324.090 134.370 325.660 134.800 ;
        RECT 324.090 79.120 324.690 134.370 ;
        RECT 324.880 134.350 325.660 134.370 ;
        RECT 425.770 134.630 426.270 134.640 ;
        RECT 425.770 134.180 426.970 134.630 ;
        RECT 425.770 78.690 425.980 134.180 ;
        RECT 426.190 134.160 426.970 134.180 ;
        RECT 87.410 70.790 88.060 77.510 ;
        RECT 189.210 76.680 189.430 77.090 ;
        RECT 87.410 69.850 88.100 70.790 ;
        RECT 87.500 19.230 88.100 69.850 ;
        RECT 189.220 22.840 189.430 76.680 ;
        RECT 323.940 70.730 324.590 77.450 ;
        RECT 425.740 76.620 425.960 77.030 ;
        RECT 323.940 69.790 324.630 70.730 ;
        RECT 87.400 7.070 88.300 19.230 ;
        RECT 188.920 7.070 189.520 22.840 ;
        RECT 324.030 19.170 324.630 69.790 ;
        RECT 425.750 22.780 425.960 76.620 ;
        RECT 87.250 6.280 189.530 7.070 ;
        RECT 323.930 7.010 324.830 19.170 ;
        RECT 425.450 7.010 426.050 22.780 ;
        RECT 87.250 6.200 96.750 6.280 ;
        RECT 139.240 6.170 189.530 6.280 ;
        RECT 323.780 6.220 426.060 7.010 ;
        RECT 139.240 6.020 160.990 6.170 ;
        RECT 189.040 -1.500 189.340 6.170 ;
        RECT 323.780 6.140 333.280 6.220 ;
        RECT 375.770 6.110 426.060 6.220 ;
        RECT 375.770 5.960 397.520 6.110 ;
        RECT 425.600 2.160 425.910 6.110 ;
        RECT 425.600 0.490 425.950 2.160 ;
        RECT 425.600 0.360 426.010 0.490 ;
        RECT 425.630 0.040 426.010 0.360 ;
        RECT 425.630 -0.020 425.950 0.040 ;
        RECT 425.600 -1.360 425.910 -1.190 ;
        RECT 189.000 -1.520 316.600 -1.500 ;
        RECT 425.600 -1.520 425.970 -1.360 ;
        RECT 189.000 -1.810 425.970 -1.520 ;
        RECT 189.000 -1.830 425.890 -1.810 ;
        RECT 189.000 -1.860 316.600 -1.830 ;
        RECT 189.040 -1.900 189.340 -1.860 ;
      LAYER mcon ;
        RECT 87.760 79.370 87.930 79.540 ;
        RECT 324.290 79.310 324.460 79.480 ;
        RECT 189.270 78.830 189.440 79.000 ;
        RECT 425.800 78.770 425.970 78.940 ;
        RECT 87.660 77.180 87.830 77.350 ;
        RECT 324.190 77.120 324.360 77.290 ;
        RECT 189.240 76.760 189.410 76.930 ;
        RECT 425.770 76.700 425.940 76.870 ;
        RECT 425.710 0.180 425.880 0.350 ;
        RECT 425.670 -1.490 425.840 -1.320 ;
        RECT 193.390 -1.750 193.560 -1.580 ;
        RECT 193.650 -1.750 193.820 -1.580 ;
        RECT 193.900 -1.750 194.070 -1.580 ;
        RECT 194.160 -1.750 194.330 -1.580 ;
      LAYER met1 ;
        RECT 87.410 76.950 88.150 79.740 ;
        RECT 189.210 76.670 189.470 79.100 ;
        RECT 323.940 76.890 324.680 79.680 ;
        RECT 425.740 76.610 426.000 79.040 ;
        RECT 425.610 0.490 425.930 0.630 ;
        RECT 425.610 0.040 426.010 0.490 ;
        RECT 425.610 -1.030 425.930 0.040 ;
        RECT 425.570 -1.360 425.930 -1.030 ;
        RECT 193.315 -15.040 194.435 -1.500 ;
        RECT 425.570 -1.810 425.970 -1.360 ;
        RECT 425.570 -1.890 425.890 -1.810 ;
      LAYER via ;
        RECT 193.450 -14.970 194.295 -14.135 ;
      LAYER met2 ;
        RECT 193.320 -19.465 194.425 -13.995 ;
        RECT 193.520 -25.310 194.100 -19.465 ;
    END
  END d5
  PIN d4
    ANTENNAGATEAREA 2.172000 ;
    PORT
      LAYER li1 ;
        RECT 71.200 198.010 71.790 198.050 ;
        RECT 72.020 198.010 72.800 198.020 ;
        RECT 71.200 197.560 72.800 198.010 ;
        RECT 307.730 197.950 308.320 197.990 ;
        RECT 308.550 197.950 309.330 197.960 ;
        RECT 71.200 197.550 71.790 197.560 ;
        RECT 72.020 197.550 72.800 197.560 ;
        RECT 172.510 197.820 173.100 197.860 ;
        RECT 173.330 197.820 174.110 197.830 ;
        RECT 71.200 165.890 71.430 197.550 ;
        RECT 172.510 197.370 174.110 197.820 ;
        RECT 172.510 197.360 173.100 197.370 ;
        RECT 173.330 197.360 174.110 197.370 ;
        RECT 307.730 197.500 309.330 197.950 ;
        RECT 307.730 197.490 308.320 197.500 ;
        RECT 308.550 197.490 309.330 197.500 ;
        RECT 409.040 197.760 409.630 197.800 ;
        RECT 409.860 197.760 410.640 197.770 ;
        RECT 71.120 165.540 71.530 165.890 ;
        RECT 172.510 165.700 172.740 197.360 ;
        RECT 307.730 165.830 307.960 197.490 ;
        RECT 409.040 197.310 410.640 197.760 ;
        RECT 409.040 197.300 409.630 197.310 ;
        RECT 409.860 197.300 410.640 197.310 ;
        RECT 172.430 165.350 172.840 165.700 ;
        RECT 307.650 165.480 308.060 165.830 ;
        RECT 409.040 165.640 409.270 197.300 ;
        RECT 408.960 165.290 409.370 165.640 ;
        RECT 71.170 163.620 71.580 163.970 ;
        RECT 71.220 110.690 71.450 163.620 ;
        RECT 172.480 163.430 172.890 163.780 ;
        RECT 307.700 163.560 308.110 163.910 ;
        RECT 71.240 109.430 71.440 110.690 ;
        RECT 172.530 110.500 172.760 163.430 ;
        RECT 307.750 110.630 307.980 163.560 ;
        RECT 409.010 163.370 409.420 163.720 ;
        RECT 71.230 109.370 71.440 109.430 ;
        RECT 71.230 107.960 71.430 109.370 ;
        RECT 172.550 109.240 172.750 110.500 ;
        RECT 307.770 109.370 307.970 110.630 ;
        RECT 409.060 110.440 409.290 163.370 ;
        RECT 71.220 107.900 71.430 107.960 ;
        RECT 172.540 109.180 172.750 109.240 ;
        RECT 307.760 109.310 307.970 109.370 ;
        RECT 71.220 105.280 71.420 107.900 ;
        RECT 172.540 107.770 172.740 109.180 ;
        RECT 307.760 107.900 307.960 109.310 ;
        RECT 409.080 109.180 409.280 110.440 ;
        RECT 172.530 107.710 172.740 107.770 ;
        RECT 307.750 107.840 307.960 107.900 ;
        RECT 409.070 109.120 409.280 109.180 ;
        RECT 71.150 104.860 71.540 105.280 ;
        RECT 172.530 105.090 172.730 107.710 ;
        RECT 307.750 105.220 307.950 107.840 ;
        RECT 409.070 107.710 409.270 109.120 ;
        RECT 409.060 107.650 409.270 107.710 ;
        RECT 172.460 104.670 172.850 105.090 ;
        RECT 307.680 104.800 308.070 105.220 ;
        RECT 409.060 105.030 409.260 107.650 ;
        RECT 408.990 104.610 409.380 105.030 ;
        RECT 71.130 103.630 71.520 104.050 ;
        RECT 71.220 101.950 71.420 103.630 ;
        RECT 172.440 103.440 172.830 103.860 ;
        RECT 307.660 103.570 308.050 103.990 ;
        RECT 71.220 101.870 71.440 101.950 ;
        RECT 71.230 77.800 71.440 101.870 ;
        RECT 172.530 101.760 172.730 103.440 ;
        RECT 307.750 101.890 307.950 103.570 ;
        RECT 408.970 103.380 409.360 103.800 ;
        RECT 307.750 101.810 307.970 101.890 ;
        RECT 172.530 101.680 172.750 101.760 ;
        RECT 172.540 77.960 172.750 101.680 ;
        RECT 70.940 77.780 71.620 77.800 ;
        RECT 70.940 77.310 72.300 77.780 ;
        RECT 172.480 77.610 172.750 77.960 ;
        RECT 307.760 77.740 307.970 101.810 ;
        RECT 409.060 101.700 409.260 103.380 ;
        RECT 409.060 101.620 409.280 101.700 ;
        RECT 409.070 77.900 409.280 101.620 ;
        RECT 307.470 77.720 308.150 77.740 ;
        RECT 172.480 77.590 172.930 77.610 ;
        RECT 70.940 77.300 71.570 77.310 ;
        RECT 70.940 77.260 71.480 77.300 ;
        RECT 70.990 58.730 71.430 77.260 ;
        RECT 70.900 52.930 71.430 58.730 ;
        RECT 172.480 77.120 173.610 77.590 ;
        RECT 307.470 77.250 308.830 77.720 ;
        RECT 409.010 77.550 409.280 77.900 ;
        RECT 409.010 77.530 409.460 77.550 ;
        RECT 307.470 77.240 308.100 77.250 ;
        RECT 307.470 77.200 308.010 77.240 ;
        RECT 172.480 77.110 172.880 77.120 ;
        RECT 70.900 49.580 71.340 52.930 ;
        RECT 70.900 46.160 71.380 49.580 ;
        RECT 172.480 49.400 172.700 77.110 ;
        RECT 307.520 58.670 307.960 77.200 ;
        RECT 70.910 45.980 71.380 46.160 ;
        RECT 172.440 48.830 172.700 49.400 ;
        RECT 307.430 52.870 307.960 58.670 ;
        RECT 409.010 77.060 410.140 77.530 ;
        RECT 409.010 77.050 409.410 77.060 ;
        RECT 307.430 49.520 307.870 52.870 ;
        RECT 172.440 45.170 172.690 48.830 ;
        RECT 307.430 46.100 307.910 49.520 ;
        RECT 409.010 49.340 409.230 77.050 ;
        RECT 307.440 45.920 307.910 46.100 ;
        RECT 408.970 48.770 409.230 49.340 ;
        RECT 408.970 45.110 409.220 48.770 ;
        RECT 70.900 32.900 71.340 43.670 ;
        RECT 172.470 43.430 172.690 43.470 ;
        RECT 172.450 43.140 172.690 43.430 ;
        RECT 70.910 32.540 71.320 32.900 ;
        RECT 70.910 31.870 71.470 32.540 ;
        RECT 70.930 17.970 71.470 31.870 ;
        RECT 70.710 16.100 71.470 17.970 ;
        RECT 70.710 4.860 71.320 16.100 ;
        RECT 172.470 14.640 172.690 43.140 ;
        RECT 307.430 32.840 307.870 43.610 ;
        RECT 409.000 43.370 409.220 43.410 ;
        RECT 408.980 43.080 409.220 43.370 ;
        RECT 307.440 32.480 307.850 32.840 ;
        RECT 307.440 31.810 308.000 32.480 ;
        RECT 307.460 17.910 308.000 31.810 ;
        RECT 172.270 14.370 172.690 14.640 ;
        RECT 307.240 16.040 308.000 17.910 ;
        RECT 172.270 13.950 172.740 14.370 ;
        RECT 172.310 11.190 172.740 13.950 ;
        RECT 172.270 10.690 172.740 11.190 ;
        RECT 172.270 7.510 172.700 10.690 ;
        RECT 171.730 5.020 172.030 5.100 ;
        RECT 169.350 4.930 172.630 5.020 ;
        RECT 103.340 4.860 172.630 4.930 ;
        RECT 70.710 4.250 172.630 4.860 ;
        RECT 70.710 4.180 104.170 4.250 ;
        RECT 169.350 4.180 172.630 4.250 ;
        RECT 307.240 4.800 307.850 16.040 ;
        RECT 409.000 14.580 409.220 43.080 ;
        RECT 408.800 14.310 409.220 14.580 ;
        RECT 408.800 13.890 409.270 14.310 ;
        RECT 408.840 11.130 409.270 13.890 ;
        RECT 408.800 10.630 409.270 11.130 ;
        RECT 408.800 7.450 409.230 10.630 ;
        RECT 408.450 4.960 408.940 5.010 ;
        RECT 405.880 4.870 409.160 4.960 ;
        RECT 339.870 4.800 409.160 4.870 ;
        RECT 307.240 4.190 409.160 4.800 ;
        RECT 171.730 -2.210 172.030 4.180 ;
        RECT 307.240 4.120 340.700 4.190 ;
        RECT 405.880 4.120 409.160 4.190 ;
        RECT 408.450 0.260 408.940 4.120 ;
        RECT 408.440 0.040 408.950 0.260 ;
        RECT 408.450 -0.240 408.940 0.040 ;
        RECT 171.750 -2.340 172.030 -2.210 ;
        RECT 408.440 -2.300 408.950 -2.100 ;
        RECT 221.400 -2.320 408.950 -2.300 ;
        RECT 196.500 -2.340 408.940 -2.320 ;
        RECT 171.750 -2.600 408.940 -2.340 ;
        RECT 171.750 -2.620 408.790 -2.600 ;
        RECT 171.750 -2.640 353.950 -2.620 ;
        RECT 171.750 -2.660 221.520 -2.640 ;
        RECT 171.750 -2.670 196.710 -2.660 ;
        RECT 172.240 -2.680 196.710 -2.670 ;
      LAYER mcon ;
        RECT 71.250 165.635 71.420 165.805 ;
        RECT 172.560 165.445 172.730 165.615 ;
        RECT 307.780 165.575 307.950 165.745 ;
        RECT 409.090 165.385 409.260 165.555 ;
        RECT 71.275 163.710 71.445 163.880 ;
        RECT 172.585 163.520 172.755 163.690 ;
        RECT 307.805 163.650 307.975 163.820 ;
        RECT 409.115 163.460 409.285 163.630 ;
        RECT 71.270 105.000 71.440 105.170 ;
        RECT 172.580 104.810 172.750 104.980 ;
        RECT 307.800 104.940 307.970 105.110 ;
        RECT 409.110 104.750 409.280 104.920 ;
        RECT 71.265 103.740 71.435 103.910 ;
        RECT 172.575 103.550 172.745 103.720 ;
        RECT 307.795 103.680 307.965 103.850 ;
        RECT 409.105 103.490 409.275 103.660 ;
        RECT 71.070 46.160 71.240 46.330 ;
        RECT 307.600 46.100 307.770 46.270 ;
        RECT 172.470 45.245 172.640 45.415 ;
        RECT 409.000 45.185 409.170 45.355 ;
        RECT 71.020 43.190 71.190 43.360 ;
        RECT 172.470 43.230 172.640 43.400 ;
        RECT 307.550 43.130 307.720 43.300 ;
        RECT 409.000 43.170 409.170 43.340 ;
        RECT 172.360 7.600 172.530 7.770 ;
        RECT 172.380 4.680 172.550 4.850 ;
        RECT 408.890 7.540 409.060 7.710 ;
        RECT 408.910 4.620 409.080 4.790 ;
        RECT 408.610 -0.090 408.780 0.080 ;
        RECT 175.665 -2.575 175.835 -2.405 ;
        RECT 175.925 -2.575 176.095 -2.405 ;
        RECT 176.175 -2.575 176.345 -2.405 ;
        RECT 176.435 -2.575 176.605 -2.405 ;
        RECT 408.620 -2.480 408.790 -2.310 ;
      LAYER met1 ;
        RECT 71.120 165.540 71.530 165.890 ;
        RECT 71.230 163.970 71.430 165.540 ;
        RECT 172.430 165.350 172.840 165.700 ;
        RECT 307.650 165.480 308.060 165.830 ;
        RECT 71.170 163.620 71.580 163.970 ;
        RECT 172.540 163.780 172.740 165.350 ;
        RECT 307.760 163.910 307.960 165.480 ;
        RECT 408.960 165.290 409.370 165.640 ;
        RECT 71.230 163.590 71.430 163.620 ;
        RECT 172.480 163.430 172.890 163.780 ;
        RECT 307.700 163.560 308.110 163.910 ;
        RECT 409.070 163.720 409.270 165.290 ;
        RECT 307.760 163.530 307.960 163.560 ;
        RECT 172.540 163.400 172.740 163.430 ;
        RECT 409.010 163.370 409.420 163.720 ;
        RECT 409.070 163.340 409.270 163.370 ;
        RECT 71.150 104.860 71.540 105.280 ;
        RECT 71.220 104.050 71.420 104.860 ;
        RECT 172.460 104.670 172.850 105.090 ;
        RECT 307.680 104.800 308.070 105.220 ;
        RECT 71.130 103.630 71.520 104.050 ;
        RECT 172.530 103.860 172.730 104.670 ;
        RECT 307.750 103.990 307.950 104.800 ;
        RECT 408.990 104.610 409.380 105.030 ;
        RECT 172.440 103.440 172.830 103.860 ;
        RECT 307.660 103.570 308.050 103.990 ;
        RECT 409.060 103.800 409.260 104.610 ;
        RECT 408.970 103.380 409.360 103.800 ;
        RECT 70.890 42.960 71.360 46.560 ;
        RECT 172.440 43.130 172.680 45.620 ;
        RECT 307.420 42.900 307.890 46.500 ;
        RECT 408.970 43.070 409.210 45.560 ;
        RECT 172.230 4.220 172.660 7.900 ;
        RECT 408.760 4.160 409.190 7.840 ;
        RECT 408.440 0.210 408.950 0.260 ;
        RECT 408.440 0.040 408.960 0.210 ;
        RECT 175.590 -15.040 176.710 -2.340 ;
        RECT 408.470 -2.670 408.960 0.040 ;
      LAYER via ;
        RECT 175.725 -14.970 176.570 -14.135 ;
      LAYER met2 ;
        RECT 175.595 -19.465 176.700 -13.995 ;
        RECT 175.845 -25.310 176.425 -19.465 ;
    END
  END d4
  PIN d3
    ANTENNAGATEAREA 4.344000 ;
    PORT
      LAYER li1 ;
        RECT 57.640 224.300 58.600 224.310 ;
        RECT 56.940 223.840 58.600 224.300 ;
        RECT 294.170 224.240 295.130 224.250 ;
        RECT 158.950 224.110 159.910 224.120 ;
        RECT 56.940 223.680 57.890 223.840 ;
        RECT 56.940 213.070 57.520 223.680 ;
        RECT 158.250 223.650 159.910 224.110 ;
        RECT 293.470 223.780 295.130 224.240 ;
        RECT 395.480 224.050 396.440 224.060 ;
        RECT 158.250 223.490 159.200 223.650 ;
        RECT 293.470 223.620 294.420 223.780 ;
        RECT 158.250 212.880 158.830 223.490 ;
        RECT 293.470 213.010 294.050 223.620 ;
        RECT 394.780 223.590 396.440 224.050 ;
        RECT 394.780 223.430 395.730 223.590 ;
        RECT 394.780 212.820 395.360 223.430 ;
        RECT 56.780 203.380 57.440 208.150 ;
        RECT 56.780 188.410 57.610 203.380 ;
        RECT 56.950 183.640 57.610 188.410 ;
        RECT 158.090 203.190 158.750 207.960 ;
        RECT 293.310 203.320 293.970 208.090 ;
        RECT 158.090 188.220 158.920 203.190 ;
        RECT 293.310 188.350 294.140 203.320 ;
        RECT 158.260 183.450 158.920 188.220 ;
        RECT 293.480 183.580 294.140 188.350 ;
        RECT 394.620 203.130 395.280 207.900 ;
        RECT 394.620 188.160 395.450 203.130 ;
        RECT 394.790 183.390 395.450 188.160 ;
        RECT 57.020 164.520 57.680 179.750 ;
        RECT 56.240 164.390 57.770 164.520 ;
        RECT 56.240 163.920 58.250 164.390 ;
        RECT 158.330 164.330 158.990 179.560 ;
        RECT 293.550 164.460 294.210 179.690 ;
        RECT 292.770 164.330 294.300 164.460 ;
        RECT 157.550 164.200 159.080 164.330 ;
        RECT 56.240 163.810 57.770 163.920 ;
        RECT 56.240 163.790 57.140 163.810 ;
        RECT 56.240 157.170 56.700 163.790 ;
        RECT 56.330 156.950 56.700 157.170 ;
        RECT 157.550 163.730 159.560 164.200 ;
        RECT 292.770 163.860 294.780 164.330 ;
        RECT 394.860 164.270 395.520 179.500 ;
        RECT 394.080 164.140 395.610 164.270 ;
        RECT 292.770 163.750 294.300 163.860 ;
        RECT 292.770 163.730 293.670 163.750 ;
        RECT 157.550 163.620 159.080 163.730 ;
        RECT 157.550 163.600 158.450 163.620 ;
        RECT 157.550 156.980 158.010 163.600 ;
        RECT 292.770 157.110 293.230 163.730 ;
        RECT 56.330 152.660 56.720 156.950 ;
        RECT 157.640 156.760 158.010 156.980 ;
        RECT 292.860 156.890 293.230 157.110 ;
        RECT 394.080 163.670 396.090 164.140 ;
        RECT 394.080 163.560 395.610 163.670 ;
        RECT 394.080 163.540 394.980 163.560 ;
        RECT 394.080 156.920 394.540 163.540 ;
        RECT 157.640 152.470 158.030 156.760 ;
        RECT 292.860 152.600 293.250 156.890 ;
        RECT 394.170 156.700 394.540 156.920 ;
        RECT 394.170 152.410 394.560 156.700 ;
        RECT 56.360 147.950 56.750 149.800 ;
        RECT 56.360 140.740 56.720 147.950 ;
        RECT 157.670 147.760 158.060 149.610 ;
        RECT 292.890 147.890 293.280 149.740 ;
        RECT 56.360 136.410 56.750 140.740 ;
        RECT 157.670 140.550 158.030 147.760 ;
        RECT 292.890 140.680 293.250 147.890 ;
        RECT 394.200 147.700 394.590 149.550 ;
        RECT 56.360 132.860 56.760 136.410 ;
        RECT 56.350 132.650 56.760 132.860 ;
        RECT 157.670 136.220 158.060 140.550 ;
        RECT 292.890 136.350 293.280 140.680 ;
        RECT 394.200 140.490 394.560 147.700 ;
        RECT 157.670 132.670 158.070 136.220 ;
        RECT 292.890 132.800 293.290 136.350 ;
        RECT 56.340 121.650 56.760 132.650 ;
        RECT 157.660 132.460 158.070 132.670 ;
        RECT 292.880 132.590 293.290 132.800 ;
        RECT 394.200 136.160 394.590 140.490 ;
        RECT 394.200 132.610 394.600 136.160 ;
        RECT 157.650 121.460 158.070 132.460 ;
        RECT 292.870 121.590 293.290 132.590 ;
        RECT 394.190 132.400 394.600 132.610 ;
        RECT 394.180 121.400 394.600 132.400 ;
        RECT 56.380 119.190 56.770 119.230 ;
        RECT 56.380 104.060 56.800 119.190 ;
        RECT 292.910 119.130 293.300 119.170 ;
        RECT 157.690 119.000 158.080 119.040 ;
        RECT 57.140 104.060 58.100 104.070 ;
        RECT 56.380 103.680 58.100 104.060 ;
        RECT 56.440 103.600 58.100 103.680 ;
        RECT 157.690 103.870 158.110 119.000 ;
        RECT 292.910 104.000 293.330 119.130 ;
        RECT 394.220 118.940 394.610 118.980 ;
        RECT 293.670 104.000 294.630 104.010 ;
        RECT 158.450 103.870 159.410 103.880 ;
        RECT 56.440 103.440 57.390 103.600 ;
        RECT 157.690 103.490 159.410 103.870 ;
        RECT 292.910 103.620 294.630 104.000 ;
        RECT 56.440 92.830 57.020 103.440 ;
        RECT 157.750 103.410 159.410 103.490 ;
        RECT 292.970 103.540 294.630 103.620 ;
        RECT 394.220 103.810 394.640 118.940 ;
        RECT 394.980 103.810 395.940 103.820 ;
        RECT 157.750 103.250 158.700 103.410 ;
        RECT 292.970 103.380 293.920 103.540 ;
        RECT 394.220 103.430 395.940 103.810 ;
        RECT 157.750 92.640 158.330 103.250 ;
        RECT 292.970 92.770 293.550 103.380 ;
        RECT 394.280 103.350 395.940 103.430 ;
        RECT 394.280 103.190 395.230 103.350 ;
        RECT 394.280 92.580 394.860 103.190 ;
        RECT 56.280 83.140 56.940 87.910 ;
        RECT 56.280 68.170 57.110 83.140 ;
        RECT 56.450 63.400 57.110 68.170 ;
        RECT 157.590 82.950 158.250 87.720 ;
        RECT 292.810 83.080 293.470 87.850 ;
        RECT 157.590 67.980 158.420 82.950 ;
        RECT 292.810 68.110 293.640 83.080 ;
        RECT 157.760 63.210 158.420 67.980 ;
        RECT 292.980 63.340 293.640 68.110 ;
        RECT 394.120 82.890 394.780 87.660 ;
        RECT 394.120 67.920 394.950 82.890 ;
        RECT 394.290 63.150 394.950 67.920 ;
        RECT 56.520 44.190 57.180 59.510 ;
        RECT 157.830 44.240 158.490 59.320 ;
        RECT 55.430 44.150 57.180 44.190 ;
        RECT 55.430 43.700 57.750 44.150 ;
        RECT 55.450 39.530 55.800 43.700 ;
        RECT 56.790 43.680 57.750 43.700 ;
        RECT 156.300 43.960 158.490 44.240 ;
        RECT 293.050 44.130 293.710 59.450 ;
        RECT 394.360 44.180 395.020 59.260 ;
        RECT 291.960 44.090 293.710 44.130 ;
        RECT 156.300 43.620 159.060 43.960 ;
        RECT 291.960 43.640 294.280 44.090 ;
        RECT 156.300 43.080 156.920 43.620 ;
        RECT 157.830 43.510 159.060 43.620 ;
        RECT 158.100 43.490 159.060 43.510 ;
        RECT 55.410 39.200 55.800 39.530 ;
        RECT 55.410 36.160 55.780 39.200 ;
        RECT 55.380 34.650 55.780 36.160 ;
        RECT 55.380 31.280 55.750 34.650 ;
        RECT 156.350 32.410 156.910 43.080 ;
        RECT 291.980 39.470 292.330 43.640 ;
        RECT 293.320 43.620 294.280 43.640 ;
        RECT 392.830 43.900 395.020 44.180 ;
        RECT 392.830 43.560 395.590 43.900 ;
        RECT 392.830 43.020 393.450 43.560 ;
        RECT 394.360 43.450 395.590 43.560 ;
        RECT 394.630 43.430 395.590 43.450 ;
        RECT 291.940 39.140 292.330 39.470 ;
        RECT 291.940 36.100 292.310 39.140 ;
        RECT 291.910 34.590 292.310 36.100 ;
        RECT 156.270 30.950 156.980 32.410 ;
        RECT 291.910 31.220 292.280 34.590 ;
        RECT 392.880 32.350 393.440 43.020 ;
        RECT 392.800 30.890 393.510 32.350 ;
        RECT 55.320 26.650 55.690 30.080 ;
        RECT 55.310 14.250 55.750 26.650 ;
        RECT 156.460 19.940 156.900 29.520 ;
        RECT 291.850 26.590 292.220 30.020 ;
        RECT 156.420 17.110 156.990 19.940 ;
        RECT 156.420 14.860 157.140 17.110 ;
        RECT 55.280 3.340 55.750 14.250 ;
        RECT 156.500 7.390 157.140 14.860 ;
        RECT 291.840 14.190 292.280 26.590 ;
        RECT 392.990 19.880 393.430 29.460 ;
        RECT 392.950 17.050 393.520 19.880 ;
        RECT 392.950 14.800 393.670 17.050 ;
        RECT 155.520 3.650 155.820 3.670 ;
        RECT 142.180 3.580 157.120 3.650 ;
        RECT 107.480 3.500 157.120 3.580 ;
        RECT 73.110 3.340 157.120 3.500 ;
        RECT 55.280 3.010 157.120 3.340 ;
        RECT 291.810 3.280 292.280 14.190 ;
        RECT 393.030 7.330 393.670 14.800 ;
        RECT 378.710 3.520 393.650 3.590 ;
        RECT 344.010 3.440 393.650 3.520 ;
        RECT 309.640 3.280 393.650 3.440 ;
        RECT 55.280 2.940 143.300 3.010 ;
        RECT 55.280 2.860 108.290 2.940 ;
        RECT 55.280 2.740 73.350 2.860 ;
        RECT 55.720 2.700 73.350 2.740 ;
        RECT 155.520 -3.180 155.820 3.010 ;
        RECT 291.810 2.950 393.650 3.280 ;
        RECT 291.810 2.880 379.830 2.950 ;
        RECT 291.810 2.800 344.820 2.880 ;
        RECT 291.810 2.680 309.880 2.800 ;
        RECT 292.250 2.640 309.880 2.680 ;
        RECT 392.710 0.250 393.190 2.950 ;
        RECT 392.700 -0.190 393.200 0.250 ;
        RECT 392.710 -0.220 393.190 -0.190 ;
        RECT 155.490 -3.220 183.420 -3.180 ;
        RECT 210.820 -3.220 287.110 -3.200 ;
        RECT 155.490 -3.240 325.260 -3.220 ;
        RECT 155.490 -3.300 363.470 -3.240 ;
        RECT 392.710 -3.300 393.190 -3.260 ;
        RECT 155.490 -3.480 393.190 -3.300 ;
        RECT 155.520 -3.520 155.820 -3.480 ;
        RECT 183.230 -3.520 393.190 -3.480 ;
        RECT 210.820 -3.560 393.190 -3.520 ;
        RECT 286.830 -3.580 393.190 -3.560 ;
        RECT 325.040 -3.600 393.190 -3.580 ;
        RECT 392.670 -3.650 393.190 -3.600 ;
      LAYER mcon ;
        RECT 57.080 213.310 57.250 213.480 ;
        RECT 158.390 213.120 158.560 213.290 ;
        RECT 293.610 213.250 293.780 213.420 ;
        RECT 394.920 213.060 395.090 213.230 ;
        RECT 57.120 207.490 57.290 207.660 ;
        RECT 158.430 207.300 158.600 207.470 ;
        RECT 293.650 207.430 293.820 207.600 ;
        RECT 394.960 207.240 395.130 207.410 ;
        RECT 57.250 184.210 57.420 184.380 ;
        RECT 158.560 184.020 158.730 184.190 ;
        RECT 293.780 184.150 293.950 184.320 ;
        RECT 395.090 183.960 395.260 184.130 ;
        RECT 57.250 179.010 57.420 179.180 ;
        RECT 158.560 178.820 158.730 178.990 ;
        RECT 293.780 178.950 293.950 179.120 ;
        RECT 395.090 178.760 395.260 178.930 ;
        RECT 56.505 152.850 56.675 153.020 ;
        RECT 157.815 152.660 157.985 152.830 ;
        RECT 293.035 152.790 293.205 152.960 ;
        RECT 394.345 152.600 394.515 152.770 ;
        RECT 56.415 149.320 56.585 149.490 ;
        RECT 157.725 149.130 157.895 149.300 ;
        RECT 292.945 149.260 293.115 149.430 ;
        RECT 394.255 149.070 394.425 149.240 ;
        RECT 56.455 121.790 56.625 121.960 ;
        RECT 157.765 121.600 157.935 121.770 ;
        RECT 292.985 121.730 293.155 121.900 ;
        RECT 394.295 121.540 394.465 121.710 ;
        RECT 56.525 118.680 56.695 118.850 ;
        RECT 157.835 118.490 158.005 118.660 ;
        RECT 293.055 118.620 293.225 118.790 ;
        RECT 394.365 118.430 394.535 118.600 ;
        RECT 56.580 93.070 56.750 93.240 ;
        RECT 157.890 92.880 158.060 93.050 ;
        RECT 293.110 93.010 293.280 93.180 ;
        RECT 394.420 92.820 394.590 92.990 ;
        RECT 56.620 87.250 56.790 87.420 ;
        RECT 157.930 87.060 158.100 87.230 ;
        RECT 293.150 87.190 293.320 87.360 ;
        RECT 394.460 87.000 394.630 87.170 ;
        RECT 56.750 63.970 56.920 64.140 ;
        RECT 158.060 63.780 158.230 63.950 ;
        RECT 293.280 63.910 293.450 64.080 ;
        RECT 394.590 63.720 394.760 63.890 ;
        RECT 56.750 58.770 56.920 58.940 ;
        RECT 158.060 58.580 158.230 58.750 ;
        RECT 293.280 58.710 293.450 58.880 ;
        RECT 394.590 58.520 394.760 58.690 ;
        RECT 55.485 31.445 55.655 31.615 ;
        RECT 156.580 31.280 156.750 31.450 ;
        RECT 292.015 31.385 292.185 31.555 ;
        RECT 393.110 31.220 393.280 31.390 ;
        RECT 55.355 29.765 55.525 29.935 ;
        RECT 291.885 29.705 292.055 29.875 ;
        RECT 156.610 29.120 156.780 29.290 ;
        RECT 393.140 29.060 393.310 29.230 ;
        RECT 156.765 7.835 156.935 8.005 ;
        RECT 156.665 3.275 156.835 3.445 ;
        RECT 393.295 7.775 393.465 7.945 ;
        RECT 393.195 3.215 393.365 3.385 ;
        RECT 392.850 -0.055 393.020 0.115 ;
        RECT 157.585 -3.415 157.755 -3.245 ;
        RECT 157.845 -3.415 158.015 -3.245 ;
        RECT 158.095 -3.415 158.265 -3.245 ;
        RECT 158.355 -3.415 158.525 -3.245 ;
        RECT 392.870 -3.545 393.040 -3.375 ;
      LAYER met1 ;
        RECT 56.860 207.130 57.400 213.900 ;
        RECT 158.170 206.940 158.710 213.710 ;
        RECT 293.390 207.070 293.930 213.840 ;
        RECT 394.700 206.880 395.240 213.650 ;
        RECT 57.060 178.390 57.600 185.160 ;
        RECT 158.370 178.200 158.910 184.970 ;
        RECT 293.590 178.330 294.130 185.100 ;
        RECT 394.900 178.140 395.440 184.910 ;
        RECT 56.330 150.020 56.720 153.420 ;
        RECT 56.360 149.960 56.720 150.020 ;
        RECT 56.360 148.060 56.750 149.960 ;
        RECT 157.640 149.830 158.030 153.230 ;
        RECT 292.860 149.960 293.250 153.360 ;
        RECT 157.670 149.770 158.030 149.830 ;
        RECT 292.890 149.900 293.250 149.960 ;
        RECT 157.670 147.870 158.060 149.770 ;
        RECT 292.890 148.000 293.280 149.900 ;
        RECT 394.170 149.770 394.560 153.170 ;
        RECT 394.200 149.710 394.560 149.770 ;
        RECT 394.200 147.810 394.590 149.710 ;
        RECT 56.340 121.590 56.810 122.350 ;
        RECT 56.330 119.640 56.810 121.590 ;
        RECT 157.650 121.400 158.120 122.160 ;
        RECT 292.870 121.530 293.340 122.290 ;
        RECT 56.330 119.190 56.770 119.640 ;
        RECT 157.640 119.450 158.120 121.400 ;
        RECT 292.860 119.580 293.340 121.530 ;
        RECT 394.180 121.340 394.650 122.100 ;
        RECT 56.330 118.370 56.800 119.190 ;
        RECT 157.640 119.000 158.080 119.450 ;
        RECT 292.860 119.130 293.300 119.580 ;
        RECT 394.170 119.390 394.650 121.340 ;
        RECT 157.640 118.180 158.110 119.000 ;
        RECT 292.860 118.310 293.330 119.130 ;
        RECT 394.170 118.940 394.610 119.390 ;
        RECT 394.170 118.120 394.640 118.940 ;
        RECT 56.360 86.890 56.900 93.660 ;
        RECT 157.670 86.700 158.210 93.470 ;
        RECT 292.890 86.830 293.430 93.600 ;
        RECT 394.200 86.640 394.740 93.410 ;
        RECT 56.560 58.150 57.100 64.920 ;
        RECT 157.870 57.960 158.410 64.730 ;
        RECT 293.090 58.090 293.630 64.860 ;
        RECT 394.400 57.900 394.940 64.670 ;
        RECT 55.270 29.680 55.700 31.830 ;
        RECT 156.330 28.920 156.950 31.710 ;
        RECT 291.800 29.620 292.230 31.770 ;
        RECT 392.860 28.860 393.480 31.650 ;
        RECT 156.500 3.990 157.140 8.270 ;
        RECT 156.500 3.010 157.120 3.990 ;
        RECT 393.030 3.930 393.670 8.210 ;
        RECT 393.030 2.950 393.650 3.930 ;
        RECT 392.700 -0.190 393.200 0.250 ;
        RECT 157.505 -15.035 158.625 -3.180 ;
        RECT 392.710 -3.460 393.190 -0.190 ;
        RECT 392.700 -3.650 393.190 -3.460 ;
      LAYER via ;
        RECT 157.640 -14.965 158.485 -14.130 ;
      LAYER met2 ;
        RECT 157.510 -19.465 158.615 -13.990 ;
        RECT 157.775 -25.310 158.355 -19.465 ;
    END
  END d3
  PIN d2
    ANTENNAGATEAREA 8.688000 ;
    PORT
      LAYER li1 ;
        RECT 40.290 240.320 41.070 240.330 ;
        RECT 39.860 239.860 41.070 240.320 ;
        RECT 276.820 240.260 277.600 240.270 ;
        RECT 141.600 240.130 142.380 240.140 ;
        RECT 39.890 233.330 40.390 239.860 ;
        RECT 141.170 239.670 142.380 240.130 ;
        RECT 276.390 239.800 277.600 240.260 ;
        RECT 378.130 240.070 378.910 240.080 ;
        RECT 141.200 233.140 141.700 239.670 ;
        RECT 276.420 233.270 276.920 239.800 ;
        RECT 377.700 239.610 378.910 240.070 ;
        RECT 377.730 233.080 378.230 239.610 ;
        RECT 39.840 228.690 40.350 230.910 ;
        RECT 39.800 227.830 40.350 228.690 ;
        RECT 141.150 228.500 141.660 230.720 ;
        RECT 276.370 228.630 276.880 230.850 ;
        RECT 39.800 223.360 40.310 227.830 ;
        RECT 141.110 227.640 141.660 228.500 ;
        RECT 276.330 227.770 276.880 228.630 ;
        RECT 377.680 228.440 378.190 230.660 ;
        RECT 39.800 222.920 40.340 223.360 ;
        RECT 39.830 217.410 40.340 222.920 ;
        RECT 141.110 223.170 141.620 227.640 ;
        RECT 276.330 223.300 276.840 227.770 ;
        RECT 377.640 227.580 378.190 228.440 ;
        RECT 141.110 222.730 141.650 223.170 ;
        RECT 276.330 222.860 276.870 223.300 ;
        RECT 141.140 217.220 141.650 222.730 ;
        RECT 276.360 217.350 276.870 222.860 ;
        RECT 377.640 223.110 378.150 227.580 ;
        RECT 377.640 222.670 378.180 223.110 ;
        RECT 377.670 217.160 378.180 222.670 ;
        RECT 39.840 210.300 40.310 215.390 ;
        RECT 39.720 210.260 40.310 210.300 ;
        RECT 39.720 209.790 41.040 210.260 ;
        RECT 141.150 210.110 141.620 215.200 ;
        RECT 276.370 210.240 276.840 215.330 ;
        RECT 141.030 210.070 141.620 210.110 ;
        RECT 276.250 210.200 276.840 210.240 ;
        RECT 39.720 203.430 40.280 209.790 ;
        RECT 141.030 209.600 142.350 210.070 ;
        RECT 276.250 209.730 277.570 210.200 ;
        RECT 377.680 210.050 378.150 215.140 ;
        RECT 377.560 210.010 378.150 210.050 ;
        RECT 141.030 203.240 141.590 209.600 ;
        RECT 276.250 203.370 276.810 209.730 ;
        RECT 377.560 209.540 378.880 210.010 ;
        RECT 377.560 203.180 378.120 209.540 ;
        RECT 39.380 191.810 40.140 200.550 ;
        RECT 39.420 188.020 39.920 191.810 ;
        RECT 140.690 191.620 141.450 200.360 ;
        RECT 275.910 191.750 276.670 200.490 ;
        RECT 140.730 187.830 141.230 191.620 ;
        RECT 275.950 187.960 276.450 191.750 ;
        RECT 377.220 191.560 377.980 200.300 ;
        RECT 377.260 187.770 377.760 191.560 ;
        RECT 39.480 180.410 39.980 184.750 ;
        RECT 39.480 180.100 40.720 180.410 ;
        RECT 39.510 179.940 40.720 180.100 ;
        RECT 140.790 180.220 141.290 184.560 ;
        RECT 276.010 180.350 276.510 184.690 ;
        RECT 39.540 173.410 40.040 179.940 ;
        RECT 140.790 179.910 142.030 180.220 ;
        RECT 276.010 180.040 277.250 180.350 ;
        RECT 140.820 179.750 142.030 179.910 ;
        RECT 276.040 179.880 277.250 180.040 ;
        RECT 377.320 180.160 377.820 184.500 ;
        RECT 140.850 173.220 141.350 179.750 ;
        RECT 276.070 173.350 276.570 179.880 ;
        RECT 377.320 179.850 378.560 180.160 ;
        RECT 377.350 179.690 378.560 179.850 ;
        RECT 377.380 173.160 377.880 179.690 ;
        RECT 39.490 168.770 40.000 170.990 ;
        RECT 39.450 167.910 40.000 168.770 ;
        RECT 140.800 168.580 141.310 170.800 ;
        RECT 276.020 168.710 276.530 170.930 ;
        RECT 39.450 163.440 39.960 167.910 ;
        RECT 140.760 167.720 141.310 168.580 ;
        RECT 275.980 167.850 276.530 168.710 ;
        RECT 377.330 168.520 377.840 170.740 ;
        RECT 39.450 163.000 39.990 163.440 ;
        RECT 39.480 157.490 39.990 163.000 ;
        RECT 140.760 163.250 141.270 167.720 ;
        RECT 275.980 163.380 276.490 167.850 ;
        RECT 377.290 167.660 377.840 168.520 ;
        RECT 140.760 162.810 141.300 163.250 ;
        RECT 275.980 162.940 276.520 163.380 ;
        RECT 140.790 157.300 141.300 162.810 ;
        RECT 276.010 157.430 276.520 162.940 ;
        RECT 377.290 163.190 377.800 167.660 ;
        RECT 377.290 162.750 377.830 163.190 ;
        RECT 377.320 157.240 377.830 162.750 ;
        RECT 39.490 150.360 39.960 155.470 ;
        RECT 39.120 150.340 39.960 150.360 ;
        RECT 39.120 149.950 40.690 150.340 ;
        RECT 140.800 150.170 141.270 155.280 ;
        RECT 276.020 150.300 276.490 155.410 ;
        RECT 39.130 149.870 40.690 149.950 ;
        RECT 140.430 150.150 141.270 150.170 ;
        RECT 275.650 150.280 276.490 150.300 ;
        RECT 39.130 149.290 39.780 149.870 ;
        RECT 140.430 149.760 142.000 150.150 ;
        RECT 275.650 149.890 277.220 150.280 ;
        RECT 377.330 150.110 377.800 155.220 ;
        RECT 140.440 149.680 142.000 149.760 ;
        RECT 275.660 149.810 277.220 149.890 ;
        RECT 376.960 150.090 377.800 150.110 ;
        RECT 39.110 144.060 39.800 149.290 ;
        RECT 140.440 149.100 141.090 149.680 ;
        RECT 275.660 149.230 276.310 149.810 ;
        RECT 376.960 149.700 378.530 150.090 ;
        RECT 376.970 149.620 378.530 149.700 ;
        RECT 140.420 143.870 141.110 149.100 ;
        RECT 275.640 144.000 276.330 149.230 ;
        RECT 376.970 149.040 377.620 149.620 ;
        RECT 376.950 143.810 377.640 149.040 ;
        RECT 39.220 131.540 39.800 140.650 ;
        RECT 39.220 127.330 39.910 131.540 ;
        RECT 140.530 131.350 141.110 140.460 ;
        RECT 275.750 131.480 276.330 140.590 ;
        RECT 140.530 127.140 141.220 131.350 ;
        RECT 275.750 127.270 276.440 131.480 ;
        RECT 377.060 131.290 377.640 140.400 ;
        RECT 377.060 127.080 377.750 131.290 ;
        RECT 39.320 120.090 39.910 124.930 ;
        RECT 39.320 119.620 40.570 120.090 ;
        RECT 140.630 119.900 141.220 124.740 ;
        RECT 275.850 120.030 276.440 124.870 ;
        RECT 39.320 119.280 39.910 119.620 ;
        RECT 140.630 119.430 141.880 119.900 ;
        RECT 275.850 119.560 277.100 120.030 ;
        RECT 377.160 119.840 377.750 124.680 ;
        RECT 39.390 113.090 39.890 119.280 ;
        RECT 140.630 119.090 141.220 119.430 ;
        RECT 275.850 119.220 276.440 119.560 ;
        RECT 377.160 119.370 378.410 119.840 ;
        RECT 140.700 112.900 141.200 119.090 ;
        RECT 275.920 113.030 276.420 119.220 ;
        RECT 377.160 119.030 377.750 119.370 ;
        RECT 377.230 112.840 377.730 119.030 ;
        RECT 39.340 108.450 39.850 110.670 ;
        RECT 39.300 107.590 39.850 108.450 ;
        RECT 140.650 108.260 141.160 110.480 ;
        RECT 275.870 108.390 276.380 110.610 ;
        RECT 39.300 103.120 39.810 107.590 ;
        RECT 140.610 107.400 141.160 108.260 ;
        RECT 275.830 107.530 276.380 108.390 ;
        RECT 377.180 108.200 377.690 110.420 ;
        RECT 39.300 102.680 39.840 103.120 ;
        RECT 39.330 97.170 39.840 102.680 ;
        RECT 140.610 102.930 141.120 107.400 ;
        RECT 275.830 103.060 276.340 107.530 ;
        RECT 377.140 107.340 377.690 108.200 ;
        RECT 140.610 102.490 141.150 102.930 ;
        RECT 275.830 102.620 276.370 103.060 ;
        RECT 140.640 96.980 141.150 102.490 ;
        RECT 275.860 97.110 276.370 102.620 ;
        RECT 377.140 102.870 377.650 107.340 ;
        RECT 377.140 102.430 377.680 102.870 ;
        RECT 377.170 96.920 377.680 102.430 ;
        RECT 39.340 90.060 39.810 95.150 ;
        RECT 39.220 90.020 39.810 90.060 ;
        RECT 39.220 89.550 40.540 90.020 ;
        RECT 140.650 89.870 141.120 94.960 ;
        RECT 275.870 90.000 276.340 95.090 ;
        RECT 140.530 89.830 141.120 89.870 ;
        RECT 275.750 89.960 276.340 90.000 ;
        RECT 39.220 83.190 39.780 89.550 ;
        RECT 140.530 89.360 141.850 89.830 ;
        RECT 275.750 89.490 277.070 89.960 ;
        RECT 377.180 89.810 377.650 94.900 ;
        RECT 377.060 89.770 377.650 89.810 ;
        RECT 140.530 83.000 141.090 89.360 ;
        RECT 275.750 83.130 276.310 89.490 ;
        RECT 377.060 89.300 378.380 89.770 ;
        RECT 377.060 82.940 377.620 89.300 ;
        RECT 38.880 71.570 39.640 80.310 ;
        RECT 38.920 67.780 39.420 71.570 ;
        RECT 140.190 71.380 140.950 80.120 ;
        RECT 275.410 71.510 276.170 80.250 ;
        RECT 140.230 67.590 140.730 71.380 ;
        RECT 275.450 67.720 275.950 71.510 ;
        RECT 376.720 71.320 377.480 80.060 ;
        RECT 376.760 67.530 377.260 71.320 ;
        RECT 38.980 60.170 39.480 64.510 ;
        RECT 38.980 59.860 40.220 60.170 ;
        RECT 39.010 59.700 40.220 59.860 ;
        RECT 140.290 59.980 140.790 64.320 ;
        RECT 275.510 60.110 276.010 64.450 ;
        RECT 39.040 53.170 39.540 59.700 ;
        RECT 140.290 59.670 141.530 59.980 ;
        RECT 275.510 59.800 276.750 60.110 ;
        RECT 140.320 59.510 141.530 59.670 ;
        RECT 275.540 59.640 276.750 59.800 ;
        RECT 376.820 59.920 377.320 64.260 ;
        RECT 140.350 52.980 140.850 59.510 ;
        RECT 275.570 53.110 276.070 59.640 ;
        RECT 376.820 59.610 378.060 59.920 ;
        RECT 376.850 59.450 378.060 59.610 ;
        RECT 376.880 52.920 377.380 59.450 ;
        RECT 38.990 48.530 39.500 50.750 ;
        RECT 38.950 47.670 39.500 48.530 ;
        RECT 140.300 48.340 140.810 50.560 ;
        RECT 275.520 48.470 276.030 50.690 ;
        RECT 38.950 43.200 39.460 47.670 ;
        RECT 140.260 47.480 140.810 48.340 ;
        RECT 275.480 47.610 276.030 48.470 ;
        RECT 376.830 48.280 377.340 50.500 ;
        RECT 38.950 42.760 39.490 43.200 ;
        RECT 38.980 37.250 39.490 42.760 ;
        RECT 140.260 43.010 140.770 47.480 ;
        RECT 275.480 43.140 275.990 47.610 ;
        RECT 376.790 47.420 377.340 48.280 ;
        RECT 140.260 42.570 140.800 43.010 ;
        RECT 275.480 42.700 276.020 43.140 ;
        RECT 140.290 37.060 140.800 42.570 ;
        RECT 275.510 37.190 276.020 42.700 ;
        RECT 376.790 42.950 377.300 47.420 ;
        RECT 376.790 42.510 377.330 42.950 ;
        RECT 376.820 37.000 377.330 42.510 ;
        RECT 38.990 30.100 39.460 35.230 ;
        RECT 38.990 30.090 40.190 30.100 ;
        RECT 38.980 30.040 40.190 30.090 ;
        RECT 38.680 29.630 40.190 30.040 ;
        RECT 140.300 29.910 140.770 35.040 ;
        RECT 275.520 30.040 275.990 35.170 ;
        RECT 275.520 30.030 276.720 30.040 ;
        RECT 275.510 29.980 276.720 30.030 ;
        RECT 140.300 29.900 141.500 29.910 ;
        RECT 140.290 29.850 141.500 29.900 ;
        RECT 38.680 29.620 39.170 29.630 ;
        RECT 38.690 26.840 38.960 29.620 ;
        RECT 140.140 29.440 141.500 29.850 ;
        RECT 275.210 29.570 276.720 29.980 ;
        RECT 376.830 29.850 377.300 34.980 ;
        RECT 376.830 29.840 378.030 29.850 ;
        RECT 376.820 29.790 378.030 29.840 ;
        RECT 275.210 29.560 275.700 29.570 ;
        RECT 38.670 22.430 38.970 26.840 ;
        RECT 140.140 22.200 140.530 29.440 ;
        RECT 275.220 26.780 275.490 29.560 ;
        RECT 376.670 29.380 378.030 29.790 ;
        RECT 275.200 22.370 275.500 26.780 ;
        RECT 376.670 22.140 377.060 29.380 ;
        RECT 38.670 17.650 38.970 21.080 ;
        RECT 38.600 17.280 38.970 17.650 ;
        RECT 38.600 14.240 38.950 17.280 ;
        RECT 38.440 2.530 39.000 14.240 ;
        RECT 140.090 13.640 140.480 20.660 ;
        RECT 275.200 17.590 275.500 21.020 ;
        RECT 275.130 17.220 275.500 17.590 ;
        RECT 275.130 14.180 275.480 17.220 ;
        RECT 139.820 13.010 140.480 13.640 ;
        RECT 139.820 7.470 140.310 13.010 ;
        RECT 38.320 2.350 39.020 2.530 ;
        RECT 274.970 2.470 275.530 14.180 ;
        RECT 376.620 13.580 377.010 20.600 ;
        RECT 376.350 12.950 377.010 13.580 ;
        RECT 376.350 7.410 376.840 12.950 ;
        RECT 58.040 2.360 59.750 2.400 ;
        RECT 58.040 2.350 124.150 2.360 ;
        RECT 38.320 2.180 124.150 2.350 ;
        RECT 274.850 2.290 275.550 2.470 ;
        RECT 294.570 2.300 296.280 2.340 ;
        RECT 294.570 2.290 360.680 2.300 ;
        RECT 138.550 2.180 138.850 2.200 ;
        RECT 38.320 1.680 140.350 2.180 ;
        RECT 274.850 2.120 360.680 2.290 ;
        RECT 38.320 1.660 124.150 1.680 ;
        RECT 38.320 1.630 58.760 1.660 ;
        RECT 38.320 1.540 39.020 1.630 ;
        RECT 138.550 -4.090 138.850 1.680 ;
        RECT 274.850 1.620 376.880 2.120 ;
        RECT 274.850 1.600 360.680 1.620 ;
        RECT 274.850 1.570 295.290 1.600 ;
        RECT 274.850 1.480 275.550 1.570 ;
        RECT 138.490 -4.110 168.640 -4.090 ;
        RECT 138.490 -4.330 376.820 -4.110 ;
        RECT 138.490 -4.380 376.810 -4.330 ;
        RECT 138.550 -4.430 138.850 -4.380 ;
        RECT 376.450 -4.420 376.810 -4.380 ;
      LAYER mcon ;
        RECT 40.060 233.490 40.230 233.660 ;
        RECT 141.370 233.300 141.540 233.470 ;
        RECT 276.590 233.430 276.760 233.600 ;
        RECT 377.900 233.240 378.070 233.410 ;
        RECT 40.010 230.470 40.180 230.640 ;
        RECT 141.320 230.280 141.490 230.450 ;
        RECT 276.540 230.410 276.710 230.580 ;
        RECT 377.850 230.220 378.020 230.390 ;
        RECT 39.990 217.590 40.160 217.760 ;
        RECT 141.300 217.400 141.470 217.570 ;
        RECT 276.520 217.530 276.690 217.700 ;
        RECT 377.830 217.340 378.000 217.510 ;
        RECT 39.960 214.960 40.130 215.130 ;
        RECT 141.270 214.770 141.440 214.940 ;
        RECT 276.490 214.900 276.660 215.070 ;
        RECT 377.800 214.710 377.970 214.880 ;
        RECT 39.810 203.545 39.980 203.715 ;
        RECT 141.120 203.355 141.290 203.525 ;
        RECT 276.340 203.485 276.510 203.655 ;
        RECT 377.650 203.295 377.820 203.465 ;
        RECT 39.850 199.975 40.020 200.145 ;
        RECT 141.160 199.785 141.330 199.955 ;
        RECT 276.380 199.915 276.550 200.085 ;
        RECT 377.690 199.725 377.860 199.895 ;
        RECT 39.560 188.285 39.730 188.455 ;
        RECT 140.870 188.095 141.040 188.265 ;
        RECT 276.090 188.225 276.260 188.395 ;
        RECT 377.400 188.035 377.570 188.205 ;
        RECT 39.640 184.265 39.810 184.435 ;
        RECT 140.950 184.075 141.120 184.245 ;
        RECT 276.170 184.205 276.340 184.375 ;
        RECT 377.480 184.015 377.650 184.185 ;
        RECT 39.710 173.570 39.880 173.740 ;
        RECT 141.020 173.380 141.190 173.550 ;
        RECT 276.240 173.510 276.410 173.680 ;
        RECT 377.550 173.320 377.720 173.490 ;
        RECT 39.660 170.550 39.830 170.720 ;
        RECT 140.970 170.360 141.140 170.530 ;
        RECT 276.190 170.490 276.360 170.660 ;
        RECT 377.500 170.300 377.670 170.470 ;
        RECT 39.640 157.670 39.810 157.840 ;
        RECT 140.950 157.480 141.120 157.650 ;
        RECT 276.170 157.610 276.340 157.780 ;
        RECT 377.480 157.420 377.650 157.590 ;
        RECT 39.610 155.040 39.780 155.210 ;
        RECT 140.920 154.850 141.090 155.020 ;
        RECT 276.140 154.980 276.310 155.150 ;
        RECT 377.450 154.790 377.620 154.960 ;
        RECT 39.350 144.250 39.520 144.420 ;
        RECT 140.660 144.060 140.830 144.230 ;
        RECT 275.880 144.190 276.050 144.360 ;
        RECT 377.190 144.000 377.360 144.170 ;
        RECT 39.420 140.010 39.590 140.180 ;
        RECT 140.730 139.820 140.900 139.990 ;
        RECT 39.540 127.540 39.710 127.710 ;
        RECT 275.950 139.950 276.120 140.120 ;
        RECT 377.260 139.760 377.430 139.930 ;
        RECT 140.850 127.350 141.020 127.520 ;
        RECT 276.070 127.480 276.240 127.650 ;
        RECT 377.380 127.290 377.550 127.460 ;
        RECT 39.550 124.520 39.720 124.690 ;
        RECT 140.860 124.330 141.030 124.500 ;
        RECT 276.080 124.460 276.250 124.630 ;
        RECT 377.390 124.270 377.560 124.440 ;
        RECT 39.560 113.250 39.730 113.420 ;
        RECT 140.870 113.060 141.040 113.230 ;
        RECT 276.090 113.190 276.260 113.360 ;
        RECT 377.400 113.000 377.570 113.170 ;
        RECT 39.510 110.230 39.680 110.400 ;
        RECT 140.820 110.040 140.990 110.210 ;
        RECT 276.040 110.170 276.210 110.340 ;
        RECT 377.350 109.980 377.520 110.150 ;
        RECT 39.490 97.350 39.660 97.520 ;
        RECT 140.800 97.160 140.970 97.330 ;
        RECT 276.020 97.290 276.190 97.460 ;
        RECT 377.330 97.100 377.500 97.270 ;
        RECT 39.460 94.720 39.630 94.890 ;
        RECT 140.770 94.530 140.940 94.700 ;
        RECT 275.990 94.660 276.160 94.830 ;
        RECT 377.300 94.470 377.470 94.640 ;
        RECT 39.310 83.305 39.480 83.475 ;
        RECT 140.620 83.115 140.790 83.285 ;
        RECT 275.840 83.245 276.010 83.415 ;
        RECT 377.150 83.055 377.320 83.225 ;
        RECT 39.350 79.735 39.520 79.905 ;
        RECT 140.660 79.545 140.830 79.715 ;
        RECT 275.880 79.675 276.050 79.845 ;
        RECT 377.190 79.485 377.360 79.655 ;
        RECT 39.060 68.045 39.230 68.215 ;
        RECT 140.370 67.855 140.540 68.025 ;
        RECT 275.590 67.985 275.760 68.155 ;
        RECT 376.900 67.795 377.070 67.965 ;
        RECT 39.140 64.025 39.310 64.195 ;
        RECT 140.450 63.835 140.620 64.005 ;
        RECT 275.670 63.965 275.840 64.135 ;
        RECT 376.980 63.775 377.150 63.945 ;
        RECT 39.210 53.330 39.380 53.500 ;
        RECT 140.520 53.140 140.690 53.310 ;
        RECT 275.740 53.270 275.910 53.440 ;
        RECT 377.050 53.080 377.220 53.250 ;
        RECT 39.160 50.310 39.330 50.480 ;
        RECT 140.470 50.120 140.640 50.290 ;
        RECT 275.690 50.250 275.860 50.420 ;
        RECT 377.000 50.060 377.170 50.230 ;
        RECT 39.140 37.430 39.310 37.600 ;
        RECT 140.450 37.240 140.620 37.410 ;
        RECT 275.670 37.370 275.840 37.540 ;
        RECT 376.980 37.180 377.150 37.350 ;
        RECT 39.110 34.800 39.280 34.970 ;
        RECT 140.420 34.610 140.590 34.780 ;
        RECT 275.640 34.740 275.810 34.910 ;
        RECT 376.950 34.550 377.120 34.720 ;
        RECT 38.725 22.685 38.895 22.855 ;
        RECT 140.275 22.530 140.445 22.700 ;
        RECT 275.255 22.625 275.425 22.795 ;
        RECT 376.805 22.470 376.975 22.640 ;
        RECT 38.725 20.805 38.895 20.975 ;
        RECT 275.255 20.745 275.425 20.915 ;
        RECT 140.185 20.170 140.355 20.340 ;
        RECT 376.715 20.110 376.885 20.280 ;
        RECT 139.925 7.650 140.095 7.820 ;
        RECT 376.455 7.590 376.625 7.760 ;
        RECT 140.005 1.850 140.175 2.020 ;
        RECT 376.535 1.790 376.705 1.960 ;
        RECT 139.255 -4.315 139.425 -4.145 ;
        RECT 139.515 -4.315 139.685 -4.145 ;
        RECT 139.765 -4.315 139.935 -4.145 ;
        RECT 140.025 -4.315 140.195 -4.145 ;
        RECT 376.555 -4.345 376.725 -4.175 ;
      LAYER met1 ;
        RECT 39.810 230.300 40.380 233.870 ;
        RECT 141.120 230.110 141.690 233.680 ;
        RECT 276.340 230.240 276.910 233.810 ;
        RECT 377.650 230.050 378.220 233.620 ;
        RECT 39.830 217.850 40.350 217.930 ;
        RECT 39.800 217.430 40.350 217.850 ;
        RECT 276.360 217.790 276.880 217.870 ;
        RECT 141.140 217.660 141.660 217.740 ;
        RECT 39.800 214.770 40.310 217.430 ;
        RECT 141.110 217.240 141.660 217.660 ;
        RECT 276.330 217.370 276.880 217.790 ;
        RECT 377.670 217.600 378.190 217.680 ;
        RECT 141.110 214.580 141.620 217.240 ;
        RECT 276.330 214.710 276.840 217.370 ;
        RECT 377.640 217.180 378.190 217.600 ;
        RECT 377.640 214.520 378.150 217.180 ;
        RECT 39.700 199.790 40.200 204.440 ;
        RECT 141.010 199.600 141.510 204.250 ;
        RECT 276.230 199.730 276.730 204.380 ;
        RECT 377.540 199.540 378.040 204.190 ;
        RECT 39.460 184.070 39.960 188.720 ;
        RECT 140.770 183.880 141.270 188.530 ;
        RECT 275.990 184.010 276.490 188.660 ;
        RECT 377.300 183.820 377.800 188.470 ;
        RECT 39.460 170.380 40.030 173.950 ;
        RECT 140.770 170.190 141.340 173.760 ;
        RECT 275.990 170.320 276.560 173.890 ;
        RECT 377.300 170.130 377.870 173.700 ;
        RECT 39.480 157.930 40.000 158.010 ;
        RECT 39.450 157.510 40.000 157.930 ;
        RECT 276.010 157.870 276.530 157.950 ;
        RECT 140.790 157.740 141.310 157.820 ;
        RECT 39.450 154.850 39.960 157.510 ;
        RECT 140.760 157.320 141.310 157.740 ;
        RECT 275.980 157.450 276.530 157.870 ;
        RECT 377.320 157.680 377.840 157.760 ;
        RECT 140.760 154.660 141.270 157.320 ;
        RECT 275.980 154.790 276.490 157.450 ;
        RECT 377.290 157.260 377.840 157.680 ;
        RECT 377.290 154.600 377.800 157.260 ;
        RECT 39.110 139.580 39.800 144.810 ;
        RECT 140.420 139.390 141.110 144.620 ;
        RECT 275.640 139.520 276.330 144.750 ;
        RECT 376.950 139.330 377.640 144.560 ;
        RECT 39.270 123.970 39.960 128.180 ;
        RECT 140.580 123.780 141.270 127.990 ;
        RECT 275.800 123.910 276.490 128.120 ;
        RECT 377.110 123.720 377.800 127.930 ;
        RECT 39.310 110.060 39.880 113.630 ;
        RECT 140.620 109.870 141.190 113.440 ;
        RECT 275.840 110.000 276.410 113.570 ;
        RECT 377.150 109.810 377.720 113.380 ;
        RECT 39.330 97.610 39.850 97.690 ;
        RECT 39.300 97.190 39.850 97.610 ;
        RECT 275.860 97.550 276.380 97.630 ;
        RECT 140.640 97.420 141.160 97.500 ;
        RECT 39.300 94.530 39.810 97.190 ;
        RECT 140.610 97.000 141.160 97.420 ;
        RECT 275.830 97.130 276.380 97.550 ;
        RECT 377.170 97.360 377.690 97.440 ;
        RECT 140.610 94.340 141.120 97.000 ;
        RECT 275.830 94.470 276.340 97.130 ;
        RECT 377.140 96.940 377.690 97.360 ;
        RECT 377.140 94.280 377.650 96.940 ;
        RECT 39.200 79.550 39.700 84.200 ;
        RECT 140.510 79.360 141.010 84.010 ;
        RECT 275.730 79.490 276.230 84.140 ;
        RECT 377.040 79.300 377.540 83.950 ;
        RECT 38.960 63.830 39.460 68.480 ;
        RECT 140.270 63.640 140.770 68.290 ;
        RECT 275.490 63.770 275.990 68.420 ;
        RECT 376.800 63.580 377.300 68.230 ;
        RECT 38.960 50.140 39.530 53.710 ;
        RECT 140.270 49.950 140.840 53.520 ;
        RECT 275.490 50.080 276.060 53.650 ;
        RECT 376.800 49.890 377.370 53.460 ;
        RECT 38.980 37.690 39.500 37.770 ;
        RECT 38.950 37.270 39.500 37.690 ;
        RECT 275.510 37.630 276.030 37.710 ;
        RECT 140.290 37.500 140.810 37.580 ;
        RECT 38.950 34.610 39.460 37.270 ;
        RECT 140.260 37.080 140.810 37.500 ;
        RECT 275.480 37.210 276.030 37.630 ;
        RECT 376.820 37.440 377.340 37.520 ;
        RECT 140.260 34.420 140.770 37.080 ;
        RECT 275.480 34.550 275.990 37.210 ;
        RECT 376.790 37.020 377.340 37.440 ;
        RECT 376.790 34.360 377.300 37.020 ;
        RECT 38.670 20.680 39.010 23.060 ;
        RECT 140.090 20.000 140.530 23.140 ;
        RECT 275.200 20.620 275.540 23.000 ;
        RECT 376.620 19.940 377.060 23.080 ;
        RECT 139.820 7.860 140.300 8.140 ;
        RECT 139.820 7.470 140.320 7.860 ;
        RECT 139.830 1.690 140.320 7.470 ;
        RECT 376.350 7.800 376.830 8.080 ;
        RECT 376.350 7.410 376.850 7.800 ;
        RECT 376.360 1.630 376.850 7.410 ;
        RECT 376.440 -3.900 376.820 1.630 ;
        RECT 139.145 -15.035 140.265 -4.090 ;
        RECT 376.440 -4.110 376.800 -3.900 ;
        RECT 376.440 -4.330 376.820 -4.110 ;
        RECT 376.440 -4.360 376.810 -4.330 ;
        RECT 376.450 -4.420 376.810 -4.360 ;
      LAYER via ;
        RECT 139.280 -14.965 140.125 -14.130 ;
      LAYER met2 ;
        RECT 139.150 -19.465 140.255 -13.990 ;
        RECT 139.380 -25.310 139.960 -19.465 ;
    END
  END d2
  PIN d1
    ANTENNAGATEAREA 17.375999 ;
    PORT
      LAYER li1 ;
        RECT 22.310 245.880 23.480 245.890 ;
        RECT 22.310 245.410 23.490 245.880 ;
        RECT 258.840 245.820 260.010 245.830 ;
        RECT 123.620 245.690 124.790 245.700 ;
        RECT 22.310 245.380 23.480 245.410 ;
        RECT 22.310 243.240 22.810 245.380 ;
        RECT 123.620 245.220 124.800 245.690 ;
        RECT 258.840 245.350 260.020 245.820 ;
        RECT 360.150 245.630 361.320 245.640 ;
        RECT 258.840 245.320 260.010 245.350 ;
        RECT 123.620 245.190 124.790 245.220 ;
        RECT 123.620 243.050 124.120 245.190 ;
        RECT 258.840 243.180 259.340 245.320 ;
        RECT 360.150 245.160 361.330 245.630 ;
        RECT 360.150 245.130 361.320 245.160 ;
        RECT 360.150 242.990 360.650 245.130 ;
        RECT 22.130 235.400 22.790 241.530 ;
        RECT 123.440 235.210 124.100 241.340 ;
        RECT 258.660 235.340 259.320 241.470 ;
        RECT 359.970 235.150 360.630 241.280 ;
        RECT 22.160 231.470 22.660 233.630 ;
        RECT 22.160 231.460 23.310 231.470 ;
        RECT 22.160 230.990 23.320 231.460 ;
        RECT 123.470 231.280 123.970 233.440 ;
        RECT 258.690 231.410 259.190 233.570 ;
        RECT 258.690 231.400 259.840 231.410 ;
        RECT 123.470 231.270 124.620 231.280 ;
        RECT 22.160 230.960 23.310 230.990 ;
        RECT 22.250 230.620 22.590 230.960 ;
        RECT 123.470 230.800 124.630 231.270 ;
        RECT 258.690 230.930 259.850 231.400 ;
        RECT 360.000 231.220 360.500 233.380 ;
        RECT 360.000 231.210 361.150 231.220 ;
        RECT 258.690 230.900 259.840 230.930 ;
        RECT 123.470 230.770 124.620 230.800 ;
        RECT 22.250 230.590 22.610 230.620 ;
        RECT 22.270 228.630 22.610 230.590 ;
        RECT 123.560 230.430 123.900 230.770 ;
        RECT 258.780 230.560 259.120 230.900 ;
        RECT 360.000 230.740 361.160 231.210 ;
        RECT 360.000 230.710 361.150 230.740 ;
        RECT 258.780 230.530 259.140 230.560 ;
        RECT 123.560 230.400 123.920 230.430 ;
        RECT 123.580 228.440 123.920 230.400 ;
        RECT 258.800 228.570 259.140 230.530 ;
        RECT 360.090 230.370 360.430 230.710 ;
        RECT 360.090 230.340 360.450 230.370 ;
        RECT 360.110 228.380 360.450 230.340 ;
        RECT 22.250 225.450 22.590 227.340 ;
        RECT 22.250 220.510 22.600 225.450 ;
        RECT 123.560 225.260 123.900 227.150 ;
        RECT 258.780 225.390 259.120 227.280 ;
        RECT 22.240 220.140 22.630 220.510 ;
        RECT 123.560 220.320 123.910 225.260 ;
        RECT 258.780 220.450 259.130 225.390 ;
        RECT 360.090 225.200 360.430 227.090 ;
        RECT 123.550 219.950 123.940 220.320 ;
        RECT 258.770 220.080 259.160 220.450 ;
        RECT 360.090 220.260 360.440 225.200 ;
        RECT 360.080 219.890 360.470 220.260 ;
        RECT 22.270 215.820 22.620 218.260 ;
        RECT 22.270 215.810 23.450 215.820 ;
        RECT 22.270 215.600 23.460 215.810 ;
        RECT 22.280 215.340 23.460 215.600 ;
        RECT 123.580 215.630 123.930 218.070 ;
        RECT 258.800 215.760 259.150 218.200 ;
        RECT 258.800 215.750 259.980 215.760 ;
        RECT 123.580 215.620 124.760 215.630 ;
        RECT 123.580 215.410 124.770 215.620 ;
        RECT 258.800 215.540 259.990 215.750 ;
        RECT 22.280 215.310 23.450 215.340 ;
        RECT 22.280 213.170 22.780 215.310 ;
        RECT 123.590 215.150 124.770 215.410 ;
        RECT 258.810 215.280 259.990 215.540 ;
        RECT 360.110 215.570 360.460 218.010 ;
        RECT 360.110 215.560 361.290 215.570 ;
        RECT 360.110 215.350 361.300 215.560 ;
        RECT 258.810 215.250 259.980 215.280 ;
        RECT 123.590 215.120 124.760 215.150 ;
        RECT 123.590 212.980 124.090 215.120 ;
        RECT 258.810 213.110 259.310 215.250 ;
        RECT 360.120 215.090 361.300 215.350 ;
        RECT 360.120 215.060 361.290 215.090 ;
        RECT 360.120 212.920 360.620 215.060 ;
        RECT 22.100 205.330 22.760 211.460 ;
        RECT 123.410 205.140 124.070 211.270 ;
        RECT 258.630 205.270 259.290 211.400 ;
        RECT 359.940 205.080 360.600 211.210 ;
        RECT 22.130 201.400 22.630 203.560 ;
        RECT 22.130 201.390 23.280 201.400 ;
        RECT 22.130 201.380 23.290 201.390 ;
        RECT 21.790 200.920 23.290 201.380 ;
        RECT 123.440 201.210 123.940 203.370 ;
        RECT 258.660 201.340 259.160 203.500 ;
        RECT 258.660 201.330 259.810 201.340 ;
        RECT 258.660 201.320 259.820 201.330 ;
        RECT 123.440 201.200 124.590 201.210 ;
        RECT 123.440 201.190 124.600 201.200 ;
        RECT 21.790 200.890 23.280 200.920 ;
        RECT 21.790 200.880 22.500 200.890 ;
        RECT 21.790 198.380 22.240 200.880 ;
        RECT 123.100 200.730 124.600 201.190 ;
        RECT 258.320 200.860 259.820 201.320 ;
        RECT 359.970 201.150 360.470 203.310 ;
        RECT 359.970 201.140 361.120 201.150 ;
        RECT 359.970 201.130 361.130 201.140 ;
        RECT 258.320 200.830 259.810 200.860 ;
        RECT 258.320 200.820 259.030 200.830 ;
        RECT 123.100 200.700 124.590 200.730 ;
        RECT 123.100 200.690 123.810 200.700 ;
        RECT 123.100 198.190 123.550 200.690 ;
        RECT 258.320 198.320 258.770 200.820 ;
        RECT 359.630 200.670 361.130 201.130 ;
        RECT 359.630 200.640 361.120 200.670 ;
        RECT 359.630 200.630 360.340 200.640 ;
        RECT 359.630 198.130 360.080 200.630 ;
        RECT 21.790 195.580 22.240 196.420 ;
        RECT 21.790 193.500 22.280 195.580 ;
        RECT 21.830 190.370 22.280 193.500 ;
        RECT 123.100 195.390 123.550 196.230 ;
        RECT 258.320 195.520 258.770 196.360 ;
        RECT 123.100 193.310 123.590 195.390 ;
        RECT 258.320 193.440 258.810 195.520 ;
        RECT 123.140 190.180 123.590 193.310 ;
        RECT 258.360 190.310 258.810 193.440 ;
        RECT 359.630 195.330 360.080 196.170 ;
        RECT 359.630 193.250 360.120 195.330 ;
        RECT 359.670 190.120 360.120 193.250 ;
        RECT 21.880 185.970 22.330 188.490 ;
        RECT 21.880 185.960 23.130 185.970 ;
        RECT 21.880 185.570 23.140 185.960 ;
        RECT 21.960 185.490 23.140 185.570 ;
        RECT 123.190 185.780 123.640 188.300 ;
        RECT 258.410 185.910 258.860 188.430 ;
        RECT 258.410 185.900 259.660 185.910 ;
        RECT 123.190 185.770 124.440 185.780 ;
        RECT 21.960 185.460 23.130 185.490 ;
        RECT 21.960 183.320 22.460 185.460 ;
        RECT 123.190 185.380 124.450 185.770 ;
        RECT 258.410 185.510 259.670 185.900 ;
        RECT 123.270 185.300 124.450 185.380 ;
        RECT 258.490 185.430 259.670 185.510 ;
        RECT 359.720 185.720 360.170 188.240 ;
        RECT 359.720 185.710 360.970 185.720 ;
        RECT 258.490 185.400 259.660 185.430 ;
        RECT 123.270 185.270 124.440 185.300 ;
        RECT 123.270 183.130 123.770 185.270 ;
        RECT 258.490 183.260 258.990 185.400 ;
        RECT 359.720 185.320 360.980 185.710 ;
        RECT 359.800 185.240 360.980 185.320 ;
        RECT 359.800 185.210 360.970 185.240 ;
        RECT 359.800 183.070 360.300 185.210 ;
        RECT 21.780 175.480 22.440 181.610 ;
        RECT 123.090 175.290 123.750 181.420 ;
        RECT 258.310 175.420 258.970 181.550 ;
        RECT 359.620 175.230 360.280 181.360 ;
        RECT 21.810 171.550 22.310 173.710 ;
        RECT 21.810 171.540 22.960 171.550 ;
        RECT 21.810 171.070 22.970 171.540 ;
        RECT 123.120 171.360 123.620 173.520 ;
        RECT 258.340 171.490 258.840 173.650 ;
        RECT 258.340 171.480 259.490 171.490 ;
        RECT 123.120 171.350 124.270 171.360 ;
        RECT 21.810 171.040 22.960 171.070 ;
        RECT 21.900 170.700 22.240 171.040 ;
        RECT 123.120 170.880 124.280 171.350 ;
        RECT 258.340 171.010 259.500 171.480 ;
        RECT 359.650 171.300 360.150 173.460 ;
        RECT 359.650 171.290 360.800 171.300 ;
        RECT 258.340 170.980 259.490 171.010 ;
        RECT 123.120 170.850 124.270 170.880 ;
        RECT 21.900 170.670 22.260 170.700 ;
        RECT 21.920 168.710 22.260 170.670 ;
        RECT 123.210 170.510 123.550 170.850 ;
        RECT 258.430 170.640 258.770 170.980 ;
        RECT 359.650 170.820 360.810 171.290 ;
        RECT 359.650 170.790 360.800 170.820 ;
        RECT 258.430 170.610 258.790 170.640 ;
        RECT 123.210 170.480 123.570 170.510 ;
        RECT 123.230 168.520 123.570 170.480 ;
        RECT 258.450 168.650 258.790 170.610 ;
        RECT 359.740 170.450 360.080 170.790 ;
        RECT 359.740 170.420 360.100 170.450 ;
        RECT 359.760 168.460 360.100 170.420 ;
        RECT 21.900 165.530 22.240 167.420 ;
        RECT 21.900 160.590 22.250 165.530 ;
        RECT 123.210 165.340 123.550 167.230 ;
        RECT 258.430 165.470 258.770 167.360 ;
        RECT 21.890 160.220 22.280 160.590 ;
        RECT 123.210 160.400 123.560 165.340 ;
        RECT 258.430 160.530 258.780 165.470 ;
        RECT 359.740 165.280 360.080 167.170 ;
        RECT 123.200 160.030 123.590 160.400 ;
        RECT 258.420 160.160 258.810 160.530 ;
        RECT 359.740 160.340 360.090 165.280 ;
        RECT 359.730 159.970 360.120 160.340 ;
        RECT 21.920 155.900 22.270 158.340 ;
        RECT 21.920 155.890 23.100 155.900 ;
        RECT 21.920 155.680 23.110 155.890 ;
        RECT 21.930 155.420 23.110 155.680 ;
        RECT 123.230 155.710 123.580 158.150 ;
        RECT 258.450 155.840 258.800 158.280 ;
        RECT 258.450 155.830 259.630 155.840 ;
        RECT 123.230 155.700 124.410 155.710 ;
        RECT 123.230 155.490 124.420 155.700 ;
        RECT 258.450 155.620 259.640 155.830 ;
        RECT 21.930 155.390 23.100 155.420 ;
        RECT 21.930 153.250 22.430 155.390 ;
        RECT 123.240 155.230 124.420 155.490 ;
        RECT 258.460 155.360 259.640 155.620 ;
        RECT 359.760 155.650 360.110 158.090 ;
        RECT 359.760 155.640 360.940 155.650 ;
        RECT 359.760 155.430 360.950 155.640 ;
        RECT 258.460 155.330 259.630 155.360 ;
        RECT 123.240 155.200 124.410 155.230 ;
        RECT 123.240 153.060 123.740 155.200 ;
        RECT 258.460 153.190 258.960 155.330 ;
        RECT 359.770 155.170 360.950 155.430 ;
        RECT 359.770 155.140 360.940 155.170 ;
        RECT 359.770 153.000 360.270 155.140 ;
        RECT 21.750 145.410 22.410 151.540 ;
        RECT 123.060 145.220 123.720 151.350 ;
        RECT 258.280 145.350 258.940 151.480 ;
        RECT 359.590 145.160 360.250 151.290 ;
        RECT 21.780 141.480 22.280 143.640 ;
        RECT 21.780 141.470 22.930 141.480 ;
        RECT 21.780 141.000 22.940 141.470 ;
        RECT 123.090 141.290 123.590 143.450 ;
        RECT 258.310 141.420 258.810 143.580 ;
        RECT 258.310 141.410 259.460 141.420 ;
        RECT 123.090 141.280 124.240 141.290 ;
        RECT 21.780 140.970 22.930 141.000 ;
        RECT 21.790 138.900 22.160 140.970 ;
        RECT 123.090 140.810 124.250 141.280 ;
        RECT 258.310 140.940 259.470 141.410 ;
        RECT 359.620 141.230 360.120 143.390 ;
        RECT 359.620 141.220 360.770 141.230 ;
        RECT 258.310 140.910 259.460 140.940 ;
        RECT 123.090 140.780 124.240 140.810 ;
        RECT 123.100 138.710 123.470 140.780 ;
        RECT 258.320 138.840 258.690 140.910 ;
        RECT 359.620 140.750 360.780 141.220 ;
        RECT 359.620 140.720 360.770 140.750 ;
        RECT 359.630 138.650 360.000 140.720 ;
        RECT 21.790 130.290 22.210 137.070 ;
        RECT 123.100 130.100 123.520 136.880 ;
        RECT 258.320 130.230 258.740 137.010 ;
        RECT 359.630 130.040 360.050 136.820 ;
        RECT 21.790 125.650 22.210 128.350 ;
        RECT 21.790 125.640 22.980 125.650 ;
        RECT 21.790 125.170 22.990 125.640 ;
        RECT 123.100 125.460 123.520 128.160 ;
        RECT 258.320 125.590 258.740 128.290 ;
        RECT 258.320 125.580 259.510 125.590 ;
        RECT 123.100 125.450 124.290 125.460 ;
        RECT 21.790 125.140 22.980 125.170 ;
        RECT 21.810 123.000 22.310 125.140 ;
        RECT 123.100 124.980 124.300 125.450 ;
        RECT 258.320 125.110 259.520 125.580 ;
        RECT 359.630 125.400 360.050 128.100 ;
        RECT 359.630 125.390 360.820 125.400 ;
        RECT 258.320 125.080 259.510 125.110 ;
        RECT 123.100 124.950 124.290 124.980 ;
        RECT 123.120 122.810 123.620 124.950 ;
        RECT 258.340 122.940 258.840 125.080 ;
        RECT 359.630 124.920 360.830 125.390 ;
        RECT 359.630 124.890 360.820 124.920 ;
        RECT 359.650 122.750 360.150 124.890 ;
        RECT 21.630 115.160 22.290 121.290 ;
        RECT 122.940 114.970 123.600 121.100 ;
        RECT 258.160 115.100 258.820 121.230 ;
        RECT 359.470 114.910 360.130 121.040 ;
        RECT 21.660 111.230 22.160 113.390 ;
        RECT 21.660 111.220 22.810 111.230 ;
        RECT 21.660 110.750 22.820 111.220 ;
        RECT 122.970 111.040 123.470 113.200 ;
        RECT 258.190 111.170 258.690 113.330 ;
        RECT 258.190 111.160 259.340 111.170 ;
        RECT 122.970 111.030 124.120 111.040 ;
        RECT 21.660 110.720 22.810 110.750 ;
        RECT 21.750 110.380 22.090 110.720 ;
        RECT 122.970 110.560 124.130 111.030 ;
        RECT 258.190 110.690 259.350 111.160 ;
        RECT 359.500 110.980 360.000 113.140 ;
        RECT 359.500 110.970 360.650 110.980 ;
        RECT 258.190 110.660 259.340 110.690 ;
        RECT 122.970 110.530 124.120 110.560 ;
        RECT 21.750 110.350 22.110 110.380 ;
        RECT 21.770 108.390 22.110 110.350 ;
        RECT 123.060 110.190 123.400 110.530 ;
        RECT 258.280 110.320 258.620 110.660 ;
        RECT 359.500 110.500 360.660 110.970 ;
        RECT 359.500 110.470 360.650 110.500 ;
        RECT 258.280 110.290 258.640 110.320 ;
        RECT 123.060 110.160 123.420 110.190 ;
        RECT 123.080 108.200 123.420 110.160 ;
        RECT 258.300 108.330 258.640 110.290 ;
        RECT 359.590 110.130 359.930 110.470 ;
        RECT 359.590 110.100 359.950 110.130 ;
        RECT 359.610 108.140 359.950 110.100 ;
        RECT 21.750 105.210 22.090 107.100 ;
        RECT 21.750 100.270 22.100 105.210 ;
        RECT 123.060 105.020 123.400 106.910 ;
        RECT 258.280 105.150 258.620 107.040 ;
        RECT 21.740 99.900 22.130 100.270 ;
        RECT 123.060 100.080 123.410 105.020 ;
        RECT 258.280 100.210 258.630 105.150 ;
        RECT 359.590 104.960 359.930 106.850 ;
        RECT 123.050 99.710 123.440 100.080 ;
        RECT 258.270 99.840 258.660 100.210 ;
        RECT 359.590 100.020 359.940 104.960 ;
        RECT 359.580 99.650 359.970 100.020 ;
        RECT 21.770 95.580 22.120 98.020 ;
        RECT 21.770 95.570 22.950 95.580 ;
        RECT 21.770 95.360 22.960 95.570 ;
        RECT 21.780 95.100 22.960 95.360 ;
        RECT 123.080 95.390 123.430 97.830 ;
        RECT 258.300 95.520 258.650 97.960 ;
        RECT 258.300 95.510 259.480 95.520 ;
        RECT 123.080 95.380 124.260 95.390 ;
        RECT 123.080 95.170 124.270 95.380 ;
        RECT 258.300 95.300 259.490 95.510 ;
        RECT 21.780 95.070 22.950 95.100 ;
        RECT 21.780 92.930 22.280 95.070 ;
        RECT 123.090 94.910 124.270 95.170 ;
        RECT 258.310 95.040 259.490 95.300 ;
        RECT 359.610 95.330 359.960 97.770 ;
        RECT 359.610 95.320 360.790 95.330 ;
        RECT 359.610 95.110 360.800 95.320 ;
        RECT 258.310 95.010 259.480 95.040 ;
        RECT 123.090 94.880 124.260 94.910 ;
        RECT 123.090 92.740 123.590 94.880 ;
        RECT 258.310 92.870 258.810 95.010 ;
        RECT 359.620 94.850 360.800 95.110 ;
        RECT 359.620 94.820 360.790 94.850 ;
        RECT 359.620 92.680 360.120 94.820 ;
        RECT 21.600 85.090 22.260 91.220 ;
        RECT 122.910 84.900 123.570 91.030 ;
        RECT 258.130 85.030 258.790 91.160 ;
        RECT 359.440 84.840 360.100 90.970 ;
        RECT 21.630 81.160 22.130 83.320 ;
        RECT 21.630 81.150 22.780 81.160 ;
        RECT 21.630 81.140 22.790 81.150 ;
        RECT 21.290 80.680 22.790 81.140 ;
        RECT 122.940 80.970 123.440 83.130 ;
        RECT 258.160 81.100 258.660 83.260 ;
        RECT 258.160 81.090 259.310 81.100 ;
        RECT 258.160 81.080 259.320 81.090 ;
        RECT 122.940 80.960 124.090 80.970 ;
        RECT 122.940 80.950 124.100 80.960 ;
        RECT 21.290 80.650 22.780 80.680 ;
        RECT 21.290 80.640 22.000 80.650 ;
        RECT 21.290 78.140 21.740 80.640 ;
        RECT 122.600 80.490 124.100 80.950 ;
        RECT 257.820 80.620 259.320 81.080 ;
        RECT 359.470 80.910 359.970 83.070 ;
        RECT 359.470 80.900 360.620 80.910 ;
        RECT 359.470 80.890 360.630 80.900 ;
        RECT 257.820 80.590 259.310 80.620 ;
        RECT 257.820 80.580 258.530 80.590 ;
        RECT 122.600 80.460 124.090 80.490 ;
        RECT 122.600 80.450 123.310 80.460 ;
        RECT 122.600 77.950 123.050 80.450 ;
        RECT 257.820 78.080 258.270 80.580 ;
        RECT 359.130 80.430 360.630 80.890 ;
        RECT 359.130 80.400 360.620 80.430 ;
        RECT 359.130 80.390 359.840 80.400 ;
        RECT 359.130 77.890 359.580 80.390 ;
        RECT 21.290 75.340 21.740 76.180 ;
        RECT 21.290 73.260 21.780 75.340 ;
        RECT 21.330 70.130 21.780 73.260 ;
        RECT 122.600 75.150 123.050 75.990 ;
        RECT 257.820 75.280 258.270 76.120 ;
        RECT 122.600 73.070 123.090 75.150 ;
        RECT 257.820 73.200 258.310 75.280 ;
        RECT 122.640 69.940 123.090 73.070 ;
        RECT 257.860 70.070 258.310 73.200 ;
        RECT 359.130 75.090 359.580 75.930 ;
        RECT 359.130 73.010 359.620 75.090 ;
        RECT 359.170 69.880 359.620 73.010 ;
        RECT 21.380 65.730 21.830 68.250 ;
        RECT 21.380 65.720 22.630 65.730 ;
        RECT 21.380 65.330 22.640 65.720 ;
        RECT 21.460 65.250 22.640 65.330 ;
        RECT 122.690 65.540 123.140 68.060 ;
        RECT 257.910 65.670 258.360 68.190 ;
        RECT 257.910 65.660 259.160 65.670 ;
        RECT 122.690 65.530 123.940 65.540 ;
        RECT 21.460 65.220 22.630 65.250 ;
        RECT 21.460 63.080 21.960 65.220 ;
        RECT 122.690 65.140 123.950 65.530 ;
        RECT 257.910 65.270 259.170 65.660 ;
        RECT 122.770 65.060 123.950 65.140 ;
        RECT 257.990 65.190 259.170 65.270 ;
        RECT 359.220 65.480 359.670 68.000 ;
        RECT 359.220 65.470 360.470 65.480 ;
        RECT 257.990 65.160 259.160 65.190 ;
        RECT 122.770 65.030 123.940 65.060 ;
        RECT 122.770 62.890 123.270 65.030 ;
        RECT 257.990 63.020 258.490 65.160 ;
        RECT 359.220 65.080 360.480 65.470 ;
        RECT 359.300 65.000 360.480 65.080 ;
        RECT 359.300 64.970 360.470 65.000 ;
        RECT 359.300 62.830 359.800 64.970 ;
        RECT 21.280 55.240 21.940 61.370 ;
        RECT 122.590 55.050 123.250 61.180 ;
        RECT 257.810 55.180 258.470 61.310 ;
        RECT 359.120 54.990 359.780 61.120 ;
        RECT 21.310 51.310 21.810 53.470 ;
        RECT 21.310 51.300 22.460 51.310 ;
        RECT 21.310 50.830 22.470 51.300 ;
        RECT 122.620 51.120 123.120 53.280 ;
        RECT 257.840 51.250 258.340 53.410 ;
        RECT 257.840 51.240 258.990 51.250 ;
        RECT 122.620 51.110 123.770 51.120 ;
        RECT 21.310 50.800 22.460 50.830 ;
        RECT 21.400 50.460 21.740 50.800 ;
        RECT 122.620 50.640 123.780 51.110 ;
        RECT 257.840 50.770 259.000 51.240 ;
        RECT 359.150 51.060 359.650 53.220 ;
        RECT 359.150 51.050 360.300 51.060 ;
        RECT 257.840 50.740 258.990 50.770 ;
        RECT 122.620 50.610 123.770 50.640 ;
        RECT 21.400 50.430 21.760 50.460 ;
        RECT 21.420 48.470 21.760 50.430 ;
        RECT 122.710 50.270 123.050 50.610 ;
        RECT 257.930 50.400 258.270 50.740 ;
        RECT 359.150 50.580 360.310 51.050 ;
        RECT 359.150 50.550 360.300 50.580 ;
        RECT 257.930 50.370 258.290 50.400 ;
        RECT 122.710 50.240 123.070 50.270 ;
        RECT 122.730 48.280 123.070 50.240 ;
        RECT 257.950 48.410 258.290 50.370 ;
        RECT 359.240 50.210 359.580 50.550 ;
        RECT 359.240 50.180 359.600 50.210 ;
        RECT 359.260 48.220 359.600 50.180 ;
        RECT 21.400 45.290 21.740 47.180 ;
        RECT 21.400 40.350 21.750 45.290 ;
        RECT 122.710 45.100 123.050 46.990 ;
        RECT 257.930 45.230 258.270 47.120 ;
        RECT 21.390 39.980 21.780 40.350 ;
        RECT 122.710 40.160 123.060 45.100 ;
        RECT 257.930 40.290 258.280 45.230 ;
        RECT 359.240 45.040 359.580 46.930 ;
        RECT 122.700 39.790 123.090 40.160 ;
        RECT 257.920 39.920 258.310 40.290 ;
        RECT 359.240 40.100 359.590 45.040 ;
        RECT 359.230 39.730 359.620 40.100 ;
        RECT 21.420 35.660 21.770 38.100 ;
        RECT 21.420 35.650 22.600 35.660 ;
        RECT 21.420 35.440 22.610 35.650 ;
        RECT 21.430 35.180 22.610 35.440 ;
        RECT 122.730 35.470 123.080 37.910 ;
        RECT 257.950 35.600 258.300 38.040 ;
        RECT 257.950 35.590 259.130 35.600 ;
        RECT 122.730 35.460 123.910 35.470 ;
        RECT 122.730 35.250 123.920 35.460 ;
        RECT 257.950 35.380 259.140 35.590 ;
        RECT 21.430 35.150 22.600 35.180 ;
        RECT 21.430 33.010 21.930 35.150 ;
        RECT 122.740 34.990 123.920 35.250 ;
        RECT 257.960 35.120 259.140 35.380 ;
        RECT 359.260 35.410 359.610 37.850 ;
        RECT 359.260 35.400 360.440 35.410 ;
        RECT 359.260 35.190 360.450 35.400 ;
        RECT 257.960 35.090 259.130 35.120 ;
        RECT 122.740 34.960 123.910 34.990 ;
        RECT 122.740 32.820 123.240 34.960 ;
        RECT 257.960 32.950 258.460 35.090 ;
        RECT 359.270 34.930 360.450 35.190 ;
        RECT 359.270 34.900 360.440 34.930 ;
        RECT 359.270 32.760 359.770 34.900 ;
        RECT 21.250 25.170 21.910 31.300 ;
        RECT 122.560 24.980 123.220 31.110 ;
        RECT 257.780 25.110 258.440 31.240 ;
        RECT 359.090 24.920 359.750 31.050 ;
        RECT 21.280 21.240 21.780 23.400 ;
        RECT 21.280 21.230 22.430 21.240 ;
        RECT 21.280 20.900 22.440 21.230 ;
        RECT 122.590 21.050 123.090 23.210 ;
        RECT 257.810 21.180 258.310 23.340 ;
        RECT 257.810 21.170 258.960 21.180 ;
        RECT 21.170 20.760 22.440 20.900 ;
        RECT 122.510 21.040 123.740 21.050 ;
        RECT 21.170 20.730 22.430 20.760 ;
        RECT 21.170 18.050 21.460 20.730 ;
        RECT 122.510 20.570 123.750 21.040 ;
        RECT 257.810 20.840 258.970 21.170 ;
        RECT 359.120 20.990 359.620 23.150 ;
        RECT 257.700 20.700 258.970 20.840 ;
        RECT 359.040 20.980 360.270 20.990 ;
        RECT 257.700 20.670 258.960 20.700 ;
        RECT 122.510 20.540 123.740 20.570 ;
        RECT 122.510 18.170 122.940 20.540 ;
        RECT 257.700 17.990 257.990 20.670 ;
        RECT 359.040 20.510 360.280 20.980 ;
        RECT 359.040 20.480 360.270 20.510 ;
        RECT 359.040 18.110 359.470 20.480 ;
        RECT 21.110 16.930 21.480 17.390 ;
        RECT 21.110 16.260 21.460 16.930 ;
        RECT 21.090 15.730 21.460 16.260 ;
        RECT 21.090 15.280 21.360 15.730 ;
        RECT 20.950 12.660 21.360 15.280 ;
        RECT 20.950 12.470 21.350 12.660 ;
        RECT 20.910 2.160 21.350 12.470 ;
        RECT 122.450 11.980 122.880 17.200 ;
        RECT 257.640 16.870 258.010 17.330 ;
        RECT 257.640 16.200 257.990 16.870 ;
        RECT 257.620 15.670 257.990 16.200 ;
        RECT 257.620 15.220 257.890 15.670 ;
        RECT 257.480 12.600 257.890 15.220 ;
        RECT 257.480 12.410 257.880 12.600 ;
        RECT 122.450 7.720 122.750 11.980 ;
        RECT 122.440 7.300 122.750 7.720 ;
        RECT 20.910 0.920 21.310 2.160 ;
        RECT 257.440 2.100 257.880 12.410 ;
        RECT 358.980 11.920 359.410 17.140 ;
        RECT 358.980 7.660 359.280 11.920 ;
        RECT 358.970 7.240 359.280 7.660 ;
        RECT 20.900 0.900 21.500 0.920 ;
        RECT 62.590 0.900 105.080 0.980 ;
        RECT 121.850 0.900 122.150 0.960 ;
        RECT 20.900 0.570 122.760 0.900 ;
        RECT 257.440 0.860 257.840 2.100 ;
        RECT 257.430 0.840 258.030 0.860 ;
        RECT 299.120 0.840 341.610 0.920 ;
        RECT 20.900 0.490 63.250 0.570 ;
        RECT 121.850 -5.130 122.150 0.570 ;
        RECT 257.430 0.510 359.290 0.840 ;
        RECT 257.430 0.430 299.780 0.510 ;
        RECT 358.970 -5.130 359.310 -5.110 ;
        RECT 121.850 -5.310 359.310 -5.130 ;
        RECT 121.850 -5.340 293.130 -5.310 ;
        RECT 121.850 -5.350 197.950 -5.340 ;
        RECT 358.970 -5.360 359.310 -5.310 ;
      LAYER mcon ;
        RECT 22.470 243.445 22.640 243.615 ;
        RECT 123.780 243.255 123.950 243.425 ;
        RECT 259.000 243.385 259.170 243.555 ;
        RECT 360.310 243.195 360.480 243.365 ;
        RECT 22.470 241.265 22.640 241.435 ;
        RECT 22.310 235.535 22.480 235.705 ;
        RECT 123.780 241.075 123.950 241.245 ;
        RECT 123.620 235.345 123.790 235.515 ;
        RECT 259.000 241.205 259.170 241.375 ;
        RECT 258.840 235.475 259.010 235.645 ;
        RECT 360.310 241.015 360.480 241.185 ;
        RECT 360.150 235.285 360.320 235.455 ;
        RECT 22.320 233.385 22.490 233.555 ;
        RECT 123.630 233.195 123.800 233.365 ;
        RECT 258.850 233.325 259.020 233.495 ;
        RECT 360.160 233.135 360.330 233.305 ;
        RECT 22.330 228.695 22.500 228.865 ;
        RECT 123.640 228.505 123.810 228.675 ;
        RECT 258.860 228.635 259.030 228.805 ;
        RECT 360.170 228.445 360.340 228.615 ;
        RECT 22.340 227.055 22.510 227.225 ;
        RECT 123.650 226.865 123.820 227.035 ;
        RECT 258.870 226.995 259.040 227.165 ;
        RECT 360.180 226.805 360.350 226.975 ;
        RECT 22.340 220.245 22.510 220.415 ;
        RECT 123.650 220.055 123.820 220.225 ;
        RECT 258.870 220.185 259.040 220.355 ;
        RECT 360.180 219.995 360.350 220.165 ;
        RECT 22.350 217.995 22.520 218.165 ;
        RECT 123.660 217.805 123.830 217.975 ;
        RECT 258.880 217.935 259.050 218.105 ;
        RECT 360.190 217.745 360.360 217.915 ;
        RECT 22.440 213.375 22.610 213.545 ;
        RECT 123.750 213.185 123.920 213.355 ;
        RECT 258.970 213.315 259.140 213.485 ;
        RECT 360.280 213.125 360.450 213.295 ;
        RECT 22.440 211.195 22.610 211.365 ;
        RECT 22.280 205.465 22.450 205.635 ;
        RECT 123.750 211.005 123.920 211.175 ;
        RECT 123.590 205.275 123.760 205.445 ;
        RECT 258.970 211.135 259.140 211.305 ;
        RECT 258.810 205.405 258.980 205.575 ;
        RECT 360.280 210.945 360.450 211.115 ;
        RECT 360.120 205.215 360.290 205.385 ;
        RECT 22.290 203.315 22.460 203.485 ;
        RECT 123.600 203.125 123.770 203.295 ;
        RECT 258.820 203.255 258.990 203.425 ;
        RECT 360.130 203.065 360.300 203.235 ;
        RECT 21.865 198.510 22.035 198.680 ;
        RECT 123.175 198.320 123.345 198.490 ;
        RECT 258.395 198.450 258.565 198.620 ;
        RECT 359.705 198.260 359.875 198.430 ;
        RECT 21.905 196.020 22.075 196.190 ;
        RECT 123.215 195.830 123.385 196.000 ;
        RECT 258.435 195.960 258.605 196.130 ;
        RECT 359.745 195.770 359.915 195.940 ;
        RECT 21.935 190.570 22.105 190.740 ;
        RECT 123.245 190.380 123.415 190.550 ;
        RECT 258.465 190.510 258.635 190.680 ;
        RECT 359.775 190.320 359.945 190.490 ;
        RECT 21.995 188.120 22.165 188.290 ;
        RECT 123.305 187.930 123.475 188.100 ;
        RECT 258.525 188.060 258.695 188.230 ;
        RECT 359.835 187.870 360.005 188.040 ;
        RECT 22.120 183.525 22.290 183.695 ;
        RECT 123.430 183.335 123.600 183.505 ;
        RECT 258.650 183.465 258.820 183.635 ;
        RECT 359.960 183.275 360.130 183.445 ;
        RECT 22.120 181.345 22.290 181.515 ;
        RECT 21.960 175.615 22.130 175.785 ;
        RECT 123.430 181.155 123.600 181.325 ;
        RECT 123.270 175.425 123.440 175.595 ;
        RECT 258.650 181.285 258.820 181.455 ;
        RECT 258.490 175.555 258.660 175.725 ;
        RECT 359.960 181.095 360.130 181.265 ;
        RECT 359.800 175.365 359.970 175.535 ;
        RECT 21.970 173.465 22.140 173.635 ;
        RECT 123.280 173.275 123.450 173.445 ;
        RECT 258.500 173.405 258.670 173.575 ;
        RECT 359.810 173.215 359.980 173.385 ;
        RECT 21.980 168.775 22.150 168.945 ;
        RECT 123.290 168.585 123.460 168.755 ;
        RECT 258.510 168.715 258.680 168.885 ;
        RECT 359.820 168.525 359.990 168.695 ;
        RECT 21.990 167.135 22.160 167.305 ;
        RECT 123.300 166.945 123.470 167.115 ;
        RECT 258.520 167.075 258.690 167.245 ;
        RECT 359.830 166.885 360.000 167.055 ;
        RECT 21.990 160.325 22.160 160.495 ;
        RECT 123.300 160.135 123.470 160.305 ;
        RECT 258.520 160.265 258.690 160.435 ;
        RECT 359.830 160.075 360.000 160.245 ;
        RECT 22.000 158.075 22.170 158.245 ;
        RECT 123.310 157.885 123.480 158.055 ;
        RECT 258.530 158.015 258.700 158.185 ;
        RECT 359.840 157.825 360.010 157.995 ;
        RECT 22.090 153.455 22.260 153.625 ;
        RECT 123.400 153.265 123.570 153.435 ;
        RECT 258.620 153.395 258.790 153.565 ;
        RECT 359.930 153.205 360.100 153.375 ;
        RECT 22.090 151.275 22.260 151.445 ;
        RECT 21.930 145.545 22.100 145.715 ;
        RECT 123.400 151.085 123.570 151.255 ;
        RECT 123.240 145.355 123.410 145.525 ;
        RECT 258.620 151.215 258.790 151.385 ;
        RECT 258.460 145.485 258.630 145.655 ;
        RECT 359.930 151.025 360.100 151.195 ;
        RECT 359.770 145.295 359.940 145.465 ;
        RECT 21.940 143.395 22.110 143.565 ;
        RECT 123.250 143.205 123.420 143.375 ;
        RECT 258.470 143.335 258.640 143.505 ;
        RECT 359.780 143.145 359.950 143.315 ;
        RECT 21.895 139.045 22.065 139.215 ;
        RECT 123.205 138.855 123.375 139.025 ;
        RECT 258.425 138.985 258.595 139.155 ;
        RECT 359.735 138.795 359.905 138.965 ;
        RECT 21.885 136.755 22.055 136.925 ;
        RECT 21.945 130.575 22.115 130.745 ;
        RECT 123.195 136.565 123.365 136.735 ;
        RECT 123.255 130.385 123.425 130.555 ;
        RECT 258.415 136.695 258.585 136.865 ;
        RECT 258.475 130.515 258.645 130.685 ;
        RECT 359.725 136.505 359.895 136.675 ;
        RECT 359.785 130.325 359.955 130.495 ;
        RECT 21.895 127.985 22.065 128.155 ;
        RECT 123.205 127.795 123.375 127.965 ;
        RECT 258.425 127.925 258.595 128.095 ;
        RECT 359.735 127.735 359.905 127.905 ;
        RECT 21.970 123.205 22.140 123.375 ;
        RECT 123.280 123.015 123.450 123.185 ;
        RECT 258.500 123.145 258.670 123.315 ;
        RECT 359.810 122.955 359.980 123.125 ;
        RECT 21.970 121.025 22.140 121.195 ;
        RECT 21.810 115.295 21.980 115.465 ;
        RECT 123.280 120.835 123.450 121.005 ;
        RECT 123.120 115.105 123.290 115.275 ;
        RECT 258.500 120.965 258.670 121.135 ;
        RECT 258.340 115.235 258.510 115.405 ;
        RECT 359.810 120.775 359.980 120.945 ;
        RECT 359.650 115.045 359.820 115.215 ;
        RECT 21.820 113.145 21.990 113.315 ;
        RECT 123.130 112.955 123.300 113.125 ;
        RECT 258.350 113.085 258.520 113.255 ;
        RECT 359.660 112.895 359.830 113.065 ;
        RECT 21.830 108.455 22.000 108.625 ;
        RECT 123.140 108.265 123.310 108.435 ;
        RECT 258.360 108.395 258.530 108.565 ;
        RECT 359.670 108.205 359.840 108.375 ;
        RECT 21.840 106.815 22.010 106.985 ;
        RECT 123.150 106.625 123.320 106.795 ;
        RECT 258.370 106.755 258.540 106.925 ;
        RECT 359.680 106.565 359.850 106.735 ;
        RECT 21.840 100.005 22.010 100.175 ;
        RECT 123.150 99.815 123.320 99.985 ;
        RECT 258.370 99.945 258.540 100.115 ;
        RECT 359.680 99.755 359.850 99.925 ;
        RECT 21.850 97.755 22.020 97.925 ;
        RECT 123.160 97.565 123.330 97.735 ;
        RECT 258.380 97.695 258.550 97.865 ;
        RECT 359.690 97.505 359.860 97.675 ;
        RECT 21.940 93.135 22.110 93.305 ;
        RECT 123.250 92.945 123.420 93.115 ;
        RECT 258.470 93.075 258.640 93.245 ;
        RECT 359.780 92.885 359.950 93.055 ;
        RECT 21.940 90.955 22.110 91.125 ;
        RECT 21.780 85.225 21.950 85.395 ;
        RECT 123.250 90.765 123.420 90.935 ;
        RECT 123.090 85.035 123.260 85.205 ;
        RECT 258.470 90.895 258.640 91.065 ;
        RECT 258.310 85.165 258.480 85.335 ;
        RECT 359.780 90.705 359.950 90.875 ;
        RECT 359.620 84.975 359.790 85.145 ;
        RECT 21.790 83.075 21.960 83.245 ;
        RECT 123.100 82.885 123.270 83.055 ;
        RECT 258.320 83.015 258.490 83.185 ;
        RECT 359.630 82.825 359.800 82.995 ;
        RECT 21.365 78.270 21.535 78.440 ;
        RECT 122.675 78.080 122.845 78.250 ;
        RECT 257.895 78.210 258.065 78.380 ;
        RECT 359.205 78.020 359.375 78.190 ;
        RECT 21.405 75.780 21.575 75.950 ;
        RECT 122.715 75.590 122.885 75.760 ;
        RECT 257.935 75.720 258.105 75.890 ;
        RECT 359.245 75.530 359.415 75.700 ;
        RECT 21.435 70.330 21.605 70.500 ;
        RECT 122.745 70.140 122.915 70.310 ;
        RECT 257.965 70.270 258.135 70.440 ;
        RECT 359.275 70.080 359.445 70.250 ;
        RECT 21.495 67.880 21.665 68.050 ;
        RECT 122.805 67.690 122.975 67.860 ;
        RECT 258.025 67.820 258.195 67.990 ;
        RECT 359.335 67.630 359.505 67.800 ;
        RECT 21.620 63.285 21.790 63.455 ;
        RECT 122.930 63.095 123.100 63.265 ;
        RECT 258.150 63.225 258.320 63.395 ;
        RECT 359.460 63.035 359.630 63.205 ;
        RECT 21.620 61.105 21.790 61.275 ;
        RECT 21.460 55.375 21.630 55.545 ;
        RECT 122.930 60.915 123.100 61.085 ;
        RECT 122.770 55.185 122.940 55.355 ;
        RECT 258.150 61.045 258.320 61.215 ;
        RECT 257.990 55.315 258.160 55.485 ;
        RECT 359.460 60.855 359.630 61.025 ;
        RECT 359.300 55.125 359.470 55.295 ;
        RECT 21.470 53.225 21.640 53.395 ;
        RECT 122.780 53.035 122.950 53.205 ;
        RECT 258.000 53.165 258.170 53.335 ;
        RECT 359.310 52.975 359.480 53.145 ;
        RECT 21.480 48.535 21.650 48.705 ;
        RECT 122.790 48.345 122.960 48.515 ;
        RECT 258.010 48.475 258.180 48.645 ;
        RECT 359.320 48.285 359.490 48.455 ;
        RECT 21.490 46.895 21.660 47.065 ;
        RECT 122.800 46.705 122.970 46.875 ;
        RECT 258.020 46.835 258.190 47.005 ;
        RECT 359.330 46.645 359.500 46.815 ;
        RECT 21.490 40.085 21.660 40.255 ;
        RECT 122.800 39.895 122.970 40.065 ;
        RECT 258.020 40.025 258.190 40.195 ;
        RECT 359.330 39.835 359.500 40.005 ;
        RECT 21.500 37.835 21.670 38.005 ;
        RECT 122.810 37.645 122.980 37.815 ;
        RECT 258.030 37.775 258.200 37.945 ;
        RECT 359.340 37.585 359.510 37.755 ;
        RECT 21.590 33.215 21.760 33.385 ;
        RECT 122.900 33.025 123.070 33.195 ;
        RECT 258.120 33.155 258.290 33.325 ;
        RECT 359.430 32.965 359.600 33.135 ;
        RECT 21.590 31.035 21.760 31.205 ;
        RECT 21.430 25.305 21.600 25.475 ;
        RECT 122.900 30.845 123.070 31.015 ;
        RECT 122.740 25.115 122.910 25.285 ;
        RECT 258.120 30.975 258.290 31.145 ;
        RECT 257.960 25.245 258.130 25.415 ;
        RECT 359.430 30.785 359.600 30.955 ;
        RECT 359.270 25.055 359.440 25.225 ;
        RECT 21.440 23.155 21.610 23.325 ;
        RECT 122.750 22.965 122.920 23.135 ;
        RECT 257.970 23.095 258.140 23.265 ;
        RECT 359.280 22.905 359.450 23.075 ;
        RECT 21.235 18.120 21.405 18.290 ;
        RECT 122.670 18.305 122.840 18.475 ;
        RECT 257.765 18.060 257.935 18.230 ;
        RECT 359.200 18.245 359.370 18.415 ;
        RECT 21.215 17.170 21.385 17.340 ;
        RECT 122.610 16.685 122.780 16.855 ;
        RECT 257.745 17.110 257.915 17.280 ;
        RECT 359.140 16.625 359.310 16.795 ;
        RECT 122.520 7.465 122.690 7.635 ;
        RECT 359.050 7.405 359.220 7.575 ;
        RECT 122.530 0.685 122.700 0.855 ;
        RECT 359.060 0.625 359.230 0.795 ;
        RECT 123.895 -5.320 124.065 -5.150 ;
        RECT 124.155 -5.320 124.325 -5.150 ;
        RECT 124.405 -5.320 124.575 -5.150 ;
        RECT 124.665 -5.320 124.835 -5.150 ;
        RECT 359.060 -5.310 359.230 -5.140 ;
      LAYER met1 ;
        RECT 22.290 241.140 22.790 243.790 ;
        RECT 123.600 240.950 124.100 243.600 ;
        RECT 258.820 241.080 259.320 243.730 ;
        RECT 360.130 240.890 360.630 243.540 ;
        RECT 22.140 233.170 22.640 235.820 ;
        RECT 123.450 232.980 123.950 235.630 ;
        RECT 258.670 233.110 259.170 235.760 ;
        RECT 359.980 232.920 360.480 235.570 ;
        RECT 22.270 228.940 22.500 229.170 ;
        RECT 22.250 226.950 22.590 228.940 ;
        RECT 123.580 228.750 123.810 228.980 ;
        RECT 258.800 228.880 259.030 229.110 ;
        RECT 123.560 226.760 123.900 228.750 ;
        RECT 258.780 226.890 259.120 228.880 ;
        RECT 360.110 228.690 360.340 228.920 ;
        RECT 360.090 226.700 360.430 228.690 ;
        RECT 22.260 220.510 22.610 220.540 ;
        RECT 22.240 220.140 22.630 220.510 ;
        RECT 258.790 220.450 259.140 220.480 ;
        RECT 123.570 220.320 123.920 220.350 ;
        RECT 22.260 217.880 22.610 220.140 ;
        RECT 123.550 219.950 123.940 220.320 ;
        RECT 258.770 220.080 259.160 220.450 ;
        RECT 360.100 220.260 360.450 220.290 ;
        RECT 123.570 217.690 123.920 219.950 ;
        RECT 258.790 217.820 259.140 220.080 ;
        RECT 360.080 219.890 360.470 220.260 ;
        RECT 360.100 217.630 360.450 219.890 ;
        RECT 22.260 211.070 22.760 213.720 ;
        RECT 123.570 210.880 124.070 213.530 ;
        RECT 258.790 211.010 259.290 213.660 ;
        RECT 360.100 210.820 360.600 213.470 ;
        RECT 22.110 203.100 22.610 205.750 ;
        RECT 123.420 202.910 123.920 205.560 ;
        RECT 258.640 203.040 259.140 205.690 ;
        RECT 359.950 202.850 360.450 205.500 ;
        RECT 21.790 195.870 22.240 198.790 ;
        RECT 123.100 195.680 123.550 198.600 ;
        RECT 258.320 195.810 258.770 198.730 ;
        RECT 359.630 195.620 360.080 198.540 ;
        RECT 21.830 187.950 22.280 190.870 ;
        RECT 123.140 187.760 123.590 190.680 ;
        RECT 258.360 187.890 258.810 190.810 ;
        RECT 359.670 187.700 360.120 190.620 ;
        RECT 21.940 181.220 22.440 183.870 ;
        RECT 123.250 181.030 123.750 183.680 ;
        RECT 258.470 181.160 258.970 183.810 ;
        RECT 359.780 180.970 360.280 183.620 ;
        RECT 21.790 173.250 22.290 175.900 ;
        RECT 123.100 173.060 123.600 175.710 ;
        RECT 258.320 173.190 258.820 175.840 ;
        RECT 359.630 173.000 360.130 175.650 ;
        RECT 21.920 169.020 22.150 169.250 ;
        RECT 21.900 167.030 22.240 169.020 ;
        RECT 123.230 168.830 123.460 169.060 ;
        RECT 258.450 168.960 258.680 169.190 ;
        RECT 123.210 166.840 123.550 168.830 ;
        RECT 258.430 166.970 258.770 168.960 ;
        RECT 359.760 168.770 359.990 169.000 ;
        RECT 359.740 166.780 360.080 168.770 ;
        RECT 21.910 160.590 22.260 160.620 ;
        RECT 21.890 160.220 22.280 160.590 ;
        RECT 258.440 160.530 258.790 160.560 ;
        RECT 123.220 160.400 123.570 160.430 ;
        RECT 21.910 157.960 22.260 160.220 ;
        RECT 123.200 160.030 123.590 160.400 ;
        RECT 258.420 160.160 258.810 160.530 ;
        RECT 359.750 160.340 360.100 160.370 ;
        RECT 123.220 157.770 123.570 160.030 ;
        RECT 258.440 157.900 258.790 160.160 ;
        RECT 359.730 159.970 360.120 160.340 ;
        RECT 359.750 157.710 360.100 159.970 ;
        RECT 21.910 151.150 22.410 153.800 ;
        RECT 123.220 150.960 123.720 153.610 ;
        RECT 258.440 151.090 258.940 153.740 ;
        RECT 359.750 150.900 360.250 153.550 ;
        RECT 21.760 143.180 22.260 145.830 ;
        RECT 123.070 142.990 123.570 145.640 ;
        RECT 258.290 143.120 258.790 145.770 ;
        RECT 359.600 142.930 360.100 145.580 ;
        RECT 21.790 136.490 22.160 139.380 ;
        RECT 123.100 136.300 123.470 139.190 ;
        RECT 258.320 136.430 258.690 139.320 ;
        RECT 359.630 136.240 360.000 139.130 ;
        RECT 21.790 127.790 22.210 131.000 ;
        RECT 123.100 127.600 123.520 130.810 ;
        RECT 258.320 127.730 258.740 130.940 ;
        RECT 359.630 127.540 360.050 130.750 ;
        RECT 21.790 120.900 22.290 123.550 ;
        RECT 123.100 120.710 123.600 123.360 ;
        RECT 258.320 120.840 258.820 123.490 ;
        RECT 359.630 120.650 360.130 123.300 ;
        RECT 21.640 112.930 22.140 115.580 ;
        RECT 122.950 112.740 123.450 115.390 ;
        RECT 258.170 112.870 258.670 115.520 ;
        RECT 359.480 112.680 359.980 115.330 ;
        RECT 21.770 108.700 22.000 108.930 ;
        RECT 21.750 106.710 22.090 108.700 ;
        RECT 123.080 108.510 123.310 108.740 ;
        RECT 258.300 108.640 258.530 108.870 ;
        RECT 123.060 106.520 123.400 108.510 ;
        RECT 258.280 106.650 258.620 108.640 ;
        RECT 359.610 108.450 359.840 108.680 ;
        RECT 359.590 106.460 359.930 108.450 ;
        RECT 21.760 100.270 22.110 100.300 ;
        RECT 21.740 99.900 22.130 100.270 ;
        RECT 258.290 100.210 258.640 100.240 ;
        RECT 123.070 100.080 123.420 100.110 ;
        RECT 21.760 97.640 22.110 99.900 ;
        RECT 123.050 99.710 123.440 100.080 ;
        RECT 258.270 99.840 258.660 100.210 ;
        RECT 359.600 100.020 359.950 100.050 ;
        RECT 123.070 97.450 123.420 99.710 ;
        RECT 258.290 97.580 258.640 99.840 ;
        RECT 359.580 99.650 359.970 100.020 ;
        RECT 359.600 97.390 359.950 99.650 ;
        RECT 21.760 90.830 22.260 93.480 ;
        RECT 123.070 90.640 123.570 93.290 ;
        RECT 258.290 90.770 258.790 93.420 ;
        RECT 359.600 90.580 360.100 93.230 ;
        RECT 21.610 82.860 22.110 85.510 ;
        RECT 122.920 82.670 123.420 85.320 ;
        RECT 258.140 82.800 258.640 85.450 ;
        RECT 359.450 82.610 359.950 85.260 ;
        RECT 21.290 75.630 21.740 78.550 ;
        RECT 122.600 75.440 123.050 78.360 ;
        RECT 257.820 75.570 258.270 78.490 ;
        RECT 359.130 75.380 359.580 78.300 ;
        RECT 21.330 67.710 21.780 70.630 ;
        RECT 122.640 67.520 123.090 70.440 ;
        RECT 257.860 67.650 258.310 70.570 ;
        RECT 359.170 67.460 359.620 70.380 ;
        RECT 21.440 60.980 21.940 63.630 ;
        RECT 122.750 60.790 123.250 63.440 ;
        RECT 257.970 60.920 258.470 63.570 ;
        RECT 359.280 60.730 359.780 63.380 ;
        RECT 21.290 53.010 21.790 55.660 ;
        RECT 122.600 52.820 123.100 55.470 ;
        RECT 257.820 52.950 258.320 55.600 ;
        RECT 359.130 52.760 359.630 55.410 ;
        RECT 21.420 48.780 21.650 49.010 ;
        RECT 21.400 46.790 21.740 48.780 ;
        RECT 122.730 48.590 122.960 48.820 ;
        RECT 257.950 48.720 258.180 48.950 ;
        RECT 122.710 46.600 123.050 48.590 ;
        RECT 257.930 46.730 258.270 48.720 ;
        RECT 359.260 48.530 359.490 48.760 ;
        RECT 359.240 46.540 359.580 48.530 ;
        RECT 21.410 40.350 21.760 40.380 ;
        RECT 21.390 39.980 21.780 40.350 ;
        RECT 257.940 40.290 258.290 40.320 ;
        RECT 122.720 40.160 123.070 40.190 ;
        RECT 21.410 37.720 21.760 39.980 ;
        RECT 122.700 39.790 123.090 40.160 ;
        RECT 257.920 39.920 258.310 40.290 ;
        RECT 359.250 40.100 359.600 40.130 ;
        RECT 122.720 37.530 123.070 39.790 ;
        RECT 257.940 37.660 258.290 39.920 ;
        RECT 359.230 39.730 359.620 40.100 ;
        RECT 359.250 37.470 359.600 39.730 ;
        RECT 21.410 30.910 21.910 33.560 ;
        RECT 122.720 30.720 123.220 33.370 ;
        RECT 257.940 30.850 258.440 33.500 ;
        RECT 359.250 30.660 359.750 33.310 ;
        RECT 21.260 22.940 21.760 25.590 ;
        RECT 122.570 22.750 123.070 25.400 ;
        RECT 257.790 22.880 258.290 25.530 ;
        RECT 359.100 22.690 359.600 25.340 ;
        RECT 21.110 17.100 21.460 18.410 ;
        RECT 122.360 16.560 122.900 18.840 ;
        RECT 257.640 17.040 257.990 18.350 ;
        RECT 358.890 16.500 359.430 18.780 ;
        RECT 122.440 0.650 122.750 7.820 ;
        RECT 122.470 0.550 122.750 0.650 ;
        RECT 358.970 0.860 359.280 7.760 ;
        RECT 358.970 0.590 359.290 0.860 ;
        RECT 123.830 -15.030 124.950 -5.100 ;
        RECT 358.990 -5.110 359.290 0.590 ;
        RECT 358.970 -5.360 359.310 -5.110 ;
      LAYER via ;
        RECT 123.965 -14.960 124.810 -14.125 ;
      LAYER met2 ;
        RECT 123.835 -19.465 124.940 -13.985 ;
        RECT 124.100 -21.310 124.675 -19.465 ;
        RECT 124.095 -25.310 124.675 -21.310 ;
    END
  END d1
  PIN d0
    ANTENNAGATEAREA 34.751999 ;
    PORT
      LAYER li1 ;
        RECT 7.030 248.280 7.810 248.300 ;
        RECT 7.010 247.830 7.810 248.280 ;
        RECT 243.560 248.220 244.340 248.240 ;
        RECT 108.340 248.090 109.120 248.110 ;
        RECT 7.010 247.040 7.250 247.830 ;
        RECT 108.320 247.640 109.120 248.090 ;
        RECT 243.540 247.770 244.340 248.220 ;
        RECT 344.870 248.030 345.650 248.050 ;
        RECT 7.010 245.830 7.260 247.040 ;
        RECT 7.030 245.630 7.260 245.830 ;
        RECT 108.320 246.850 108.560 247.640 ;
        RECT 243.540 246.980 243.780 247.770 ;
        RECT 344.850 247.580 345.650 248.030 ;
        RECT 108.320 245.640 108.570 246.850 ;
        RECT 243.540 245.770 243.790 246.980 ;
        RECT 7.030 245.610 7.250 245.630 ;
        RECT 7.020 245.050 7.250 245.610 ;
        RECT 108.340 245.440 108.570 245.640 ;
        RECT 243.560 245.570 243.790 245.770 ;
        RECT 344.850 246.790 345.090 247.580 ;
        RECT 344.850 245.580 345.100 246.790 ;
        RECT 243.560 245.550 243.780 245.570 ;
        RECT 108.340 245.420 108.560 245.440 ;
        RECT 7.020 244.860 7.260 245.050 ;
        RECT 108.330 244.860 108.560 245.420 ;
        RECT 243.550 244.990 243.780 245.550 ;
        RECT 344.870 245.380 345.100 245.580 ;
        RECT 344.870 245.360 345.090 245.380 ;
        RECT 7.020 244.390 7.250 244.860 ;
        RECT 6.650 244.170 7.250 244.390 ;
        RECT 108.330 244.670 108.570 244.860 ;
        RECT 243.550 244.800 243.790 244.990 ;
        RECT 344.860 244.800 345.090 245.360 ;
        RECT 108.330 244.200 108.560 244.670 ;
        RECT 243.550 244.330 243.780 244.800 ;
        RECT 7.010 241.900 7.250 244.170 ;
        RECT 107.960 243.980 108.560 244.200 ;
        RECT 243.180 244.110 243.780 244.330 ;
        RECT 344.860 244.610 345.100 244.800 ;
        RECT 344.860 244.140 345.090 244.610 ;
        RECT 7.010 241.660 7.970 241.900 ;
        RECT 6.830 241.430 7.970 241.660 ;
        RECT 108.320 241.710 108.560 243.980 ;
        RECT 243.540 241.840 243.780 244.110 ;
        RECT 344.490 243.920 345.090 244.140 ;
        RECT 108.320 241.470 109.280 241.710 ;
        RECT 243.540 241.600 244.500 241.840 ;
        RECT 6.830 239.810 7.310 241.430 ;
        RECT 108.140 241.240 109.280 241.470 ;
        RECT 243.360 241.370 244.500 241.600 ;
        RECT 344.850 241.650 345.090 243.920 ;
        RECT 344.850 241.410 345.810 241.650 ;
        RECT 108.140 239.620 108.620 241.240 ;
        RECT 243.360 239.750 243.840 241.370 ;
        RECT 344.670 241.180 345.810 241.410 ;
        RECT 344.670 239.560 345.150 241.180 ;
        RECT 6.850 235.700 7.310 236.440 ;
        RECT 6.850 233.880 7.330 235.700 ;
        RECT 108.160 235.510 108.620 236.250 ;
        RECT 243.380 235.640 243.840 236.380 ;
        RECT 6.850 233.860 7.640 233.880 ;
        RECT 6.840 233.410 7.640 233.860 ;
        RECT 108.160 233.690 108.640 235.510 ;
        RECT 243.380 233.820 243.860 235.640 ;
        RECT 344.690 235.450 345.150 236.190 ;
        RECT 243.380 233.800 244.170 233.820 ;
        RECT 108.160 233.670 108.950 233.690 ;
        RECT 6.840 232.620 7.080 233.410 ;
        RECT 108.150 233.220 108.950 233.670 ;
        RECT 243.370 233.350 244.170 233.800 ;
        RECT 344.690 233.630 345.170 235.450 ;
        RECT 344.690 233.610 345.480 233.630 ;
        RECT 6.840 231.410 7.090 232.620 ;
        RECT 6.860 231.210 7.090 231.410 ;
        RECT 108.150 232.430 108.390 233.220 ;
        RECT 243.370 232.560 243.610 233.350 ;
        RECT 344.680 233.160 345.480 233.610 ;
        RECT 108.150 231.220 108.400 232.430 ;
        RECT 243.370 231.350 243.620 232.560 ;
        RECT 6.860 231.190 7.080 231.210 ;
        RECT 6.850 230.630 7.080 231.190 ;
        RECT 108.170 231.020 108.400 231.220 ;
        RECT 243.390 231.150 243.620 231.350 ;
        RECT 344.680 232.370 344.920 233.160 ;
        RECT 344.680 231.160 344.930 232.370 ;
        RECT 243.390 231.130 243.610 231.150 ;
        RECT 108.170 231.000 108.390 231.020 ;
        RECT 6.850 230.440 7.090 230.630 ;
        RECT 108.160 230.440 108.390 231.000 ;
        RECT 243.380 230.570 243.610 231.130 ;
        RECT 344.700 230.960 344.930 231.160 ;
        RECT 344.700 230.940 344.920 230.960 ;
        RECT 6.850 229.970 7.080 230.440 ;
        RECT 6.480 229.750 7.080 229.970 ;
        RECT 108.160 230.250 108.400 230.440 ;
        RECT 243.380 230.380 243.620 230.570 ;
        RECT 344.690 230.380 344.920 230.940 ;
        RECT 108.160 229.780 108.390 230.250 ;
        RECT 243.380 229.910 243.610 230.380 ;
        RECT 6.840 227.480 7.080 229.750 ;
        RECT 107.790 229.560 108.390 229.780 ;
        RECT 243.010 229.690 243.610 229.910 ;
        RECT 344.690 230.190 344.930 230.380 ;
        RECT 344.690 229.720 344.920 230.190 ;
        RECT 6.840 227.040 7.800 227.480 ;
        RECT 6.850 227.010 7.800 227.040 ;
        RECT 108.150 227.290 108.390 229.560 ;
        RECT 243.370 227.420 243.610 229.690 ;
        RECT 344.320 229.500 344.920 229.720 ;
        RECT 6.850 225.860 7.070 227.010 ;
        RECT 108.150 226.850 109.110 227.290 ;
        RECT 243.370 226.980 244.330 227.420 ;
        RECT 108.160 226.820 109.110 226.850 ;
        RECT 243.380 226.950 244.330 226.980 ;
        RECT 344.680 227.230 344.920 229.500 ;
        RECT 6.790 225.640 7.110 225.860 ;
        RECT 108.160 225.670 108.380 226.820 ;
        RECT 243.380 225.800 243.600 226.950 ;
        RECT 344.680 226.790 345.640 227.230 ;
        RECT 344.690 226.760 345.640 226.790 ;
        RECT 108.100 225.450 108.420 225.670 ;
        RECT 243.320 225.580 243.640 225.800 ;
        RECT 344.690 225.610 344.910 226.760 ;
        RECT 344.630 225.390 344.950 225.610 ;
        RECT 6.820 224.450 7.140 224.690 ;
        RECT 6.850 222.040 7.080 224.450 ;
        RECT 108.130 224.260 108.450 224.500 ;
        RECT 243.350 224.390 243.670 224.630 ;
        RECT 6.790 221.990 7.170 222.040 ;
        RECT 6.790 221.720 7.180 221.990 ;
        RECT 108.160 221.850 108.390 224.260 ;
        RECT 243.380 221.980 243.610 224.390 ;
        RECT 344.660 224.200 344.980 224.440 ;
        RECT 243.320 221.930 243.700 221.980 ;
        RECT 6.800 221.670 7.180 221.720 ;
        RECT 108.100 221.800 108.480 221.850 ;
        RECT 108.100 221.530 108.490 221.800 ;
        RECT 243.320 221.660 243.710 221.930 ;
        RECT 344.690 221.790 344.920 224.200 ;
        RECT 243.330 221.610 243.710 221.660 ;
        RECT 344.630 221.740 345.010 221.790 ;
        RECT 108.110 221.480 108.490 221.530 ;
        RECT 344.630 221.470 345.020 221.740 ;
        RECT 344.640 221.420 345.020 221.470 ;
        RECT 6.780 220.560 7.150 220.930 ;
        RECT 6.840 219.750 7.070 220.560 ;
        RECT 108.090 220.370 108.460 220.740 ;
        RECT 243.310 220.500 243.680 220.870 ;
        RECT 6.830 218.310 7.080 219.750 ;
        RECT 108.150 219.560 108.380 220.370 ;
        RECT 243.370 219.690 243.600 220.500 ;
        RECT 344.620 220.310 344.990 220.680 ;
        RECT 6.830 218.230 7.210 218.310 ;
        RECT 6.830 218.170 7.780 218.230 ;
        RECT 6.840 217.990 7.780 218.170 ;
        RECT 6.980 217.760 7.780 217.990 ;
        RECT 108.140 218.120 108.390 219.560 ;
        RECT 243.360 218.250 243.610 219.690 ;
        RECT 344.680 219.500 344.910 220.310 ;
        RECT 243.360 218.170 243.740 218.250 ;
        RECT 108.140 218.040 108.520 218.120 ;
        RECT 243.360 218.110 244.310 218.170 ;
        RECT 108.140 217.980 109.090 218.040 ;
        RECT 108.150 217.800 109.090 217.980 ;
        RECT 243.370 217.930 244.310 218.110 ;
        RECT 6.980 216.970 7.220 217.760 ;
        RECT 108.290 217.570 109.090 217.800 ;
        RECT 243.510 217.700 244.310 217.930 ;
        RECT 344.670 218.060 344.920 219.500 ;
        RECT 344.670 217.980 345.050 218.060 ;
        RECT 344.670 217.920 345.620 217.980 ;
        RECT 344.680 217.740 345.620 217.920 ;
        RECT 6.980 215.760 7.230 216.970 ;
        RECT 7.000 215.560 7.230 215.760 ;
        RECT 108.290 216.780 108.530 217.570 ;
        RECT 243.510 216.910 243.750 217.700 ;
        RECT 344.820 217.510 345.620 217.740 ;
        RECT 108.290 215.570 108.540 216.780 ;
        RECT 243.510 215.700 243.760 216.910 ;
        RECT 7.000 215.540 7.220 215.560 ;
        RECT 6.990 214.980 7.220 215.540 ;
        RECT 108.310 215.370 108.540 215.570 ;
        RECT 243.530 215.500 243.760 215.700 ;
        RECT 344.820 216.720 345.060 217.510 ;
        RECT 344.820 215.510 345.070 216.720 ;
        RECT 243.530 215.480 243.750 215.500 ;
        RECT 108.310 215.350 108.530 215.370 ;
        RECT 6.990 214.790 7.230 214.980 ;
        RECT 108.300 214.790 108.530 215.350 ;
        RECT 243.520 214.920 243.750 215.480 ;
        RECT 344.840 215.310 345.070 215.510 ;
        RECT 344.840 215.290 345.060 215.310 ;
        RECT 6.990 214.320 7.220 214.790 ;
        RECT 6.620 214.100 7.220 214.320 ;
        RECT 108.300 214.600 108.540 214.790 ;
        RECT 243.520 214.730 243.760 214.920 ;
        RECT 344.830 214.730 345.060 215.290 ;
        RECT 108.300 214.130 108.530 214.600 ;
        RECT 243.520 214.260 243.750 214.730 ;
        RECT 6.980 211.830 7.220 214.100 ;
        RECT 107.930 213.910 108.530 214.130 ;
        RECT 243.150 214.040 243.750 214.260 ;
        RECT 344.830 214.540 345.070 214.730 ;
        RECT 344.830 214.070 345.060 214.540 ;
        RECT 6.980 211.590 7.940 211.830 ;
        RECT 6.800 211.360 7.940 211.590 ;
        RECT 108.290 211.640 108.530 213.910 ;
        RECT 243.510 211.770 243.750 214.040 ;
        RECT 344.460 213.850 345.060 214.070 ;
        RECT 108.290 211.400 109.250 211.640 ;
        RECT 243.510 211.530 244.470 211.770 ;
        RECT 6.800 209.740 7.280 211.360 ;
        RECT 108.110 211.170 109.250 211.400 ;
        RECT 243.330 211.300 244.470 211.530 ;
        RECT 344.820 211.580 345.060 213.850 ;
        RECT 344.820 211.340 345.780 211.580 ;
        RECT 108.110 209.550 108.590 211.170 ;
        RECT 243.330 209.680 243.810 211.300 ;
        RECT 344.640 211.110 345.780 211.340 ;
        RECT 344.640 209.490 345.120 211.110 ;
        RECT 6.820 205.630 7.280 206.370 ;
        RECT 6.820 203.810 7.300 205.630 ;
        RECT 108.130 205.440 108.590 206.180 ;
        RECT 243.350 205.570 243.810 206.310 ;
        RECT 6.820 203.790 7.610 203.810 ;
        RECT 6.810 203.340 7.610 203.790 ;
        RECT 108.130 203.620 108.610 205.440 ;
        RECT 243.350 203.750 243.830 205.570 ;
        RECT 344.660 205.380 345.120 206.120 ;
        RECT 243.350 203.730 244.140 203.750 ;
        RECT 108.130 203.600 108.920 203.620 ;
        RECT 6.810 202.550 7.050 203.340 ;
        RECT 108.120 203.150 108.920 203.600 ;
        RECT 243.340 203.280 244.140 203.730 ;
        RECT 344.660 203.560 345.140 205.380 ;
        RECT 344.660 203.540 345.450 203.560 ;
        RECT 6.810 201.340 7.060 202.550 ;
        RECT 6.830 201.140 7.060 201.340 ;
        RECT 108.120 202.360 108.360 203.150 ;
        RECT 243.340 202.490 243.580 203.280 ;
        RECT 344.650 203.090 345.450 203.540 ;
        RECT 108.120 201.150 108.370 202.360 ;
        RECT 243.340 201.280 243.590 202.490 ;
        RECT 6.830 201.120 7.050 201.140 ;
        RECT 6.820 200.560 7.050 201.120 ;
        RECT 108.140 200.950 108.370 201.150 ;
        RECT 243.360 201.080 243.590 201.280 ;
        RECT 344.650 202.300 344.890 203.090 ;
        RECT 344.650 201.090 344.900 202.300 ;
        RECT 243.360 201.060 243.580 201.080 ;
        RECT 108.140 200.930 108.360 200.950 ;
        RECT 6.820 200.370 7.060 200.560 ;
        RECT 108.130 200.370 108.360 200.930 ;
        RECT 243.350 200.500 243.580 201.060 ;
        RECT 344.670 200.890 344.900 201.090 ;
        RECT 344.670 200.870 344.890 200.890 ;
        RECT 6.820 199.900 7.050 200.370 ;
        RECT 6.450 199.680 7.050 199.900 ;
        RECT 108.130 200.180 108.370 200.370 ;
        RECT 243.350 200.310 243.590 200.500 ;
        RECT 344.660 200.310 344.890 200.870 ;
        RECT 108.130 199.710 108.360 200.180 ;
        RECT 243.350 199.840 243.580 200.310 ;
        RECT 6.810 197.420 7.050 199.680 ;
        RECT 107.760 199.490 108.360 199.710 ;
        RECT 242.980 199.620 243.580 199.840 ;
        RECT 344.660 200.120 344.900 200.310 ;
        RECT 344.660 199.650 344.890 200.120 ;
        RECT 6.590 197.410 7.050 197.420 ;
        RECT 6.590 196.940 7.770 197.410 ;
        RECT 108.120 197.230 108.360 199.490 ;
        RECT 243.340 197.360 243.580 199.620 ;
        RECT 344.290 199.430 344.890 199.650 ;
        RECT 107.900 197.220 108.360 197.230 ;
        RECT 243.120 197.350 243.580 197.360 ;
        RECT 6.590 195.470 6.930 196.940 ;
        RECT 107.900 196.750 109.080 197.220 ;
        RECT 243.120 196.880 244.300 197.350 ;
        RECT 344.650 197.170 344.890 199.430 ;
        RECT 344.430 197.160 344.890 197.170 ;
        RECT 107.900 195.280 108.240 196.750 ;
        RECT 243.120 195.410 243.460 196.880 ;
        RECT 344.430 196.690 345.610 197.160 ;
        RECT 344.430 195.220 344.770 196.690 ;
        RECT 6.650 192.030 6.990 194.170 ;
        RECT 107.960 191.840 108.300 193.980 ;
        RECT 243.180 191.970 243.520 194.110 ;
        RECT 344.490 191.780 344.830 193.920 ;
        RECT 6.630 188.380 6.990 190.870 ;
        RECT 6.630 188.090 7.460 188.380 ;
        RECT 6.660 187.910 7.460 188.090 ;
        RECT 107.940 188.190 108.300 190.680 ;
        RECT 243.160 188.320 243.520 190.810 ;
        RECT 6.660 187.120 6.900 187.910 ;
        RECT 107.940 187.900 108.770 188.190 ;
        RECT 243.160 188.030 243.990 188.320 ;
        RECT 107.970 187.720 108.770 187.900 ;
        RECT 243.190 187.850 243.990 188.030 ;
        RECT 344.470 188.130 344.830 190.620 ;
        RECT 6.660 185.910 6.910 187.120 ;
        RECT 6.680 185.710 6.910 185.910 ;
        RECT 107.970 186.930 108.210 187.720 ;
        RECT 243.190 187.060 243.430 187.850 ;
        RECT 344.470 187.840 345.300 188.130 ;
        RECT 344.500 187.660 345.300 187.840 ;
        RECT 107.970 185.720 108.220 186.930 ;
        RECT 243.190 185.850 243.440 187.060 ;
        RECT 6.680 185.690 6.900 185.710 ;
        RECT 6.670 185.130 6.900 185.690 ;
        RECT 107.990 185.520 108.220 185.720 ;
        RECT 243.210 185.650 243.440 185.850 ;
        RECT 344.500 186.870 344.740 187.660 ;
        RECT 344.500 185.660 344.750 186.870 ;
        RECT 243.210 185.630 243.430 185.650 ;
        RECT 107.990 185.500 108.210 185.520 ;
        RECT 6.670 184.940 6.910 185.130 ;
        RECT 107.980 184.940 108.210 185.500 ;
        RECT 243.200 185.070 243.430 185.630 ;
        RECT 344.520 185.460 344.750 185.660 ;
        RECT 344.520 185.440 344.740 185.460 ;
        RECT 6.670 184.470 6.900 184.940 ;
        RECT 6.300 184.250 6.900 184.470 ;
        RECT 107.980 184.750 108.220 184.940 ;
        RECT 243.200 184.880 243.440 185.070 ;
        RECT 344.510 184.880 344.740 185.440 ;
        RECT 107.980 184.280 108.210 184.750 ;
        RECT 243.200 184.410 243.430 184.880 ;
        RECT 6.660 181.980 6.900 184.250 ;
        RECT 107.610 184.060 108.210 184.280 ;
        RECT 242.830 184.190 243.430 184.410 ;
        RECT 344.510 184.690 344.750 184.880 ;
        RECT 344.510 184.220 344.740 184.690 ;
        RECT 6.660 181.740 7.620 181.980 ;
        RECT 6.480 181.510 7.620 181.740 ;
        RECT 107.970 181.790 108.210 184.060 ;
        RECT 243.190 181.920 243.430 184.190 ;
        RECT 344.140 184.000 344.740 184.220 ;
        RECT 107.970 181.550 108.930 181.790 ;
        RECT 243.190 181.680 244.150 181.920 ;
        RECT 6.480 179.890 6.960 181.510 ;
        RECT 107.790 181.320 108.930 181.550 ;
        RECT 243.010 181.450 244.150 181.680 ;
        RECT 344.500 181.730 344.740 184.000 ;
        RECT 344.500 181.490 345.460 181.730 ;
        RECT 107.790 179.700 108.270 181.320 ;
        RECT 243.010 179.830 243.490 181.450 ;
        RECT 344.320 181.260 345.460 181.490 ;
        RECT 344.320 179.640 344.800 181.260 ;
        RECT 6.500 175.780 6.960 176.520 ;
        RECT 6.500 173.960 6.980 175.780 ;
        RECT 107.810 175.590 108.270 176.330 ;
        RECT 243.030 175.720 243.490 176.460 ;
        RECT 6.500 173.940 7.290 173.960 ;
        RECT 6.490 173.490 7.290 173.940 ;
        RECT 107.810 173.770 108.290 175.590 ;
        RECT 243.030 173.900 243.510 175.720 ;
        RECT 344.340 175.530 344.800 176.270 ;
        RECT 243.030 173.880 243.820 173.900 ;
        RECT 107.810 173.750 108.600 173.770 ;
        RECT 6.490 172.700 6.730 173.490 ;
        RECT 107.800 173.300 108.600 173.750 ;
        RECT 243.020 173.430 243.820 173.880 ;
        RECT 344.340 173.710 344.820 175.530 ;
        RECT 344.340 173.690 345.130 173.710 ;
        RECT 6.490 171.490 6.740 172.700 ;
        RECT 6.510 171.290 6.740 171.490 ;
        RECT 107.800 172.510 108.040 173.300 ;
        RECT 243.020 172.640 243.260 173.430 ;
        RECT 344.330 173.240 345.130 173.690 ;
        RECT 107.800 171.300 108.050 172.510 ;
        RECT 243.020 171.430 243.270 172.640 ;
        RECT 6.510 171.270 6.730 171.290 ;
        RECT 6.500 170.710 6.730 171.270 ;
        RECT 107.820 171.100 108.050 171.300 ;
        RECT 243.040 171.230 243.270 171.430 ;
        RECT 344.330 172.450 344.570 173.240 ;
        RECT 344.330 171.240 344.580 172.450 ;
        RECT 243.040 171.210 243.260 171.230 ;
        RECT 107.820 171.080 108.040 171.100 ;
        RECT 6.500 170.520 6.740 170.710 ;
        RECT 107.810 170.520 108.040 171.080 ;
        RECT 243.030 170.650 243.260 171.210 ;
        RECT 344.350 171.040 344.580 171.240 ;
        RECT 344.350 171.020 344.570 171.040 ;
        RECT 6.500 170.050 6.730 170.520 ;
        RECT 6.130 169.830 6.730 170.050 ;
        RECT 107.810 170.330 108.050 170.520 ;
        RECT 243.030 170.460 243.270 170.650 ;
        RECT 344.340 170.460 344.570 171.020 ;
        RECT 107.810 169.860 108.040 170.330 ;
        RECT 243.030 169.990 243.260 170.460 ;
        RECT 6.490 167.560 6.730 169.830 ;
        RECT 107.440 169.640 108.040 169.860 ;
        RECT 242.660 169.770 243.260 169.990 ;
        RECT 344.340 170.270 344.580 170.460 ;
        RECT 344.340 169.800 344.570 170.270 ;
        RECT 6.490 167.120 7.450 167.560 ;
        RECT 6.500 167.090 7.450 167.120 ;
        RECT 107.800 167.370 108.040 169.640 ;
        RECT 243.020 167.500 243.260 169.770 ;
        RECT 343.970 169.580 344.570 169.800 ;
        RECT 6.500 165.940 6.720 167.090 ;
        RECT 107.800 166.930 108.760 167.370 ;
        RECT 243.020 167.060 243.980 167.500 ;
        RECT 107.810 166.900 108.760 166.930 ;
        RECT 243.030 167.030 243.980 167.060 ;
        RECT 344.330 167.310 344.570 169.580 ;
        RECT 6.440 165.720 6.760 165.940 ;
        RECT 107.810 165.750 108.030 166.900 ;
        RECT 243.030 165.880 243.250 167.030 ;
        RECT 344.330 166.870 345.290 167.310 ;
        RECT 344.340 166.840 345.290 166.870 ;
        RECT 107.750 165.530 108.070 165.750 ;
        RECT 242.970 165.660 243.290 165.880 ;
        RECT 344.340 165.690 344.560 166.840 ;
        RECT 344.280 165.470 344.600 165.690 ;
        RECT 6.470 164.530 6.790 164.770 ;
        RECT 6.500 162.120 6.730 164.530 ;
        RECT 107.780 164.340 108.100 164.580 ;
        RECT 243.000 164.470 243.320 164.710 ;
        RECT 6.440 162.070 6.820 162.120 ;
        RECT 6.440 161.800 6.830 162.070 ;
        RECT 107.810 161.930 108.040 164.340 ;
        RECT 243.030 162.060 243.260 164.470 ;
        RECT 344.310 164.280 344.630 164.520 ;
        RECT 242.970 162.010 243.350 162.060 ;
        RECT 6.450 161.750 6.830 161.800 ;
        RECT 107.750 161.880 108.130 161.930 ;
        RECT 107.750 161.610 108.140 161.880 ;
        RECT 242.970 161.740 243.360 162.010 ;
        RECT 344.340 161.870 344.570 164.280 ;
        RECT 242.980 161.690 243.360 161.740 ;
        RECT 344.280 161.820 344.660 161.870 ;
        RECT 107.760 161.560 108.140 161.610 ;
        RECT 344.280 161.550 344.670 161.820 ;
        RECT 344.290 161.500 344.670 161.550 ;
        RECT 6.430 160.640 6.800 161.010 ;
        RECT 6.490 159.830 6.720 160.640 ;
        RECT 107.740 160.450 108.110 160.820 ;
        RECT 242.960 160.580 243.330 160.950 ;
        RECT 6.480 158.390 6.730 159.830 ;
        RECT 107.800 159.640 108.030 160.450 ;
        RECT 243.020 159.770 243.250 160.580 ;
        RECT 344.270 160.390 344.640 160.760 ;
        RECT 6.480 158.310 6.860 158.390 ;
        RECT 6.480 158.250 7.430 158.310 ;
        RECT 6.490 158.070 7.430 158.250 ;
        RECT 6.630 157.840 7.430 158.070 ;
        RECT 107.790 158.200 108.040 159.640 ;
        RECT 243.010 158.330 243.260 159.770 ;
        RECT 344.330 159.580 344.560 160.390 ;
        RECT 243.010 158.250 243.390 158.330 ;
        RECT 107.790 158.120 108.170 158.200 ;
        RECT 243.010 158.190 243.960 158.250 ;
        RECT 107.790 158.060 108.740 158.120 ;
        RECT 107.800 157.880 108.740 158.060 ;
        RECT 243.020 158.010 243.960 158.190 ;
        RECT 6.630 157.050 6.870 157.840 ;
        RECT 107.940 157.650 108.740 157.880 ;
        RECT 243.160 157.780 243.960 158.010 ;
        RECT 344.320 158.140 344.570 159.580 ;
        RECT 344.320 158.060 344.700 158.140 ;
        RECT 344.320 158.000 345.270 158.060 ;
        RECT 344.330 157.820 345.270 158.000 ;
        RECT 6.630 155.840 6.880 157.050 ;
        RECT 6.650 155.640 6.880 155.840 ;
        RECT 107.940 156.860 108.180 157.650 ;
        RECT 243.160 156.990 243.400 157.780 ;
        RECT 344.470 157.590 345.270 157.820 ;
        RECT 107.940 155.650 108.190 156.860 ;
        RECT 243.160 155.780 243.410 156.990 ;
        RECT 6.650 155.620 6.870 155.640 ;
        RECT 6.640 155.060 6.870 155.620 ;
        RECT 107.960 155.450 108.190 155.650 ;
        RECT 243.180 155.580 243.410 155.780 ;
        RECT 344.470 156.800 344.710 157.590 ;
        RECT 344.470 155.590 344.720 156.800 ;
        RECT 243.180 155.560 243.400 155.580 ;
        RECT 107.960 155.430 108.180 155.450 ;
        RECT 6.640 154.870 6.880 155.060 ;
        RECT 107.950 154.870 108.180 155.430 ;
        RECT 243.170 155.000 243.400 155.560 ;
        RECT 344.490 155.390 344.720 155.590 ;
        RECT 344.490 155.370 344.710 155.390 ;
        RECT 6.640 154.400 6.870 154.870 ;
        RECT 6.270 154.180 6.870 154.400 ;
        RECT 107.950 154.680 108.190 154.870 ;
        RECT 243.170 154.810 243.410 155.000 ;
        RECT 344.480 154.810 344.710 155.370 ;
        RECT 107.950 154.210 108.180 154.680 ;
        RECT 243.170 154.340 243.400 154.810 ;
        RECT 6.630 151.910 6.870 154.180 ;
        RECT 107.580 153.990 108.180 154.210 ;
        RECT 242.800 154.120 243.400 154.340 ;
        RECT 344.480 154.620 344.720 154.810 ;
        RECT 344.480 154.150 344.710 154.620 ;
        RECT 6.630 151.670 7.590 151.910 ;
        RECT 6.450 151.440 7.590 151.670 ;
        RECT 107.940 151.720 108.180 153.990 ;
        RECT 243.160 151.850 243.400 154.120 ;
        RECT 344.110 153.930 344.710 154.150 ;
        RECT 107.940 151.480 108.900 151.720 ;
        RECT 243.160 151.610 244.120 151.850 ;
        RECT 6.450 149.820 6.930 151.440 ;
        RECT 107.760 151.250 108.900 151.480 ;
        RECT 242.980 151.380 244.120 151.610 ;
        RECT 344.470 151.660 344.710 153.930 ;
        RECT 344.470 151.420 345.430 151.660 ;
        RECT 107.760 149.630 108.240 151.250 ;
        RECT 242.980 149.760 243.460 151.380 ;
        RECT 344.290 151.190 345.430 151.420 ;
        RECT 344.290 149.570 344.770 151.190 ;
        RECT 6.470 145.710 6.930 146.450 ;
        RECT 6.470 143.890 6.950 145.710 ;
        RECT 107.780 145.520 108.240 146.260 ;
        RECT 243.000 145.650 243.460 146.390 ;
        RECT 6.470 143.870 7.260 143.890 ;
        RECT 6.460 143.420 7.260 143.870 ;
        RECT 107.780 143.700 108.260 145.520 ;
        RECT 243.000 143.830 243.480 145.650 ;
        RECT 344.310 145.460 344.770 146.200 ;
        RECT 243.000 143.810 243.790 143.830 ;
        RECT 107.780 143.680 108.570 143.700 ;
        RECT 6.460 142.630 6.700 143.420 ;
        RECT 107.770 143.230 108.570 143.680 ;
        RECT 242.990 143.360 243.790 143.810 ;
        RECT 344.310 143.640 344.790 145.460 ;
        RECT 344.310 143.620 345.100 143.640 ;
        RECT 6.460 141.420 6.710 142.630 ;
        RECT 6.480 141.220 6.710 141.420 ;
        RECT 107.770 142.440 108.010 143.230 ;
        RECT 242.990 142.570 243.230 143.360 ;
        RECT 344.300 143.170 345.100 143.620 ;
        RECT 107.770 141.230 108.020 142.440 ;
        RECT 242.990 141.360 243.240 142.570 ;
        RECT 6.480 141.200 6.700 141.220 ;
        RECT 6.470 140.640 6.700 141.200 ;
        RECT 107.790 141.030 108.020 141.230 ;
        RECT 243.010 141.160 243.240 141.360 ;
        RECT 344.300 142.380 344.540 143.170 ;
        RECT 344.300 141.170 344.550 142.380 ;
        RECT 243.010 141.140 243.230 141.160 ;
        RECT 107.790 141.010 108.010 141.030 ;
        RECT 6.470 140.450 6.710 140.640 ;
        RECT 107.780 140.450 108.010 141.010 ;
        RECT 243.000 140.580 243.230 141.140 ;
        RECT 344.320 140.970 344.550 141.170 ;
        RECT 344.320 140.950 344.540 140.970 ;
        RECT 6.470 139.980 6.700 140.450 ;
        RECT 6.100 139.760 6.700 139.980 ;
        RECT 107.780 140.260 108.020 140.450 ;
        RECT 243.000 140.390 243.240 140.580 ;
        RECT 344.310 140.390 344.540 140.950 ;
        RECT 107.780 139.790 108.010 140.260 ;
        RECT 243.000 139.920 243.230 140.390 ;
        RECT 6.460 137.490 6.700 139.760 ;
        RECT 107.410 139.570 108.010 139.790 ;
        RECT 242.630 139.700 243.230 139.920 ;
        RECT 344.310 140.200 344.550 140.390 ;
        RECT 344.310 139.730 344.540 140.200 ;
        RECT 6.460 137.050 7.420 137.490 ;
        RECT 6.500 137.020 7.420 137.050 ;
        RECT 107.770 137.300 108.010 139.570 ;
        RECT 242.990 137.430 243.230 139.700 ;
        RECT 343.940 139.510 344.540 139.730 ;
        RECT 6.510 135.360 6.800 137.020 ;
        RECT 107.770 136.860 108.730 137.300 ;
        RECT 242.990 136.990 243.950 137.430 ;
        RECT 243.030 136.960 243.950 136.990 ;
        RECT 344.300 137.240 344.540 139.510 ;
        RECT 107.810 136.830 108.730 136.860 ;
        RECT 107.820 135.170 108.110 136.830 ;
        RECT 243.040 135.300 243.330 136.960 ;
        RECT 344.300 136.800 345.260 137.240 ;
        RECT 344.340 136.770 345.260 136.800 ;
        RECT 344.350 135.110 344.640 136.770 ;
        RECT 6.510 131.850 6.800 134.640 ;
        RECT 107.820 131.660 108.110 134.450 ;
        RECT 243.040 131.790 243.330 134.580 ;
        RECT 344.350 131.600 344.640 134.390 ;
        RECT 6.500 128.060 6.790 130.600 ;
        RECT 6.500 127.740 7.310 128.060 ;
        RECT 6.510 127.590 7.310 127.740 ;
        RECT 107.810 127.870 108.100 130.410 ;
        RECT 243.030 128.000 243.320 130.540 ;
        RECT 6.510 126.800 6.750 127.590 ;
        RECT 107.810 127.550 108.620 127.870 ;
        RECT 243.030 127.680 243.840 128.000 ;
        RECT 107.820 127.400 108.620 127.550 ;
        RECT 243.040 127.530 243.840 127.680 ;
        RECT 344.340 127.810 344.630 130.350 ;
        RECT 6.510 125.590 6.760 126.800 ;
        RECT 6.530 125.390 6.760 125.590 ;
        RECT 107.820 126.610 108.060 127.400 ;
        RECT 243.040 126.740 243.280 127.530 ;
        RECT 344.340 127.490 345.150 127.810 ;
        RECT 344.350 127.340 345.150 127.490 ;
        RECT 107.820 125.400 108.070 126.610 ;
        RECT 243.040 125.530 243.290 126.740 ;
        RECT 6.530 125.370 6.750 125.390 ;
        RECT 6.520 124.810 6.750 125.370 ;
        RECT 107.840 125.200 108.070 125.400 ;
        RECT 243.060 125.330 243.290 125.530 ;
        RECT 344.350 126.550 344.590 127.340 ;
        RECT 344.350 125.340 344.600 126.550 ;
        RECT 243.060 125.310 243.280 125.330 ;
        RECT 107.840 125.180 108.060 125.200 ;
        RECT 6.520 124.620 6.760 124.810 ;
        RECT 107.830 124.620 108.060 125.180 ;
        RECT 243.050 124.750 243.280 125.310 ;
        RECT 344.370 125.140 344.600 125.340 ;
        RECT 344.370 125.120 344.590 125.140 ;
        RECT 6.520 124.150 6.750 124.620 ;
        RECT 6.150 123.930 6.750 124.150 ;
        RECT 107.830 124.430 108.070 124.620 ;
        RECT 243.050 124.560 243.290 124.750 ;
        RECT 344.360 124.560 344.590 125.120 ;
        RECT 107.830 123.960 108.060 124.430 ;
        RECT 243.050 124.090 243.280 124.560 ;
        RECT 6.510 121.660 6.750 123.930 ;
        RECT 107.460 123.740 108.060 123.960 ;
        RECT 242.680 123.870 243.280 124.090 ;
        RECT 344.360 124.370 344.600 124.560 ;
        RECT 344.360 123.900 344.590 124.370 ;
        RECT 6.510 121.420 7.470 121.660 ;
        RECT 6.330 121.190 7.470 121.420 ;
        RECT 107.820 121.470 108.060 123.740 ;
        RECT 243.040 121.600 243.280 123.870 ;
        RECT 343.990 123.680 344.590 123.900 ;
        RECT 107.820 121.230 108.780 121.470 ;
        RECT 243.040 121.360 244.000 121.600 ;
        RECT 6.330 119.570 6.810 121.190 ;
        RECT 107.640 121.000 108.780 121.230 ;
        RECT 242.860 121.130 244.000 121.360 ;
        RECT 344.350 121.410 344.590 123.680 ;
        RECT 344.350 121.170 345.310 121.410 ;
        RECT 107.640 119.380 108.120 121.000 ;
        RECT 242.860 119.510 243.340 121.130 ;
        RECT 344.170 120.940 345.310 121.170 ;
        RECT 344.170 119.320 344.650 120.940 ;
        RECT 6.350 115.460 6.810 116.200 ;
        RECT 6.350 113.640 6.830 115.460 ;
        RECT 107.660 115.270 108.120 116.010 ;
        RECT 242.880 115.400 243.340 116.140 ;
        RECT 6.350 113.620 7.140 113.640 ;
        RECT 6.340 113.170 7.140 113.620 ;
        RECT 107.660 113.450 108.140 115.270 ;
        RECT 242.880 113.580 243.360 115.400 ;
        RECT 344.190 115.210 344.650 115.950 ;
        RECT 242.880 113.560 243.670 113.580 ;
        RECT 107.660 113.430 108.450 113.450 ;
        RECT 6.340 112.380 6.580 113.170 ;
        RECT 107.650 112.980 108.450 113.430 ;
        RECT 242.870 113.110 243.670 113.560 ;
        RECT 344.190 113.390 344.670 115.210 ;
        RECT 344.190 113.370 344.980 113.390 ;
        RECT 6.340 111.170 6.590 112.380 ;
        RECT 6.360 110.970 6.590 111.170 ;
        RECT 107.650 112.190 107.890 112.980 ;
        RECT 242.870 112.320 243.110 113.110 ;
        RECT 344.180 112.920 344.980 113.370 ;
        RECT 107.650 110.980 107.900 112.190 ;
        RECT 242.870 111.110 243.120 112.320 ;
        RECT 6.360 110.950 6.580 110.970 ;
        RECT 6.350 110.390 6.580 110.950 ;
        RECT 107.670 110.780 107.900 110.980 ;
        RECT 242.890 110.910 243.120 111.110 ;
        RECT 344.180 112.130 344.420 112.920 ;
        RECT 344.180 110.920 344.430 112.130 ;
        RECT 242.890 110.890 243.110 110.910 ;
        RECT 107.670 110.760 107.890 110.780 ;
        RECT 6.350 110.200 6.590 110.390 ;
        RECT 107.660 110.200 107.890 110.760 ;
        RECT 242.880 110.330 243.110 110.890 ;
        RECT 344.200 110.720 344.430 110.920 ;
        RECT 344.200 110.700 344.420 110.720 ;
        RECT 6.350 109.730 6.580 110.200 ;
        RECT 5.980 109.510 6.580 109.730 ;
        RECT 107.660 110.010 107.900 110.200 ;
        RECT 242.880 110.140 243.120 110.330 ;
        RECT 344.190 110.140 344.420 110.700 ;
        RECT 107.660 109.540 107.890 110.010 ;
        RECT 242.880 109.670 243.110 110.140 ;
        RECT 6.340 107.240 6.580 109.510 ;
        RECT 107.290 109.320 107.890 109.540 ;
        RECT 242.510 109.450 243.110 109.670 ;
        RECT 344.190 109.950 344.430 110.140 ;
        RECT 344.190 109.480 344.420 109.950 ;
        RECT 6.340 106.800 7.300 107.240 ;
        RECT 6.350 106.770 7.300 106.800 ;
        RECT 107.650 107.050 107.890 109.320 ;
        RECT 242.870 107.180 243.110 109.450 ;
        RECT 343.820 109.260 344.420 109.480 ;
        RECT 6.350 105.620 6.570 106.770 ;
        RECT 107.650 106.610 108.610 107.050 ;
        RECT 242.870 106.740 243.830 107.180 ;
        RECT 107.660 106.580 108.610 106.610 ;
        RECT 242.880 106.710 243.830 106.740 ;
        RECT 344.180 106.990 344.420 109.260 ;
        RECT 6.290 105.400 6.610 105.620 ;
        RECT 107.660 105.430 107.880 106.580 ;
        RECT 242.880 105.560 243.100 106.710 ;
        RECT 344.180 106.550 345.140 106.990 ;
        RECT 344.190 106.520 345.140 106.550 ;
        RECT 107.600 105.210 107.920 105.430 ;
        RECT 242.820 105.340 243.140 105.560 ;
        RECT 344.190 105.370 344.410 106.520 ;
        RECT 344.130 105.150 344.450 105.370 ;
        RECT 6.320 104.210 6.640 104.450 ;
        RECT 6.350 101.800 6.580 104.210 ;
        RECT 107.630 104.020 107.950 104.260 ;
        RECT 242.850 104.150 243.170 104.390 ;
        RECT 6.290 101.750 6.670 101.800 ;
        RECT 6.290 101.480 6.680 101.750 ;
        RECT 107.660 101.610 107.890 104.020 ;
        RECT 242.880 101.740 243.110 104.150 ;
        RECT 344.160 103.960 344.480 104.200 ;
        RECT 242.820 101.690 243.200 101.740 ;
        RECT 6.300 101.430 6.680 101.480 ;
        RECT 107.600 101.560 107.980 101.610 ;
        RECT 107.600 101.290 107.990 101.560 ;
        RECT 242.820 101.420 243.210 101.690 ;
        RECT 344.190 101.550 344.420 103.960 ;
        RECT 242.830 101.370 243.210 101.420 ;
        RECT 344.130 101.500 344.510 101.550 ;
        RECT 107.610 101.240 107.990 101.290 ;
        RECT 344.130 101.230 344.520 101.500 ;
        RECT 344.140 101.180 344.520 101.230 ;
        RECT 6.280 100.320 6.650 100.690 ;
        RECT 6.340 99.510 6.570 100.320 ;
        RECT 107.590 100.130 107.960 100.500 ;
        RECT 242.810 100.260 243.180 100.630 ;
        RECT 6.330 98.070 6.580 99.510 ;
        RECT 107.650 99.320 107.880 100.130 ;
        RECT 242.870 99.450 243.100 100.260 ;
        RECT 344.120 100.070 344.490 100.440 ;
        RECT 6.330 97.990 6.710 98.070 ;
        RECT 6.330 97.930 7.280 97.990 ;
        RECT 6.340 97.750 7.280 97.930 ;
        RECT 6.480 97.520 7.280 97.750 ;
        RECT 107.640 97.880 107.890 99.320 ;
        RECT 242.860 98.010 243.110 99.450 ;
        RECT 344.180 99.260 344.410 100.070 ;
        RECT 242.860 97.930 243.240 98.010 ;
        RECT 107.640 97.800 108.020 97.880 ;
        RECT 242.860 97.870 243.810 97.930 ;
        RECT 107.640 97.740 108.590 97.800 ;
        RECT 107.650 97.560 108.590 97.740 ;
        RECT 242.870 97.690 243.810 97.870 ;
        RECT 6.480 96.730 6.720 97.520 ;
        RECT 107.790 97.330 108.590 97.560 ;
        RECT 243.010 97.460 243.810 97.690 ;
        RECT 344.170 97.820 344.420 99.260 ;
        RECT 344.170 97.740 344.550 97.820 ;
        RECT 344.170 97.680 345.120 97.740 ;
        RECT 344.180 97.500 345.120 97.680 ;
        RECT 6.480 95.520 6.730 96.730 ;
        RECT 6.500 95.320 6.730 95.520 ;
        RECT 107.790 96.540 108.030 97.330 ;
        RECT 243.010 96.670 243.250 97.460 ;
        RECT 344.320 97.270 345.120 97.500 ;
        RECT 107.790 95.330 108.040 96.540 ;
        RECT 243.010 95.460 243.260 96.670 ;
        RECT 6.500 95.300 6.720 95.320 ;
        RECT 6.490 94.740 6.720 95.300 ;
        RECT 107.810 95.130 108.040 95.330 ;
        RECT 243.030 95.260 243.260 95.460 ;
        RECT 344.320 96.480 344.560 97.270 ;
        RECT 344.320 95.270 344.570 96.480 ;
        RECT 243.030 95.240 243.250 95.260 ;
        RECT 107.810 95.110 108.030 95.130 ;
        RECT 6.490 94.550 6.730 94.740 ;
        RECT 107.800 94.550 108.030 95.110 ;
        RECT 243.020 94.680 243.250 95.240 ;
        RECT 344.340 95.070 344.570 95.270 ;
        RECT 344.340 95.050 344.560 95.070 ;
        RECT 6.490 94.080 6.720 94.550 ;
        RECT 6.120 93.860 6.720 94.080 ;
        RECT 107.800 94.360 108.040 94.550 ;
        RECT 243.020 94.490 243.260 94.680 ;
        RECT 344.330 94.490 344.560 95.050 ;
        RECT 107.800 93.890 108.030 94.360 ;
        RECT 243.020 94.020 243.250 94.490 ;
        RECT 6.480 91.590 6.720 93.860 ;
        RECT 107.430 93.670 108.030 93.890 ;
        RECT 242.650 93.800 243.250 94.020 ;
        RECT 344.330 94.300 344.570 94.490 ;
        RECT 344.330 93.830 344.560 94.300 ;
        RECT 6.480 91.350 7.440 91.590 ;
        RECT 6.300 91.120 7.440 91.350 ;
        RECT 107.790 91.400 108.030 93.670 ;
        RECT 243.010 91.530 243.250 93.800 ;
        RECT 343.960 93.610 344.560 93.830 ;
        RECT 107.790 91.160 108.750 91.400 ;
        RECT 243.010 91.290 243.970 91.530 ;
        RECT 6.300 89.500 6.780 91.120 ;
        RECT 107.610 90.930 108.750 91.160 ;
        RECT 242.830 91.060 243.970 91.290 ;
        RECT 344.320 91.340 344.560 93.610 ;
        RECT 344.320 91.100 345.280 91.340 ;
        RECT 107.610 89.310 108.090 90.930 ;
        RECT 242.830 89.440 243.310 91.060 ;
        RECT 344.140 90.870 345.280 91.100 ;
        RECT 344.140 89.250 344.620 90.870 ;
        RECT 6.320 85.390 6.780 86.130 ;
        RECT 6.320 83.570 6.800 85.390 ;
        RECT 107.630 85.200 108.090 85.940 ;
        RECT 242.850 85.330 243.310 86.070 ;
        RECT 6.320 83.550 7.110 83.570 ;
        RECT 6.310 83.100 7.110 83.550 ;
        RECT 107.630 83.380 108.110 85.200 ;
        RECT 242.850 83.510 243.330 85.330 ;
        RECT 344.160 85.140 344.620 85.880 ;
        RECT 242.850 83.490 243.640 83.510 ;
        RECT 107.630 83.360 108.420 83.380 ;
        RECT 6.310 82.310 6.550 83.100 ;
        RECT 107.620 82.910 108.420 83.360 ;
        RECT 242.840 83.040 243.640 83.490 ;
        RECT 344.160 83.320 344.640 85.140 ;
        RECT 344.160 83.300 344.950 83.320 ;
        RECT 6.310 81.100 6.560 82.310 ;
        RECT 6.330 80.900 6.560 81.100 ;
        RECT 107.620 82.120 107.860 82.910 ;
        RECT 242.840 82.250 243.080 83.040 ;
        RECT 344.150 82.850 344.950 83.300 ;
        RECT 107.620 80.910 107.870 82.120 ;
        RECT 242.840 81.040 243.090 82.250 ;
        RECT 6.330 80.880 6.550 80.900 ;
        RECT 6.320 80.320 6.550 80.880 ;
        RECT 107.640 80.710 107.870 80.910 ;
        RECT 242.860 80.840 243.090 81.040 ;
        RECT 344.150 82.060 344.390 82.850 ;
        RECT 344.150 80.850 344.400 82.060 ;
        RECT 242.860 80.820 243.080 80.840 ;
        RECT 107.640 80.690 107.860 80.710 ;
        RECT 6.320 80.130 6.560 80.320 ;
        RECT 107.630 80.130 107.860 80.690 ;
        RECT 242.850 80.260 243.080 80.820 ;
        RECT 344.170 80.650 344.400 80.850 ;
        RECT 344.170 80.630 344.390 80.650 ;
        RECT 6.320 79.660 6.550 80.130 ;
        RECT 5.950 79.440 6.550 79.660 ;
        RECT 107.630 79.940 107.870 80.130 ;
        RECT 242.850 80.070 243.090 80.260 ;
        RECT 344.160 80.070 344.390 80.630 ;
        RECT 107.630 79.470 107.860 79.940 ;
        RECT 242.850 79.600 243.080 80.070 ;
        RECT 6.310 77.180 6.550 79.440 ;
        RECT 107.260 79.250 107.860 79.470 ;
        RECT 242.480 79.380 243.080 79.600 ;
        RECT 344.160 79.880 344.400 80.070 ;
        RECT 344.160 79.410 344.390 79.880 ;
        RECT 6.090 77.170 6.550 77.180 ;
        RECT 6.090 76.700 7.270 77.170 ;
        RECT 107.620 76.990 107.860 79.250 ;
        RECT 242.840 77.120 243.080 79.380 ;
        RECT 343.790 79.190 344.390 79.410 ;
        RECT 107.400 76.980 107.860 76.990 ;
        RECT 242.620 77.110 243.080 77.120 ;
        RECT 6.090 75.230 6.430 76.700 ;
        RECT 107.400 76.510 108.580 76.980 ;
        RECT 242.620 76.640 243.800 77.110 ;
        RECT 344.150 76.930 344.390 79.190 ;
        RECT 343.930 76.920 344.390 76.930 ;
        RECT 107.400 75.040 107.740 76.510 ;
        RECT 242.620 75.170 242.960 76.640 ;
        RECT 343.930 76.450 345.110 76.920 ;
        RECT 343.930 74.980 344.270 76.450 ;
        RECT 6.150 71.790 6.490 73.930 ;
        RECT 107.460 71.600 107.800 73.740 ;
        RECT 242.680 71.730 243.020 73.870 ;
        RECT 343.990 71.540 344.330 73.680 ;
        RECT 6.130 68.140 6.490 70.630 ;
        RECT 6.130 67.850 6.960 68.140 ;
        RECT 6.160 67.670 6.960 67.850 ;
        RECT 107.440 67.950 107.800 70.440 ;
        RECT 242.660 68.080 243.020 70.570 ;
        RECT 6.160 66.880 6.400 67.670 ;
        RECT 107.440 67.660 108.270 67.950 ;
        RECT 242.660 67.790 243.490 68.080 ;
        RECT 107.470 67.480 108.270 67.660 ;
        RECT 242.690 67.610 243.490 67.790 ;
        RECT 343.970 67.890 344.330 70.380 ;
        RECT 6.160 65.670 6.410 66.880 ;
        RECT 6.180 65.470 6.410 65.670 ;
        RECT 107.470 66.690 107.710 67.480 ;
        RECT 242.690 66.820 242.930 67.610 ;
        RECT 343.970 67.600 344.800 67.890 ;
        RECT 344.000 67.420 344.800 67.600 ;
        RECT 107.470 65.480 107.720 66.690 ;
        RECT 242.690 65.610 242.940 66.820 ;
        RECT 6.180 65.450 6.400 65.470 ;
        RECT 6.170 64.890 6.400 65.450 ;
        RECT 107.490 65.280 107.720 65.480 ;
        RECT 242.710 65.410 242.940 65.610 ;
        RECT 344.000 66.630 344.240 67.420 ;
        RECT 344.000 65.420 344.250 66.630 ;
        RECT 242.710 65.390 242.930 65.410 ;
        RECT 107.490 65.260 107.710 65.280 ;
        RECT 6.170 64.700 6.410 64.890 ;
        RECT 107.480 64.700 107.710 65.260 ;
        RECT 242.700 64.830 242.930 65.390 ;
        RECT 344.020 65.220 344.250 65.420 ;
        RECT 344.020 65.200 344.240 65.220 ;
        RECT 6.170 64.230 6.400 64.700 ;
        RECT 5.800 64.010 6.400 64.230 ;
        RECT 107.480 64.510 107.720 64.700 ;
        RECT 242.700 64.640 242.940 64.830 ;
        RECT 344.010 64.640 344.240 65.200 ;
        RECT 107.480 64.040 107.710 64.510 ;
        RECT 242.700 64.170 242.930 64.640 ;
        RECT 6.160 61.740 6.400 64.010 ;
        RECT 107.110 63.820 107.710 64.040 ;
        RECT 242.330 63.950 242.930 64.170 ;
        RECT 344.010 64.450 344.250 64.640 ;
        RECT 344.010 63.980 344.240 64.450 ;
        RECT 6.160 61.500 7.120 61.740 ;
        RECT 5.980 61.270 7.120 61.500 ;
        RECT 107.470 61.550 107.710 63.820 ;
        RECT 242.690 61.680 242.930 63.950 ;
        RECT 343.640 63.760 344.240 63.980 ;
        RECT 107.470 61.310 108.430 61.550 ;
        RECT 242.690 61.440 243.650 61.680 ;
        RECT 5.980 59.650 6.460 61.270 ;
        RECT 107.290 61.080 108.430 61.310 ;
        RECT 242.510 61.210 243.650 61.440 ;
        RECT 344.000 61.490 344.240 63.760 ;
        RECT 344.000 61.250 344.960 61.490 ;
        RECT 107.290 59.460 107.770 61.080 ;
        RECT 242.510 59.590 242.990 61.210 ;
        RECT 343.820 61.020 344.960 61.250 ;
        RECT 343.820 59.400 344.300 61.020 ;
        RECT 6.000 55.540 6.460 56.280 ;
        RECT 6.000 53.720 6.480 55.540 ;
        RECT 107.310 55.350 107.770 56.090 ;
        RECT 242.530 55.480 242.990 56.220 ;
        RECT 6.000 53.700 6.790 53.720 ;
        RECT 5.990 53.250 6.790 53.700 ;
        RECT 107.310 53.530 107.790 55.350 ;
        RECT 242.530 53.660 243.010 55.480 ;
        RECT 343.840 55.290 344.300 56.030 ;
        RECT 242.530 53.640 243.320 53.660 ;
        RECT 107.310 53.510 108.100 53.530 ;
        RECT 5.990 52.460 6.230 53.250 ;
        RECT 107.300 53.060 108.100 53.510 ;
        RECT 242.520 53.190 243.320 53.640 ;
        RECT 343.840 53.470 344.320 55.290 ;
        RECT 343.840 53.450 344.630 53.470 ;
        RECT 5.990 51.250 6.240 52.460 ;
        RECT 6.010 51.050 6.240 51.250 ;
        RECT 107.300 52.270 107.540 53.060 ;
        RECT 242.520 52.400 242.760 53.190 ;
        RECT 343.830 53.000 344.630 53.450 ;
        RECT 107.300 51.060 107.550 52.270 ;
        RECT 242.520 51.190 242.770 52.400 ;
        RECT 6.010 51.030 6.230 51.050 ;
        RECT 6.000 50.470 6.230 51.030 ;
        RECT 107.320 50.860 107.550 51.060 ;
        RECT 242.540 50.990 242.770 51.190 ;
        RECT 343.830 52.210 344.070 53.000 ;
        RECT 343.830 51.000 344.080 52.210 ;
        RECT 242.540 50.970 242.760 50.990 ;
        RECT 107.320 50.840 107.540 50.860 ;
        RECT 6.000 50.280 6.240 50.470 ;
        RECT 107.310 50.280 107.540 50.840 ;
        RECT 242.530 50.410 242.760 50.970 ;
        RECT 343.850 50.800 344.080 51.000 ;
        RECT 343.850 50.780 344.070 50.800 ;
        RECT 6.000 49.810 6.230 50.280 ;
        RECT 5.630 49.590 6.230 49.810 ;
        RECT 107.310 50.090 107.550 50.280 ;
        RECT 242.530 50.220 242.770 50.410 ;
        RECT 343.840 50.220 344.070 50.780 ;
        RECT 107.310 49.620 107.540 50.090 ;
        RECT 242.530 49.750 242.760 50.220 ;
        RECT 5.990 47.320 6.230 49.590 ;
        RECT 106.940 49.400 107.540 49.620 ;
        RECT 242.160 49.530 242.760 49.750 ;
        RECT 343.840 50.030 344.080 50.220 ;
        RECT 343.840 49.560 344.070 50.030 ;
        RECT 5.990 46.880 6.950 47.320 ;
        RECT 6.000 46.850 6.950 46.880 ;
        RECT 107.300 47.130 107.540 49.400 ;
        RECT 242.520 47.260 242.760 49.530 ;
        RECT 343.470 49.340 344.070 49.560 ;
        RECT 6.000 45.700 6.220 46.850 ;
        RECT 107.300 46.690 108.260 47.130 ;
        RECT 242.520 46.820 243.480 47.260 ;
        RECT 107.310 46.660 108.260 46.690 ;
        RECT 242.530 46.790 243.480 46.820 ;
        RECT 343.830 47.070 344.070 49.340 ;
        RECT 5.940 45.480 6.260 45.700 ;
        RECT 107.310 45.510 107.530 46.660 ;
        RECT 242.530 45.640 242.750 46.790 ;
        RECT 343.830 46.630 344.790 47.070 ;
        RECT 343.840 46.600 344.790 46.630 ;
        RECT 107.250 45.290 107.570 45.510 ;
        RECT 242.470 45.420 242.790 45.640 ;
        RECT 343.840 45.450 344.060 46.600 ;
        RECT 343.780 45.230 344.100 45.450 ;
        RECT 5.970 44.290 6.290 44.530 ;
        RECT 6.000 41.880 6.230 44.290 ;
        RECT 107.280 44.100 107.600 44.340 ;
        RECT 242.500 44.230 242.820 44.470 ;
        RECT 5.940 41.830 6.320 41.880 ;
        RECT 5.940 41.560 6.330 41.830 ;
        RECT 107.310 41.690 107.540 44.100 ;
        RECT 242.530 41.820 242.760 44.230 ;
        RECT 343.810 44.040 344.130 44.280 ;
        RECT 242.470 41.770 242.850 41.820 ;
        RECT 5.950 41.510 6.330 41.560 ;
        RECT 107.250 41.640 107.630 41.690 ;
        RECT 107.250 41.370 107.640 41.640 ;
        RECT 242.470 41.500 242.860 41.770 ;
        RECT 343.840 41.630 344.070 44.040 ;
        RECT 242.480 41.450 242.860 41.500 ;
        RECT 343.780 41.580 344.160 41.630 ;
        RECT 107.260 41.320 107.640 41.370 ;
        RECT 343.780 41.310 344.170 41.580 ;
        RECT 343.790 41.260 344.170 41.310 ;
        RECT 5.930 40.400 6.300 40.770 ;
        RECT 5.990 39.590 6.220 40.400 ;
        RECT 107.240 40.210 107.610 40.580 ;
        RECT 242.460 40.340 242.830 40.710 ;
        RECT 5.980 38.150 6.230 39.590 ;
        RECT 107.300 39.400 107.530 40.210 ;
        RECT 242.520 39.530 242.750 40.340 ;
        RECT 343.770 40.150 344.140 40.520 ;
        RECT 5.980 38.070 6.360 38.150 ;
        RECT 5.980 38.010 6.930 38.070 ;
        RECT 5.990 37.830 6.930 38.010 ;
        RECT 6.130 37.600 6.930 37.830 ;
        RECT 107.290 37.960 107.540 39.400 ;
        RECT 242.510 38.090 242.760 39.530 ;
        RECT 343.830 39.340 344.060 40.150 ;
        RECT 242.510 38.010 242.890 38.090 ;
        RECT 107.290 37.880 107.670 37.960 ;
        RECT 242.510 37.950 243.460 38.010 ;
        RECT 107.290 37.820 108.240 37.880 ;
        RECT 107.300 37.640 108.240 37.820 ;
        RECT 242.520 37.770 243.460 37.950 ;
        RECT 6.130 36.810 6.370 37.600 ;
        RECT 107.440 37.410 108.240 37.640 ;
        RECT 242.660 37.540 243.460 37.770 ;
        RECT 343.820 37.900 344.070 39.340 ;
        RECT 343.820 37.820 344.200 37.900 ;
        RECT 343.820 37.760 344.770 37.820 ;
        RECT 343.830 37.580 344.770 37.760 ;
        RECT 6.130 35.600 6.380 36.810 ;
        RECT 6.150 35.400 6.380 35.600 ;
        RECT 107.440 36.620 107.680 37.410 ;
        RECT 242.660 36.750 242.900 37.540 ;
        RECT 343.970 37.350 344.770 37.580 ;
        RECT 107.440 35.410 107.690 36.620 ;
        RECT 242.660 35.540 242.910 36.750 ;
        RECT 6.150 35.380 6.370 35.400 ;
        RECT 6.140 34.820 6.370 35.380 ;
        RECT 107.460 35.210 107.690 35.410 ;
        RECT 242.680 35.340 242.910 35.540 ;
        RECT 343.970 36.560 344.210 37.350 ;
        RECT 343.970 35.350 344.220 36.560 ;
        RECT 242.680 35.320 242.900 35.340 ;
        RECT 107.460 35.190 107.680 35.210 ;
        RECT 6.140 34.630 6.380 34.820 ;
        RECT 107.450 34.630 107.680 35.190 ;
        RECT 242.670 34.760 242.900 35.320 ;
        RECT 343.990 35.150 344.220 35.350 ;
        RECT 343.990 35.130 344.210 35.150 ;
        RECT 6.140 34.160 6.370 34.630 ;
        RECT 5.770 33.940 6.370 34.160 ;
        RECT 107.450 34.440 107.690 34.630 ;
        RECT 242.670 34.570 242.910 34.760 ;
        RECT 343.980 34.570 344.210 35.130 ;
        RECT 107.450 33.970 107.680 34.440 ;
        RECT 242.670 34.100 242.900 34.570 ;
        RECT 6.130 31.670 6.370 33.940 ;
        RECT 107.080 33.750 107.680 33.970 ;
        RECT 242.300 33.880 242.900 34.100 ;
        RECT 343.980 34.380 344.220 34.570 ;
        RECT 343.980 33.910 344.210 34.380 ;
        RECT 6.130 31.430 7.090 31.670 ;
        RECT 5.950 31.200 7.090 31.430 ;
        RECT 107.440 31.480 107.680 33.750 ;
        RECT 242.660 31.610 242.900 33.880 ;
        RECT 343.610 33.690 344.210 33.910 ;
        RECT 107.440 31.240 108.400 31.480 ;
        RECT 242.660 31.370 243.620 31.610 ;
        RECT 5.950 29.580 6.430 31.200 ;
        RECT 107.260 31.010 108.400 31.240 ;
        RECT 242.480 31.140 243.620 31.370 ;
        RECT 343.970 31.420 344.210 33.690 ;
        RECT 343.970 31.180 344.930 31.420 ;
        RECT 107.260 29.390 107.740 31.010 ;
        RECT 242.480 29.520 242.960 31.140 ;
        RECT 343.790 30.950 344.930 31.180 ;
        RECT 343.790 29.330 344.270 30.950 ;
        RECT 5.970 25.470 6.430 26.210 ;
        RECT 5.970 23.650 6.450 25.470 ;
        RECT 107.280 25.280 107.740 26.020 ;
        RECT 242.500 25.410 242.960 26.150 ;
        RECT 5.970 23.630 6.760 23.650 ;
        RECT 5.960 23.180 6.760 23.630 ;
        RECT 107.280 23.460 107.760 25.280 ;
        RECT 242.500 23.590 242.980 25.410 ;
        RECT 343.810 25.220 344.270 25.960 ;
        RECT 242.500 23.570 243.290 23.590 ;
        RECT 107.280 23.440 108.070 23.460 ;
        RECT 5.960 22.390 6.200 23.180 ;
        RECT 107.270 22.990 108.070 23.440 ;
        RECT 242.490 23.120 243.290 23.570 ;
        RECT 343.810 23.400 344.290 25.220 ;
        RECT 343.810 23.380 344.600 23.400 ;
        RECT 5.960 21.180 6.210 22.390 ;
        RECT 5.980 20.980 6.210 21.180 ;
        RECT 107.270 22.200 107.510 22.990 ;
        RECT 242.490 22.330 242.730 23.120 ;
        RECT 343.800 22.930 344.600 23.380 ;
        RECT 107.270 20.990 107.520 22.200 ;
        RECT 242.490 21.120 242.740 22.330 ;
        RECT 5.980 20.960 6.200 20.980 ;
        RECT 5.970 20.400 6.200 20.960 ;
        RECT 107.290 20.790 107.520 20.990 ;
        RECT 242.510 20.920 242.740 21.120 ;
        RECT 343.800 22.140 344.040 22.930 ;
        RECT 343.800 20.930 344.050 22.140 ;
        RECT 242.510 20.900 242.730 20.920 ;
        RECT 107.290 20.770 107.510 20.790 ;
        RECT 5.970 20.210 6.210 20.400 ;
        RECT 107.280 20.210 107.510 20.770 ;
        RECT 242.500 20.340 242.730 20.900 ;
        RECT 343.820 20.730 344.050 20.930 ;
        RECT 343.820 20.710 344.040 20.730 ;
        RECT 5.970 19.740 6.200 20.210 ;
        RECT 5.600 19.520 6.200 19.740 ;
        RECT 107.280 20.020 107.520 20.210 ;
        RECT 242.500 20.150 242.740 20.340 ;
        RECT 343.810 20.150 344.040 20.710 ;
        RECT 107.280 19.550 107.510 20.020 ;
        RECT 242.500 19.680 242.730 20.150 ;
        RECT 5.960 17.250 6.200 19.520 ;
        RECT 106.910 19.330 107.510 19.550 ;
        RECT 242.130 19.460 242.730 19.680 ;
        RECT 343.810 19.960 344.050 20.150 ;
        RECT 343.810 19.490 344.040 19.960 ;
        RECT 5.960 16.810 6.920 17.250 ;
        RECT 107.270 17.060 107.510 19.330 ;
        RECT 242.490 17.190 242.730 19.460 ;
        RECT 343.440 19.270 344.040 19.490 ;
        RECT 107.270 16.880 108.230 17.060 ;
        RECT 5.970 16.780 6.920 16.810 ;
        RECT 5.970 15.780 6.320 16.780 ;
        RECT 107.250 16.590 108.230 16.880 ;
        RECT 242.490 16.750 243.450 17.190 ;
        RECT 343.800 17.000 344.040 19.270 ;
        RECT 343.800 16.820 344.760 17.000 ;
        RECT 242.500 16.720 243.450 16.750 ;
        RECT 5.970 15.740 6.310 15.780 ;
        RECT 5.980 15.450 6.310 15.740 ;
        RECT 5.980 15.300 6.300 15.450 ;
        RECT 5.940 15.030 6.300 15.300 ;
        RECT 107.250 14.920 107.580 16.590 ;
        RECT 242.500 15.720 242.850 16.720 ;
        RECT 343.780 16.530 344.760 16.820 ;
        RECT 242.500 15.680 242.840 15.720 ;
        RECT 242.510 15.390 242.840 15.680 ;
        RECT 242.510 15.240 242.830 15.390 ;
        RECT 242.470 14.970 242.830 15.240 ;
        RECT 107.290 14.910 107.470 14.920 ;
        RECT 343.780 14.860 344.110 16.530 ;
        RECT 343.820 14.850 344.000 14.860 ;
        RECT 5.980 14.340 6.320 14.370 ;
        RECT 5.980 14.100 6.350 14.340 ;
        RECT 242.510 14.280 242.850 14.310 ;
        RECT 5.980 14.070 6.310 14.100 ;
        RECT 6.000 13.730 6.310 14.070 ;
        RECT 6.000 13.120 6.320 13.730 ;
        RECT 5.980 12.140 6.320 13.120 ;
        RECT 107.210 12.620 107.540 14.150 ;
        RECT 242.510 14.040 242.880 14.280 ;
        RECT 242.510 14.010 242.840 14.040 ;
        RECT 242.530 13.670 242.840 14.010 ;
        RECT 242.530 13.060 242.850 13.670 ;
        RECT 107.210 12.190 107.550 12.620 ;
        RECT 5.940 4.440 6.320 12.140 ;
        RECT 107.320 7.520 107.550 12.190 ;
        RECT 242.510 12.080 242.850 13.060 ;
        RECT 343.740 12.560 344.070 14.090 ;
        RECT 343.740 12.130 344.080 12.560 ;
        RECT 107.290 7.250 107.600 7.520 ;
        RECT 5.940 2.580 6.330 4.440 ;
        RECT 242.470 4.380 242.850 12.080 ;
        RECT 343.850 7.460 344.080 12.130 ;
        RECT 343.820 7.190 344.130 7.460 ;
        RECT 5.940 0.300 6.340 2.580 ;
        RECT 242.470 2.520 242.860 4.380 ;
        RECT 5.970 0.290 6.340 0.300 ;
        RECT 107.260 0.290 107.560 0.330 ;
        RECT 5.970 0.280 21.690 0.290 ;
        RECT 99.280 0.280 107.560 0.290 ;
        RECT 5.970 0.040 107.560 0.280 ;
        RECT 242.470 0.240 242.870 2.520 ;
        RECT 5.970 0.010 99.970 0.040 ;
        RECT 5.970 0.000 6.340 0.010 ;
        RECT 21.560 0.000 99.970 0.010 ;
        RECT 106.460 -5.850 106.760 0.040 ;
        RECT 107.260 0.020 107.560 0.040 ;
        RECT 242.500 0.230 242.870 0.240 ;
        RECT 343.790 0.230 344.090 0.270 ;
        RECT 242.500 0.220 258.220 0.230 ;
        RECT 335.810 0.220 344.090 0.230 ;
        RECT 242.500 -0.020 344.090 0.220 ;
        RECT 242.500 -0.050 336.500 -0.020 ;
        RECT 343.790 -0.040 344.090 -0.020 ;
        RECT 242.500 -0.060 242.870 -0.050 ;
        RECT 258.090 -0.060 336.500 -0.050 ;
        RECT 234.980 -5.850 242.870 -5.800 ;
        RECT 106.430 -5.860 138.760 -5.850 ;
        RECT 203.130 -5.860 242.870 -5.850 ;
        RECT 106.430 -6.120 242.870 -5.860 ;
        RECT 106.430 -6.150 235.460 -6.120 ;
        RECT 107.120 -6.160 132.250 -6.150 ;
        RECT 138.670 -6.160 203.250 -6.150 ;
      LAYER mcon ;
        RECT 6.960 239.995 7.130 240.165 ;
        RECT 108.270 239.805 108.440 239.975 ;
        RECT 243.490 239.935 243.660 240.105 ;
        RECT 344.800 239.745 344.970 239.915 ;
        RECT 7.000 236.155 7.170 236.325 ;
        RECT 108.310 235.965 108.480 236.135 ;
        RECT 243.530 236.095 243.700 236.265 ;
        RECT 344.840 235.905 345.010 236.075 ;
        RECT 6.875 225.670 7.045 225.840 ;
        RECT 108.185 225.480 108.355 225.650 ;
        RECT 243.405 225.610 243.575 225.780 ;
        RECT 344.715 225.420 344.885 225.590 ;
        RECT 6.890 224.480 7.060 224.650 ;
        RECT 108.200 224.290 108.370 224.460 ;
        RECT 243.420 224.420 243.590 224.590 ;
        RECT 6.895 221.765 7.065 221.935 ;
        RECT 344.730 224.230 344.900 224.400 ;
        RECT 108.205 221.575 108.375 221.745 ;
        RECT 243.425 221.705 243.595 221.875 ;
        RECT 344.735 221.515 344.905 221.685 ;
        RECT 6.880 220.655 7.050 220.825 ;
        RECT 108.190 220.465 108.360 220.635 ;
        RECT 243.410 220.595 243.580 220.765 ;
        RECT 344.720 220.405 344.890 220.575 ;
        RECT 6.930 209.925 7.100 210.095 ;
        RECT 108.240 209.735 108.410 209.905 ;
        RECT 243.460 209.865 243.630 210.035 ;
        RECT 344.770 209.675 344.940 209.845 ;
        RECT 6.970 206.085 7.140 206.255 ;
        RECT 108.280 205.895 108.450 206.065 ;
        RECT 243.500 206.025 243.670 206.195 ;
        RECT 344.810 205.835 344.980 206.005 ;
        RECT 6.710 195.625 6.880 195.795 ;
        RECT 108.020 195.435 108.190 195.605 ;
        RECT 243.240 195.565 243.410 195.735 ;
        RECT 344.550 195.375 344.720 195.545 ;
        RECT 6.700 193.925 6.870 194.095 ;
        RECT 6.750 192.175 6.920 192.345 ;
        RECT 108.010 193.735 108.180 193.905 ;
        RECT 108.060 191.985 108.230 192.155 ;
        RECT 243.230 193.865 243.400 194.035 ;
        RECT 243.280 192.115 243.450 192.285 ;
        RECT 344.540 193.675 344.710 193.845 ;
        RECT 344.590 191.925 344.760 192.095 ;
        RECT 6.730 190.485 6.900 190.655 ;
        RECT 108.040 190.295 108.210 190.465 ;
        RECT 243.260 190.425 243.430 190.595 ;
        RECT 344.570 190.235 344.740 190.405 ;
        RECT 6.610 180.075 6.780 180.245 ;
        RECT 107.920 179.885 108.090 180.055 ;
        RECT 243.140 180.015 243.310 180.185 ;
        RECT 344.450 179.825 344.620 179.995 ;
        RECT 6.650 176.235 6.820 176.405 ;
        RECT 107.960 176.045 108.130 176.215 ;
        RECT 243.180 176.175 243.350 176.345 ;
        RECT 344.490 175.985 344.660 176.155 ;
        RECT 6.525 165.750 6.695 165.920 ;
        RECT 107.835 165.560 108.005 165.730 ;
        RECT 243.055 165.690 243.225 165.860 ;
        RECT 344.365 165.500 344.535 165.670 ;
        RECT 6.540 164.560 6.710 164.730 ;
        RECT 107.850 164.370 108.020 164.540 ;
        RECT 243.070 164.500 243.240 164.670 ;
        RECT 6.545 161.845 6.715 162.015 ;
        RECT 344.380 164.310 344.550 164.480 ;
        RECT 107.855 161.655 108.025 161.825 ;
        RECT 243.075 161.785 243.245 161.955 ;
        RECT 344.385 161.595 344.555 161.765 ;
        RECT 6.530 160.735 6.700 160.905 ;
        RECT 107.840 160.545 108.010 160.715 ;
        RECT 243.060 160.675 243.230 160.845 ;
        RECT 344.370 160.485 344.540 160.655 ;
        RECT 6.580 150.005 6.750 150.175 ;
        RECT 107.890 149.815 108.060 149.985 ;
        RECT 243.110 149.945 243.280 150.115 ;
        RECT 344.420 149.755 344.590 149.925 ;
        RECT 6.620 146.165 6.790 146.335 ;
        RECT 107.930 145.975 108.100 146.145 ;
        RECT 243.150 146.105 243.320 146.275 ;
        RECT 344.460 145.915 344.630 146.085 ;
        RECT 6.585 135.415 6.755 135.585 ;
        RECT 107.895 135.225 108.065 135.395 ;
        RECT 243.115 135.355 243.285 135.525 ;
        RECT 344.425 135.165 344.595 135.335 ;
        RECT 6.560 134.395 6.730 134.565 ;
        RECT 6.565 131.890 6.735 132.060 ;
        RECT 107.870 134.205 108.040 134.375 ;
        RECT 107.875 131.700 108.045 131.870 ;
        RECT 243.090 134.335 243.260 134.505 ;
        RECT 243.095 131.830 243.265 132.000 ;
        RECT 344.400 134.145 344.570 134.315 ;
        RECT 344.405 131.640 344.575 131.810 ;
        RECT 6.565 130.290 6.735 130.460 ;
        RECT 107.875 130.100 108.045 130.270 ;
        RECT 243.095 130.230 243.265 130.400 ;
        RECT 344.405 130.040 344.575 130.210 ;
        RECT 6.460 119.755 6.630 119.925 ;
        RECT 107.770 119.565 107.940 119.735 ;
        RECT 242.990 119.695 243.160 119.865 ;
        RECT 344.300 119.505 344.470 119.675 ;
        RECT 6.500 115.915 6.670 116.085 ;
        RECT 107.810 115.725 107.980 115.895 ;
        RECT 243.030 115.855 243.200 116.025 ;
        RECT 344.340 115.665 344.510 115.835 ;
        RECT 6.375 105.430 6.545 105.600 ;
        RECT 107.685 105.240 107.855 105.410 ;
        RECT 242.905 105.370 243.075 105.540 ;
        RECT 344.215 105.180 344.385 105.350 ;
        RECT 6.390 104.240 6.560 104.410 ;
        RECT 107.700 104.050 107.870 104.220 ;
        RECT 242.920 104.180 243.090 104.350 ;
        RECT 6.395 101.525 6.565 101.695 ;
        RECT 344.230 103.990 344.400 104.160 ;
        RECT 107.705 101.335 107.875 101.505 ;
        RECT 242.925 101.465 243.095 101.635 ;
        RECT 344.235 101.275 344.405 101.445 ;
        RECT 6.380 100.415 6.550 100.585 ;
        RECT 107.690 100.225 107.860 100.395 ;
        RECT 242.910 100.355 243.080 100.525 ;
        RECT 344.220 100.165 344.390 100.335 ;
        RECT 6.430 89.685 6.600 89.855 ;
        RECT 107.740 89.495 107.910 89.665 ;
        RECT 242.960 89.625 243.130 89.795 ;
        RECT 344.270 89.435 344.440 89.605 ;
        RECT 6.470 85.845 6.640 86.015 ;
        RECT 107.780 85.655 107.950 85.825 ;
        RECT 243.000 85.785 243.170 85.955 ;
        RECT 344.310 85.595 344.480 85.765 ;
        RECT 6.210 75.385 6.380 75.555 ;
        RECT 107.520 75.195 107.690 75.365 ;
        RECT 242.740 75.325 242.910 75.495 ;
        RECT 344.050 75.135 344.220 75.305 ;
        RECT 6.200 73.685 6.370 73.855 ;
        RECT 6.250 71.935 6.420 72.105 ;
        RECT 107.510 73.495 107.680 73.665 ;
        RECT 107.560 71.745 107.730 71.915 ;
        RECT 242.730 73.625 242.900 73.795 ;
        RECT 242.780 71.875 242.950 72.045 ;
        RECT 344.040 73.435 344.210 73.605 ;
        RECT 344.090 71.685 344.260 71.855 ;
        RECT 6.230 70.245 6.400 70.415 ;
        RECT 107.540 70.055 107.710 70.225 ;
        RECT 242.760 70.185 242.930 70.355 ;
        RECT 344.070 69.995 344.240 70.165 ;
        RECT 6.110 59.835 6.280 60.005 ;
        RECT 107.420 59.645 107.590 59.815 ;
        RECT 242.640 59.775 242.810 59.945 ;
        RECT 343.950 59.585 344.120 59.755 ;
        RECT 6.150 55.995 6.320 56.165 ;
        RECT 107.460 55.805 107.630 55.975 ;
        RECT 242.680 55.935 242.850 56.105 ;
        RECT 343.990 55.745 344.160 55.915 ;
        RECT 6.025 45.510 6.195 45.680 ;
        RECT 107.335 45.320 107.505 45.490 ;
        RECT 242.555 45.450 242.725 45.620 ;
        RECT 343.865 45.260 344.035 45.430 ;
        RECT 6.040 44.320 6.210 44.490 ;
        RECT 107.350 44.130 107.520 44.300 ;
        RECT 242.570 44.260 242.740 44.430 ;
        RECT 6.045 41.605 6.215 41.775 ;
        RECT 343.880 44.070 344.050 44.240 ;
        RECT 107.355 41.415 107.525 41.585 ;
        RECT 242.575 41.545 242.745 41.715 ;
        RECT 343.885 41.355 344.055 41.525 ;
        RECT 6.030 40.495 6.200 40.665 ;
        RECT 107.340 40.305 107.510 40.475 ;
        RECT 242.560 40.435 242.730 40.605 ;
        RECT 343.870 40.245 344.040 40.415 ;
        RECT 6.080 29.765 6.250 29.935 ;
        RECT 107.390 29.575 107.560 29.745 ;
        RECT 242.610 29.705 242.780 29.875 ;
        RECT 343.920 29.515 344.090 29.685 ;
        RECT 6.120 25.925 6.290 26.095 ;
        RECT 107.430 25.735 107.600 25.905 ;
        RECT 242.650 25.865 242.820 26.035 ;
        RECT 343.960 25.675 344.130 25.845 ;
        RECT 6.025 15.090 6.195 15.260 ;
        RECT 107.295 14.950 107.465 15.120 ;
        RECT 242.555 15.030 242.725 15.200 ;
        RECT 343.825 14.890 343.995 15.060 ;
        RECT 6.075 14.140 6.245 14.310 ;
        RECT 107.295 13.900 107.465 14.070 ;
        RECT 242.605 14.080 242.775 14.250 ;
        RECT 343.825 13.840 343.995 14.010 ;
        RECT 107.340 7.280 107.510 7.450 ;
        RECT 343.870 7.220 344.040 7.390 ;
        RECT 107.315 0.085 107.485 0.255 ;
        RECT 242.615 0.025 242.785 0.195 ;
        RECT 343.845 0.025 344.015 0.195 ;
        RECT 106.530 -6.080 106.700 -5.910 ;
        RECT 106.790 -6.080 106.960 -5.910 ;
        RECT 107.040 -6.080 107.210 -5.910 ;
        RECT 107.300 -6.080 107.470 -5.910 ;
        RECT 242.605 -6.055 242.775 -5.885 ;
      LAYER met1 ;
        RECT 6.830 236.040 7.320 240.270 ;
        RECT 108.140 235.850 108.630 240.080 ;
        RECT 243.360 235.980 243.850 240.210 ;
        RECT 344.670 235.790 345.160 240.020 ;
        RECT 6.840 225.870 7.070 226.030 ;
        RECT 6.840 225.860 7.080 225.870 ;
        RECT 6.790 225.640 7.110 225.860 ;
        RECT 108.150 225.680 108.380 225.840 ;
        RECT 243.370 225.810 243.600 225.970 ;
        RECT 243.370 225.800 243.610 225.810 ;
        RECT 108.150 225.670 108.390 225.680 ;
        RECT 6.850 224.690 7.080 225.640 ;
        RECT 108.100 225.450 108.420 225.670 ;
        RECT 243.320 225.580 243.640 225.800 ;
        RECT 344.680 225.620 344.910 225.780 ;
        RECT 344.680 225.610 344.920 225.620 ;
        RECT 6.820 224.450 7.140 224.690 ;
        RECT 108.160 224.500 108.390 225.450 ;
        RECT 243.380 224.630 243.610 225.580 ;
        RECT 344.630 225.390 344.950 225.610 ;
        RECT 108.130 224.260 108.450 224.500 ;
        RECT 243.350 224.390 243.670 224.630 ;
        RECT 344.690 224.440 344.920 225.390 ;
        RECT 344.660 224.200 344.980 224.440 ;
        RECT 6.790 221.990 7.170 222.040 ;
        RECT 6.790 221.720 7.180 221.990 ;
        RECT 243.320 221.930 243.700 221.980 ;
        RECT 6.800 221.670 7.180 221.720 ;
        RECT 108.100 221.800 108.480 221.850 ;
        RECT 6.850 220.930 7.080 221.670 ;
        RECT 108.100 221.530 108.490 221.800 ;
        RECT 243.320 221.660 243.710 221.930 ;
        RECT 243.330 221.610 243.710 221.660 ;
        RECT 344.630 221.740 345.010 221.790 ;
        RECT 108.110 221.480 108.490 221.530 ;
        RECT 6.780 220.560 7.150 220.930 ;
        RECT 108.160 220.740 108.390 221.480 ;
        RECT 243.380 220.870 243.610 221.610 ;
        RECT 344.630 221.470 345.020 221.740 ;
        RECT 344.640 221.420 345.020 221.470 ;
        RECT 108.090 220.370 108.460 220.740 ;
        RECT 243.310 220.500 243.680 220.870 ;
        RECT 344.690 220.680 344.920 221.420 ;
        RECT 344.620 220.310 344.990 220.680 ;
        RECT 6.800 205.970 7.290 210.200 ;
        RECT 108.110 205.780 108.600 210.010 ;
        RECT 243.330 205.910 243.820 210.140 ;
        RECT 344.640 205.720 345.130 209.950 ;
        RECT 6.630 193.810 6.970 195.950 ;
        RECT 107.940 193.620 108.280 195.760 ;
        RECT 243.160 193.750 243.500 195.890 ;
        RECT 344.470 193.560 344.810 195.700 ;
        RECT 6.630 190.280 6.970 192.420 ;
        RECT 107.940 190.090 108.280 192.230 ;
        RECT 243.160 190.220 243.500 192.360 ;
        RECT 344.470 190.030 344.810 192.170 ;
        RECT 6.480 176.120 6.970 180.350 ;
        RECT 107.790 175.930 108.280 180.160 ;
        RECT 243.010 176.060 243.500 180.290 ;
        RECT 344.320 175.870 344.810 180.100 ;
        RECT 6.490 165.950 6.720 166.110 ;
        RECT 6.490 165.940 6.730 165.950 ;
        RECT 6.440 165.720 6.760 165.940 ;
        RECT 107.800 165.760 108.030 165.920 ;
        RECT 243.020 165.890 243.250 166.050 ;
        RECT 243.020 165.880 243.260 165.890 ;
        RECT 107.800 165.750 108.040 165.760 ;
        RECT 6.500 164.770 6.730 165.720 ;
        RECT 107.750 165.530 108.070 165.750 ;
        RECT 242.970 165.660 243.290 165.880 ;
        RECT 344.330 165.700 344.560 165.860 ;
        RECT 344.330 165.690 344.570 165.700 ;
        RECT 6.470 164.530 6.790 164.770 ;
        RECT 107.810 164.580 108.040 165.530 ;
        RECT 243.030 164.710 243.260 165.660 ;
        RECT 344.280 165.470 344.600 165.690 ;
        RECT 107.780 164.340 108.100 164.580 ;
        RECT 243.000 164.470 243.320 164.710 ;
        RECT 344.340 164.520 344.570 165.470 ;
        RECT 344.310 164.280 344.630 164.520 ;
        RECT 6.440 162.070 6.820 162.120 ;
        RECT 6.440 161.800 6.830 162.070 ;
        RECT 242.970 162.010 243.350 162.060 ;
        RECT 6.450 161.750 6.830 161.800 ;
        RECT 107.750 161.880 108.130 161.930 ;
        RECT 6.500 161.010 6.730 161.750 ;
        RECT 107.750 161.610 108.140 161.880 ;
        RECT 242.970 161.740 243.360 162.010 ;
        RECT 242.980 161.690 243.360 161.740 ;
        RECT 344.280 161.820 344.660 161.870 ;
        RECT 107.760 161.560 108.140 161.610 ;
        RECT 6.430 160.640 6.800 161.010 ;
        RECT 107.810 160.820 108.040 161.560 ;
        RECT 243.030 160.950 243.260 161.690 ;
        RECT 344.280 161.550 344.670 161.820 ;
        RECT 344.290 161.500 344.670 161.550 ;
        RECT 107.740 160.450 108.110 160.820 ;
        RECT 242.960 160.580 243.330 160.950 ;
        RECT 344.340 160.760 344.570 161.500 ;
        RECT 344.270 160.390 344.640 160.760 ;
        RECT 6.450 146.050 6.940 150.280 ;
        RECT 107.760 145.860 108.250 150.090 ;
        RECT 242.980 145.990 243.470 150.220 ;
        RECT 344.290 145.800 344.780 150.030 ;
        RECT 6.500 135.380 6.820 135.700 ;
        RECT 6.520 134.670 6.810 135.380 ;
        RECT 107.810 135.190 108.130 135.510 ;
        RECT 243.030 135.320 243.350 135.640 ;
        RECT 6.510 134.570 6.810 134.670 ;
        RECT 6.500 134.380 6.810 134.570 ;
        RECT 107.830 134.480 108.120 135.190 ;
        RECT 243.050 134.610 243.340 135.320 ;
        RECT 344.340 135.130 344.660 135.450 ;
        RECT 243.040 134.510 243.340 134.610 ;
        RECT 107.820 134.380 108.120 134.480 ;
        RECT 6.500 134.360 6.780 134.380 ;
        RECT 6.510 134.260 6.780 134.360 ;
        RECT 107.810 134.190 108.120 134.380 ;
        RECT 243.030 134.320 243.340 134.510 ;
        RECT 344.360 134.420 344.650 135.130 ;
        RECT 344.350 134.320 344.650 134.420 ;
        RECT 243.030 134.300 243.310 134.320 ;
        RECT 243.040 134.200 243.310 134.300 ;
        RECT 107.810 134.170 108.090 134.190 ;
        RECT 107.820 134.070 108.090 134.170 ;
        RECT 344.340 134.130 344.650 134.320 ;
        RECT 344.340 134.110 344.620 134.130 ;
        RECT 344.350 134.010 344.620 134.110 ;
        RECT 6.500 131.980 6.810 132.130 ;
        RECT 6.510 130.160 6.800 131.980 ;
        RECT 107.810 131.790 108.120 131.940 ;
        RECT 243.030 131.920 243.340 132.070 ;
        RECT 107.820 129.970 108.110 131.790 ;
        RECT 243.040 130.100 243.330 131.920 ;
        RECT 344.340 131.730 344.650 131.880 ;
        RECT 344.350 129.910 344.640 131.730 ;
        RECT 6.330 115.800 6.820 120.030 ;
        RECT 107.640 115.610 108.130 119.840 ;
        RECT 242.860 115.740 243.350 119.970 ;
        RECT 344.170 115.550 344.660 119.780 ;
        RECT 6.340 105.630 6.570 105.790 ;
        RECT 6.340 105.620 6.580 105.630 ;
        RECT 6.290 105.400 6.610 105.620 ;
        RECT 107.650 105.440 107.880 105.600 ;
        RECT 242.870 105.570 243.100 105.730 ;
        RECT 242.870 105.560 243.110 105.570 ;
        RECT 107.650 105.430 107.890 105.440 ;
        RECT 6.350 104.450 6.580 105.400 ;
        RECT 107.600 105.210 107.920 105.430 ;
        RECT 242.820 105.340 243.140 105.560 ;
        RECT 344.180 105.380 344.410 105.540 ;
        RECT 344.180 105.370 344.420 105.380 ;
        RECT 6.320 104.210 6.640 104.450 ;
        RECT 107.660 104.260 107.890 105.210 ;
        RECT 242.880 104.390 243.110 105.340 ;
        RECT 344.130 105.150 344.450 105.370 ;
        RECT 107.630 104.020 107.950 104.260 ;
        RECT 242.850 104.150 243.170 104.390 ;
        RECT 344.190 104.200 344.420 105.150 ;
        RECT 344.160 103.960 344.480 104.200 ;
        RECT 6.290 101.750 6.670 101.800 ;
        RECT 6.290 101.480 6.680 101.750 ;
        RECT 242.820 101.690 243.200 101.740 ;
        RECT 6.300 101.430 6.680 101.480 ;
        RECT 107.600 101.560 107.980 101.610 ;
        RECT 6.350 100.690 6.580 101.430 ;
        RECT 107.600 101.290 107.990 101.560 ;
        RECT 242.820 101.420 243.210 101.690 ;
        RECT 242.830 101.370 243.210 101.420 ;
        RECT 344.130 101.500 344.510 101.550 ;
        RECT 107.610 101.240 107.990 101.290 ;
        RECT 6.280 100.320 6.650 100.690 ;
        RECT 107.660 100.500 107.890 101.240 ;
        RECT 242.880 100.630 243.110 101.370 ;
        RECT 344.130 101.230 344.520 101.500 ;
        RECT 344.140 101.180 344.520 101.230 ;
        RECT 107.590 100.130 107.960 100.500 ;
        RECT 242.810 100.260 243.180 100.630 ;
        RECT 344.190 100.440 344.420 101.180 ;
        RECT 344.120 100.070 344.490 100.440 ;
        RECT 6.300 85.730 6.790 89.960 ;
        RECT 107.610 85.540 108.100 89.770 ;
        RECT 242.830 85.670 243.320 89.900 ;
        RECT 344.140 85.480 344.630 89.710 ;
        RECT 6.130 73.570 6.470 75.710 ;
        RECT 107.440 73.380 107.780 75.520 ;
        RECT 242.660 73.510 243.000 75.650 ;
        RECT 343.970 73.320 344.310 75.460 ;
        RECT 6.130 70.040 6.470 72.180 ;
        RECT 107.440 69.850 107.780 71.990 ;
        RECT 242.660 69.980 243.000 72.120 ;
        RECT 343.970 69.790 344.310 71.930 ;
        RECT 5.980 55.880 6.470 60.110 ;
        RECT 107.290 55.690 107.780 59.920 ;
        RECT 242.510 55.820 243.000 60.050 ;
        RECT 343.820 55.630 344.310 59.860 ;
        RECT 5.990 45.710 6.220 45.870 ;
        RECT 5.990 45.700 6.230 45.710 ;
        RECT 5.940 45.480 6.260 45.700 ;
        RECT 107.300 45.520 107.530 45.680 ;
        RECT 242.520 45.650 242.750 45.810 ;
        RECT 242.520 45.640 242.760 45.650 ;
        RECT 107.300 45.510 107.540 45.520 ;
        RECT 6.000 44.530 6.230 45.480 ;
        RECT 107.250 45.290 107.570 45.510 ;
        RECT 242.470 45.420 242.790 45.640 ;
        RECT 343.830 45.460 344.060 45.620 ;
        RECT 343.830 45.450 344.070 45.460 ;
        RECT 5.970 44.290 6.290 44.530 ;
        RECT 107.310 44.340 107.540 45.290 ;
        RECT 242.530 44.470 242.760 45.420 ;
        RECT 343.780 45.230 344.100 45.450 ;
        RECT 107.280 44.100 107.600 44.340 ;
        RECT 242.500 44.230 242.820 44.470 ;
        RECT 343.840 44.280 344.070 45.230 ;
        RECT 343.810 44.040 344.130 44.280 ;
        RECT 5.940 41.830 6.320 41.880 ;
        RECT 5.940 41.560 6.330 41.830 ;
        RECT 242.470 41.770 242.850 41.820 ;
        RECT 5.950 41.510 6.330 41.560 ;
        RECT 107.250 41.640 107.630 41.690 ;
        RECT 6.000 40.770 6.230 41.510 ;
        RECT 107.250 41.370 107.640 41.640 ;
        RECT 242.470 41.500 242.860 41.770 ;
        RECT 242.480 41.450 242.860 41.500 ;
        RECT 343.780 41.580 344.160 41.630 ;
        RECT 107.260 41.320 107.640 41.370 ;
        RECT 5.930 40.400 6.300 40.770 ;
        RECT 107.310 40.580 107.540 41.320 ;
        RECT 242.530 40.710 242.760 41.450 ;
        RECT 343.780 41.310 344.170 41.580 ;
        RECT 343.790 41.260 344.170 41.310 ;
        RECT 107.240 40.210 107.610 40.580 ;
        RECT 242.460 40.340 242.830 40.710 ;
        RECT 343.840 40.520 344.070 41.260 ;
        RECT 343.770 40.150 344.140 40.520 ;
        RECT 5.950 25.810 6.440 30.040 ;
        RECT 107.260 25.620 107.750 29.850 ;
        RECT 242.480 25.750 242.970 29.980 ;
        RECT 343.790 25.560 344.280 29.790 ;
        RECT 5.980 15.300 6.300 15.350 ;
        RECT 5.940 14.910 6.300 15.300 ;
        RECT 242.510 15.240 242.830 15.290 ;
        RECT 5.940 14.870 6.310 14.910 ;
        RECT 5.920 14.650 6.360 14.870 ;
        RECT 5.920 14.630 6.320 14.650 ;
        RECT 6.010 14.400 6.320 14.630 ;
        RECT 5.980 14.340 6.320 14.400 ;
        RECT 5.980 14.100 6.350 14.340 ;
        RECT 5.980 14.090 6.310 14.100 ;
        RECT 107.200 13.840 107.570 15.240 ;
        RECT 242.470 14.850 242.830 15.240 ;
        RECT 242.470 14.810 242.840 14.850 ;
        RECT 242.450 14.590 242.890 14.810 ;
        RECT 242.450 14.570 242.850 14.590 ;
        RECT 242.540 14.340 242.850 14.570 ;
        RECT 242.510 14.280 242.850 14.340 ;
        RECT 242.510 14.040 242.880 14.280 ;
        RECT 242.510 14.030 242.840 14.040 ;
        RECT 107.200 13.810 107.560 13.840 ;
        RECT 343.730 13.780 344.100 15.180 ;
        RECT 343.730 13.750 344.090 13.780 ;
        RECT 107.290 7.250 107.600 7.520 ;
        RECT 107.300 0.330 107.480 7.250 ;
        RECT 343.820 7.190 344.130 7.460 ;
        RECT 107.260 0.020 107.560 0.330 ;
        RECT 343.830 0.270 344.010 7.190 ;
        RECT 242.510 0.230 242.860 0.270 ;
        RECT 242.510 -0.050 242.870 0.230 ;
        RECT 343.790 -0.040 344.090 0.270 ;
        RECT 242.560 -5.810 242.870 -0.050 ;
        RECT 106.435 -15.030 107.555 -5.850 ;
        RECT 242.530 -6.120 242.870 -5.810 ;
      LAYER via ;
        RECT 106.570 -14.960 107.415 -14.125 ;
      LAYER met2 ;
        RECT 106.440 -19.465 107.545 -13.985 ;
        RECT 106.715 -21.310 107.290 -19.465 ;
        RECT 106.710 -25.310 107.290 -21.310 ;
    END
  END d0
  PIN vdd
    ANTENNADIFFAREA 566.099976 ;
    PORT
      LAYER nwell ;
        RECT 7.950 250.020 11.280 251.100 ;
        RECT 7.950 248.350 11.250 250.020 ;
        RECT 109.260 249.830 112.590 250.910 ;
        RECT 244.480 249.960 247.810 251.040 ;
        RECT 23.630 247.600 26.960 248.680 ;
        RECT 109.260 248.160 112.560 249.830 ;
        RECT 23.630 245.930 26.930 247.600 ;
        RECT 124.940 247.410 128.270 248.490 ;
        RECT 244.480 248.290 247.780 249.960 ;
        RECT 345.790 249.770 349.120 250.850 ;
        RECT 260.160 247.540 263.490 248.620 ;
        RECT 345.790 248.100 349.090 249.770 ;
        RECT 124.940 245.740 128.240 247.410 ;
        RECT 260.160 245.870 263.460 247.540 ;
        RECT 361.470 247.350 364.800 248.430 ;
        RECT 361.470 245.680 364.770 247.350 ;
        RECT 8.110 243.620 11.440 244.700 ;
        RECT 8.110 241.950 11.410 243.620 ;
        RECT 109.420 243.430 112.750 244.510 ;
        RECT 244.640 243.560 247.970 244.640 ;
        RECT 41.210 242.050 44.540 243.130 ;
        RECT 41.210 240.380 44.510 242.050 ;
        RECT 109.420 241.760 112.720 243.430 ;
        RECT 142.520 241.860 145.850 242.940 ;
        RECT 244.640 241.890 247.940 243.560 ;
        RECT 345.950 243.370 349.280 244.450 ;
        RECT 277.740 241.990 281.070 243.070 ;
        RECT 142.520 240.190 145.820 241.860 ;
        RECT 277.740 240.320 281.040 241.990 ;
        RECT 345.950 241.700 349.250 243.370 ;
        RECT 379.050 241.800 382.380 242.880 ;
        RECT 379.050 240.130 382.350 241.800 ;
        RECT 7.780 235.600 11.110 236.680 ;
        RECT 7.780 233.930 11.080 235.600 ;
        RECT 109.090 235.410 112.420 236.490 ;
        RECT 244.310 235.540 247.640 236.620 ;
        RECT 23.460 233.180 26.790 234.260 ;
        RECT 109.090 233.740 112.390 235.410 ;
        RECT 23.460 231.510 26.760 233.180 ;
        RECT 124.770 232.990 128.100 234.070 ;
        RECT 244.310 233.870 247.610 235.540 ;
        RECT 345.620 235.350 348.950 236.430 ;
        RECT 259.990 233.120 263.320 234.200 ;
        RECT 345.620 233.680 348.920 235.350 ;
        RECT 124.770 231.320 128.070 232.990 ;
        RECT 259.990 231.450 263.290 233.120 ;
        RECT 361.300 232.930 364.630 234.010 ;
        RECT 361.300 231.260 364.600 232.930 ;
        RECT 7.940 229.200 11.270 230.280 ;
        RECT 7.940 227.530 11.240 229.200 ;
        RECT 109.250 229.010 112.580 230.090 ;
        RECT 244.470 229.140 247.800 230.220 ;
        RECT 109.250 227.340 112.550 229.010 ;
        RECT 244.470 227.470 247.770 229.140 ;
        RECT 345.780 228.950 349.110 230.030 ;
        RECT 345.780 227.280 349.080 228.950 ;
        RECT 58.740 226.030 62.070 227.110 ;
        RECT 58.740 224.360 62.040 226.030 ;
        RECT 160.050 225.840 163.380 226.920 ;
        RECT 295.270 225.970 298.600 227.050 ;
        RECT 160.050 224.170 163.350 225.840 ;
        RECT 295.270 224.300 298.570 225.970 ;
        RECT 396.580 225.780 399.910 226.860 ;
        RECT 396.580 224.110 399.880 225.780 ;
        RECT 7.920 219.950 11.250 221.030 ;
        RECT 7.920 218.280 11.220 219.950 ;
        RECT 109.230 219.760 112.560 220.840 ;
        RECT 244.450 219.890 247.780 220.970 ;
        RECT 23.600 217.530 26.930 218.610 ;
        RECT 109.230 218.090 112.530 219.760 ;
        RECT 23.600 215.860 26.900 217.530 ;
        RECT 124.910 217.340 128.240 218.420 ;
        RECT 244.450 218.220 247.750 219.890 ;
        RECT 345.760 219.700 349.090 220.780 ;
        RECT 260.130 217.470 263.460 218.550 ;
        RECT 345.760 218.030 349.060 219.700 ;
        RECT 124.910 215.670 128.210 217.340 ;
        RECT 260.130 215.800 263.430 217.470 ;
        RECT 361.440 217.280 364.770 218.360 ;
        RECT 361.440 215.610 364.740 217.280 ;
        RECT 8.080 213.550 11.410 214.630 ;
        RECT 8.080 211.880 11.380 213.550 ;
        RECT 109.390 213.360 112.720 214.440 ;
        RECT 244.610 213.490 247.940 214.570 ;
        RECT 41.180 211.980 44.510 213.060 ;
        RECT 41.180 210.310 44.480 211.980 ;
        RECT 109.390 211.690 112.690 213.360 ;
        RECT 142.490 211.790 145.820 212.870 ;
        RECT 244.610 211.820 247.910 213.490 ;
        RECT 345.920 213.300 349.250 214.380 ;
        RECT 277.710 211.920 281.040 213.000 ;
        RECT 142.490 210.120 145.790 211.790 ;
        RECT 277.710 210.250 281.010 211.920 ;
        RECT 345.920 211.630 349.220 213.300 ;
        RECT 379.020 211.730 382.350 212.810 ;
        RECT 379.020 210.060 382.320 211.730 ;
        RECT 7.750 205.530 11.080 206.610 ;
        RECT 7.750 203.860 11.050 205.530 ;
        RECT 109.060 205.340 112.390 206.420 ;
        RECT 244.280 205.470 247.610 206.550 ;
        RECT 23.430 203.110 26.760 204.190 ;
        RECT 109.060 203.670 112.360 205.340 ;
        RECT 23.430 201.440 26.730 203.110 ;
        RECT 124.740 202.920 128.070 204.000 ;
        RECT 244.280 203.800 247.580 205.470 ;
        RECT 345.590 205.280 348.920 206.360 ;
        RECT 259.960 203.050 263.290 204.130 ;
        RECT 345.590 203.610 348.890 205.280 ;
        RECT 124.740 201.250 128.040 202.920 ;
        RECT 259.960 201.380 263.260 203.050 ;
        RECT 361.270 202.860 364.600 203.940 ;
        RECT 361.270 201.190 364.570 202.860 ;
        RECT 7.910 199.130 11.240 200.210 ;
        RECT 72.940 199.740 76.270 200.820 ;
        RECT 7.910 197.460 11.210 199.130 ;
        RECT 72.940 198.070 76.240 199.740 ;
        RECT 109.220 198.940 112.550 200.020 ;
        RECT 174.250 199.550 177.580 200.630 ;
        RECT 109.220 197.270 112.520 198.940 ;
        RECT 174.250 197.880 177.550 199.550 ;
        RECT 244.440 199.070 247.770 200.150 ;
        RECT 309.470 199.680 312.800 200.760 ;
        RECT 244.440 197.400 247.740 199.070 ;
        RECT 309.470 198.010 312.770 199.680 ;
        RECT 345.750 198.880 349.080 199.960 ;
        RECT 410.780 199.490 414.110 200.570 ;
        RECT 345.750 197.210 349.050 198.880 ;
        RECT 410.780 197.820 414.080 199.490 ;
        RECT 7.600 190.100 10.930 191.180 ;
        RECT 7.600 188.430 10.900 190.100 ;
        RECT 108.910 189.910 112.240 190.990 ;
        RECT 244.130 190.040 247.460 191.120 ;
        RECT 23.280 187.680 26.610 188.760 ;
        RECT 108.910 188.240 112.210 189.910 ;
        RECT 23.280 186.010 26.580 187.680 ;
        RECT 124.590 187.490 127.920 188.570 ;
        RECT 244.130 188.370 247.430 190.040 ;
        RECT 345.440 189.850 348.770 190.930 ;
        RECT 259.810 187.620 263.140 188.700 ;
        RECT 345.440 188.180 348.740 189.850 ;
        RECT 124.590 185.820 127.890 187.490 ;
        RECT 259.810 185.950 263.110 187.620 ;
        RECT 361.120 187.430 364.450 188.510 ;
        RECT 361.120 185.760 364.420 187.430 ;
        RECT 7.760 183.700 11.090 184.780 ;
        RECT 7.760 182.030 11.060 183.700 ;
        RECT 109.070 183.510 112.400 184.590 ;
        RECT 244.290 183.640 247.620 184.720 ;
        RECT 40.860 182.130 44.190 183.210 ;
        RECT 40.860 180.460 44.160 182.130 ;
        RECT 109.070 181.840 112.370 183.510 ;
        RECT 142.170 181.940 145.500 183.020 ;
        RECT 244.290 181.970 247.590 183.640 ;
        RECT 345.600 183.450 348.930 184.530 ;
        RECT 277.390 182.070 280.720 183.150 ;
        RECT 142.170 180.270 145.470 181.940 ;
        RECT 277.390 180.400 280.690 182.070 ;
        RECT 345.600 181.780 348.900 183.450 ;
        RECT 378.700 181.880 382.030 182.960 ;
        RECT 378.700 180.210 382.000 181.880 ;
        RECT 7.430 175.680 10.760 176.760 ;
        RECT 7.430 174.010 10.730 175.680 ;
        RECT 108.740 175.490 112.070 176.570 ;
        RECT 243.960 175.620 247.290 176.700 ;
        RECT 23.110 173.260 26.440 174.340 ;
        RECT 108.740 173.820 112.040 175.490 ;
        RECT 23.110 171.590 26.410 173.260 ;
        RECT 124.420 173.070 127.750 174.150 ;
        RECT 243.960 173.950 247.260 175.620 ;
        RECT 345.270 175.430 348.600 176.510 ;
        RECT 259.640 173.200 262.970 174.280 ;
        RECT 345.270 173.760 348.570 175.430 ;
        RECT 124.420 171.400 127.720 173.070 ;
        RECT 259.640 171.530 262.940 173.200 ;
        RECT 360.950 173.010 364.280 174.090 ;
        RECT 360.950 171.340 364.250 173.010 ;
        RECT 7.590 169.280 10.920 170.360 ;
        RECT 7.590 167.610 10.890 169.280 ;
        RECT 108.900 169.090 112.230 170.170 ;
        RECT 244.120 169.220 247.450 170.300 ;
        RECT 108.900 167.420 112.200 169.090 ;
        RECT 244.120 167.550 247.420 169.220 ;
        RECT 345.430 169.030 348.760 170.110 ;
        RECT 345.430 167.360 348.730 169.030 ;
        RECT 58.390 166.110 61.720 167.190 ;
        RECT 58.390 164.440 61.690 166.110 ;
        RECT 159.700 165.920 163.030 167.000 ;
        RECT 294.920 166.050 298.250 167.130 ;
        RECT 159.700 164.250 163.000 165.920 ;
        RECT 294.920 164.380 298.220 166.050 ;
        RECT 396.230 165.860 399.560 166.940 ;
        RECT 396.230 164.190 399.530 165.860 ;
        RECT 7.570 160.030 10.900 161.110 ;
        RECT 7.570 158.360 10.870 160.030 ;
        RECT 108.880 159.840 112.210 160.920 ;
        RECT 244.100 159.970 247.430 161.050 ;
        RECT 23.250 157.610 26.580 158.690 ;
        RECT 108.880 158.170 112.180 159.840 ;
        RECT 23.250 155.940 26.550 157.610 ;
        RECT 124.560 157.420 127.890 158.500 ;
        RECT 244.100 158.300 247.400 159.970 ;
        RECT 345.410 159.780 348.740 160.860 ;
        RECT 259.780 157.550 263.110 158.630 ;
        RECT 345.410 158.110 348.710 159.780 ;
        RECT 124.560 155.750 127.860 157.420 ;
        RECT 259.780 155.880 263.080 157.550 ;
        RECT 361.090 157.360 364.420 158.440 ;
        RECT 361.090 155.690 364.390 157.360 ;
        RECT 7.730 153.630 11.060 154.710 ;
        RECT 7.730 151.960 11.030 153.630 ;
        RECT 109.040 153.440 112.370 154.520 ;
        RECT 244.260 153.570 247.590 154.650 ;
        RECT 40.830 152.060 44.160 153.140 ;
        RECT 40.830 150.390 44.130 152.060 ;
        RECT 109.040 151.770 112.340 153.440 ;
        RECT 142.140 151.870 145.470 152.950 ;
        RECT 244.260 151.900 247.560 153.570 ;
        RECT 345.570 153.380 348.900 154.460 ;
        RECT 277.360 152.000 280.690 153.080 ;
        RECT 142.140 150.200 145.440 151.870 ;
        RECT 277.360 150.330 280.660 152.000 ;
        RECT 345.570 151.710 348.870 153.380 ;
        RECT 378.670 151.810 382.000 152.890 ;
        RECT 378.670 150.140 381.970 151.810 ;
        RECT 7.400 145.610 10.730 146.690 ;
        RECT 7.400 143.940 10.700 145.610 ;
        RECT 108.710 145.420 112.040 146.500 ;
        RECT 243.930 145.550 247.260 146.630 ;
        RECT 23.080 143.190 26.410 144.270 ;
        RECT 108.710 143.750 112.010 145.420 ;
        RECT 23.080 141.520 26.380 143.190 ;
        RECT 124.390 143.000 127.720 144.080 ;
        RECT 243.930 143.880 247.230 145.550 ;
        RECT 345.240 145.360 348.570 146.440 ;
        RECT 259.610 143.130 262.940 144.210 ;
        RECT 345.240 143.690 348.540 145.360 ;
        RECT 124.390 141.330 127.690 143.000 ;
        RECT 259.610 141.460 262.910 143.130 ;
        RECT 360.920 142.940 364.250 144.020 ;
        RECT 360.920 141.270 364.220 142.940 ;
        RECT 7.560 139.210 10.890 140.290 ;
        RECT 7.560 137.540 10.860 139.210 ;
        RECT 108.870 139.020 112.200 140.100 ;
        RECT 89.270 136.600 92.600 137.680 ;
        RECT 108.870 137.350 112.170 139.020 ;
        RECT 216.860 138.740 220.190 139.820 ;
        RECT 244.090 139.150 247.420 140.230 ;
        RECT 89.270 134.930 92.570 136.600 ;
        RECT 190.580 136.410 193.910 137.490 ;
        RECT 216.860 137.070 220.160 138.740 ;
        RECT 244.090 137.480 247.390 139.150 ;
        RECT 345.400 138.960 348.730 140.040 ;
        RECT 325.800 136.540 329.130 137.620 ;
        RECT 345.400 137.290 348.700 138.960 ;
        RECT 453.390 138.680 456.720 139.760 ;
        RECT 190.580 134.740 193.880 136.410 ;
        RECT 325.800 134.870 329.100 136.540 ;
        RECT 427.110 136.350 430.440 137.430 ;
        RECT 453.390 137.010 456.690 138.680 ;
        RECT 427.110 134.680 430.410 136.350 ;
        RECT 470.690 136.330 474.020 137.410 ;
        RECT 470.690 134.660 473.990 136.330 ;
        RECT 7.450 129.780 10.780 130.860 ;
        RECT 7.450 128.110 10.750 129.780 ;
        RECT 108.760 129.590 112.090 130.670 ;
        RECT 243.980 129.720 247.310 130.800 ;
        RECT 23.130 127.360 26.460 128.440 ;
        RECT 108.760 127.920 112.060 129.590 ;
        RECT 23.130 125.690 26.430 127.360 ;
        RECT 124.440 127.170 127.770 128.250 ;
        RECT 243.980 128.050 247.280 129.720 ;
        RECT 345.290 129.530 348.620 130.610 ;
        RECT 259.660 127.300 262.990 128.380 ;
        RECT 345.290 127.860 348.590 129.530 ;
        RECT 124.440 125.500 127.740 127.170 ;
        RECT 259.660 125.630 262.960 127.300 ;
        RECT 360.970 127.110 364.300 128.190 ;
        RECT 360.970 125.440 364.270 127.110 ;
        RECT 7.610 123.380 10.940 124.460 ;
        RECT 7.610 121.710 10.910 123.380 ;
        RECT 108.920 123.190 112.250 124.270 ;
        RECT 244.140 123.320 247.470 124.400 ;
        RECT 40.710 121.810 44.040 122.890 ;
        RECT 40.710 120.140 44.010 121.810 ;
        RECT 108.920 121.520 112.220 123.190 ;
        RECT 142.020 121.620 145.350 122.700 ;
        RECT 244.140 121.650 247.440 123.320 ;
        RECT 345.450 123.130 348.780 124.210 ;
        RECT 277.240 121.750 280.570 122.830 ;
        RECT 142.020 119.950 145.320 121.620 ;
        RECT 277.240 120.080 280.540 121.750 ;
        RECT 345.450 121.460 348.750 123.130 ;
        RECT 378.550 121.560 381.880 122.640 ;
        RECT 378.550 119.890 381.850 121.560 ;
        RECT 7.280 115.360 10.610 116.440 ;
        RECT 7.280 113.690 10.580 115.360 ;
        RECT 108.590 115.170 111.920 116.250 ;
        RECT 243.810 115.300 247.140 116.380 ;
        RECT 22.960 112.940 26.290 114.020 ;
        RECT 108.590 113.500 111.890 115.170 ;
        RECT 22.960 111.270 26.260 112.940 ;
        RECT 124.270 112.750 127.600 113.830 ;
        RECT 243.810 113.630 247.110 115.300 ;
        RECT 345.120 115.110 348.450 116.190 ;
        RECT 259.490 112.880 262.820 113.960 ;
        RECT 345.120 113.440 348.420 115.110 ;
        RECT 124.270 111.080 127.570 112.750 ;
        RECT 259.490 111.210 262.790 112.880 ;
        RECT 360.800 112.690 364.130 113.770 ;
        RECT 360.800 111.020 364.100 112.690 ;
        RECT 7.440 108.960 10.770 110.040 ;
        RECT 7.440 107.290 10.740 108.960 ;
        RECT 108.750 108.770 112.080 109.850 ;
        RECT 243.970 108.900 247.300 109.980 ;
        RECT 108.750 107.100 112.050 108.770 ;
        RECT 243.970 107.230 247.270 108.900 ;
        RECT 345.280 108.710 348.610 109.790 ;
        RECT 345.280 107.040 348.580 108.710 ;
        RECT 58.240 105.790 61.570 106.870 ;
        RECT 58.240 104.120 61.540 105.790 ;
        RECT 159.550 105.600 162.880 106.680 ;
        RECT 294.770 105.730 298.100 106.810 ;
        RECT 159.550 103.930 162.850 105.600 ;
        RECT 294.770 104.060 298.070 105.730 ;
        RECT 396.080 105.540 399.410 106.620 ;
        RECT 396.080 103.870 399.380 105.540 ;
        RECT 7.420 99.710 10.750 100.790 ;
        RECT 7.420 98.040 10.720 99.710 ;
        RECT 108.730 99.520 112.060 100.600 ;
        RECT 243.950 99.650 247.280 100.730 ;
        RECT 23.100 97.290 26.430 98.370 ;
        RECT 108.730 97.850 112.030 99.520 ;
        RECT 23.100 95.620 26.400 97.290 ;
        RECT 124.410 97.100 127.740 98.180 ;
        RECT 243.950 97.980 247.250 99.650 ;
        RECT 345.260 99.460 348.590 100.540 ;
        RECT 259.630 97.230 262.960 98.310 ;
        RECT 345.260 97.790 348.560 99.460 ;
        RECT 124.410 95.430 127.710 97.100 ;
        RECT 259.630 95.560 262.930 97.230 ;
        RECT 360.940 97.040 364.270 98.120 ;
        RECT 360.940 95.370 364.240 97.040 ;
        RECT 7.580 93.310 10.910 94.390 ;
        RECT 7.580 91.640 10.880 93.310 ;
        RECT 108.890 93.120 112.220 94.200 ;
        RECT 244.110 93.250 247.440 94.330 ;
        RECT 40.680 91.740 44.010 92.820 ;
        RECT 40.680 90.070 43.980 91.740 ;
        RECT 108.890 91.450 112.190 93.120 ;
        RECT 141.990 91.550 145.320 92.630 ;
        RECT 244.110 91.580 247.410 93.250 ;
        RECT 345.420 93.060 348.750 94.140 ;
        RECT 277.210 91.680 280.540 92.760 ;
        RECT 141.990 89.880 145.290 91.550 ;
        RECT 277.210 90.010 280.510 91.680 ;
        RECT 345.420 91.390 348.720 93.060 ;
        RECT 378.520 91.490 381.850 92.570 ;
        RECT 378.520 89.820 381.820 91.490 ;
        RECT 7.250 85.290 10.580 86.370 ;
        RECT 7.250 83.620 10.550 85.290 ;
        RECT 108.560 85.100 111.890 86.180 ;
        RECT 243.780 85.230 247.110 86.310 ;
        RECT 22.930 82.870 26.260 83.950 ;
        RECT 108.560 83.430 111.860 85.100 ;
        RECT 22.930 81.200 26.230 82.870 ;
        RECT 124.240 82.680 127.570 83.760 ;
        RECT 243.780 83.560 247.080 85.230 ;
        RECT 345.090 85.040 348.420 86.120 ;
        RECT 259.460 82.810 262.790 83.890 ;
        RECT 345.090 83.370 348.390 85.040 ;
        RECT 124.240 81.010 127.540 82.680 ;
        RECT 259.460 81.140 262.760 82.810 ;
        RECT 360.770 82.620 364.100 83.700 ;
        RECT 360.770 80.950 364.070 82.620 ;
        RECT 7.410 78.890 10.740 79.970 ;
        RECT 72.440 79.500 75.770 80.580 ;
        RECT 7.410 77.220 10.710 78.890 ;
        RECT 72.440 77.830 75.740 79.500 ;
        RECT 108.720 78.700 112.050 79.780 ;
        RECT 173.750 79.310 177.080 80.390 ;
        RECT 108.720 77.030 112.020 78.700 ;
        RECT 173.750 77.640 177.050 79.310 ;
        RECT 243.940 78.830 247.270 79.910 ;
        RECT 308.970 79.440 312.300 80.520 ;
        RECT 243.940 77.160 247.240 78.830 ;
        RECT 308.970 77.770 312.270 79.440 ;
        RECT 345.250 78.640 348.580 79.720 ;
        RECT 410.280 79.250 413.610 80.330 ;
        RECT 345.250 76.970 348.550 78.640 ;
        RECT 410.280 77.580 413.580 79.250 ;
        RECT 7.100 69.860 10.430 70.940 ;
        RECT 7.100 68.190 10.400 69.860 ;
        RECT 108.410 69.670 111.740 70.750 ;
        RECT 243.630 69.800 246.960 70.880 ;
        RECT 22.780 67.440 26.110 68.520 ;
        RECT 108.410 68.000 111.710 69.670 ;
        RECT 22.780 65.770 26.080 67.440 ;
        RECT 124.090 67.250 127.420 68.330 ;
        RECT 243.630 68.130 246.930 69.800 ;
        RECT 344.940 69.610 348.270 70.690 ;
        RECT 259.310 67.380 262.640 68.460 ;
        RECT 344.940 67.940 348.240 69.610 ;
        RECT 124.090 65.580 127.390 67.250 ;
        RECT 259.310 65.710 262.610 67.380 ;
        RECT 360.620 67.190 363.950 68.270 ;
        RECT 360.620 65.520 363.920 67.190 ;
        RECT 7.260 63.460 10.590 64.540 ;
        RECT 7.260 61.790 10.560 63.460 ;
        RECT 108.570 63.270 111.900 64.350 ;
        RECT 243.790 63.400 247.120 64.480 ;
        RECT 40.360 61.890 43.690 62.970 ;
        RECT 40.360 60.220 43.660 61.890 ;
        RECT 108.570 61.600 111.870 63.270 ;
        RECT 141.670 61.700 145.000 62.780 ;
        RECT 243.790 61.730 247.090 63.400 ;
        RECT 345.100 63.210 348.430 64.290 ;
        RECT 276.890 61.830 280.220 62.910 ;
        RECT 141.670 60.030 144.970 61.700 ;
        RECT 276.890 60.160 280.190 61.830 ;
        RECT 345.100 61.540 348.400 63.210 ;
        RECT 378.200 61.640 381.530 62.720 ;
        RECT 378.200 59.970 381.500 61.640 ;
        RECT 6.930 55.440 10.260 56.520 ;
        RECT 6.930 53.770 10.230 55.440 ;
        RECT 108.240 55.250 111.570 56.330 ;
        RECT 243.460 55.380 246.790 56.460 ;
        RECT 22.610 53.020 25.940 54.100 ;
        RECT 108.240 53.580 111.540 55.250 ;
        RECT 22.610 51.350 25.910 53.020 ;
        RECT 123.920 52.830 127.250 53.910 ;
        RECT 243.460 53.710 246.760 55.380 ;
        RECT 344.770 55.190 348.100 56.270 ;
        RECT 259.140 52.960 262.470 54.040 ;
        RECT 344.770 53.520 348.070 55.190 ;
        RECT 123.920 51.160 127.220 52.830 ;
        RECT 259.140 51.290 262.440 52.960 ;
        RECT 360.450 52.770 363.780 53.850 ;
        RECT 360.450 51.100 363.750 52.770 ;
        RECT 7.090 49.040 10.420 50.120 ;
        RECT 7.090 47.370 10.390 49.040 ;
        RECT 108.400 48.850 111.730 49.930 ;
        RECT 243.620 48.980 246.950 50.060 ;
        RECT 108.400 47.180 111.700 48.850 ;
        RECT 243.620 47.310 246.920 48.980 ;
        RECT 344.930 48.790 348.260 49.870 ;
        RECT 344.930 47.120 348.230 48.790 ;
        RECT 57.890 45.870 61.220 46.950 ;
        RECT 57.890 44.200 61.190 45.870 ;
        RECT 159.200 45.680 162.530 46.760 ;
        RECT 294.420 45.810 297.750 46.890 ;
        RECT 159.200 44.010 162.500 45.680 ;
        RECT 294.420 44.140 297.720 45.810 ;
        RECT 395.730 45.620 399.060 46.700 ;
        RECT 395.730 43.950 399.030 45.620 ;
        RECT 7.070 39.790 10.400 40.870 ;
        RECT 7.070 38.120 10.370 39.790 ;
        RECT 108.380 39.600 111.710 40.680 ;
        RECT 243.600 39.730 246.930 40.810 ;
        RECT 22.750 37.370 26.080 38.450 ;
        RECT 108.380 37.930 111.680 39.600 ;
        RECT 22.750 35.700 26.050 37.370 ;
        RECT 124.060 37.180 127.390 38.260 ;
        RECT 243.600 38.060 246.900 39.730 ;
        RECT 344.910 39.540 348.240 40.620 ;
        RECT 259.280 37.310 262.610 38.390 ;
        RECT 344.910 37.870 348.210 39.540 ;
        RECT 124.060 35.510 127.360 37.180 ;
        RECT 259.280 35.640 262.580 37.310 ;
        RECT 360.590 37.120 363.920 38.200 ;
        RECT 360.590 35.450 363.890 37.120 ;
        RECT 7.230 33.390 10.560 34.470 ;
        RECT 7.230 31.720 10.530 33.390 ;
        RECT 108.540 33.200 111.870 34.280 ;
        RECT 243.760 33.330 247.090 34.410 ;
        RECT 40.330 31.820 43.660 32.900 ;
        RECT 40.330 30.150 43.630 31.820 ;
        RECT 108.540 31.530 111.840 33.200 ;
        RECT 141.640 31.630 144.970 32.710 ;
        RECT 243.760 31.660 247.060 33.330 ;
        RECT 345.070 33.140 348.400 34.220 ;
        RECT 276.860 31.760 280.190 32.840 ;
        RECT 141.640 29.960 144.940 31.630 ;
        RECT 276.860 30.090 280.160 31.760 ;
        RECT 345.070 31.470 348.370 33.140 ;
        RECT 378.170 31.570 381.500 32.650 ;
        RECT 378.170 29.900 381.470 31.570 ;
        RECT 6.900 25.370 10.230 26.450 ;
        RECT 6.900 23.700 10.200 25.370 ;
        RECT 108.210 25.180 111.540 26.260 ;
        RECT 243.430 25.310 246.760 26.390 ;
        RECT 22.580 22.950 25.910 24.030 ;
        RECT 108.210 23.510 111.510 25.180 ;
        RECT 22.580 21.280 25.880 22.950 ;
        RECT 123.890 22.760 127.220 23.840 ;
        RECT 243.430 23.640 246.730 25.310 ;
        RECT 344.740 25.120 348.070 26.200 ;
        RECT 259.110 22.890 262.440 23.970 ;
        RECT 344.740 23.450 348.040 25.120 ;
        RECT 123.890 21.090 127.190 22.760 ;
        RECT 259.110 21.220 262.410 22.890 ;
        RECT 360.420 22.700 363.750 23.780 ;
        RECT 360.420 21.030 363.720 22.700 ;
        RECT 7.060 18.970 10.390 20.050 ;
        RECT 7.060 17.300 10.360 18.970 ;
        RECT 108.370 18.780 111.700 19.860 ;
        RECT 243.590 18.910 246.920 19.990 ;
        RECT 108.370 17.110 111.670 18.780 ;
        RECT 243.590 17.240 246.890 18.910 ;
        RECT 344.900 18.720 348.230 19.800 ;
        RECT 344.900 17.050 348.200 18.720 ;
      LAYER li1 ;
        RECT 8.000 250.200 11.190 250.950 ;
        RECT 8.000 250.190 9.300 250.200 ;
        RECT 9.890 250.190 11.190 250.200 ;
        RECT 8.200 249.860 8.450 250.190 ;
        RECT 10.090 249.860 10.340 250.190 ;
        RECT 109.310 250.010 112.500 250.760 ;
        RECT 244.530 250.140 247.720 250.890 ;
        RECT 244.530 250.130 245.830 250.140 ;
        RECT 246.420 250.130 247.720 250.140 ;
        RECT 109.310 250.000 110.610 250.010 ;
        RECT 111.200 250.000 112.500 250.010 ;
        RECT 8.200 248.640 8.460 249.860 ;
        RECT 10.090 248.640 10.350 249.860 ;
        RECT 109.510 249.670 109.760 250.000 ;
        RECT 111.400 249.670 111.650 250.000 ;
        RECT 244.730 249.800 244.980 250.130 ;
        RECT 246.620 249.800 246.870 250.130 ;
        RECT 345.840 249.950 349.030 250.700 ;
        RECT 345.840 249.940 347.140 249.950 ;
        RECT 347.730 249.940 349.030 249.950 ;
        RECT 23.680 247.780 26.870 248.530 ;
        RECT 109.510 248.450 109.770 249.670 ;
        RECT 111.400 248.450 111.660 249.670 ;
        RECT 244.730 248.580 244.990 249.800 ;
        RECT 246.620 248.580 246.880 249.800 ;
        RECT 346.040 249.610 346.290 249.940 ;
        RECT 347.930 249.610 348.180 249.940 ;
        RECT 23.680 247.770 24.980 247.780 ;
        RECT 25.570 247.770 26.870 247.780 ;
        RECT 23.880 247.440 24.130 247.770 ;
        RECT 25.770 247.440 26.020 247.770 ;
        RECT 124.990 247.590 128.180 248.340 ;
        RECT 260.210 247.720 263.400 248.470 ;
        RECT 346.040 248.390 346.300 249.610 ;
        RECT 347.930 248.390 348.190 249.610 ;
        RECT 260.210 247.710 261.510 247.720 ;
        RECT 262.100 247.710 263.400 247.720 ;
        RECT 124.990 247.580 126.290 247.590 ;
        RECT 126.880 247.580 128.180 247.590 ;
        RECT 23.880 246.220 24.140 247.440 ;
        RECT 25.770 246.220 26.030 247.440 ;
        RECT 125.190 247.250 125.440 247.580 ;
        RECT 127.080 247.250 127.330 247.580 ;
        RECT 260.410 247.380 260.660 247.710 ;
        RECT 262.300 247.380 262.550 247.710 ;
        RECT 361.520 247.530 364.710 248.280 ;
        RECT 361.520 247.520 362.820 247.530 ;
        RECT 363.410 247.520 364.710 247.530 ;
        RECT 125.190 246.030 125.450 247.250 ;
        RECT 127.080 246.030 127.340 247.250 ;
        RECT 260.410 246.160 260.670 247.380 ;
        RECT 262.300 246.160 262.560 247.380 ;
        RECT 361.720 247.190 361.970 247.520 ;
        RECT 363.610 247.190 363.860 247.520 ;
        RECT 361.720 245.970 361.980 247.190 ;
        RECT 363.610 245.970 363.870 247.190 ;
        RECT 8.160 243.800 11.350 244.550 ;
        RECT 8.160 243.790 9.460 243.800 ;
        RECT 10.050 243.790 11.350 243.800 ;
        RECT 8.360 243.460 8.610 243.790 ;
        RECT 10.250 243.460 10.500 243.790 ;
        RECT 109.470 243.610 112.660 244.360 ;
        RECT 244.690 243.740 247.880 244.490 ;
        RECT 244.690 243.730 245.990 243.740 ;
        RECT 246.580 243.730 247.880 243.740 ;
        RECT 109.470 243.600 110.770 243.610 ;
        RECT 111.360 243.600 112.660 243.610 ;
        RECT 8.360 242.240 8.620 243.460 ;
        RECT 10.250 242.240 10.510 243.460 ;
        RECT 109.670 243.270 109.920 243.600 ;
        RECT 111.560 243.270 111.810 243.600 ;
        RECT 244.890 243.400 245.140 243.730 ;
        RECT 246.780 243.400 247.030 243.730 ;
        RECT 346.000 243.550 349.190 244.300 ;
        RECT 346.000 243.540 347.300 243.550 ;
        RECT 347.890 243.540 349.190 243.550 ;
        RECT 41.260 242.230 44.450 242.980 ;
        RECT 41.260 242.220 42.560 242.230 ;
        RECT 43.150 242.220 44.450 242.230 ;
        RECT 41.460 241.890 41.710 242.220 ;
        RECT 43.350 241.890 43.600 242.220 ;
        RECT 109.670 242.050 109.930 243.270 ;
        RECT 111.560 242.050 111.820 243.270 ;
        RECT 142.570 242.040 145.760 242.790 ;
        RECT 244.890 242.180 245.150 243.400 ;
        RECT 246.780 242.180 247.040 243.400 ;
        RECT 346.200 243.210 346.450 243.540 ;
        RECT 348.090 243.210 348.340 243.540 ;
        RECT 277.790 242.170 280.980 242.920 ;
        RECT 277.790 242.160 279.090 242.170 ;
        RECT 279.680 242.160 280.980 242.170 ;
        RECT 142.570 242.030 143.870 242.040 ;
        RECT 144.460 242.030 145.760 242.040 ;
        RECT 41.460 240.670 41.720 241.890 ;
        RECT 43.350 240.670 43.610 241.890 ;
        RECT 142.770 241.700 143.020 242.030 ;
        RECT 144.660 241.700 144.910 242.030 ;
        RECT 277.990 241.830 278.240 242.160 ;
        RECT 279.880 241.830 280.130 242.160 ;
        RECT 346.200 241.990 346.460 243.210 ;
        RECT 348.090 241.990 348.350 243.210 ;
        RECT 379.100 241.980 382.290 242.730 ;
        RECT 379.100 241.970 380.400 241.980 ;
        RECT 380.990 241.970 382.290 241.980 ;
        RECT 142.770 240.480 143.030 241.700 ;
        RECT 144.660 240.480 144.920 241.700 ;
        RECT 277.990 240.610 278.250 241.830 ;
        RECT 279.880 240.610 280.140 241.830 ;
        RECT 379.300 241.640 379.550 241.970 ;
        RECT 381.190 241.640 381.440 241.970 ;
        RECT 379.300 240.420 379.560 241.640 ;
        RECT 381.190 240.420 381.450 241.640 ;
        RECT 7.830 235.780 11.020 236.530 ;
        RECT 7.830 235.770 9.130 235.780 ;
        RECT 9.720 235.770 11.020 235.780 ;
        RECT 8.030 235.440 8.280 235.770 ;
        RECT 9.920 235.440 10.170 235.770 ;
        RECT 109.140 235.590 112.330 236.340 ;
        RECT 244.360 235.720 247.550 236.470 ;
        RECT 244.360 235.710 245.660 235.720 ;
        RECT 246.250 235.710 247.550 235.720 ;
        RECT 109.140 235.580 110.440 235.590 ;
        RECT 111.030 235.580 112.330 235.590 ;
        RECT 8.030 234.220 8.290 235.440 ;
        RECT 9.920 234.220 10.180 235.440 ;
        RECT 109.340 235.250 109.590 235.580 ;
        RECT 111.230 235.250 111.480 235.580 ;
        RECT 244.560 235.380 244.810 235.710 ;
        RECT 246.450 235.380 246.700 235.710 ;
        RECT 345.670 235.530 348.860 236.280 ;
        RECT 345.670 235.520 346.970 235.530 ;
        RECT 347.560 235.520 348.860 235.530 ;
        RECT 23.510 233.360 26.700 234.110 ;
        RECT 109.340 234.030 109.600 235.250 ;
        RECT 111.230 234.030 111.490 235.250 ;
        RECT 244.560 234.160 244.820 235.380 ;
        RECT 246.450 234.160 246.710 235.380 ;
        RECT 345.870 235.190 346.120 235.520 ;
        RECT 347.760 235.190 348.010 235.520 ;
        RECT 23.510 233.350 24.810 233.360 ;
        RECT 25.400 233.350 26.700 233.360 ;
        RECT 23.710 233.020 23.960 233.350 ;
        RECT 25.600 233.020 25.850 233.350 ;
        RECT 124.820 233.170 128.010 233.920 ;
        RECT 260.040 233.300 263.230 234.050 ;
        RECT 345.870 233.970 346.130 235.190 ;
        RECT 347.760 233.970 348.020 235.190 ;
        RECT 260.040 233.290 261.340 233.300 ;
        RECT 261.930 233.290 263.230 233.300 ;
        RECT 124.820 233.160 126.120 233.170 ;
        RECT 126.710 233.160 128.010 233.170 ;
        RECT 23.710 231.800 23.970 233.020 ;
        RECT 25.600 231.800 25.860 233.020 ;
        RECT 125.020 232.830 125.270 233.160 ;
        RECT 126.910 232.830 127.160 233.160 ;
        RECT 260.240 232.960 260.490 233.290 ;
        RECT 262.130 232.960 262.380 233.290 ;
        RECT 361.350 233.110 364.540 233.860 ;
        RECT 361.350 233.100 362.650 233.110 ;
        RECT 363.240 233.100 364.540 233.110 ;
        RECT 125.020 231.610 125.280 232.830 ;
        RECT 126.910 231.610 127.170 232.830 ;
        RECT 260.240 231.740 260.500 232.960 ;
        RECT 262.130 231.740 262.390 232.960 ;
        RECT 361.550 232.770 361.800 233.100 ;
        RECT 363.440 232.770 363.690 233.100 ;
        RECT 361.550 231.550 361.810 232.770 ;
        RECT 363.440 231.550 363.700 232.770 ;
        RECT 7.990 229.380 11.180 230.130 ;
        RECT 7.990 229.370 9.290 229.380 ;
        RECT 9.880 229.370 11.180 229.380 ;
        RECT 8.190 229.040 8.440 229.370 ;
        RECT 10.080 229.040 10.330 229.370 ;
        RECT 109.300 229.190 112.490 229.940 ;
        RECT 244.520 229.320 247.710 230.070 ;
        RECT 244.520 229.310 245.820 229.320 ;
        RECT 246.410 229.310 247.710 229.320 ;
        RECT 109.300 229.180 110.600 229.190 ;
        RECT 111.190 229.180 112.490 229.190 ;
        RECT 8.190 227.820 8.450 229.040 ;
        RECT 10.080 227.820 10.340 229.040 ;
        RECT 109.500 228.850 109.750 229.180 ;
        RECT 111.390 228.850 111.640 229.180 ;
        RECT 244.720 228.980 244.970 229.310 ;
        RECT 246.610 228.980 246.860 229.310 ;
        RECT 345.830 229.130 349.020 229.880 ;
        RECT 345.830 229.120 347.130 229.130 ;
        RECT 347.720 229.120 349.020 229.130 ;
        RECT 109.500 227.630 109.760 228.850 ;
        RECT 111.390 227.630 111.650 228.850 ;
        RECT 244.720 227.760 244.980 228.980 ;
        RECT 246.610 227.760 246.870 228.980 ;
        RECT 346.030 228.790 346.280 229.120 ;
        RECT 347.920 228.790 348.170 229.120 ;
        RECT 346.030 227.570 346.290 228.790 ;
        RECT 347.920 227.570 348.180 228.790 ;
        RECT 58.790 226.210 61.980 226.960 ;
        RECT 58.790 226.200 60.090 226.210 ;
        RECT 60.680 226.200 61.980 226.210 ;
        RECT 58.990 225.870 59.240 226.200 ;
        RECT 60.880 225.870 61.130 226.200 ;
        RECT 160.100 226.020 163.290 226.770 ;
        RECT 295.320 226.150 298.510 226.900 ;
        RECT 295.320 226.140 296.620 226.150 ;
        RECT 297.210 226.140 298.510 226.150 ;
        RECT 160.100 226.010 161.400 226.020 ;
        RECT 161.990 226.010 163.290 226.020 ;
        RECT 58.990 224.650 59.250 225.870 ;
        RECT 60.880 224.650 61.140 225.870 ;
        RECT 160.300 225.680 160.550 226.010 ;
        RECT 162.190 225.680 162.440 226.010 ;
        RECT 295.520 225.810 295.770 226.140 ;
        RECT 297.410 225.810 297.660 226.140 ;
        RECT 396.630 225.960 399.820 226.710 ;
        RECT 396.630 225.950 397.930 225.960 ;
        RECT 398.520 225.950 399.820 225.960 ;
        RECT 160.300 224.460 160.560 225.680 ;
        RECT 162.190 224.460 162.450 225.680 ;
        RECT 295.520 224.590 295.780 225.810 ;
        RECT 297.410 224.590 297.670 225.810 ;
        RECT 396.830 225.620 397.080 225.950 ;
        RECT 398.720 225.620 398.970 225.950 ;
        RECT 396.830 224.400 397.090 225.620 ;
        RECT 398.720 224.400 398.980 225.620 ;
        RECT 7.970 220.130 11.160 220.880 ;
        RECT 7.970 220.120 9.270 220.130 ;
        RECT 9.860 220.120 11.160 220.130 ;
        RECT 8.170 219.790 8.420 220.120 ;
        RECT 10.060 219.790 10.310 220.120 ;
        RECT 109.280 219.940 112.470 220.690 ;
        RECT 244.500 220.070 247.690 220.820 ;
        RECT 244.500 220.060 245.800 220.070 ;
        RECT 246.390 220.060 247.690 220.070 ;
        RECT 109.280 219.930 110.580 219.940 ;
        RECT 111.170 219.930 112.470 219.940 ;
        RECT 8.170 218.570 8.430 219.790 ;
        RECT 10.060 218.570 10.320 219.790 ;
        RECT 109.480 219.600 109.730 219.930 ;
        RECT 111.370 219.600 111.620 219.930 ;
        RECT 244.700 219.730 244.950 220.060 ;
        RECT 246.590 219.730 246.840 220.060 ;
        RECT 345.810 219.880 349.000 220.630 ;
        RECT 345.810 219.870 347.110 219.880 ;
        RECT 347.700 219.870 349.000 219.880 ;
        RECT 23.650 217.710 26.840 218.460 ;
        RECT 109.480 218.380 109.740 219.600 ;
        RECT 111.370 218.380 111.630 219.600 ;
        RECT 244.700 218.510 244.960 219.730 ;
        RECT 246.590 218.510 246.850 219.730 ;
        RECT 346.010 219.540 346.260 219.870 ;
        RECT 347.900 219.540 348.150 219.870 ;
        RECT 23.650 217.700 24.950 217.710 ;
        RECT 25.540 217.700 26.840 217.710 ;
        RECT 23.850 217.370 24.100 217.700 ;
        RECT 25.740 217.370 25.990 217.700 ;
        RECT 124.960 217.520 128.150 218.270 ;
        RECT 260.180 217.650 263.370 218.400 ;
        RECT 346.010 218.320 346.270 219.540 ;
        RECT 347.900 218.320 348.160 219.540 ;
        RECT 260.180 217.640 261.480 217.650 ;
        RECT 262.070 217.640 263.370 217.650 ;
        RECT 124.960 217.510 126.260 217.520 ;
        RECT 126.850 217.510 128.150 217.520 ;
        RECT 23.850 216.150 24.110 217.370 ;
        RECT 25.740 216.150 26.000 217.370 ;
        RECT 125.160 217.180 125.410 217.510 ;
        RECT 127.050 217.180 127.300 217.510 ;
        RECT 260.380 217.310 260.630 217.640 ;
        RECT 262.270 217.310 262.520 217.640 ;
        RECT 361.490 217.460 364.680 218.210 ;
        RECT 361.490 217.450 362.790 217.460 ;
        RECT 363.380 217.450 364.680 217.460 ;
        RECT 125.160 215.960 125.420 217.180 ;
        RECT 127.050 215.960 127.310 217.180 ;
        RECT 260.380 216.090 260.640 217.310 ;
        RECT 262.270 216.090 262.530 217.310 ;
        RECT 361.690 217.120 361.940 217.450 ;
        RECT 363.580 217.120 363.830 217.450 ;
        RECT 361.690 215.900 361.950 217.120 ;
        RECT 363.580 215.900 363.840 217.120 ;
        RECT 8.130 213.730 11.320 214.480 ;
        RECT 8.130 213.720 9.430 213.730 ;
        RECT 10.020 213.720 11.320 213.730 ;
        RECT 8.330 213.390 8.580 213.720 ;
        RECT 10.220 213.390 10.470 213.720 ;
        RECT 109.440 213.540 112.630 214.290 ;
        RECT 244.660 213.670 247.850 214.420 ;
        RECT 244.660 213.660 245.960 213.670 ;
        RECT 246.550 213.660 247.850 213.670 ;
        RECT 109.440 213.530 110.740 213.540 ;
        RECT 111.330 213.530 112.630 213.540 ;
        RECT 8.330 212.170 8.590 213.390 ;
        RECT 10.220 212.170 10.480 213.390 ;
        RECT 109.640 213.200 109.890 213.530 ;
        RECT 111.530 213.200 111.780 213.530 ;
        RECT 244.860 213.330 245.110 213.660 ;
        RECT 246.750 213.330 247.000 213.660 ;
        RECT 345.970 213.480 349.160 214.230 ;
        RECT 345.970 213.470 347.270 213.480 ;
        RECT 347.860 213.470 349.160 213.480 ;
        RECT 41.230 212.160 44.420 212.910 ;
        RECT 41.230 212.150 42.530 212.160 ;
        RECT 43.120 212.150 44.420 212.160 ;
        RECT 41.430 211.820 41.680 212.150 ;
        RECT 43.320 211.820 43.570 212.150 ;
        RECT 109.640 211.980 109.900 213.200 ;
        RECT 111.530 211.980 111.790 213.200 ;
        RECT 142.540 211.970 145.730 212.720 ;
        RECT 244.860 212.110 245.120 213.330 ;
        RECT 246.750 212.110 247.010 213.330 ;
        RECT 346.170 213.140 346.420 213.470 ;
        RECT 348.060 213.140 348.310 213.470 ;
        RECT 277.760 212.100 280.950 212.850 ;
        RECT 277.760 212.090 279.060 212.100 ;
        RECT 279.650 212.090 280.950 212.100 ;
        RECT 142.540 211.960 143.840 211.970 ;
        RECT 144.430 211.960 145.730 211.970 ;
        RECT 41.430 210.600 41.690 211.820 ;
        RECT 43.320 210.600 43.580 211.820 ;
        RECT 142.740 211.630 142.990 211.960 ;
        RECT 144.630 211.630 144.880 211.960 ;
        RECT 277.960 211.760 278.210 212.090 ;
        RECT 279.850 211.760 280.100 212.090 ;
        RECT 346.170 211.920 346.430 213.140 ;
        RECT 348.060 211.920 348.320 213.140 ;
        RECT 379.070 211.910 382.260 212.660 ;
        RECT 379.070 211.900 380.370 211.910 ;
        RECT 380.960 211.900 382.260 211.910 ;
        RECT 142.740 210.410 143.000 211.630 ;
        RECT 144.630 210.410 144.890 211.630 ;
        RECT 277.960 210.540 278.220 211.760 ;
        RECT 279.850 210.540 280.110 211.760 ;
        RECT 379.270 211.570 379.520 211.900 ;
        RECT 381.160 211.570 381.410 211.900 ;
        RECT 379.270 210.350 379.530 211.570 ;
        RECT 381.160 210.350 381.420 211.570 ;
        RECT 7.800 205.710 10.990 206.460 ;
        RECT 7.800 205.700 9.100 205.710 ;
        RECT 9.690 205.700 10.990 205.710 ;
        RECT 8.000 205.370 8.250 205.700 ;
        RECT 9.890 205.370 10.140 205.700 ;
        RECT 109.110 205.520 112.300 206.270 ;
        RECT 244.330 205.650 247.520 206.400 ;
        RECT 244.330 205.640 245.630 205.650 ;
        RECT 246.220 205.640 247.520 205.650 ;
        RECT 109.110 205.510 110.410 205.520 ;
        RECT 111.000 205.510 112.300 205.520 ;
        RECT 8.000 204.150 8.260 205.370 ;
        RECT 9.890 204.150 10.150 205.370 ;
        RECT 109.310 205.180 109.560 205.510 ;
        RECT 111.200 205.180 111.450 205.510 ;
        RECT 244.530 205.310 244.780 205.640 ;
        RECT 246.420 205.310 246.670 205.640 ;
        RECT 345.640 205.460 348.830 206.210 ;
        RECT 345.640 205.450 346.940 205.460 ;
        RECT 347.530 205.450 348.830 205.460 ;
        RECT 23.480 203.290 26.670 204.040 ;
        RECT 109.310 203.960 109.570 205.180 ;
        RECT 111.200 203.960 111.460 205.180 ;
        RECT 244.530 204.090 244.790 205.310 ;
        RECT 246.420 204.090 246.680 205.310 ;
        RECT 345.840 205.120 346.090 205.450 ;
        RECT 347.730 205.120 347.980 205.450 ;
        RECT 23.480 203.280 24.780 203.290 ;
        RECT 25.370 203.280 26.670 203.290 ;
        RECT 23.680 202.950 23.930 203.280 ;
        RECT 25.570 202.950 25.820 203.280 ;
        RECT 124.790 203.100 127.980 203.850 ;
        RECT 260.010 203.230 263.200 203.980 ;
        RECT 345.840 203.900 346.100 205.120 ;
        RECT 347.730 203.900 347.990 205.120 ;
        RECT 260.010 203.220 261.310 203.230 ;
        RECT 261.900 203.220 263.200 203.230 ;
        RECT 124.790 203.090 126.090 203.100 ;
        RECT 126.680 203.090 127.980 203.100 ;
        RECT 23.680 201.730 23.940 202.950 ;
        RECT 25.570 201.730 25.830 202.950 ;
        RECT 124.990 202.760 125.240 203.090 ;
        RECT 126.880 202.760 127.130 203.090 ;
        RECT 260.210 202.890 260.460 203.220 ;
        RECT 262.100 202.890 262.350 203.220 ;
        RECT 361.320 203.040 364.510 203.790 ;
        RECT 361.320 203.030 362.620 203.040 ;
        RECT 363.210 203.030 364.510 203.040 ;
        RECT 124.990 201.540 125.250 202.760 ;
        RECT 126.880 201.540 127.140 202.760 ;
        RECT 260.210 201.670 260.470 202.890 ;
        RECT 262.100 201.670 262.360 202.890 ;
        RECT 361.520 202.700 361.770 203.030 ;
        RECT 363.410 202.700 363.660 203.030 ;
        RECT 361.520 201.480 361.780 202.700 ;
        RECT 363.410 201.480 363.670 202.700 ;
        RECT 7.960 199.310 11.150 200.060 ;
        RECT 72.990 199.920 76.180 200.670 ;
        RECT 72.990 199.910 74.290 199.920 ;
        RECT 74.880 199.910 76.180 199.920 ;
        RECT 7.960 199.300 9.260 199.310 ;
        RECT 9.850 199.300 11.150 199.310 ;
        RECT 73.190 199.580 73.440 199.910 ;
        RECT 75.080 199.580 75.330 199.910 ;
        RECT 8.160 198.970 8.410 199.300 ;
        RECT 10.050 198.970 10.300 199.300 ;
        RECT 8.160 197.750 8.420 198.970 ;
        RECT 10.050 197.750 10.310 198.970 ;
        RECT 73.190 198.360 73.450 199.580 ;
        RECT 75.080 198.360 75.340 199.580 ;
        RECT 109.270 199.120 112.460 199.870 ;
        RECT 174.300 199.730 177.490 200.480 ;
        RECT 174.300 199.720 175.600 199.730 ;
        RECT 176.190 199.720 177.490 199.730 ;
        RECT 109.270 199.110 110.570 199.120 ;
        RECT 111.160 199.110 112.460 199.120 ;
        RECT 174.500 199.390 174.750 199.720 ;
        RECT 176.390 199.390 176.640 199.720 ;
        RECT 109.470 198.780 109.720 199.110 ;
        RECT 111.360 198.780 111.610 199.110 ;
        RECT 109.470 197.560 109.730 198.780 ;
        RECT 111.360 197.560 111.620 198.780 ;
        RECT 174.500 198.170 174.760 199.390 ;
        RECT 176.390 198.170 176.650 199.390 ;
        RECT 244.490 199.250 247.680 200.000 ;
        RECT 309.520 199.860 312.710 200.610 ;
        RECT 309.520 199.850 310.820 199.860 ;
        RECT 311.410 199.850 312.710 199.860 ;
        RECT 244.490 199.240 245.790 199.250 ;
        RECT 246.380 199.240 247.680 199.250 ;
        RECT 309.720 199.520 309.970 199.850 ;
        RECT 311.610 199.520 311.860 199.850 ;
        RECT 244.690 198.910 244.940 199.240 ;
        RECT 246.580 198.910 246.830 199.240 ;
        RECT 244.690 197.690 244.950 198.910 ;
        RECT 246.580 197.690 246.840 198.910 ;
        RECT 309.720 198.300 309.980 199.520 ;
        RECT 311.610 198.300 311.870 199.520 ;
        RECT 345.800 199.060 348.990 199.810 ;
        RECT 410.830 199.670 414.020 200.420 ;
        RECT 410.830 199.660 412.130 199.670 ;
        RECT 412.720 199.660 414.020 199.670 ;
        RECT 345.800 199.050 347.100 199.060 ;
        RECT 347.690 199.050 348.990 199.060 ;
        RECT 411.030 199.330 411.280 199.660 ;
        RECT 412.920 199.330 413.170 199.660 ;
        RECT 346.000 198.720 346.250 199.050 ;
        RECT 347.890 198.720 348.140 199.050 ;
        RECT 346.000 197.500 346.260 198.720 ;
        RECT 347.890 197.500 348.150 198.720 ;
        RECT 411.030 198.110 411.290 199.330 ;
        RECT 412.920 198.110 413.180 199.330 ;
        RECT 7.650 190.280 10.840 191.030 ;
        RECT 7.650 190.270 8.950 190.280 ;
        RECT 9.540 190.270 10.840 190.280 ;
        RECT 7.850 189.940 8.100 190.270 ;
        RECT 9.740 189.940 9.990 190.270 ;
        RECT 108.960 190.090 112.150 190.840 ;
        RECT 244.180 190.220 247.370 190.970 ;
        RECT 244.180 190.210 245.480 190.220 ;
        RECT 246.070 190.210 247.370 190.220 ;
        RECT 108.960 190.080 110.260 190.090 ;
        RECT 110.850 190.080 112.150 190.090 ;
        RECT 7.850 188.720 8.110 189.940 ;
        RECT 9.740 188.720 10.000 189.940 ;
        RECT 109.160 189.750 109.410 190.080 ;
        RECT 111.050 189.750 111.300 190.080 ;
        RECT 244.380 189.880 244.630 190.210 ;
        RECT 246.270 189.880 246.520 190.210 ;
        RECT 345.490 190.030 348.680 190.780 ;
        RECT 345.490 190.020 346.790 190.030 ;
        RECT 347.380 190.020 348.680 190.030 ;
        RECT 23.330 187.860 26.520 188.610 ;
        RECT 109.160 188.530 109.420 189.750 ;
        RECT 111.050 188.530 111.310 189.750 ;
        RECT 244.380 188.660 244.640 189.880 ;
        RECT 246.270 188.660 246.530 189.880 ;
        RECT 345.690 189.690 345.940 190.020 ;
        RECT 347.580 189.690 347.830 190.020 ;
        RECT 23.330 187.850 24.630 187.860 ;
        RECT 25.220 187.850 26.520 187.860 ;
        RECT 23.530 187.520 23.780 187.850 ;
        RECT 25.420 187.520 25.670 187.850 ;
        RECT 124.640 187.670 127.830 188.420 ;
        RECT 259.860 187.800 263.050 188.550 ;
        RECT 345.690 188.470 345.950 189.690 ;
        RECT 347.580 188.470 347.840 189.690 ;
        RECT 259.860 187.790 261.160 187.800 ;
        RECT 261.750 187.790 263.050 187.800 ;
        RECT 124.640 187.660 125.940 187.670 ;
        RECT 126.530 187.660 127.830 187.670 ;
        RECT 23.530 186.300 23.790 187.520 ;
        RECT 25.420 186.300 25.680 187.520 ;
        RECT 124.840 187.330 125.090 187.660 ;
        RECT 126.730 187.330 126.980 187.660 ;
        RECT 260.060 187.460 260.310 187.790 ;
        RECT 261.950 187.460 262.200 187.790 ;
        RECT 361.170 187.610 364.360 188.360 ;
        RECT 361.170 187.600 362.470 187.610 ;
        RECT 363.060 187.600 364.360 187.610 ;
        RECT 124.840 186.110 125.100 187.330 ;
        RECT 126.730 186.110 126.990 187.330 ;
        RECT 260.060 186.240 260.320 187.460 ;
        RECT 261.950 186.240 262.210 187.460 ;
        RECT 361.370 187.270 361.620 187.600 ;
        RECT 363.260 187.270 363.510 187.600 ;
        RECT 361.370 186.050 361.630 187.270 ;
        RECT 363.260 186.050 363.520 187.270 ;
        RECT 7.810 183.880 11.000 184.630 ;
        RECT 7.810 183.870 9.110 183.880 ;
        RECT 9.700 183.870 11.000 183.880 ;
        RECT 8.010 183.540 8.260 183.870 ;
        RECT 9.900 183.540 10.150 183.870 ;
        RECT 109.120 183.690 112.310 184.440 ;
        RECT 244.340 183.820 247.530 184.570 ;
        RECT 244.340 183.810 245.640 183.820 ;
        RECT 246.230 183.810 247.530 183.820 ;
        RECT 109.120 183.680 110.420 183.690 ;
        RECT 111.010 183.680 112.310 183.690 ;
        RECT 8.010 182.320 8.270 183.540 ;
        RECT 9.900 182.320 10.160 183.540 ;
        RECT 109.320 183.350 109.570 183.680 ;
        RECT 111.210 183.350 111.460 183.680 ;
        RECT 244.540 183.480 244.790 183.810 ;
        RECT 246.430 183.480 246.680 183.810 ;
        RECT 345.650 183.630 348.840 184.380 ;
        RECT 345.650 183.620 346.950 183.630 ;
        RECT 347.540 183.620 348.840 183.630 ;
        RECT 40.910 182.310 44.100 183.060 ;
        RECT 40.910 182.300 42.210 182.310 ;
        RECT 42.800 182.300 44.100 182.310 ;
        RECT 41.110 181.970 41.360 182.300 ;
        RECT 43.000 181.970 43.250 182.300 ;
        RECT 109.320 182.130 109.580 183.350 ;
        RECT 111.210 182.130 111.470 183.350 ;
        RECT 142.220 182.120 145.410 182.870 ;
        RECT 244.540 182.260 244.800 183.480 ;
        RECT 246.430 182.260 246.690 183.480 ;
        RECT 345.850 183.290 346.100 183.620 ;
        RECT 347.740 183.290 347.990 183.620 ;
        RECT 277.440 182.250 280.630 183.000 ;
        RECT 277.440 182.240 278.740 182.250 ;
        RECT 279.330 182.240 280.630 182.250 ;
        RECT 142.220 182.110 143.520 182.120 ;
        RECT 144.110 182.110 145.410 182.120 ;
        RECT 41.110 180.750 41.370 181.970 ;
        RECT 43.000 180.750 43.260 181.970 ;
        RECT 142.420 181.780 142.670 182.110 ;
        RECT 144.310 181.780 144.560 182.110 ;
        RECT 277.640 181.910 277.890 182.240 ;
        RECT 279.530 181.910 279.780 182.240 ;
        RECT 345.850 182.070 346.110 183.290 ;
        RECT 347.740 182.070 348.000 183.290 ;
        RECT 378.750 182.060 381.940 182.810 ;
        RECT 378.750 182.050 380.050 182.060 ;
        RECT 380.640 182.050 381.940 182.060 ;
        RECT 142.420 180.560 142.680 181.780 ;
        RECT 144.310 180.560 144.570 181.780 ;
        RECT 277.640 180.690 277.900 181.910 ;
        RECT 279.530 180.690 279.790 181.910 ;
        RECT 378.950 181.720 379.200 182.050 ;
        RECT 380.840 181.720 381.090 182.050 ;
        RECT 378.950 180.500 379.210 181.720 ;
        RECT 380.840 180.500 381.100 181.720 ;
        RECT 7.480 175.860 10.670 176.610 ;
        RECT 7.480 175.850 8.780 175.860 ;
        RECT 9.370 175.850 10.670 175.860 ;
        RECT 7.680 175.520 7.930 175.850 ;
        RECT 9.570 175.520 9.820 175.850 ;
        RECT 108.790 175.670 111.980 176.420 ;
        RECT 244.010 175.800 247.200 176.550 ;
        RECT 244.010 175.790 245.310 175.800 ;
        RECT 245.900 175.790 247.200 175.800 ;
        RECT 108.790 175.660 110.090 175.670 ;
        RECT 110.680 175.660 111.980 175.670 ;
        RECT 7.680 174.300 7.940 175.520 ;
        RECT 9.570 174.300 9.830 175.520 ;
        RECT 108.990 175.330 109.240 175.660 ;
        RECT 110.880 175.330 111.130 175.660 ;
        RECT 244.210 175.460 244.460 175.790 ;
        RECT 246.100 175.460 246.350 175.790 ;
        RECT 345.320 175.610 348.510 176.360 ;
        RECT 345.320 175.600 346.620 175.610 ;
        RECT 347.210 175.600 348.510 175.610 ;
        RECT 23.160 173.440 26.350 174.190 ;
        RECT 108.990 174.110 109.250 175.330 ;
        RECT 110.880 174.110 111.140 175.330 ;
        RECT 244.210 174.240 244.470 175.460 ;
        RECT 246.100 174.240 246.360 175.460 ;
        RECT 345.520 175.270 345.770 175.600 ;
        RECT 347.410 175.270 347.660 175.600 ;
        RECT 23.160 173.430 24.460 173.440 ;
        RECT 25.050 173.430 26.350 173.440 ;
        RECT 23.360 173.100 23.610 173.430 ;
        RECT 25.250 173.100 25.500 173.430 ;
        RECT 124.470 173.250 127.660 174.000 ;
        RECT 259.690 173.380 262.880 174.130 ;
        RECT 345.520 174.050 345.780 175.270 ;
        RECT 347.410 174.050 347.670 175.270 ;
        RECT 259.690 173.370 260.990 173.380 ;
        RECT 261.580 173.370 262.880 173.380 ;
        RECT 124.470 173.240 125.770 173.250 ;
        RECT 126.360 173.240 127.660 173.250 ;
        RECT 23.360 171.880 23.620 173.100 ;
        RECT 25.250 171.880 25.510 173.100 ;
        RECT 124.670 172.910 124.920 173.240 ;
        RECT 126.560 172.910 126.810 173.240 ;
        RECT 259.890 173.040 260.140 173.370 ;
        RECT 261.780 173.040 262.030 173.370 ;
        RECT 361.000 173.190 364.190 173.940 ;
        RECT 361.000 173.180 362.300 173.190 ;
        RECT 362.890 173.180 364.190 173.190 ;
        RECT 124.670 171.690 124.930 172.910 ;
        RECT 126.560 171.690 126.820 172.910 ;
        RECT 259.890 171.820 260.150 173.040 ;
        RECT 261.780 171.820 262.040 173.040 ;
        RECT 361.200 172.850 361.450 173.180 ;
        RECT 363.090 172.850 363.340 173.180 ;
        RECT 361.200 171.630 361.460 172.850 ;
        RECT 363.090 171.630 363.350 172.850 ;
        RECT 7.640 169.460 10.830 170.210 ;
        RECT 7.640 169.450 8.940 169.460 ;
        RECT 9.530 169.450 10.830 169.460 ;
        RECT 7.840 169.120 8.090 169.450 ;
        RECT 9.730 169.120 9.980 169.450 ;
        RECT 108.950 169.270 112.140 170.020 ;
        RECT 244.170 169.400 247.360 170.150 ;
        RECT 244.170 169.390 245.470 169.400 ;
        RECT 246.060 169.390 247.360 169.400 ;
        RECT 108.950 169.260 110.250 169.270 ;
        RECT 110.840 169.260 112.140 169.270 ;
        RECT 7.840 167.900 8.100 169.120 ;
        RECT 9.730 167.900 9.990 169.120 ;
        RECT 109.150 168.930 109.400 169.260 ;
        RECT 111.040 168.930 111.290 169.260 ;
        RECT 244.370 169.060 244.620 169.390 ;
        RECT 246.260 169.060 246.510 169.390 ;
        RECT 345.480 169.210 348.670 169.960 ;
        RECT 345.480 169.200 346.780 169.210 ;
        RECT 347.370 169.200 348.670 169.210 ;
        RECT 109.150 167.710 109.410 168.930 ;
        RECT 111.040 167.710 111.300 168.930 ;
        RECT 244.370 167.840 244.630 169.060 ;
        RECT 246.260 167.840 246.520 169.060 ;
        RECT 345.680 168.870 345.930 169.200 ;
        RECT 347.570 168.870 347.820 169.200 ;
        RECT 345.680 167.650 345.940 168.870 ;
        RECT 347.570 167.650 347.830 168.870 ;
        RECT 58.440 166.290 61.630 167.040 ;
        RECT 58.440 166.280 59.740 166.290 ;
        RECT 60.330 166.280 61.630 166.290 ;
        RECT 58.640 165.950 58.890 166.280 ;
        RECT 60.530 165.950 60.780 166.280 ;
        RECT 159.750 166.100 162.940 166.850 ;
        RECT 294.970 166.230 298.160 166.980 ;
        RECT 294.970 166.220 296.270 166.230 ;
        RECT 296.860 166.220 298.160 166.230 ;
        RECT 159.750 166.090 161.050 166.100 ;
        RECT 161.640 166.090 162.940 166.100 ;
        RECT 58.640 164.730 58.900 165.950 ;
        RECT 60.530 164.730 60.790 165.950 ;
        RECT 159.950 165.760 160.200 166.090 ;
        RECT 161.840 165.760 162.090 166.090 ;
        RECT 295.170 165.890 295.420 166.220 ;
        RECT 297.060 165.890 297.310 166.220 ;
        RECT 396.280 166.040 399.470 166.790 ;
        RECT 396.280 166.030 397.580 166.040 ;
        RECT 398.170 166.030 399.470 166.040 ;
        RECT 159.950 164.540 160.210 165.760 ;
        RECT 161.840 164.540 162.100 165.760 ;
        RECT 295.170 164.670 295.430 165.890 ;
        RECT 297.060 164.670 297.320 165.890 ;
        RECT 396.480 165.700 396.730 166.030 ;
        RECT 398.370 165.700 398.620 166.030 ;
        RECT 396.480 164.480 396.740 165.700 ;
        RECT 398.370 164.480 398.630 165.700 ;
        RECT 7.620 160.210 10.810 160.960 ;
        RECT 7.620 160.200 8.920 160.210 ;
        RECT 9.510 160.200 10.810 160.210 ;
        RECT 7.820 159.870 8.070 160.200 ;
        RECT 9.710 159.870 9.960 160.200 ;
        RECT 108.930 160.020 112.120 160.770 ;
        RECT 244.150 160.150 247.340 160.900 ;
        RECT 244.150 160.140 245.450 160.150 ;
        RECT 246.040 160.140 247.340 160.150 ;
        RECT 108.930 160.010 110.230 160.020 ;
        RECT 110.820 160.010 112.120 160.020 ;
        RECT 7.820 158.650 8.080 159.870 ;
        RECT 9.710 158.650 9.970 159.870 ;
        RECT 109.130 159.680 109.380 160.010 ;
        RECT 111.020 159.680 111.270 160.010 ;
        RECT 244.350 159.810 244.600 160.140 ;
        RECT 246.240 159.810 246.490 160.140 ;
        RECT 345.460 159.960 348.650 160.710 ;
        RECT 345.460 159.950 346.760 159.960 ;
        RECT 347.350 159.950 348.650 159.960 ;
        RECT 23.300 157.790 26.490 158.540 ;
        RECT 109.130 158.460 109.390 159.680 ;
        RECT 111.020 158.460 111.280 159.680 ;
        RECT 244.350 158.590 244.610 159.810 ;
        RECT 246.240 158.590 246.500 159.810 ;
        RECT 345.660 159.620 345.910 159.950 ;
        RECT 347.550 159.620 347.800 159.950 ;
        RECT 23.300 157.780 24.600 157.790 ;
        RECT 25.190 157.780 26.490 157.790 ;
        RECT 23.500 157.450 23.750 157.780 ;
        RECT 25.390 157.450 25.640 157.780 ;
        RECT 124.610 157.600 127.800 158.350 ;
        RECT 259.830 157.730 263.020 158.480 ;
        RECT 345.660 158.400 345.920 159.620 ;
        RECT 347.550 158.400 347.810 159.620 ;
        RECT 259.830 157.720 261.130 157.730 ;
        RECT 261.720 157.720 263.020 157.730 ;
        RECT 124.610 157.590 125.910 157.600 ;
        RECT 126.500 157.590 127.800 157.600 ;
        RECT 23.500 156.230 23.760 157.450 ;
        RECT 25.390 156.230 25.650 157.450 ;
        RECT 124.810 157.260 125.060 157.590 ;
        RECT 126.700 157.260 126.950 157.590 ;
        RECT 260.030 157.390 260.280 157.720 ;
        RECT 261.920 157.390 262.170 157.720 ;
        RECT 361.140 157.540 364.330 158.290 ;
        RECT 361.140 157.530 362.440 157.540 ;
        RECT 363.030 157.530 364.330 157.540 ;
        RECT 124.810 156.040 125.070 157.260 ;
        RECT 126.700 156.040 126.960 157.260 ;
        RECT 260.030 156.170 260.290 157.390 ;
        RECT 261.920 156.170 262.180 157.390 ;
        RECT 361.340 157.200 361.590 157.530 ;
        RECT 363.230 157.200 363.480 157.530 ;
        RECT 361.340 155.980 361.600 157.200 ;
        RECT 363.230 155.980 363.490 157.200 ;
        RECT 7.780 153.810 10.970 154.560 ;
        RECT 7.780 153.800 9.080 153.810 ;
        RECT 9.670 153.800 10.970 153.810 ;
        RECT 7.980 153.470 8.230 153.800 ;
        RECT 9.870 153.470 10.120 153.800 ;
        RECT 109.090 153.620 112.280 154.370 ;
        RECT 244.310 153.750 247.500 154.500 ;
        RECT 244.310 153.740 245.610 153.750 ;
        RECT 246.200 153.740 247.500 153.750 ;
        RECT 109.090 153.610 110.390 153.620 ;
        RECT 110.980 153.610 112.280 153.620 ;
        RECT 7.980 152.250 8.240 153.470 ;
        RECT 9.870 152.250 10.130 153.470 ;
        RECT 109.290 153.280 109.540 153.610 ;
        RECT 111.180 153.280 111.430 153.610 ;
        RECT 244.510 153.410 244.760 153.740 ;
        RECT 246.400 153.410 246.650 153.740 ;
        RECT 345.620 153.560 348.810 154.310 ;
        RECT 345.620 153.550 346.920 153.560 ;
        RECT 347.510 153.550 348.810 153.560 ;
        RECT 40.880 152.240 44.070 152.990 ;
        RECT 40.880 152.230 42.180 152.240 ;
        RECT 42.770 152.230 44.070 152.240 ;
        RECT 41.080 151.900 41.330 152.230 ;
        RECT 42.970 151.900 43.220 152.230 ;
        RECT 109.290 152.060 109.550 153.280 ;
        RECT 111.180 152.060 111.440 153.280 ;
        RECT 142.190 152.050 145.380 152.800 ;
        RECT 244.510 152.190 244.770 153.410 ;
        RECT 246.400 152.190 246.660 153.410 ;
        RECT 345.820 153.220 346.070 153.550 ;
        RECT 347.710 153.220 347.960 153.550 ;
        RECT 277.410 152.180 280.600 152.930 ;
        RECT 277.410 152.170 278.710 152.180 ;
        RECT 279.300 152.170 280.600 152.180 ;
        RECT 142.190 152.040 143.490 152.050 ;
        RECT 144.080 152.040 145.380 152.050 ;
        RECT 41.080 150.680 41.340 151.900 ;
        RECT 42.970 150.680 43.230 151.900 ;
        RECT 142.390 151.710 142.640 152.040 ;
        RECT 144.280 151.710 144.530 152.040 ;
        RECT 277.610 151.840 277.860 152.170 ;
        RECT 279.500 151.840 279.750 152.170 ;
        RECT 345.820 152.000 346.080 153.220 ;
        RECT 347.710 152.000 347.970 153.220 ;
        RECT 378.720 151.990 381.910 152.740 ;
        RECT 378.720 151.980 380.020 151.990 ;
        RECT 380.610 151.980 381.910 151.990 ;
        RECT 142.390 150.490 142.650 151.710 ;
        RECT 144.280 150.490 144.540 151.710 ;
        RECT 277.610 150.620 277.870 151.840 ;
        RECT 279.500 150.620 279.760 151.840 ;
        RECT 378.920 151.650 379.170 151.980 ;
        RECT 380.810 151.650 381.060 151.980 ;
        RECT 378.920 150.430 379.180 151.650 ;
        RECT 380.810 150.430 381.070 151.650 ;
        RECT 7.450 145.790 10.640 146.540 ;
        RECT 7.450 145.780 8.750 145.790 ;
        RECT 9.340 145.780 10.640 145.790 ;
        RECT 7.650 145.450 7.900 145.780 ;
        RECT 9.540 145.450 9.790 145.780 ;
        RECT 108.760 145.600 111.950 146.350 ;
        RECT 243.980 145.730 247.170 146.480 ;
        RECT 243.980 145.720 245.280 145.730 ;
        RECT 245.870 145.720 247.170 145.730 ;
        RECT 108.760 145.590 110.060 145.600 ;
        RECT 110.650 145.590 111.950 145.600 ;
        RECT 7.650 144.230 7.910 145.450 ;
        RECT 9.540 144.230 9.800 145.450 ;
        RECT 108.960 145.260 109.210 145.590 ;
        RECT 110.850 145.260 111.100 145.590 ;
        RECT 244.180 145.390 244.430 145.720 ;
        RECT 246.070 145.390 246.320 145.720 ;
        RECT 345.290 145.540 348.480 146.290 ;
        RECT 345.290 145.530 346.590 145.540 ;
        RECT 347.180 145.530 348.480 145.540 ;
        RECT 23.130 143.370 26.320 144.120 ;
        RECT 108.960 144.040 109.220 145.260 ;
        RECT 110.850 144.040 111.110 145.260 ;
        RECT 244.180 144.170 244.440 145.390 ;
        RECT 246.070 144.170 246.330 145.390 ;
        RECT 345.490 145.200 345.740 145.530 ;
        RECT 347.380 145.200 347.630 145.530 ;
        RECT 23.130 143.360 24.430 143.370 ;
        RECT 25.020 143.360 26.320 143.370 ;
        RECT 23.330 143.030 23.580 143.360 ;
        RECT 25.220 143.030 25.470 143.360 ;
        RECT 124.440 143.180 127.630 143.930 ;
        RECT 259.660 143.310 262.850 144.060 ;
        RECT 345.490 143.980 345.750 145.200 ;
        RECT 347.380 143.980 347.640 145.200 ;
        RECT 259.660 143.300 260.960 143.310 ;
        RECT 261.550 143.300 262.850 143.310 ;
        RECT 124.440 143.170 125.740 143.180 ;
        RECT 126.330 143.170 127.630 143.180 ;
        RECT 23.330 141.810 23.590 143.030 ;
        RECT 25.220 141.810 25.480 143.030 ;
        RECT 124.640 142.840 124.890 143.170 ;
        RECT 126.530 142.840 126.780 143.170 ;
        RECT 259.860 142.970 260.110 143.300 ;
        RECT 261.750 142.970 262.000 143.300 ;
        RECT 360.970 143.120 364.160 143.870 ;
        RECT 360.970 143.110 362.270 143.120 ;
        RECT 362.860 143.110 364.160 143.120 ;
        RECT 124.640 141.620 124.900 142.840 ;
        RECT 126.530 141.620 126.790 142.840 ;
        RECT 259.860 141.750 260.120 142.970 ;
        RECT 261.750 141.750 262.010 142.970 ;
        RECT 361.170 142.780 361.420 143.110 ;
        RECT 363.060 142.780 363.310 143.110 ;
        RECT 361.170 141.560 361.430 142.780 ;
        RECT 363.060 141.560 363.320 142.780 ;
        RECT 7.610 139.390 10.800 140.140 ;
        RECT 7.610 139.380 8.910 139.390 ;
        RECT 9.500 139.380 10.800 139.390 ;
        RECT 7.810 139.050 8.060 139.380 ;
        RECT 9.700 139.050 9.950 139.380 ;
        RECT 108.920 139.200 112.110 139.950 ;
        RECT 108.920 139.190 110.220 139.200 ;
        RECT 110.810 139.190 112.110 139.200 ;
        RECT 7.810 137.830 8.070 139.050 ;
        RECT 9.700 137.830 9.960 139.050 ;
        RECT 109.120 138.860 109.370 139.190 ;
        RECT 111.010 138.860 111.260 139.190 ;
        RECT 216.910 138.920 220.100 139.670 ;
        RECT 244.140 139.330 247.330 140.080 ;
        RECT 244.140 139.320 245.440 139.330 ;
        RECT 246.030 139.320 247.330 139.330 ;
        RECT 216.910 138.910 218.210 138.920 ;
        RECT 218.800 138.910 220.100 138.920 ;
        RECT 244.340 138.990 244.590 139.320 ;
        RECT 246.230 138.990 246.480 139.320 ;
        RECT 345.450 139.140 348.640 139.890 ;
        RECT 345.450 139.130 346.750 139.140 ;
        RECT 347.340 139.130 348.640 139.140 ;
        RECT 109.120 137.640 109.380 138.860 ;
        RECT 111.010 137.640 111.270 138.860 ;
        RECT 217.110 138.580 217.360 138.910 ;
        RECT 219.000 138.580 219.250 138.910 ;
        RECT 89.320 136.780 92.510 137.530 ;
        RECT 217.110 137.360 217.370 138.580 ;
        RECT 219.000 137.360 219.260 138.580 ;
        RECT 244.340 137.770 244.600 138.990 ;
        RECT 246.230 137.770 246.490 138.990 ;
        RECT 345.650 138.800 345.900 139.130 ;
        RECT 347.540 138.800 347.790 139.130 ;
        RECT 453.440 138.860 456.630 139.610 ;
        RECT 453.440 138.850 454.740 138.860 ;
        RECT 455.330 138.850 456.630 138.860 ;
        RECT 345.650 137.580 345.910 138.800 ;
        RECT 347.540 137.580 347.800 138.800 ;
        RECT 453.640 138.520 453.890 138.850 ;
        RECT 455.530 138.520 455.780 138.850 ;
        RECT 89.320 136.770 90.620 136.780 ;
        RECT 91.210 136.770 92.510 136.780 ;
        RECT 89.520 136.440 89.770 136.770 ;
        RECT 91.410 136.440 91.660 136.770 ;
        RECT 190.630 136.590 193.820 137.340 ;
        RECT 325.850 136.720 329.040 137.470 ;
        RECT 453.640 137.300 453.900 138.520 ;
        RECT 455.530 137.300 455.790 138.520 ;
        RECT 325.850 136.710 327.150 136.720 ;
        RECT 327.740 136.710 329.040 136.720 ;
        RECT 190.630 136.580 191.930 136.590 ;
        RECT 192.520 136.580 193.820 136.590 ;
        RECT 89.520 135.220 89.780 136.440 ;
        RECT 91.410 135.220 91.670 136.440 ;
        RECT 190.830 136.250 191.080 136.580 ;
        RECT 192.720 136.250 192.970 136.580 ;
        RECT 326.050 136.380 326.300 136.710 ;
        RECT 327.940 136.380 328.190 136.710 ;
        RECT 427.160 136.530 430.350 137.280 ;
        RECT 427.160 136.520 428.460 136.530 ;
        RECT 429.050 136.520 430.350 136.530 ;
        RECT 190.830 135.030 191.090 136.250 ;
        RECT 192.720 135.030 192.980 136.250 ;
        RECT 326.050 135.160 326.310 136.380 ;
        RECT 327.940 135.160 328.200 136.380 ;
        RECT 427.360 136.190 427.610 136.520 ;
        RECT 429.250 136.190 429.500 136.520 ;
        RECT 470.740 136.510 473.930 137.260 ;
        RECT 470.740 136.500 472.040 136.510 ;
        RECT 472.630 136.500 473.930 136.510 ;
        RECT 427.360 134.970 427.620 136.190 ;
        RECT 429.250 134.970 429.510 136.190 ;
        RECT 470.940 136.170 471.190 136.500 ;
        RECT 472.830 136.170 473.080 136.500 ;
        RECT 470.940 134.950 471.200 136.170 ;
        RECT 472.830 134.950 473.090 136.170 ;
        RECT 7.500 129.960 10.690 130.710 ;
        RECT 7.500 129.950 8.800 129.960 ;
        RECT 9.390 129.950 10.690 129.960 ;
        RECT 7.700 129.620 7.950 129.950 ;
        RECT 9.590 129.620 9.840 129.950 ;
        RECT 108.810 129.770 112.000 130.520 ;
        RECT 244.030 129.900 247.220 130.650 ;
        RECT 244.030 129.890 245.330 129.900 ;
        RECT 245.920 129.890 247.220 129.900 ;
        RECT 108.810 129.760 110.110 129.770 ;
        RECT 110.700 129.760 112.000 129.770 ;
        RECT 7.700 128.400 7.960 129.620 ;
        RECT 9.590 128.400 9.850 129.620 ;
        RECT 109.010 129.430 109.260 129.760 ;
        RECT 110.900 129.430 111.150 129.760 ;
        RECT 244.230 129.560 244.480 129.890 ;
        RECT 246.120 129.560 246.370 129.890 ;
        RECT 345.340 129.710 348.530 130.460 ;
        RECT 345.340 129.700 346.640 129.710 ;
        RECT 347.230 129.700 348.530 129.710 ;
        RECT 23.180 127.540 26.370 128.290 ;
        RECT 109.010 128.210 109.270 129.430 ;
        RECT 110.900 128.210 111.160 129.430 ;
        RECT 244.230 128.340 244.490 129.560 ;
        RECT 246.120 128.340 246.380 129.560 ;
        RECT 345.540 129.370 345.790 129.700 ;
        RECT 347.430 129.370 347.680 129.700 ;
        RECT 23.180 127.530 24.480 127.540 ;
        RECT 25.070 127.530 26.370 127.540 ;
        RECT 23.380 127.200 23.630 127.530 ;
        RECT 25.270 127.200 25.520 127.530 ;
        RECT 124.490 127.350 127.680 128.100 ;
        RECT 259.710 127.480 262.900 128.230 ;
        RECT 345.540 128.150 345.800 129.370 ;
        RECT 347.430 128.150 347.690 129.370 ;
        RECT 259.710 127.470 261.010 127.480 ;
        RECT 261.600 127.470 262.900 127.480 ;
        RECT 124.490 127.340 125.790 127.350 ;
        RECT 126.380 127.340 127.680 127.350 ;
        RECT 23.380 125.980 23.640 127.200 ;
        RECT 25.270 125.980 25.530 127.200 ;
        RECT 124.690 127.010 124.940 127.340 ;
        RECT 126.580 127.010 126.830 127.340 ;
        RECT 259.910 127.140 260.160 127.470 ;
        RECT 261.800 127.140 262.050 127.470 ;
        RECT 361.020 127.290 364.210 128.040 ;
        RECT 361.020 127.280 362.320 127.290 ;
        RECT 362.910 127.280 364.210 127.290 ;
        RECT 124.690 125.790 124.950 127.010 ;
        RECT 126.580 125.790 126.840 127.010 ;
        RECT 259.910 125.920 260.170 127.140 ;
        RECT 261.800 125.920 262.060 127.140 ;
        RECT 361.220 126.950 361.470 127.280 ;
        RECT 363.110 126.950 363.360 127.280 ;
        RECT 361.220 125.730 361.480 126.950 ;
        RECT 363.110 125.730 363.370 126.950 ;
        RECT 7.660 123.560 10.850 124.310 ;
        RECT 7.660 123.550 8.960 123.560 ;
        RECT 9.550 123.550 10.850 123.560 ;
        RECT 7.860 123.220 8.110 123.550 ;
        RECT 9.750 123.220 10.000 123.550 ;
        RECT 108.970 123.370 112.160 124.120 ;
        RECT 244.190 123.500 247.380 124.250 ;
        RECT 244.190 123.490 245.490 123.500 ;
        RECT 246.080 123.490 247.380 123.500 ;
        RECT 108.970 123.360 110.270 123.370 ;
        RECT 110.860 123.360 112.160 123.370 ;
        RECT 7.860 122.000 8.120 123.220 ;
        RECT 9.750 122.000 10.010 123.220 ;
        RECT 109.170 123.030 109.420 123.360 ;
        RECT 111.060 123.030 111.310 123.360 ;
        RECT 244.390 123.160 244.640 123.490 ;
        RECT 246.280 123.160 246.530 123.490 ;
        RECT 345.500 123.310 348.690 124.060 ;
        RECT 345.500 123.300 346.800 123.310 ;
        RECT 347.390 123.300 348.690 123.310 ;
        RECT 40.760 121.990 43.950 122.740 ;
        RECT 40.760 121.980 42.060 121.990 ;
        RECT 42.650 121.980 43.950 121.990 ;
        RECT 40.960 121.650 41.210 121.980 ;
        RECT 42.850 121.650 43.100 121.980 ;
        RECT 109.170 121.810 109.430 123.030 ;
        RECT 111.060 121.810 111.320 123.030 ;
        RECT 142.070 121.800 145.260 122.550 ;
        RECT 244.390 121.940 244.650 123.160 ;
        RECT 246.280 121.940 246.540 123.160 ;
        RECT 345.700 122.970 345.950 123.300 ;
        RECT 347.590 122.970 347.840 123.300 ;
        RECT 277.290 121.930 280.480 122.680 ;
        RECT 277.290 121.920 278.590 121.930 ;
        RECT 279.180 121.920 280.480 121.930 ;
        RECT 142.070 121.790 143.370 121.800 ;
        RECT 143.960 121.790 145.260 121.800 ;
        RECT 40.960 120.430 41.220 121.650 ;
        RECT 42.850 120.430 43.110 121.650 ;
        RECT 142.270 121.460 142.520 121.790 ;
        RECT 144.160 121.460 144.410 121.790 ;
        RECT 277.490 121.590 277.740 121.920 ;
        RECT 279.380 121.590 279.630 121.920 ;
        RECT 345.700 121.750 345.960 122.970 ;
        RECT 347.590 121.750 347.850 122.970 ;
        RECT 378.600 121.740 381.790 122.490 ;
        RECT 378.600 121.730 379.900 121.740 ;
        RECT 380.490 121.730 381.790 121.740 ;
        RECT 142.270 120.240 142.530 121.460 ;
        RECT 144.160 120.240 144.420 121.460 ;
        RECT 277.490 120.370 277.750 121.590 ;
        RECT 279.380 120.370 279.640 121.590 ;
        RECT 378.800 121.400 379.050 121.730 ;
        RECT 380.690 121.400 380.940 121.730 ;
        RECT 378.800 120.180 379.060 121.400 ;
        RECT 380.690 120.180 380.950 121.400 ;
        RECT 7.330 115.540 10.520 116.290 ;
        RECT 7.330 115.530 8.630 115.540 ;
        RECT 9.220 115.530 10.520 115.540 ;
        RECT 7.530 115.200 7.780 115.530 ;
        RECT 9.420 115.200 9.670 115.530 ;
        RECT 108.640 115.350 111.830 116.100 ;
        RECT 243.860 115.480 247.050 116.230 ;
        RECT 243.860 115.470 245.160 115.480 ;
        RECT 245.750 115.470 247.050 115.480 ;
        RECT 108.640 115.340 109.940 115.350 ;
        RECT 110.530 115.340 111.830 115.350 ;
        RECT 7.530 113.980 7.790 115.200 ;
        RECT 9.420 113.980 9.680 115.200 ;
        RECT 108.840 115.010 109.090 115.340 ;
        RECT 110.730 115.010 110.980 115.340 ;
        RECT 244.060 115.140 244.310 115.470 ;
        RECT 245.950 115.140 246.200 115.470 ;
        RECT 345.170 115.290 348.360 116.040 ;
        RECT 345.170 115.280 346.470 115.290 ;
        RECT 347.060 115.280 348.360 115.290 ;
        RECT 23.010 113.120 26.200 113.870 ;
        RECT 108.840 113.790 109.100 115.010 ;
        RECT 110.730 113.790 110.990 115.010 ;
        RECT 244.060 113.920 244.320 115.140 ;
        RECT 245.950 113.920 246.210 115.140 ;
        RECT 345.370 114.950 345.620 115.280 ;
        RECT 347.260 114.950 347.510 115.280 ;
        RECT 23.010 113.110 24.310 113.120 ;
        RECT 24.900 113.110 26.200 113.120 ;
        RECT 23.210 112.780 23.460 113.110 ;
        RECT 25.100 112.780 25.350 113.110 ;
        RECT 124.320 112.930 127.510 113.680 ;
        RECT 259.540 113.060 262.730 113.810 ;
        RECT 345.370 113.730 345.630 114.950 ;
        RECT 347.260 113.730 347.520 114.950 ;
        RECT 259.540 113.050 260.840 113.060 ;
        RECT 261.430 113.050 262.730 113.060 ;
        RECT 124.320 112.920 125.620 112.930 ;
        RECT 126.210 112.920 127.510 112.930 ;
        RECT 23.210 111.560 23.470 112.780 ;
        RECT 25.100 111.560 25.360 112.780 ;
        RECT 124.520 112.590 124.770 112.920 ;
        RECT 126.410 112.590 126.660 112.920 ;
        RECT 259.740 112.720 259.990 113.050 ;
        RECT 261.630 112.720 261.880 113.050 ;
        RECT 360.850 112.870 364.040 113.620 ;
        RECT 360.850 112.860 362.150 112.870 ;
        RECT 362.740 112.860 364.040 112.870 ;
        RECT 124.520 111.370 124.780 112.590 ;
        RECT 126.410 111.370 126.670 112.590 ;
        RECT 259.740 111.500 260.000 112.720 ;
        RECT 261.630 111.500 261.890 112.720 ;
        RECT 361.050 112.530 361.300 112.860 ;
        RECT 362.940 112.530 363.190 112.860 ;
        RECT 361.050 111.310 361.310 112.530 ;
        RECT 362.940 111.310 363.200 112.530 ;
        RECT 7.490 109.140 10.680 109.890 ;
        RECT 7.490 109.130 8.790 109.140 ;
        RECT 9.380 109.130 10.680 109.140 ;
        RECT 7.690 108.800 7.940 109.130 ;
        RECT 9.580 108.800 9.830 109.130 ;
        RECT 108.800 108.950 111.990 109.700 ;
        RECT 244.020 109.080 247.210 109.830 ;
        RECT 244.020 109.070 245.320 109.080 ;
        RECT 245.910 109.070 247.210 109.080 ;
        RECT 108.800 108.940 110.100 108.950 ;
        RECT 110.690 108.940 111.990 108.950 ;
        RECT 7.690 107.580 7.950 108.800 ;
        RECT 9.580 107.580 9.840 108.800 ;
        RECT 109.000 108.610 109.250 108.940 ;
        RECT 110.890 108.610 111.140 108.940 ;
        RECT 244.220 108.740 244.470 109.070 ;
        RECT 246.110 108.740 246.360 109.070 ;
        RECT 345.330 108.890 348.520 109.640 ;
        RECT 345.330 108.880 346.630 108.890 ;
        RECT 347.220 108.880 348.520 108.890 ;
        RECT 109.000 107.390 109.260 108.610 ;
        RECT 110.890 107.390 111.150 108.610 ;
        RECT 244.220 107.520 244.480 108.740 ;
        RECT 246.110 107.520 246.370 108.740 ;
        RECT 345.530 108.550 345.780 108.880 ;
        RECT 347.420 108.550 347.670 108.880 ;
        RECT 345.530 107.330 345.790 108.550 ;
        RECT 347.420 107.330 347.680 108.550 ;
        RECT 58.290 105.970 61.480 106.720 ;
        RECT 58.290 105.960 59.590 105.970 ;
        RECT 60.180 105.960 61.480 105.970 ;
        RECT 58.490 105.630 58.740 105.960 ;
        RECT 60.380 105.630 60.630 105.960 ;
        RECT 159.600 105.780 162.790 106.530 ;
        RECT 294.820 105.910 298.010 106.660 ;
        RECT 294.820 105.900 296.120 105.910 ;
        RECT 296.710 105.900 298.010 105.910 ;
        RECT 159.600 105.770 160.900 105.780 ;
        RECT 161.490 105.770 162.790 105.780 ;
        RECT 58.490 104.410 58.750 105.630 ;
        RECT 60.380 104.410 60.640 105.630 ;
        RECT 159.800 105.440 160.050 105.770 ;
        RECT 161.690 105.440 161.940 105.770 ;
        RECT 295.020 105.570 295.270 105.900 ;
        RECT 296.910 105.570 297.160 105.900 ;
        RECT 396.130 105.720 399.320 106.470 ;
        RECT 396.130 105.710 397.430 105.720 ;
        RECT 398.020 105.710 399.320 105.720 ;
        RECT 159.800 104.220 160.060 105.440 ;
        RECT 161.690 104.220 161.950 105.440 ;
        RECT 295.020 104.350 295.280 105.570 ;
        RECT 296.910 104.350 297.170 105.570 ;
        RECT 396.330 105.380 396.580 105.710 ;
        RECT 398.220 105.380 398.470 105.710 ;
        RECT 396.330 104.160 396.590 105.380 ;
        RECT 398.220 104.160 398.480 105.380 ;
        RECT 7.470 99.890 10.660 100.640 ;
        RECT 7.470 99.880 8.770 99.890 ;
        RECT 9.360 99.880 10.660 99.890 ;
        RECT 7.670 99.550 7.920 99.880 ;
        RECT 9.560 99.550 9.810 99.880 ;
        RECT 108.780 99.700 111.970 100.450 ;
        RECT 244.000 99.830 247.190 100.580 ;
        RECT 244.000 99.820 245.300 99.830 ;
        RECT 245.890 99.820 247.190 99.830 ;
        RECT 108.780 99.690 110.080 99.700 ;
        RECT 110.670 99.690 111.970 99.700 ;
        RECT 7.670 98.330 7.930 99.550 ;
        RECT 9.560 98.330 9.820 99.550 ;
        RECT 108.980 99.360 109.230 99.690 ;
        RECT 110.870 99.360 111.120 99.690 ;
        RECT 244.200 99.490 244.450 99.820 ;
        RECT 246.090 99.490 246.340 99.820 ;
        RECT 345.310 99.640 348.500 100.390 ;
        RECT 345.310 99.630 346.610 99.640 ;
        RECT 347.200 99.630 348.500 99.640 ;
        RECT 23.150 97.470 26.340 98.220 ;
        RECT 108.980 98.140 109.240 99.360 ;
        RECT 110.870 98.140 111.130 99.360 ;
        RECT 244.200 98.270 244.460 99.490 ;
        RECT 246.090 98.270 246.350 99.490 ;
        RECT 345.510 99.300 345.760 99.630 ;
        RECT 347.400 99.300 347.650 99.630 ;
        RECT 23.150 97.460 24.450 97.470 ;
        RECT 25.040 97.460 26.340 97.470 ;
        RECT 23.350 97.130 23.600 97.460 ;
        RECT 25.240 97.130 25.490 97.460 ;
        RECT 124.460 97.280 127.650 98.030 ;
        RECT 259.680 97.410 262.870 98.160 ;
        RECT 345.510 98.080 345.770 99.300 ;
        RECT 347.400 98.080 347.660 99.300 ;
        RECT 259.680 97.400 260.980 97.410 ;
        RECT 261.570 97.400 262.870 97.410 ;
        RECT 124.460 97.270 125.760 97.280 ;
        RECT 126.350 97.270 127.650 97.280 ;
        RECT 23.350 95.910 23.610 97.130 ;
        RECT 25.240 95.910 25.500 97.130 ;
        RECT 124.660 96.940 124.910 97.270 ;
        RECT 126.550 96.940 126.800 97.270 ;
        RECT 259.880 97.070 260.130 97.400 ;
        RECT 261.770 97.070 262.020 97.400 ;
        RECT 360.990 97.220 364.180 97.970 ;
        RECT 360.990 97.210 362.290 97.220 ;
        RECT 362.880 97.210 364.180 97.220 ;
        RECT 124.660 95.720 124.920 96.940 ;
        RECT 126.550 95.720 126.810 96.940 ;
        RECT 259.880 95.850 260.140 97.070 ;
        RECT 261.770 95.850 262.030 97.070 ;
        RECT 361.190 96.880 361.440 97.210 ;
        RECT 363.080 96.880 363.330 97.210 ;
        RECT 361.190 95.660 361.450 96.880 ;
        RECT 363.080 95.660 363.340 96.880 ;
        RECT 7.630 93.490 10.820 94.240 ;
        RECT 7.630 93.480 8.930 93.490 ;
        RECT 9.520 93.480 10.820 93.490 ;
        RECT 7.830 93.150 8.080 93.480 ;
        RECT 9.720 93.150 9.970 93.480 ;
        RECT 108.940 93.300 112.130 94.050 ;
        RECT 244.160 93.430 247.350 94.180 ;
        RECT 244.160 93.420 245.460 93.430 ;
        RECT 246.050 93.420 247.350 93.430 ;
        RECT 108.940 93.290 110.240 93.300 ;
        RECT 110.830 93.290 112.130 93.300 ;
        RECT 7.830 91.930 8.090 93.150 ;
        RECT 9.720 91.930 9.980 93.150 ;
        RECT 109.140 92.960 109.390 93.290 ;
        RECT 111.030 92.960 111.280 93.290 ;
        RECT 244.360 93.090 244.610 93.420 ;
        RECT 246.250 93.090 246.500 93.420 ;
        RECT 345.470 93.240 348.660 93.990 ;
        RECT 345.470 93.230 346.770 93.240 ;
        RECT 347.360 93.230 348.660 93.240 ;
        RECT 40.730 91.920 43.920 92.670 ;
        RECT 40.730 91.910 42.030 91.920 ;
        RECT 42.620 91.910 43.920 91.920 ;
        RECT 40.930 91.580 41.180 91.910 ;
        RECT 42.820 91.580 43.070 91.910 ;
        RECT 109.140 91.740 109.400 92.960 ;
        RECT 111.030 91.740 111.290 92.960 ;
        RECT 142.040 91.730 145.230 92.480 ;
        RECT 244.360 91.870 244.620 93.090 ;
        RECT 246.250 91.870 246.510 93.090 ;
        RECT 345.670 92.900 345.920 93.230 ;
        RECT 347.560 92.900 347.810 93.230 ;
        RECT 277.260 91.860 280.450 92.610 ;
        RECT 277.260 91.850 278.560 91.860 ;
        RECT 279.150 91.850 280.450 91.860 ;
        RECT 142.040 91.720 143.340 91.730 ;
        RECT 143.930 91.720 145.230 91.730 ;
        RECT 40.930 90.360 41.190 91.580 ;
        RECT 42.820 90.360 43.080 91.580 ;
        RECT 142.240 91.390 142.490 91.720 ;
        RECT 144.130 91.390 144.380 91.720 ;
        RECT 277.460 91.520 277.710 91.850 ;
        RECT 279.350 91.520 279.600 91.850 ;
        RECT 345.670 91.680 345.930 92.900 ;
        RECT 347.560 91.680 347.820 92.900 ;
        RECT 378.570 91.670 381.760 92.420 ;
        RECT 378.570 91.660 379.870 91.670 ;
        RECT 380.460 91.660 381.760 91.670 ;
        RECT 142.240 90.170 142.500 91.390 ;
        RECT 144.130 90.170 144.390 91.390 ;
        RECT 277.460 90.300 277.720 91.520 ;
        RECT 279.350 90.300 279.610 91.520 ;
        RECT 378.770 91.330 379.020 91.660 ;
        RECT 380.660 91.330 380.910 91.660 ;
        RECT 378.770 90.110 379.030 91.330 ;
        RECT 380.660 90.110 380.920 91.330 ;
        RECT 7.300 85.470 10.490 86.220 ;
        RECT 7.300 85.460 8.600 85.470 ;
        RECT 9.190 85.460 10.490 85.470 ;
        RECT 7.500 85.130 7.750 85.460 ;
        RECT 9.390 85.130 9.640 85.460 ;
        RECT 108.610 85.280 111.800 86.030 ;
        RECT 243.830 85.410 247.020 86.160 ;
        RECT 243.830 85.400 245.130 85.410 ;
        RECT 245.720 85.400 247.020 85.410 ;
        RECT 108.610 85.270 109.910 85.280 ;
        RECT 110.500 85.270 111.800 85.280 ;
        RECT 7.500 83.910 7.760 85.130 ;
        RECT 9.390 83.910 9.650 85.130 ;
        RECT 108.810 84.940 109.060 85.270 ;
        RECT 110.700 84.940 110.950 85.270 ;
        RECT 244.030 85.070 244.280 85.400 ;
        RECT 245.920 85.070 246.170 85.400 ;
        RECT 345.140 85.220 348.330 85.970 ;
        RECT 345.140 85.210 346.440 85.220 ;
        RECT 347.030 85.210 348.330 85.220 ;
        RECT 22.980 83.050 26.170 83.800 ;
        RECT 108.810 83.720 109.070 84.940 ;
        RECT 110.700 83.720 110.960 84.940 ;
        RECT 244.030 83.850 244.290 85.070 ;
        RECT 245.920 83.850 246.180 85.070 ;
        RECT 345.340 84.880 345.590 85.210 ;
        RECT 347.230 84.880 347.480 85.210 ;
        RECT 22.980 83.040 24.280 83.050 ;
        RECT 24.870 83.040 26.170 83.050 ;
        RECT 23.180 82.710 23.430 83.040 ;
        RECT 25.070 82.710 25.320 83.040 ;
        RECT 124.290 82.860 127.480 83.610 ;
        RECT 259.510 82.990 262.700 83.740 ;
        RECT 345.340 83.660 345.600 84.880 ;
        RECT 347.230 83.660 347.490 84.880 ;
        RECT 259.510 82.980 260.810 82.990 ;
        RECT 261.400 82.980 262.700 82.990 ;
        RECT 124.290 82.850 125.590 82.860 ;
        RECT 126.180 82.850 127.480 82.860 ;
        RECT 23.180 81.490 23.440 82.710 ;
        RECT 25.070 81.490 25.330 82.710 ;
        RECT 124.490 82.520 124.740 82.850 ;
        RECT 126.380 82.520 126.630 82.850 ;
        RECT 259.710 82.650 259.960 82.980 ;
        RECT 261.600 82.650 261.850 82.980 ;
        RECT 360.820 82.800 364.010 83.550 ;
        RECT 360.820 82.790 362.120 82.800 ;
        RECT 362.710 82.790 364.010 82.800 ;
        RECT 124.490 81.300 124.750 82.520 ;
        RECT 126.380 81.300 126.640 82.520 ;
        RECT 259.710 81.430 259.970 82.650 ;
        RECT 261.600 81.430 261.860 82.650 ;
        RECT 361.020 82.460 361.270 82.790 ;
        RECT 362.910 82.460 363.160 82.790 ;
        RECT 361.020 81.240 361.280 82.460 ;
        RECT 362.910 81.240 363.170 82.460 ;
        RECT 7.460 79.070 10.650 79.820 ;
        RECT 72.490 79.680 75.680 80.430 ;
        RECT 72.490 79.670 73.790 79.680 ;
        RECT 74.380 79.670 75.680 79.680 ;
        RECT 7.460 79.060 8.760 79.070 ;
        RECT 9.350 79.060 10.650 79.070 ;
        RECT 72.690 79.340 72.940 79.670 ;
        RECT 74.580 79.340 74.830 79.670 ;
        RECT 7.660 78.730 7.910 79.060 ;
        RECT 9.550 78.730 9.800 79.060 ;
        RECT 7.660 77.510 7.920 78.730 ;
        RECT 9.550 77.510 9.810 78.730 ;
        RECT 72.690 78.120 72.950 79.340 ;
        RECT 74.580 78.120 74.840 79.340 ;
        RECT 108.770 78.880 111.960 79.630 ;
        RECT 173.800 79.490 176.990 80.240 ;
        RECT 173.800 79.480 175.100 79.490 ;
        RECT 175.690 79.480 176.990 79.490 ;
        RECT 108.770 78.870 110.070 78.880 ;
        RECT 110.660 78.870 111.960 78.880 ;
        RECT 174.000 79.150 174.250 79.480 ;
        RECT 175.890 79.150 176.140 79.480 ;
        RECT 108.970 78.540 109.220 78.870 ;
        RECT 110.860 78.540 111.110 78.870 ;
        RECT 108.970 77.320 109.230 78.540 ;
        RECT 110.860 77.320 111.120 78.540 ;
        RECT 174.000 77.930 174.260 79.150 ;
        RECT 175.890 77.930 176.150 79.150 ;
        RECT 243.990 79.010 247.180 79.760 ;
        RECT 309.020 79.620 312.210 80.370 ;
        RECT 309.020 79.610 310.320 79.620 ;
        RECT 310.910 79.610 312.210 79.620 ;
        RECT 243.990 79.000 245.290 79.010 ;
        RECT 245.880 79.000 247.180 79.010 ;
        RECT 309.220 79.280 309.470 79.610 ;
        RECT 311.110 79.280 311.360 79.610 ;
        RECT 244.190 78.670 244.440 79.000 ;
        RECT 246.080 78.670 246.330 79.000 ;
        RECT 244.190 77.450 244.450 78.670 ;
        RECT 246.080 77.450 246.340 78.670 ;
        RECT 309.220 78.060 309.480 79.280 ;
        RECT 311.110 78.060 311.370 79.280 ;
        RECT 345.300 78.820 348.490 79.570 ;
        RECT 410.330 79.430 413.520 80.180 ;
        RECT 410.330 79.420 411.630 79.430 ;
        RECT 412.220 79.420 413.520 79.430 ;
        RECT 345.300 78.810 346.600 78.820 ;
        RECT 347.190 78.810 348.490 78.820 ;
        RECT 410.530 79.090 410.780 79.420 ;
        RECT 412.420 79.090 412.670 79.420 ;
        RECT 345.500 78.480 345.750 78.810 ;
        RECT 347.390 78.480 347.640 78.810 ;
        RECT 345.500 77.260 345.760 78.480 ;
        RECT 347.390 77.260 347.650 78.480 ;
        RECT 410.530 77.870 410.790 79.090 ;
        RECT 412.420 77.870 412.680 79.090 ;
        RECT 7.150 70.040 10.340 70.790 ;
        RECT 7.150 70.030 8.450 70.040 ;
        RECT 9.040 70.030 10.340 70.040 ;
        RECT 7.350 69.700 7.600 70.030 ;
        RECT 9.240 69.700 9.490 70.030 ;
        RECT 108.460 69.850 111.650 70.600 ;
        RECT 243.680 69.980 246.870 70.730 ;
        RECT 243.680 69.970 244.980 69.980 ;
        RECT 245.570 69.970 246.870 69.980 ;
        RECT 108.460 69.840 109.760 69.850 ;
        RECT 110.350 69.840 111.650 69.850 ;
        RECT 7.350 68.480 7.610 69.700 ;
        RECT 9.240 68.480 9.500 69.700 ;
        RECT 108.660 69.510 108.910 69.840 ;
        RECT 110.550 69.510 110.800 69.840 ;
        RECT 243.880 69.640 244.130 69.970 ;
        RECT 245.770 69.640 246.020 69.970 ;
        RECT 344.990 69.790 348.180 70.540 ;
        RECT 344.990 69.780 346.290 69.790 ;
        RECT 346.880 69.780 348.180 69.790 ;
        RECT 22.830 67.620 26.020 68.370 ;
        RECT 108.660 68.290 108.920 69.510 ;
        RECT 110.550 68.290 110.810 69.510 ;
        RECT 243.880 68.420 244.140 69.640 ;
        RECT 245.770 68.420 246.030 69.640 ;
        RECT 345.190 69.450 345.440 69.780 ;
        RECT 347.080 69.450 347.330 69.780 ;
        RECT 22.830 67.610 24.130 67.620 ;
        RECT 24.720 67.610 26.020 67.620 ;
        RECT 23.030 67.280 23.280 67.610 ;
        RECT 24.920 67.280 25.170 67.610 ;
        RECT 124.140 67.430 127.330 68.180 ;
        RECT 259.360 67.560 262.550 68.310 ;
        RECT 345.190 68.230 345.450 69.450 ;
        RECT 347.080 68.230 347.340 69.450 ;
        RECT 259.360 67.550 260.660 67.560 ;
        RECT 261.250 67.550 262.550 67.560 ;
        RECT 124.140 67.420 125.440 67.430 ;
        RECT 126.030 67.420 127.330 67.430 ;
        RECT 23.030 66.060 23.290 67.280 ;
        RECT 24.920 66.060 25.180 67.280 ;
        RECT 124.340 67.090 124.590 67.420 ;
        RECT 126.230 67.090 126.480 67.420 ;
        RECT 259.560 67.220 259.810 67.550 ;
        RECT 261.450 67.220 261.700 67.550 ;
        RECT 360.670 67.370 363.860 68.120 ;
        RECT 360.670 67.360 361.970 67.370 ;
        RECT 362.560 67.360 363.860 67.370 ;
        RECT 124.340 65.870 124.600 67.090 ;
        RECT 126.230 65.870 126.490 67.090 ;
        RECT 259.560 66.000 259.820 67.220 ;
        RECT 261.450 66.000 261.710 67.220 ;
        RECT 360.870 67.030 361.120 67.360 ;
        RECT 362.760 67.030 363.010 67.360 ;
        RECT 360.870 65.810 361.130 67.030 ;
        RECT 362.760 65.810 363.020 67.030 ;
        RECT 7.310 63.640 10.500 64.390 ;
        RECT 7.310 63.630 8.610 63.640 ;
        RECT 9.200 63.630 10.500 63.640 ;
        RECT 7.510 63.300 7.760 63.630 ;
        RECT 9.400 63.300 9.650 63.630 ;
        RECT 108.620 63.450 111.810 64.200 ;
        RECT 243.840 63.580 247.030 64.330 ;
        RECT 243.840 63.570 245.140 63.580 ;
        RECT 245.730 63.570 247.030 63.580 ;
        RECT 108.620 63.440 109.920 63.450 ;
        RECT 110.510 63.440 111.810 63.450 ;
        RECT 7.510 62.080 7.770 63.300 ;
        RECT 9.400 62.080 9.660 63.300 ;
        RECT 108.820 63.110 109.070 63.440 ;
        RECT 110.710 63.110 110.960 63.440 ;
        RECT 244.040 63.240 244.290 63.570 ;
        RECT 245.930 63.240 246.180 63.570 ;
        RECT 345.150 63.390 348.340 64.140 ;
        RECT 345.150 63.380 346.450 63.390 ;
        RECT 347.040 63.380 348.340 63.390 ;
        RECT 40.410 62.070 43.600 62.820 ;
        RECT 40.410 62.060 41.710 62.070 ;
        RECT 42.300 62.060 43.600 62.070 ;
        RECT 40.610 61.730 40.860 62.060 ;
        RECT 42.500 61.730 42.750 62.060 ;
        RECT 108.820 61.890 109.080 63.110 ;
        RECT 110.710 61.890 110.970 63.110 ;
        RECT 141.720 61.880 144.910 62.630 ;
        RECT 244.040 62.020 244.300 63.240 ;
        RECT 245.930 62.020 246.190 63.240 ;
        RECT 345.350 63.050 345.600 63.380 ;
        RECT 347.240 63.050 347.490 63.380 ;
        RECT 276.940 62.010 280.130 62.760 ;
        RECT 276.940 62.000 278.240 62.010 ;
        RECT 278.830 62.000 280.130 62.010 ;
        RECT 141.720 61.870 143.020 61.880 ;
        RECT 143.610 61.870 144.910 61.880 ;
        RECT 40.610 60.510 40.870 61.730 ;
        RECT 42.500 60.510 42.760 61.730 ;
        RECT 141.920 61.540 142.170 61.870 ;
        RECT 143.810 61.540 144.060 61.870 ;
        RECT 277.140 61.670 277.390 62.000 ;
        RECT 279.030 61.670 279.280 62.000 ;
        RECT 345.350 61.830 345.610 63.050 ;
        RECT 347.240 61.830 347.500 63.050 ;
        RECT 378.250 61.820 381.440 62.570 ;
        RECT 378.250 61.810 379.550 61.820 ;
        RECT 380.140 61.810 381.440 61.820 ;
        RECT 141.920 60.320 142.180 61.540 ;
        RECT 143.810 60.320 144.070 61.540 ;
        RECT 277.140 60.450 277.400 61.670 ;
        RECT 279.030 60.450 279.290 61.670 ;
        RECT 378.450 61.480 378.700 61.810 ;
        RECT 380.340 61.480 380.590 61.810 ;
        RECT 378.450 60.260 378.710 61.480 ;
        RECT 380.340 60.260 380.600 61.480 ;
        RECT 6.980 55.620 10.170 56.370 ;
        RECT 6.980 55.610 8.280 55.620 ;
        RECT 8.870 55.610 10.170 55.620 ;
        RECT 7.180 55.280 7.430 55.610 ;
        RECT 9.070 55.280 9.320 55.610 ;
        RECT 108.290 55.430 111.480 56.180 ;
        RECT 243.510 55.560 246.700 56.310 ;
        RECT 243.510 55.550 244.810 55.560 ;
        RECT 245.400 55.550 246.700 55.560 ;
        RECT 108.290 55.420 109.590 55.430 ;
        RECT 110.180 55.420 111.480 55.430 ;
        RECT 7.180 54.060 7.440 55.280 ;
        RECT 9.070 54.060 9.330 55.280 ;
        RECT 108.490 55.090 108.740 55.420 ;
        RECT 110.380 55.090 110.630 55.420 ;
        RECT 243.710 55.220 243.960 55.550 ;
        RECT 245.600 55.220 245.850 55.550 ;
        RECT 344.820 55.370 348.010 56.120 ;
        RECT 344.820 55.360 346.120 55.370 ;
        RECT 346.710 55.360 348.010 55.370 ;
        RECT 22.660 53.200 25.850 53.950 ;
        RECT 108.490 53.870 108.750 55.090 ;
        RECT 110.380 53.870 110.640 55.090 ;
        RECT 243.710 54.000 243.970 55.220 ;
        RECT 245.600 54.000 245.860 55.220 ;
        RECT 345.020 55.030 345.270 55.360 ;
        RECT 346.910 55.030 347.160 55.360 ;
        RECT 22.660 53.190 23.960 53.200 ;
        RECT 24.550 53.190 25.850 53.200 ;
        RECT 22.860 52.860 23.110 53.190 ;
        RECT 24.750 52.860 25.000 53.190 ;
        RECT 123.970 53.010 127.160 53.760 ;
        RECT 259.190 53.140 262.380 53.890 ;
        RECT 345.020 53.810 345.280 55.030 ;
        RECT 346.910 53.810 347.170 55.030 ;
        RECT 259.190 53.130 260.490 53.140 ;
        RECT 261.080 53.130 262.380 53.140 ;
        RECT 123.970 53.000 125.270 53.010 ;
        RECT 125.860 53.000 127.160 53.010 ;
        RECT 22.860 51.640 23.120 52.860 ;
        RECT 24.750 51.640 25.010 52.860 ;
        RECT 124.170 52.670 124.420 53.000 ;
        RECT 126.060 52.670 126.310 53.000 ;
        RECT 259.390 52.800 259.640 53.130 ;
        RECT 261.280 52.800 261.530 53.130 ;
        RECT 360.500 52.950 363.690 53.700 ;
        RECT 360.500 52.940 361.800 52.950 ;
        RECT 362.390 52.940 363.690 52.950 ;
        RECT 124.170 51.450 124.430 52.670 ;
        RECT 126.060 51.450 126.320 52.670 ;
        RECT 259.390 51.580 259.650 52.800 ;
        RECT 261.280 51.580 261.540 52.800 ;
        RECT 360.700 52.610 360.950 52.940 ;
        RECT 362.590 52.610 362.840 52.940 ;
        RECT 360.700 51.390 360.960 52.610 ;
        RECT 362.590 51.390 362.850 52.610 ;
        RECT 7.140 49.220 10.330 49.970 ;
        RECT 7.140 49.210 8.440 49.220 ;
        RECT 9.030 49.210 10.330 49.220 ;
        RECT 7.340 48.880 7.590 49.210 ;
        RECT 9.230 48.880 9.480 49.210 ;
        RECT 108.450 49.030 111.640 49.780 ;
        RECT 243.670 49.160 246.860 49.910 ;
        RECT 243.670 49.150 244.970 49.160 ;
        RECT 245.560 49.150 246.860 49.160 ;
        RECT 108.450 49.020 109.750 49.030 ;
        RECT 110.340 49.020 111.640 49.030 ;
        RECT 7.340 47.660 7.600 48.880 ;
        RECT 9.230 47.660 9.490 48.880 ;
        RECT 108.650 48.690 108.900 49.020 ;
        RECT 110.540 48.690 110.790 49.020 ;
        RECT 243.870 48.820 244.120 49.150 ;
        RECT 245.760 48.820 246.010 49.150 ;
        RECT 344.980 48.970 348.170 49.720 ;
        RECT 344.980 48.960 346.280 48.970 ;
        RECT 346.870 48.960 348.170 48.970 ;
        RECT 108.650 47.470 108.910 48.690 ;
        RECT 110.540 47.470 110.800 48.690 ;
        RECT 243.870 47.600 244.130 48.820 ;
        RECT 245.760 47.600 246.020 48.820 ;
        RECT 345.180 48.630 345.430 48.960 ;
        RECT 347.070 48.630 347.320 48.960 ;
        RECT 345.180 47.410 345.440 48.630 ;
        RECT 347.070 47.410 347.330 48.630 ;
        RECT 57.940 46.050 61.130 46.800 ;
        RECT 57.940 46.040 59.240 46.050 ;
        RECT 59.830 46.040 61.130 46.050 ;
        RECT 58.140 45.710 58.390 46.040 ;
        RECT 60.030 45.710 60.280 46.040 ;
        RECT 159.250 45.860 162.440 46.610 ;
        RECT 294.470 45.990 297.660 46.740 ;
        RECT 294.470 45.980 295.770 45.990 ;
        RECT 296.360 45.980 297.660 45.990 ;
        RECT 159.250 45.850 160.550 45.860 ;
        RECT 161.140 45.850 162.440 45.860 ;
        RECT 58.140 44.490 58.400 45.710 ;
        RECT 60.030 44.490 60.290 45.710 ;
        RECT 159.450 45.520 159.700 45.850 ;
        RECT 161.340 45.520 161.590 45.850 ;
        RECT 294.670 45.650 294.920 45.980 ;
        RECT 296.560 45.650 296.810 45.980 ;
        RECT 395.780 45.800 398.970 46.550 ;
        RECT 395.780 45.790 397.080 45.800 ;
        RECT 397.670 45.790 398.970 45.800 ;
        RECT 159.450 44.300 159.710 45.520 ;
        RECT 161.340 44.300 161.600 45.520 ;
        RECT 294.670 44.430 294.930 45.650 ;
        RECT 296.560 44.430 296.820 45.650 ;
        RECT 395.980 45.460 396.230 45.790 ;
        RECT 397.870 45.460 398.120 45.790 ;
        RECT 395.980 44.240 396.240 45.460 ;
        RECT 397.870 44.240 398.130 45.460 ;
        RECT 7.120 39.970 10.310 40.720 ;
        RECT 7.120 39.960 8.420 39.970 ;
        RECT 9.010 39.960 10.310 39.970 ;
        RECT 7.320 39.630 7.570 39.960 ;
        RECT 9.210 39.630 9.460 39.960 ;
        RECT 108.430 39.780 111.620 40.530 ;
        RECT 243.650 39.910 246.840 40.660 ;
        RECT 243.650 39.900 244.950 39.910 ;
        RECT 245.540 39.900 246.840 39.910 ;
        RECT 108.430 39.770 109.730 39.780 ;
        RECT 110.320 39.770 111.620 39.780 ;
        RECT 7.320 38.410 7.580 39.630 ;
        RECT 9.210 38.410 9.470 39.630 ;
        RECT 108.630 39.440 108.880 39.770 ;
        RECT 110.520 39.440 110.770 39.770 ;
        RECT 243.850 39.570 244.100 39.900 ;
        RECT 245.740 39.570 245.990 39.900 ;
        RECT 344.960 39.720 348.150 40.470 ;
        RECT 344.960 39.710 346.260 39.720 ;
        RECT 346.850 39.710 348.150 39.720 ;
        RECT 22.800 37.550 25.990 38.300 ;
        RECT 108.630 38.220 108.890 39.440 ;
        RECT 110.520 38.220 110.780 39.440 ;
        RECT 243.850 38.350 244.110 39.570 ;
        RECT 245.740 38.350 246.000 39.570 ;
        RECT 345.160 39.380 345.410 39.710 ;
        RECT 347.050 39.380 347.300 39.710 ;
        RECT 22.800 37.540 24.100 37.550 ;
        RECT 24.690 37.540 25.990 37.550 ;
        RECT 23.000 37.210 23.250 37.540 ;
        RECT 24.890 37.210 25.140 37.540 ;
        RECT 124.110 37.360 127.300 38.110 ;
        RECT 259.330 37.490 262.520 38.240 ;
        RECT 345.160 38.160 345.420 39.380 ;
        RECT 347.050 38.160 347.310 39.380 ;
        RECT 259.330 37.480 260.630 37.490 ;
        RECT 261.220 37.480 262.520 37.490 ;
        RECT 124.110 37.350 125.410 37.360 ;
        RECT 126.000 37.350 127.300 37.360 ;
        RECT 23.000 35.990 23.260 37.210 ;
        RECT 24.890 35.990 25.150 37.210 ;
        RECT 124.310 37.020 124.560 37.350 ;
        RECT 126.200 37.020 126.450 37.350 ;
        RECT 259.530 37.150 259.780 37.480 ;
        RECT 261.420 37.150 261.670 37.480 ;
        RECT 360.640 37.300 363.830 38.050 ;
        RECT 360.640 37.290 361.940 37.300 ;
        RECT 362.530 37.290 363.830 37.300 ;
        RECT 124.310 35.800 124.570 37.020 ;
        RECT 126.200 35.800 126.460 37.020 ;
        RECT 259.530 35.930 259.790 37.150 ;
        RECT 261.420 35.930 261.680 37.150 ;
        RECT 360.840 36.960 361.090 37.290 ;
        RECT 362.730 36.960 362.980 37.290 ;
        RECT 360.840 35.740 361.100 36.960 ;
        RECT 362.730 35.740 362.990 36.960 ;
        RECT 7.280 33.570 10.470 34.320 ;
        RECT 7.280 33.560 8.580 33.570 ;
        RECT 9.170 33.560 10.470 33.570 ;
        RECT 7.480 33.230 7.730 33.560 ;
        RECT 9.370 33.230 9.620 33.560 ;
        RECT 108.590 33.380 111.780 34.130 ;
        RECT 243.810 33.510 247.000 34.260 ;
        RECT 243.810 33.500 245.110 33.510 ;
        RECT 245.700 33.500 247.000 33.510 ;
        RECT 108.590 33.370 109.890 33.380 ;
        RECT 110.480 33.370 111.780 33.380 ;
        RECT 7.480 32.010 7.740 33.230 ;
        RECT 9.370 32.010 9.630 33.230 ;
        RECT 108.790 33.040 109.040 33.370 ;
        RECT 110.680 33.040 110.930 33.370 ;
        RECT 244.010 33.170 244.260 33.500 ;
        RECT 245.900 33.170 246.150 33.500 ;
        RECT 345.120 33.320 348.310 34.070 ;
        RECT 345.120 33.310 346.420 33.320 ;
        RECT 347.010 33.310 348.310 33.320 ;
        RECT 40.380 32.000 43.570 32.750 ;
        RECT 40.380 31.990 41.680 32.000 ;
        RECT 42.270 31.990 43.570 32.000 ;
        RECT 40.580 31.660 40.830 31.990 ;
        RECT 42.470 31.660 42.720 31.990 ;
        RECT 108.790 31.820 109.050 33.040 ;
        RECT 110.680 31.820 110.940 33.040 ;
        RECT 141.690 31.810 144.880 32.560 ;
        RECT 244.010 31.950 244.270 33.170 ;
        RECT 245.900 31.950 246.160 33.170 ;
        RECT 345.320 32.980 345.570 33.310 ;
        RECT 347.210 32.980 347.460 33.310 ;
        RECT 276.910 31.940 280.100 32.690 ;
        RECT 276.910 31.930 278.210 31.940 ;
        RECT 278.800 31.930 280.100 31.940 ;
        RECT 141.690 31.800 142.990 31.810 ;
        RECT 143.580 31.800 144.880 31.810 ;
        RECT 40.580 30.440 40.840 31.660 ;
        RECT 42.470 30.440 42.730 31.660 ;
        RECT 141.890 31.470 142.140 31.800 ;
        RECT 143.780 31.470 144.030 31.800 ;
        RECT 277.110 31.600 277.360 31.930 ;
        RECT 279.000 31.600 279.250 31.930 ;
        RECT 345.320 31.760 345.580 32.980 ;
        RECT 347.210 31.760 347.470 32.980 ;
        RECT 378.220 31.750 381.410 32.500 ;
        RECT 378.220 31.740 379.520 31.750 ;
        RECT 380.110 31.740 381.410 31.750 ;
        RECT 141.890 30.250 142.150 31.470 ;
        RECT 143.780 30.250 144.040 31.470 ;
        RECT 277.110 30.380 277.370 31.600 ;
        RECT 279.000 30.380 279.260 31.600 ;
        RECT 378.420 31.410 378.670 31.740 ;
        RECT 380.310 31.410 380.560 31.740 ;
        RECT 378.420 30.190 378.680 31.410 ;
        RECT 380.310 30.190 380.570 31.410 ;
        RECT 6.950 25.550 10.140 26.300 ;
        RECT 6.950 25.540 8.250 25.550 ;
        RECT 8.840 25.540 10.140 25.550 ;
        RECT 7.150 25.210 7.400 25.540 ;
        RECT 9.040 25.210 9.290 25.540 ;
        RECT 108.260 25.360 111.450 26.110 ;
        RECT 243.480 25.490 246.670 26.240 ;
        RECT 243.480 25.480 244.780 25.490 ;
        RECT 245.370 25.480 246.670 25.490 ;
        RECT 108.260 25.350 109.560 25.360 ;
        RECT 110.150 25.350 111.450 25.360 ;
        RECT 7.150 23.990 7.410 25.210 ;
        RECT 9.040 23.990 9.300 25.210 ;
        RECT 108.460 25.020 108.710 25.350 ;
        RECT 110.350 25.020 110.600 25.350 ;
        RECT 243.680 25.150 243.930 25.480 ;
        RECT 245.570 25.150 245.820 25.480 ;
        RECT 344.790 25.300 347.980 26.050 ;
        RECT 344.790 25.290 346.090 25.300 ;
        RECT 346.680 25.290 347.980 25.300 ;
        RECT 22.630 23.130 25.820 23.880 ;
        RECT 108.460 23.800 108.720 25.020 ;
        RECT 110.350 23.800 110.610 25.020 ;
        RECT 243.680 23.930 243.940 25.150 ;
        RECT 245.570 23.930 245.830 25.150 ;
        RECT 344.990 24.960 345.240 25.290 ;
        RECT 346.880 24.960 347.130 25.290 ;
        RECT 22.630 23.120 23.930 23.130 ;
        RECT 24.520 23.120 25.820 23.130 ;
        RECT 22.830 22.790 23.080 23.120 ;
        RECT 24.720 22.790 24.970 23.120 ;
        RECT 123.940 22.940 127.130 23.690 ;
        RECT 259.160 23.070 262.350 23.820 ;
        RECT 344.990 23.740 345.250 24.960 ;
        RECT 346.880 23.740 347.140 24.960 ;
        RECT 259.160 23.060 260.460 23.070 ;
        RECT 261.050 23.060 262.350 23.070 ;
        RECT 123.940 22.930 125.240 22.940 ;
        RECT 125.830 22.930 127.130 22.940 ;
        RECT 22.830 21.570 23.090 22.790 ;
        RECT 24.720 21.570 24.980 22.790 ;
        RECT 124.140 22.600 124.390 22.930 ;
        RECT 126.030 22.600 126.280 22.930 ;
        RECT 259.360 22.730 259.610 23.060 ;
        RECT 261.250 22.730 261.500 23.060 ;
        RECT 360.470 22.880 363.660 23.630 ;
        RECT 360.470 22.870 361.770 22.880 ;
        RECT 362.360 22.870 363.660 22.880 ;
        RECT 124.140 21.380 124.400 22.600 ;
        RECT 126.030 21.380 126.290 22.600 ;
        RECT 259.360 21.510 259.620 22.730 ;
        RECT 261.250 21.510 261.510 22.730 ;
        RECT 360.670 22.540 360.920 22.870 ;
        RECT 362.560 22.540 362.810 22.870 ;
        RECT 360.670 21.320 360.930 22.540 ;
        RECT 362.560 21.320 362.820 22.540 ;
        RECT 7.110 19.150 10.300 19.900 ;
        RECT 7.110 19.140 8.410 19.150 ;
        RECT 9.000 19.140 10.300 19.150 ;
        RECT 7.310 18.810 7.560 19.140 ;
        RECT 9.200 18.810 9.450 19.140 ;
        RECT 108.420 18.960 111.610 19.710 ;
        RECT 243.640 19.090 246.830 19.840 ;
        RECT 243.640 19.080 244.940 19.090 ;
        RECT 245.530 19.080 246.830 19.090 ;
        RECT 108.420 18.950 109.720 18.960 ;
        RECT 110.310 18.950 111.610 18.960 ;
        RECT 7.310 17.590 7.570 18.810 ;
        RECT 9.200 17.590 9.460 18.810 ;
        RECT 108.620 18.620 108.870 18.950 ;
        RECT 110.510 18.620 110.760 18.950 ;
        RECT 243.840 18.750 244.090 19.080 ;
        RECT 245.730 18.750 245.980 19.080 ;
        RECT 344.950 18.900 348.140 19.650 ;
        RECT 344.950 18.890 346.250 18.900 ;
        RECT 346.840 18.890 348.140 18.900 ;
        RECT 108.620 17.400 108.880 18.620 ;
        RECT 110.510 17.400 110.770 18.620 ;
        RECT 243.840 17.530 244.100 18.750 ;
        RECT 245.730 17.530 245.990 18.750 ;
        RECT 345.150 18.560 345.400 18.890 ;
        RECT 347.040 18.560 347.290 18.890 ;
        RECT 345.150 17.340 345.410 18.560 ;
        RECT 347.040 17.340 347.300 18.560 ;
      LAYER mcon ;
        RECT 8.155 250.305 8.325 250.475 ;
        RECT 9.015 250.305 9.185 250.475 ;
        RECT 10.045 250.305 10.215 250.475 ;
        RECT 10.905 250.305 11.075 250.475 ;
        RECT 109.465 250.115 109.635 250.285 ;
        RECT 110.325 250.115 110.495 250.285 ;
        RECT 111.355 250.115 111.525 250.285 ;
        RECT 112.215 250.115 112.385 250.285 ;
        RECT 244.685 250.245 244.855 250.415 ;
        RECT 245.545 250.245 245.715 250.415 ;
        RECT 246.575 250.245 246.745 250.415 ;
        RECT 247.435 250.245 247.605 250.415 ;
        RECT 345.995 250.055 346.165 250.225 ;
        RECT 346.855 250.055 347.025 250.225 ;
        RECT 347.885 250.055 348.055 250.225 ;
        RECT 348.745 250.055 348.915 250.225 ;
        RECT 23.835 247.885 24.005 248.055 ;
        RECT 24.695 247.885 24.865 248.055 ;
        RECT 25.725 247.885 25.895 248.055 ;
        RECT 26.585 247.885 26.755 248.055 ;
        RECT 125.145 247.695 125.315 247.865 ;
        RECT 126.005 247.695 126.175 247.865 ;
        RECT 127.035 247.695 127.205 247.865 ;
        RECT 127.895 247.695 128.065 247.865 ;
        RECT 260.365 247.825 260.535 247.995 ;
        RECT 261.225 247.825 261.395 247.995 ;
        RECT 262.255 247.825 262.425 247.995 ;
        RECT 263.115 247.825 263.285 247.995 ;
        RECT 361.675 247.635 361.845 247.805 ;
        RECT 362.535 247.635 362.705 247.805 ;
        RECT 363.565 247.635 363.735 247.805 ;
        RECT 364.425 247.635 364.595 247.805 ;
        RECT 8.315 243.905 8.485 244.075 ;
        RECT 9.175 243.905 9.345 244.075 ;
        RECT 10.205 243.905 10.375 244.075 ;
        RECT 11.065 243.905 11.235 244.075 ;
        RECT 109.625 243.715 109.795 243.885 ;
        RECT 110.485 243.715 110.655 243.885 ;
        RECT 111.515 243.715 111.685 243.885 ;
        RECT 112.375 243.715 112.545 243.885 ;
        RECT 244.845 243.845 245.015 244.015 ;
        RECT 245.705 243.845 245.875 244.015 ;
        RECT 246.735 243.845 246.905 244.015 ;
        RECT 247.595 243.845 247.765 244.015 ;
        RECT 346.155 243.655 346.325 243.825 ;
        RECT 347.015 243.655 347.185 243.825 ;
        RECT 348.045 243.655 348.215 243.825 ;
        RECT 348.905 243.655 349.075 243.825 ;
        RECT 41.415 242.335 41.585 242.505 ;
        RECT 42.275 242.335 42.445 242.505 ;
        RECT 43.305 242.335 43.475 242.505 ;
        RECT 44.165 242.335 44.335 242.505 ;
        RECT 142.725 242.145 142.895 242.315 ;
        RECT 143.585 242.145 143.755 242.315 ;
        RECT 144.615 242.145 144.785 242.315 ;
        RECT 145.475 242.145 145.645 242.315 ;
        RECT 277.945 242.275 278.115 242.445 ;
        RECT 278.805 242.275 278.975 242.445 ;
        RECT 279.835 242.275 280.005 242.445 ;
        RECT 280.695 242.275 280.865 242.445 ;
        RECT 379.255 242.085 379.425 242.255 ;
        RECT 380.115 242.085 380.285 242.255 ;
        RECT 381.145 242.085 381.315 242.255 ;
        RECT 382.005 242.085 382.175 242.255 ;
        RECT 7.985 235.885 8.155 236.055 ;
        RECT 8.845 235.885 9.015 236.055 ;
        RECT 9.875 235.885 10.045 236.055 ;
        RECT 10.735 235.885 10.905 236.055 ;
        RECT 109.295 235.695 109.465 235.865 ;
        RECT 110.155 235.695 110.325 235.865 ;
        RECT 111.185 235.695 111.355 235.865 ;
        RECT 112.045 235.695 112.215 235.865 ;
        RECT 244.515 235.825 244.685 235.995 ;
        RECT 245.375 235.825 245.545 235.995 ;
        RECT 246.405 235.825 246.575 235.995 ;
        RECT 247.265 235.825 247.435 235.995 ;
        RECT 345.825 235.635 345.995 235.805 ;
        RECT 346.685 235.635 346.855 235.805 ;
        RECT 347.715 235.635 347.885 235.805 ;
        RECT 348.575 235.635 348.745 235.805 ;
        RECT 23.665 233.465 23.835 233.635 ;
        RECT 24.525 233.465 24.695 233.635 ;
        RECT 25.555 233.465 25.725 233.635 ;
        RECT 26.415 233.465 26.585 233.635 ;
        RECT 124.975 233.275 125.145 233.445 ;
        RECT 125.835 233.275 126.005 233.445 ;
        RECT 126.865 233.275 127.035 233.445 ;
        RECT 127.725 233.275 127.895 233.445 ;
        RECT 260.195 233.405 260.365 233.575 ;
        RECT 261.055 233.405 261.225 233.575 ;
        RECT 262.085 233.405 262.255 233.575 ;
        RECT 262.945 233.405 263.115 233.575 ;
        RECT 361.505 233.215 361.675 233.385 ;
        RECT 362.365 233.215 362.535 233.385 ;
        RECT 363.395 233.215 363.565 233.385 ;
        RECT 364.255 233.215 364.425 233.385 ;
        RECT 8.145 229.485 8.315 229.655 ;
        RECT 9.005 229.485 9.175 229.655 ;
        RECT 10.035 229.485 10.205 229.655 ;
        RECT 10.895 229.485 11.065 229.655 ;
        RECT 109.455 229.295 109.625 229.465 ;
        RECT 110.315 229.295 110.485 229.465 ;
        RECT 111.345 229.295 111.515 229.465 ;
        RECT 112.205 229.295 112.375 229.465 ;
        RECT 244.675 229.425 244.845 229.595 ;
        RECT 245.535 229.425 245.705 229.595 ;
        RECT 246.565 229.425 246.735 229.595 ;
        RECT 247.425 229.425 247.595 229.595 ;
        RECT 345.985 229.235 346.155 229.405 ;
        RECT 346.845 229.235 347.015 229.405 ;
        RECT 347.875 229.235 348.045 229.405 ;
        RECT 348.735 229.235 348.905 229.405 ;
        RECT 58.945 226.315 59.115 226.485 ;
        RECT 59.805 226.315 59.975 226.485 ;
        RECT 60.835 226.315 61.005 226.485 ;
        RECT 61.695 226.315 61.865 226.485 ;
        RECT 160.255 226.125 160.425 226.295 ;
        RECT 161.115 226.125 161.285 226.295 ;
        RECT 162.145 226.125 162.315 226.295 ;
        RECT 163.005 226.125 163.175 226.295 ;
        RECT 295.475 226.255 295.645 226.425 ;
        RECT 296.335 226.255 296.505 226.425 ;
        RECT 297.365 226.255 297.535 226.425 ;
        RECT 298.225 226.255 298.395 226.425 ;
        RECT 396.785 226.065 396.955 226.235 ;
        RECT 397.645 226.065 397.815 226.235 ;
        RECT 398.675 226.065 398.845 226.235 ;
        RECT 399.535 226.065 399.705 226.235 ;
        RECT 8.125 220.235 8.295 220.405 ;
        RECT 8.985 220.235 9.155 220.405 ;
        RECT 10.015 220.235 10.185 220.405 ;
        RECT 10.875 220.235 11.045 220.405 ;
        RECT 109.435 220.045 109.605 220.215 ;
        RECT 110.295 220.045 110.465 220.215 ;
        RECT 111.325 220.045 111.495 220.215 ;
        RECT 112.185 220.045 112.355 220.215 ;
        RECT 244.655 220.175 244.825 220.345 ;
        RECT 245.515 220.175 245.685 220.345 ;
        RECT 246.545 220.175 246.715 220.345 ;
        RECT 247.405 220.175 247.575 220.345 ;
        RECT 345.965 219.985 346.135 220.155 ;
        RECT 346.825 219.985 346.995 220.155 ;
        RECT 347.855 219.985 348.025 220.155 ;
        RECT 348.715 219.985 348.885 220.155 ;
        RECT 23.805 217.815 23.975 217.985 ;
        RECT 24.665 217.815 24.835 217.985 ;
        RECT 25.695 217.815 25.865 217.985 ;
        RECT 26.555 217.815 26.725 217.985 ;
        RECT 125.115 217.625 125.285 217.795 ;
        RECT 125.975 217.625 126.145 217.795 ;
        RECT 127.005 217.625 127.175 217.795 ;
        RECT 127.865 217.625 128.035 217.795 ;
        RECT 260.335 217.755 260.505 217.925 ;
        RECT 261.195 217.755 261.365 217.925 ;
        RECT 262.225 217.755 262.395 217.925 ;
        RECT 263.085 217.755 263.255 217.925 ;
        RECT 361.645 217.565 361.815 217.735 ;
        RECT 362.505 217.565 362.675 217.735 ;
        RECT 363.535 217.565 363.705 217.735 ;
        RECT 364.395 217.565 364.565 217.735 ;
        RECT 8.285 213.835 8.455 214.005 ;
        RECT 9.145 213.835 9.315 214.005 ;
        RECT 10.175 213.835 10.345 214.005 ;
        RECT 11.035 213.835 11.205 214.005 ;
        RECT 109.595 213.645 109.765 213.815 ;
        RECT 110.455 213.645 110.625 213.815 ;
        RECT 111.485 213.645 111.655 213.815 ;
        RECT 112.345 213.645 112.515 213.815 ;
        RECT 244.815 213.775 244.985 213.945 ;
        RECT 245.675 213.775 245.845 213.945 ;
        RECT 246.705 213.775 246.875 213.945 ;
        RECT 247.565 213.775 247.735 213.945 ;
        RECT 346.125 213.585 346.295 213.755 ;
        RECT 346.985 213.585 347.155 213.755 ;
        RECT 348.015 213.585 348.185 213.755 ;
        RECT 348.875 213.585 349.045 213.755 ;
        RECT 41.385 212.265 41.555 212.435 ;
        RECT 42.245 212.265 42.415 212.435 ;
        RECT 43.275 212.265 43.445 212.435 ;
        RECT 44.135 212.265 44.305 212.435 ;
        RECT 142.695 212.075 142.865 212.245 ;
        RECT 143.555 212.075 143.725 212.245 ;
        RECT 144.585 212.075 144.755 212.245 ;
        RECT 145.445 212.075 145.615 212.245 ;
        RECT 277.915 212.205 278.085 212.375 ;
        RECT 278.775 212.205 278.945 212.375 ;
        RECT 279.805 212.205 279.975 212.375 ;
        RECT 280.665 212.205 280.835 212.375 ;
        RECT 379.225 212.015 379.395 212.185 ;
        RECT 380.085 212.015 380.255 212.185 ;
        RECT 381.115 212.015 381.285 212.185 ;
        RECT 381.975 212.015 382.145 212.185 ;
        RECT 7.955 205.815 8.125 205.985 ;
        RECT 8.815 205.815 8.985 205.985 ;
        RECT 9.845 205.815 10.015 205.985 ;
        RECT 10.705 205.815 10.875 205.985 ;
        RECT 109.265 205.625 109.435 205.795 ;
        RECT 110.125 205.625 110.295 205.795 ;
        RECT 111.155 205.625 111.325 205.795 ;
        RECT 112.015 205.625 112.185 205.795 ;
        RECT 244.485 205.755 244.655 205.925 ;
        RECT 245.345 205.755 245.515 205.925 ;
        RECT 246.375 205.755 246.545 205.925 ;
        RECT 247.235 205.755 247.405 205.925 ;
        RECT 345.795 205.565 345.965 205.735 ;
        RECT 346.655 205.565 346.825 205.735 ;
        RECT 347.685 205.565 347.855 205.735 ;
        RECT 348.545 205.565 348.715 205.735 ;
        RECT 23.635 203.395 23.805 203.565 ;
        RECT 24.495 203.395 24.665 203.565 ;
        RECT 25.525 203.395 25.695 203.565 ;
        RECT 26.385 203.395 26.555 203.565 ;
        RECT 124.945 203.205 125.115 203.375 ;
        RECT 125.805 203.205 125.975 203.375 ;
        RECT 126.835 203.205 127.005 203.375 ;
        RECT 127.695 203.205 127.865 203.375 ;
        RECT 260.165 203.335 260.335 203.505 ;
        RECT 261.025 203.335 261.195 203.505 ;
        RECT 262.055 203.335 262.225 203.505 ;
        RECT 262.915 203.335 263.085 203.505 ;
        RECT 361.475 203.145 361.645 203.315 ;
        RECT 362.335 203.145 362.505 203.315 ;
        RECT 363.365 203.145 363.535 203.315 ;
        RECT 364.225 203.145 364.395 203.315 ;
        RECT 73.145 200.025 73.315 200.195 ;
        RECT 74.005 200.025 74.175 200.195 ;
        RECT 75.035 200.025 75.205 200.195 ;
        RECT 75.895 200.025 76.065 200.195 ;
        RECT 8.115 199.415 8.285 199.585 ;
        RECT 8.975 199.415 9.145 199.585 ;
        RECT 10.005 199.415 10.175 199.585 ;
        RECT 10.865 199.415 11.035 199.585 ;
        RECT 174.455 199.835 174.625 200.005 ;
        RECT 175.315 199.835 175.485 200.005 ;
        RECT 176.345 199.835 176.515 200.005 ;
        RECT 177.205 199.835 177.375 200.005 ;
        RECT 109.425 199.225 109.595 199.395 ;
        RECT 110.285 199.225 110.455 199.395 ;
        RECT 111.315 199.225 111.485 199.395 ;
        RECT 112.175 199.225 112.345 199.395 ;
        RECT 309.675 199.965 309.845 200.135 ;
        RECT 310.535 199.965 310.705 200.135 ;
        RECT 311.565 199.965 311.735 200.135 ;
        RECT 312.425 199.965 312.595 200.135 ;
        RECT 244.645 199.355 244.815 199.525 ;
        RECT 245.505 199.355 245.675 199.525 ;
        RECT 246.535 199.355 246.705 199.525 ;
        RECT 247.395 199.355 247.565 199.525 ;
        RECT 410.985 199.775 411.155 199.945 ;
        RECT 411.845 199.775 412.015 199.945 ;
        RECT 412.875 199.775 413.045 199.945 ;
        RECT 413.735 199.775 413.905 199.945 ;
        RECT 345.955 199.165 346.125 199.335 ;
        RECT 346.815 199.165 346.985 199.335 ;
        RECT 347.845 199.165 348.015 199.335 ;
        RECT 348.705 199.165 348.875 199.335 ;
        RECT 7.805 190.385 7.975 190.555 ;
        RECT 8.665 190.385 8.835 190.555 ;
        RECT 9.695 190.385 9.865 190.555 ;
        RECT 10.555 190.385 10.725 190.555 ;
        RECT 109.115 190.195 109.285 190.365 ;
        RECT 109.975 190.195 110.145 190.365 ;
        RECT 111.005 190.195 111.175 190.365 ;
        RECT 111.865 190.195 112.035 190.365 ;
        RECT 244.335 190.325 244.505 190.495 ;
        RECT 245.195 190.325 245.365 190.495 ;
        RECT 246.225 190.325 246.395 190.495 ;
        RECT 247.085 190.325 247.255 190.495 ;
        RECT 345.645 190.135 345.815 190.305 ;
        RECT 346.505 190.135 346.675 190.305 ;
        RECT 347.535 190.135 347.705 190.305 ;
        RECT 348.395 190.135 348.565 190.305 ;
        RECT 23.485 187.965 23.655 188.135 ;
        RECT 24.345 187.965 24.515 188.135 ;
        RECT 25.375 187.965 25.545 188.135 ;
        RECT 26.235 187.965 26.405 188.135 ;
        RECT 124.795 187.775 124.965 187.945 ;
        RECT 125.655 187.775 125.825 187.945 ;
        RECT 126.685 187.775 126.855 187.945 ;
        RECT 127.545 187.775 127.715 187.945 ;
        RECT 260.015 187.905 260.185 188.075 ;
        RECT 260.875 187.905 261.045 188.075 ;
        RECT 261.905 187.905 262.075 188.075 ;
        RECT 262.765 187.905 262.935 188.075 ;
        RECT 361.325 187.715 361.495 187.885 ;
        RECT 362.185 187.715 362.355 187.885 ;
        RECT 363.215 187.715 363.385 187.885 ;
        RECT 364.075 187.715 364.245 187.885 ;
        RECT 7.965 183.985 8.135 184.155 ;
        RECT 8.825 183.985 8.995 184.155 ;
        RECT 9.855 183.985 10.025 184.155 ;
        RECT 10.715 183.985 10.885 184.155 ;
        RECT 109.275 183.795 109.445 183.965 ;
        RECT 110.135 183.795 110.305 183.965 ;
        RECT 111.165 183.795 111.335 183.965 ;
        RECT 112.025 183.795 112.195 183.965 ;
        RECT 244.495 183.925 244.665 184.095 ;
        RECT 245.355 183.925 245.525 184.095 ;
        RECT 246.385 183.925 246.555 184.095 ;
        RECT 247.245 183.925 247.415 184.095 ;
        RECT 345.805 183.735 345.975 183.905 ;
        RECT 346.665 183.735 346.835 183.905 ;
        RECT 347.695 183.735 347.865 183.905 ;
        RECT 348.555 183.735 348.725 183.905 ;
        RECT 41.065 182.415 41.235 182.585 ;
        RECT 41.925 182.415 42.095 182.585 ;
        RECT 42.955 182.415 43.125 182.585 ;
        RECT 43.815 182.415 43.985 182.585 ;
        RECT 142.375 182.225 142.545 182.395 ;
        RECT 143.235 182.225 143.405 182.395 ;
        RECT 144.265 182.225 144.435 182.395 ;
        RECT 145.125 182.225 145.295 182.395 ;
        RECT 277.595 182.355 277.765 182.525 ;
        RECT 278.455 182.355 278.625 182.525 ;
        RECT 279.485 182.355 279.655 182.525 ;
        RECT 280.345 182.355 280.515 182.525 ;
        RECT 378.905 182.165 379.075 182.335 ;
        RECT 379.765 182.165 379.935 182.335 ;
        RECT 380.795 182.165 380.965 182.335 ;
        RECT 381.655 182.165 381.825 182.335 ;
        RECT 7.635 175.965 7.805 176.135 ;
        RECT 8.495 175.965 8.665 176.135 ;
        RECT 9.525 175.965 9.695 176.135 ;
        RECT 10.385 175.965 10.555 176.135 ;
        RECT 108.945 175.775 109.115 175.945 ;
        RECT 109.805 175.775 109.975 175.945 ;
        RECT 110.835 175.775 111.005 175.945 ;
        RECT 111.695 175.775 111.865 175.945 ;
        RECT 244.165 175.905 244.335 176.075 ;
        RECT 245.025 175.905 245.195 176.075 ;
        RECT 246.055 175.905 246.225 176.075 ;
        RECT 246.915 175.905 247.085 176.075 ;
        RECT 345.475 175.715 345.645 175.885 ;
        RECT 346.335 175.715 346.505 175.885 ;
        RECT 347.365 175.715 347.535 175.885 ;
        RECT 348.225 175.715 348.395 175.885 ;
        RECT 23.315 173.545 23.485 173.715 ;
        RECT 24.175 173.545 24.345 173.715 ;
        RECT 25.205 173.545 25.375 173.715 ;
        RECT 26.065 173.545 26.235 173.715 ;
        RECT 124.625 173.355 124.795 173.525 ;
        RECT 125.485 173.355 125.655 173.525 ;
        RECT 126.515 173.355 126.685 173.525 ;
        RECT 127.375 173.355 127.545 173.525 ;
        RECT 259.845 173.485 260.015 173.655 ;
        RECT 260.705 173.485 260.875 173.655 ;
        RECT 261.735 173.485 261.905 173.655 ;
        RECT 262.595 173.485 262.765 173.655 ;
        RECT 361.155 173.295 361.325 173.465 ;
        RECT 362.015 173.295 362.185 173.465 ;
        RECT 363.045 173.295 363.215 173.465 ;
        RECT 363.905 173.295 364.075 173.465 ;
        RECT 7.795 169.565 7.965 169.735 ;
        RECT 8.655 169.565 8.825 169.735 ;
        RECT 9.685 169.565 9.855 169.735 ;
        RECT 10.545 169.565 10.715 169.735 ;
        RECT 109.105 169.375 109.275 169.545 ;
        RECT 109.965 169.375 110.135 169.545 ;
        RECT 110.995 169.375 111.165 169.545 ;
        RECT 111.855 169.375 112.025 169.545 ;
        RECT 244.325 169.505 244.495 169.675 ;
        RECT 245.185 169.505 245.355 169.675 ;
        RECT 246.215 169.505 246.385 169.675 ;
        RECT 247.075 169.505 247.245 169.675 ;
        RECT 345.635 169.315 345.805 169.485 ;
        RECT 346.495 169.315 346.665 169.485 ;
        RECT 347.525 169.315 347.695 169.485 ;
        RECT 348.385 169.315 348.555 169.485 ;
        RECT 58.595 166.395 58.765 166.565 ;
        RECT 59.455 166.395 59.625 166.565 ;
        RECT 60.485 166.395 60.655 166.565 ;
        RECT 61.345 166.395 61.515 166.565 ;
        RECT 159.905 166.205 160.075 166.375 ;
        RECT 160.765 166.205 160.935 166.375 ;
        RECT 161.795 166.205 161.965 166.375 ;
        RECT 162.655 166.205 162.825 166.375 ;
        RECT 295.125 166.335 295.295 166.505 ;
        RECT 295.985 166.335 296.155 166.505 ;
        RECT 297.015 166.335 297.185 166.505 ;
        RECT 297.875 166.335 298.045 166.505 ;
        RECT 396.435 166.145 396.605 166.315 ;
        RECT 397.295 166.145 397.465 166.315 ;
        RECT 398.325 166.145 398.495 166.315 ;
        RECT 399.185 166.145 399.355 166.315 ;
        RECT 7.775 160.315 7.945 160.485 ;
        RECT 8.635 160.315 8.805 160.485 ;
        RECT 9.665 160.315 9.835 160.485 ;
        RECT 10.525 160.315 10.695 160.485 ;
        RECT 109.085 160.125 109.255 160.295 ;
        RECT 109.945 160.125 110.115 160.295 ;
        RECT 110.975 160.125 111.145 160.295 ;
        RECT 111.835 160.125 112.005 160.295 ;
        RECT 244.305 160.255 244.475 160.425 ;
        RECT 245.165 160.255 245.335 160.425 ;
        RECT 246.195 160.255 246.365 160.425 ;
        RECT 247.055 160.255 247.225 160.425 ;
        RECT 345.615 160.065 345.785 160.235 ;
        RECT 346.475 160.065 346.645 160.235 ;
        RECT 347.505 160.065 347.675 160.235 ;
        RECT 348.365 160.065 348.535 160.235 ;
        RECT 23.455 157.895 23.625 158.065 ;
        RECT 24.315 157.895 24.485 158.065 ;
        RECT 25.345 157.895 25.515 158.065 ;
        RECT 26.205 157.895 26.375 158.065 ;
        RECT 124.765 157.705 124.935 157.875 ;
        RECT 125.625 157.705 125.795 157.875 ;
        RECT 126.655 157.705 126.825 157.875 ;
        RECT 127.515 157.705 127.685 157.875 ;
        RECT 259.985 157.835 260.155 158.005 ;
        RECT 260.845 157.835 261.015 158.005 ;
        RECT 261.875 157.835 262.045 158.005 ;
        RECT 262.735 157.835 262.905 158.005 ;
        RECT 361.295 157.645 361.465 157.815 ;
        RECT 362.155 157.645 362.325 157.815 ;
        RECT 363.185 157.645 363.355 157.815 ;
        RECT 364.045 157.645 364.215 157.815 ;
        RECT 7.935 153.915 8.105 154.085 ;
        RECT 8.795 153.915 8.965 154.085 ;
        RECT 9.825 153.915 9.995 154.085 ;
        RECT 10.685 153.915 10.855 154.085 ;
        RECT 109.245 153.725 109.415 153.895 ;
        RECT 110.105 153.725 110.275 153.895 ;
        RECT 111.135 153.725 111.305 153.895 ;
        RECT 111.995 153.725 112.165 153.895 ;
        RECT 244.465 153.855 244.635 154.025 ;
        RECT 245.325 153.855 245.495 154.025 ;
        RECT 246.355 153.855 246.525 154.025 ;
        RECT 247.215 153.855 247.385 154.025 ;
        RECT 345.775 153.665 345.945 153.835 ;
        RECT 346.635 153.665 346.805 153.835 ;
        RECT 347.665 153.665 347.835 153.835 ;
        RECT 348.525 153.665 348.695 153.835 ;
        RECT 41.035 152.345 41.205 152.515 ;
        RECT 41.895 152.345 42.065 152.515 ;
        RECT 42.925 152.345 43.095 152.515 ;
        RECT 43.785 152.345 43.955 152.515 ;
        RECT 142.345 152.155 142.515 152.325 ;
        RECT 143.205 152.155 143.375 152.325 ;
        RECT 144.235 152.155 144.405 152.325 ;
        RECT 145.095 152.155 145.265 152.325 ;
        RECT 277.565 152.285 277.735 152.455 ;
        RECT 278.425 152.285 278.595 152.455 ;
        RECT 279.455 152.285 279.625 152.455 ;
        RECT 280.315 152.285 280.485 152.455 ;
        RECT 378.875 152.095 379.045 152.265 ;
        RECT 379.735 152.095 379.905 152.265 ;
        RECT 380.765 152.095 380.935 152.265 ;
        RECT 381.625 152.095 381.795 152.265 ;
        RECT 7.605 145.895 7.775 146.065 ;
        RECT 8.465 145.895 8.635 146.065 ;
        RECT 9.495 145.895 9.665 146.065 ;
        RECT 10.355 145.895 10.525 146.065 ;
        RECT 108.915 145.705 109.085 145.875 ;
        RECT 109.775 145.705 109.945 145.875 ;
        RECT 110.805 145.705 110.975 145.875 ;
        RECT 111.665 145.705 111.835 145.875 ;
        RECT 244.135 145.835 244.305 146.005 ;
        RECT 244.995 145.835 245.165 146.005 ;
        RECT 246.025 145.835 246.195 146.005 ;
        RECT 246.885 145.835 247.055 146.005 ;
        RECT 345.445 145.645 345.615 145.815 ;
        RECT 346.305 145.645 346.475 145.815 ;
        RECT 347.335 145.645 347.505 145.815 ;
        RECT 348.195 145.645 348.365 145.815 ;
        RECT 23.285 143.475 23.455 143.645 ;
        RECT 24.145 143.475 24.315 143.645 ;
        RECT 25.175 143.475 25.345 143.645 ;
        RECT 26.035 143.475 26.205 143.645 ;
        RECT 124.595 143.285 124.765 143.455 ;
        RECT 125.455 143.285 125.625 143.455 ;
        RECT 126.485 143.285 126.655 143.455 ;
        RECT 127.345 143.285 127.515 143.455 ;
        RECT 259.815 143.415 259.985 143.585 ;
        RECT 260.675 143.415 260.845 143.585 ;
        RECT 261.705 143.415 261.875 143.585 ;
        RECT 262.565 143.415 262.735 143.585 ;
        RECT 361.125 143.225 361.295 143.395 ;
        RECT 361.985 143.225 362.155 143.395 ;
        RECT 363.015 143.225 363.185 143.395 ;
        RECT 363.875 143.225 364.045 143.395 ;
        RECT 7.765 139.495 7.935 139.665 ;
        RECT 8.625 139.495 8.795 139.665 ;
        RECT 9.655 139.495 9.825 139.665 ;
        RECT 10.515 139.495 10.685 139.665 ;
        RECT 109.075 139.305 109.245 139.475 ;
        RECT 109.935 139.305 110.105 139.475 ;
        RECT 110.965 139.305 111.135 139.475 ;
        RECT 111.825 139.305 111.995 139.475 ;
        RECT 244.295 139.435 244.465 139.605 ;
        RECT 245.155 139.435 245.325 139.605 ;
        RECT 246.185 139.435 246.355 139.605 ;
        RECT 247.045 139.435 247.215 139.605 ;
        RECT 217.065 139.025 217.235 139.195 ;
        RECT 217.925 139.025 218.095 139.195 ;
        RECT 218.955 139.025 219.125 139.195 ;
        RECT 219.815 139.025 219.985 139.195 ;
        RECT 345.605 139.245 345.775 139.415 ;
        RECT 346.465 139.245 346.635 139.415 ;
        RECT 347.495 139.245 347.665 139.415 ;
        RECT 348.355 139.245 348.525 139.415 ;
        RECT 453.595 138.965 453.765 139.135 ;
        RECT 454.455 138.965 454.625 139.135 ;
        RECT 455.485 138.965 455.655 139.135 ;
        RECT 456.345 138.965 456.515 139.135 ;
        RECT 89.475 136.885 89.645 137.055 ;
        RECT 90.335 136.885 90.505 137.055 ;
        RECT 91.365 136.885 91.535 137.055 ;
        RECT 92.225 136.885 92.395 137.055 ;
        RECT 190.785 136.695 190.955 136.865 ;
        RECT 191.645 136.695 191.815 136.865 ;
        RECT 192.675 136.695 192.845 136.865 ;
        RECT 193.535 136.695 193.705 136.865 ;
        RECT 326.005 136.825 326.175 136.995 ;
        RECT 326.865 136.825 327.035 136.995 ;
        RECT 327.895 136.825 328.065 136.995 ;
        RECT 328.755 136.825 328.925 136.995 ;
        RECT 427.315 136.635 427.485 136.805 ;
        RECT 428.175 136.635 428.345 136.805 ;
        RECT 429.205 136.635 429.375 136.805 ;
        RECT 430.065 136.635 430.235 136.805 ;
        RECT 470.895 136.615 471.065 136.785 ;
        RECT 471.755 136.615 471.925 136.785 ;
        RECT 472.785 136.615 472.955 136.785 ;
        RECT 473.645 136.615 473.815 136.785 ;
        RECT 7.655 130.065 7.825 130.235 ;
        RECT 8.515 130.065 8.685 130.235 ;
        RECT 9.545 130.065 9.715 130.235 ;
        RECT 10.405 130.065 10.575 130.235 ;
        RECT 108.965 129.875 109.135 130.045 ;
        RECT 109.825 129.875 109.995 130.045 ;
        RECT 110.855 129.875 111.025 130.045 ;
        RECT 111.715 129.875 111.885 130.045 ;
        RECT 244.185 130.005 244.355 130.175 ;
        RECT 245.045 130.005 245.215 130.175 ;
        RECT 246.075 130.005 246.245 130.175 ;
        RECT 246.935 130.005 247.105 130.175 ;
        RECT 345.495 129.815 345.665 129.985 ;
        RECT 346.355 129.815 346.525 129.985 ;
        RECT 347.385 129.815 347.555 129.985 ;
        RECT 348.245 129.815 348.415 129.985 ;
        RECT 23.335 127.645 23.505 127.815 ;
        RECT 24.195 127.645 24.365 127.815 ;
        RECT 25.225 127.645 25.395 127.815 ;
        RECT 26.085 127.645 26.255 127.815 ;
        RECT 124.645 127.455 124.815 127.625 ;
        RECT 125.505 127.455 125.675 127.625 ;
        RECT 126.535 127.455 126.705 127.625 ;
        RECT 127.395 127.455 127.565 127.625 ;
        RECT 259.865 127.585 260.035 127.755 ;
        RECT 260.725 127.585 260.895 127.755 ;
        RECT 261.755 127.585 261.925 127.755 ;
        RECT 262.615 127.585 262.785 127.755 ;
        RECT 361.175 127.395 361.345 127.565 ;
        RECT 362.035 127.395 362.205 127.565 ;
        RECT 363.065 127.395 363.235 127.565 ;
        RECT 363.925 127.395 364.095 127.565 ;
        RECT 7.815 123.665 7.985 123.835 ;
        RECT 8.675 123.665 8.845 123.835 ;
        RECT 9.705 123.665 9.875 123.835 ;
        RECT 10.565 123.665 10.735 123.835 ;
        RECT 109.125 123.475 109.295 123.645 ;
        RECT 109.985 123.475 110.155 123.645 ;
        RECT 111.015 123.475 111.185 123.645 ;
        RECT 111.875 123.475 112.045 123.645 ;
        RECT 244.345 123.605 244.515 123.775 ;
        RECT 245.205 123.605 245.375 123.775 ;
        RECT 246.235 123.605 246.405 123.775 ;
        RECT 247.095 123.605 247.265 123.775 ;
        RECT 345.655 123.415 345.825 123.585 ;
        RECT 346.515 123.415 346.685 123.585 ;
        RECT 347.545 123.415 347.715 123.585 ;
        RECT 348.405 123.415 348.575 123.585 ;
        RECT 40.915 122.095 41.085 122.265 ;
        RECT 41.775 122.095 41.945 122.265 ;
        RECT 42.805 122.095 42.975 122.265 ;
        RECT 43.665 122.095 43.835 122.265 ;
        RECT 142.225 121.905 142.395 122.075 ;
        RECT 143.085 121.905 143.255 122.075 ;
        RECT 144.115 121.905 144.285 122.075 ;
        RECT 144.975 121.905 145.145 122.075 ;
        RECT 277.445 122.035 277.615 122.205 ;
        RECT 278.305 122.035 278.475 122.205 ;
        RECT 279.335 122.035 279.505 122.205 ;
        RECT 280.195 122.035 280.365 122.205 ;
        RECT 378.755 121.845 378.925 122.015 ;
        RECT 379.615 121.845 379.785 122.015 ;
        RECT 380.645 121.845 380.815 122.015 ;
        RECT 381.505 121.845 381.675 122.015 ;
        RECT 7.485 115.645 7.655 115.815 ;
        RECT 8.345 115.645 8.515 115.815 ;
        RECT 9.375 115.645 9.545 115.815 ;
        RECT 10.235 115.645 10.405 115.815 ;
        RECT 108.795 115.455 108.965 115.625 ;
        RECT 109.655 115.455 109.825 115.625 ;
        RECT 110.685 115.455 110.855 115.625 ;
        RECT 111.545 115.455 111.715 115.625 ;
        RECT 244.015 115.585 244.185 115.755 ;
        RECT 244.875 115.585 245.045 115.755 ;
        RECT 245.905 115.585 246.075 115.755 ;
        RECT 246.765 115.585 246.935 115.755 ;
        RECT 345.325 115.395 345.495 115.565 ;
        RECT 346.185 115.395 346.355 115.565 ;
        RECT 347.215 115.395 347.385 115.565 ;
        RECT 348.075 115.395 348.245 115.565 ;
        RECT 23.165 113.225 23.335 113.395 ;
        RECT 24.025 113.225 24.195 113.395 ;
        RECT 25.055 113.225 25.225 113.395 ;
        RECT 25.915 113.225 26.085 113.395 ;
        RECT 124.475 113.035 124.645 113.205 ;
        RECT 125.335 113.035 125.505 113.205 ;
        RECT 126.365 113.035 126.535 113.205 ;
        RECT 127.225 113.035 127.395 113.205 ;
        RECT 259.695 113.165 259.865 113.335 ;
        RECT 260.555 113.165 260.725 113.335 ;
        RECT 261.585 113.165 261.755 113.335 ;
        RECT 262.445 113.165 262.615 113.335 ;
        RECT 361.005 112.975 361.175 113.145 ;
        RECT 361.865 112.975 362.035 113.145 ;
        RECT 362.895 112.975 363.065 113.145 ;
        RECT 363.755 112.975 363.925 113.145 ;
        RECT 7.645 109.245 7.815 109.415 ;
        RECT 8.505 109.245 8.675 109.415 ;
        RECT 9.535 109.245 9.705 109.415 ;
        RECT 10.395 109.245 10.565 109.415 ;
        RECT 108.955 109.055 109.125 109.225 ;
        RECT 109.815 109.055 109.985 109.225 ;
        RECT 110.845 109.055 111.015 109.225 ;
        RECT 111.705 109.055 111.875 109.225 ;
        RECT 244.175 109.185 244.345 109.355 ;
        RECT 245.035 109.185 245.205 109.355 ;
        RECT 246.065 109.185 246.235 109.355 ;
        RECT 246.925 109.185 247.095 109.355 ;
        RECT 345.485 108.995 345.655 109.165 ;
        RECT 346.345 108.995 346.515 109.165 ;
        RECT 347.375 108.995 347.545 109.165 ;
        RECT 348.235 108.995 348.405 109.165 ;
        RECT 58.445 106.075 58.615 106.245 ;
        RECT 59.305 106.075 59.475 106.245 ;
        RECT 60.335 106.075 60.505 106.245 ;
        RECT 61.195 106.075 61.365 106.245 ;
        RECT 159.755 105.885 159.925 106.055 ;
        RECT 160.615 105.885 160.785 106.055 ;
        RECT 161.645 105.885 161.815 106.055 ;
        RECT 162.505 105.885 162.675 106.055 ;
        RECT 294.975 106.015 295.145 106.185 ;
        RECT 295.835 106.015 296.005 106.185 ;
        RECT 296.865 106.015 297.035 106.185 ;
        RECT 297.725 106.015 297.895 106.185 ;
        RECT 396.285 105.825 396.455 105.995 ;
        RECT 397.145 105.825 397.315 105.995 ;
        RECT 398.175 105.825 398.345 105.995 ;
        RECT 399.035 105.825 399.205 105.995 ;
        RECT 7.625 99.995 7.795 100.165 ;
        RECT 8.485 99.995 8.655 100.165 ;
        RECT 9.515 99.995 9.685 100.165 ;
        RECT 10.375 99.995 10.545 100.165 ;
        RECT 108.935 99.805 109.105 99.975 ;
        RECT 109.795 99.805 109.965 99.975 ;
        RECT 110.825 99.805 110.995 99.975 ;
        RECT 111.685 99.805 111.855 99.975 ;
        RECT 244.155 99.935 244.325 100.105 ;
        RECT 245.015 99.935 245.185 100.105 ;
        RECT 246.045 99.935 246.215 100.105 ;
        RECT 246.905 99.935 247.075 100.105 ;
        RECT 345.465 99.745 345.635 99.915 ;
        RECT 346.325 99.745 346.495 99.915 ;
        RECT 347.355 99.745 347.525 99.915 ;
        RECT 348.215 99.745 348.385 99.915 ;
        RECT 23.305 97.575 23.475 97.745 ;
        RECT 24.165 97.575 24.335 97.745 ;
        RECT 25.195 97.575 25.365 97.745 ;
        RECT 26.055 97.575 26.225 97.745 ;
        RECT 124.615 97.385 124.785 97.555 ;
        RECT 125.475 97.385 125.645 97.555 ;
        RECT 126.505 97.385 126.675 97.555 ;
        RECT 127.365 97.385 127.535 97.555 ;
        RECT 259.835 97.515 260.005 97.685 ;
        RECT 260.695 97.515 260.865 97.685 ;
        RECT 261.725 97.515 261.895 97.685 ;
        RECT 262.585 97.515 262.755 97.685 ;
        RECT 361.145 97.325 361.315 97.495 ;
        RECT 362.005 97.325 362.175 97.495 ;
        RECT 363.035 97.325 363.205 97.495 ;
        RECT 363.895 97.325 364.065 97.495 ;
        RECT 7.785 93.595 7.955 93.765 ;
        RECT 8.645 93.595 8.815 93.765 ;
        RECT 9.675 93.595 9.845 93.765 ;
        RECT 10.535 93.595 10.705 93.765 ;
        RECT 109.095 93.405 109.265 93.575 ;
        RECT 109.955 93.405 110.125 93.575 ;
        RECT 110.985 93.405 111.155 93.575 ;
        RECT 111.845 93.405 112.015 93.575 ;
        RECT 244.315 93.535 244.485 93.705 ;
        RECT 245.175 93.535 245.345 93.705 ;
        RECT 246.205 93.535 246.375 93.705 ;
        RECT 247.065 93.535 247.235 93.705 ;
        RECT 345.625 93.345 345.795 93.515 ;
        RECT 346.485 93.345 346.655 93.515 ;
        RECT 347.515 93.345 347.685 93.515 ;
        RECT 348.375 93.345 348.545 93.515 ;
        RECT 40.885 92.025 41.055 92.195 ;
        RECT 41.745 92.025 41.915 92.195 ;
        RECT 42.775 92.025 42.945 92.195 ;
        RECT 43.635 92.025 43.805 92.195 ;
        RECT 142.195 91.835 142.365 92.005 ;
        RECT 143.055 91.835 143.225 92.005 ;
        RECT 144.085 91.835 144.255 92.005 ;
        RECT 144.945 91.835 145.115 92.005 ;
        RECT 277.415 91.965 277.585 92.135 ;
        RECT 278.275 91.965 278.445 92.135 ;
        RECT 279.305 91.965 279.475 92.135 ;
        RECT 280.165 91.965 280.335 92.135 ;
        RECT 378.725 91.775 378.895 91.945 ;
        RECT 379.585 91.775 379.755 91.945 ;
        RECT 380.615 91.775 380.785 91.945 ;
        RECT 381.475 91.775 381.645 91.945 ;
        RECT 7.455 85.575 7.625 85.745 ;
        RECT 8.315 85.575 8.485 85.745 ;
        RECT 9.345 85.575 9.515 85.745 ;
        RECT 10.205 85.575 10.375 85.745 ;
        RECT 108.765 85.385 108.935 85.555 ;
        RECT 109.625 85.385 109.795 85.555 ;
        RECT 110.655 85.385 110.825 85.555 ;
        RECT 111.515 85.385 111.685 85.555 ;
        RECT 243.985 85.515 244.155 85.685 ;
        RECT 244.845 85.515 245.015 85.685 ;
        RECT 245.875 85.515 246.045 85.685 ;
        RECT 246.735 85.515 246.905 85.685 ;
        RECT 345.295 85.325 345.465 85.495 ;
        RECT 346.155 85.325 346.325 85.495 ;
        RECT 347.185 85.325 347.355 85.495 ;
        RECT 348.045 85.325 348.215 85.495 ;
        RECT 23.135 83.155 23.305 83.325 ;
        RECT 23.995 83.155 24.165 83.325 ;
        RECT 25.025 83.155 25.195 83.325 ;
        RECT 25.885 83.155 26.055 83.325 ;
        RECT 124.445 82.965 124.615 83.135 ;
        RECT 125.305 82.965 125.475 83.135 ;
        RECT 126.335 82.965 126.505 83.135 ;
        RECT 127.195 82.965 127.365 83.135 ;
        RECT 259.665 83.095 259.835 83.265 ;
        RECT 260.525 83.095 260.695 83.265 ;
        RECT 261.555 83.095 261.725 83.265 ;
        RECT 262.415 83.095 262.585 83.265 ;
        RECT 360.975 82.905 361.145 83.075 ;
        RECT 361.835 82.905 362.005 83.075 ;
        RECT 362.865 82.905 363.035 83.075 ;
        RECT 363.725 82.905 363.895 83.075 ;
        RECT 72.645 79.785 72.815 79.955 ;
        RECT 73.505 79.785 73.675 79.955 ;
        RECT 74.535 79.785 74.705 79.955 ;
        RECT 75.395 79.785 75.565 79.955 ;
        RECT 7.615 79.175 7.785 79.345 ;
        RECT 8.475 79.175 8.645 79.345 ;
        RECT 9.505 79.175 9.675 79.345 ;
        RECT 10.365 79.175 10.535 79.345 ;
        RECT 173.955 79.595 174.125 79.765 ;
        RECT 174.815 79.595 174.985 79.765 ;
        RECT 175.845 79.595 176.015 79.765 ;
        RECT 176.705 79.595 176.875 79.765 ;
        RECT 108.925 78.985 109.095 79.155 ;
        RECT 109.785 78.985 109.955 79.155 ;
        RECT 110.815 78.985 110.985 79.155 ;
        RECT 111.675 78.985 111.845 79.155 ;
        RECT 309.175 79.725 309.345 79.895 ;
        RECT 310.035 79.725 310.205 79.895 ;
        RECT 311.065 79.725 311.235 79.895 ;
        RECT 311.925 79.725 312.095 79.895 ;
        RECT 244.145 79.115 244.315 79.285 ;
        RECT 245.005 79.115 245.175 79.285 ;
        RECT 246.035 79.115 246.205 79.285 ;
        RECT 246.895 79.115 247.065 79.285 ;
        RECT 410.485 79.535 410.655 79.705 ;
        RECT 411.345 79.535 411.515 79.705 ;
        RECT 412.375 79.535 412.545 79.705 ;
        RECT 413.235 79.535 413.405 79.705 ;
        RECT 345.455 78.925 345.625 79.095 ;
        RECT 346.315 78.925 346.485 79.095 ;
        RECT 347.345 78.925 347.515 79.095 ;
        RECT 348.205 78.925 348.375 79.095 ;
        RECT 7.305 70.145 7.475 70.315 ;
        RECT 8.165 70.145 8.335 70.315 ;
        RECT 9.195 70.145 9.365 70.315 ;
        RECT 10.055 70.145 10.225 70.315 ;
        RECT 108.615 69.955 108.785 70.125 ;
        RECT 109.475 69.955 109.645 70.125 ;
        RECT 110.505 69.955 110.675 70.125 ;
        RECT 111.365 69.955 111.535 70.125 ;
        RECT 243.835 70.085 244.005 70.255 ;
        RECT 244.695 70.085 244.865 70.255 ;
        RECT 245.725 70.085 245.895 70.255 ;
        RECT 246.585 70.085 246.755 70.255 ;
        RECT 345.145 69.895 345.315 70.065 ;
        RECT 346.005 69.895 346.175 70.065 ;
        RECT 347.035 69.895 347.205 70.065 ;
        RECT 347.895 69.895 348.065 70.065 ;
        RECT 22.985 67.725 23.155 67.895 ;
        RECT 23.845 67.725 24.015 67.895 ;
        RECT 24.875 67.725 25.045 67.895 ;
        RECT 25.735 67.725 25.905 67.895 ;
        RECT 124.295 67.535 124.465 67.705 ;
        RECT 125.155 67.535 125.325 67.705 ;
        RECT 126.185 67.535 126.355 67.705 ;
        RECT 127.045 67.535 127.215 67.705 ;
        RECT 259.515 67.665 259.685 67.835 ;
        RECT 260.375 67.665 260.545 67.835 ;
        RECT 261.405 67.665 261.575 67.835 ;
        RECT 262.265 67.665 262.435 67.835 ;
        RECT 360.825 67.475 360.995 67.645 ;
        RECT 361.685 67.475 361.855 67.645 ;
        RECT 362.715 67.475 362.885 67.645 ;
        RECT 363.575 67.475 363.745 67.645 ;
        RECT 7.465 63.745 7.635 63.915 ;
        RECT 8.325 63.745 8.495 63.915 ;
        RECT 9.355 63.745 9.525 63.915 ;
        RECT 10.215 63.745 10.385 63.915 ;
        RECT 108.775 63.555 108.945 63.725 ;
        RECT 109.635 63.555 109.805 63.725 ;
        RECT 110.665 63.555 110.835 63.725 ;
        RECT 111.525 63.555 111.695 63.725 ;
        RECT 243.995 63.685 244.165 63.855 ;
        RECT 244.855 63.685 245.025 63.855 ;
        RECT 245.885 63.685 246.055 63.855 ;
        RECT 246.745 63.685 246.915 63.855 ;
        RECT 345.305 63.495 345.475 63.665 ;
        RECT 346.165 63.495 346.335 63.665 ;
        RECT 347.195 63.495 347.365 63.665 ;
        RECT 348.055 63.495 348.225 63.665 ;
        RECT 40.565 62.175 40.735 62.345 ;
        RECT 41.425 62.175 41.595 62.345 ;
        RECT 42.455 62.175 42.625 62.345 ;
        RECT 43.315 62.175 43.485 62.345 ;
        RECT 141.875 61.985 142.045 62.155 ;
        RECT 142.735 61.985 142.905 62.155 ;
        RECT 143.765 61.985 143.935 62.155 ;
        RECT 144.625 61.985 144.795 62.155 ;
        RECT 277.095 62.115 277.265 62.285 ;
        RECT 277.955 62.115 278.125 62.285 ;
        RECT 278.985 62.115 279.155 62.285 ;
        RECT 279.845 62.115 280.015 62.285 ;
        RECT 378.405 61.925 378.575 62.095 ;
        RECT 379.265 61.925 379.435 62.095 ;
        RECT 380.295 61.925 380.465 62.095 ;
        RECT 381.155 61.925 381.325 62.095 ;
        RECT 7.135 55.725 7.305 55.895 ;
        RECT 7.995 55.725 8.165 55.895 ;
        RECT 9.025 55.725 9.195 55.895 ;
        RECT 9.885 55.725 10.055 55.895 ;
        RECT 108.445 55.535 108.615 55.705 ;
        RECT 109.305 55.535 109.475 55.705 ;
        RECT 110.335 55.535 110.505 55.705 ;
        RECT 111.195 55.535 111.365 55.705 ;
        RECT 243.665 55.665 243.835 55.835 ;
        RECT 244.525 55.665 244.695 55.835 ;
        RECT 245.555 55.665 245.725 55.835 ;
        RECT 246.415 55.665 246.585 55.835 ;
        RECT 344.975 55.475 345.145 55.645 ;
        RECT 345.835 55.475 346.005 55.645 ;
        RECT 346.865 55.475 347.035 55.645 ;
        RECT 347.725 55.475 347.895 55.645 ;
        RECT 22.815 53.305 22.985 53.475 ;
        RECT 23.675 53.305 23.845 53.475 ;
        RECT 24.705 53.305 24.875 53.475 ;
        RECT 25.565 53.305 25.735 53.475 ;
        RECT 124.125 53.115 124.295 53.285 ;
        RECT 124.985 53.115 125.155 53.285 ;
        RECT 126.015 53.115 126.185 53.285 ;
        RECT 126.875 53.115 127.045 53.285 ;
        RECT 259.345 53.245 259.515 53.415 ;
        RECT 260.205 53.245 260.375 53.415 ;
        RECT 261.235 53.245 261.405 53.415 ;
        RECT 262.095 53.245 262.265 53.415 ;
        RECT 360.655 53.055 360.825 53.225 ;
        RECT 361.515 53.055 361.685 53.225 ;
        RECT 362.545 53.055 362.715 53.225 ;
        RECT 363.405 53.055 363.575 53.225 ;
        RECT 7.295 49.325 7.465 49.495 ;
        RECT 8.155 49.325 8.325 49.495 ;
        RECT 9.185 49.325 9.355 49.495 ;
        RECT 10.045 49.325 10.215 49.495 ;
        RECT 108.605 49.135 108.775 49.305 ;
        RECT 109.465 49.135 109.635 49.305 ;
        RECT 110.495 49.135 110.665 49.305 ;
        RECT 111.355 49.135 111.525 49.305 ;
        RECT 243.825 49.265 243.995 49.435 ;
        RECT 244.685 49.265 244.855 49.435 ;
        RECT 245.715 49.265 245.885 49.435 ;
        RECT 246.575 49.265 246.745 49.435 ;
        RECT 345.135 49.075 345.305 49.245 ;
        RECT 345.995 49.075 346.165 49.245 ;
        RECT 347.025 49.075 347.195 49.245 ;
        RECT 347.885 49.075 348.055 49.245 ;
        RECT 58.095 46.155 58.265 46.325 ;
        RECT 58.955 46.155 59.125 46.325 ;
        RECT 59.985 46.155 60.155 46.325 ;
        RECT 60.845 46.155 61.015 46.325 ;
        RECT 159.405 45.965 159.575 46.135 ;
        RECT 160.265 45.965 160.435 46.135 ;
        RECT 161.295 45.965 161.465 46.135 ;
        RECT 162.155 45.965 162.325 46.135 ;
        RECT 294.625 46.095 294.795 46.265 ;
        RECT 295.485 46.095 295.655 46.265 ;
        RECT 296.515 46.095 296.685 46.265 ;
        RECT 297.375 46.095 297.545 46.265 ;
        RECT 395.935 45.905 396.105 46.075 ;
        RECT 396.795 45.905 396.965 46.075 ;
        RECT 397.825 45.905 397.995 46.075 ;
        RECT 398.685 45.905 398.855 46.075 ;
        RECT 7.275 40.075 7.445 40.245 ;
        RECT 8.135 40.075 8.305 40.245 ;
        RECT 9.165 40.075 9.335 40.245 ;
        RECT 10.025 40.075 10.195 40.245 ;
        RECT 108.585 39.885 108.755 40.055 ;
        RECT 109.445 39.885 109.615 40.055 ;
        RECT 110.475 39.885 110.645 40.055 ;
        RECT 111.335 39.885 111.505 40.055 ;
        RECT 243.805 40.015 243.975 40.185 ;
        RECT 244.665 40.015 244.835 40.185 ;
        RECT 245.695 40.015 245.865 40.185 ;
        RECT 246.555 40.015 246.725 40.185 ;
        RECT 345.115 39.825 345.285 39.995 ;
        RECT 345.975 39.825 346.145 39.995 ;
        RECT 347.005 39.825 347.175 39.995 ;
        RECT 347.865 39.825 348.035 39.995 ;
        RECT 22.955 37.655 23.125 37.825 ;
        RECT 23.815 37.655 23.985 37.825 ;
        RECT 24.845 37.655 25.015 37.825 ;
        RECT 25.705 37.655 25.875 37.825 ;
        RECT 124.265 37.465 124.435 37.635 ;
        RECT 125.125 37.465 125.295 37.635 ;
        RECT 126.155 37.465 126.325 37.635 ;
        RECT 127.015 37.465 127.185 37.635 ;
        RECT 259.485 37.595 259.655 37.765 ;
        RECT 260.345 37.595 260.515 37.765 ;
        RECT 261.375 37.595 261.545 37.765 ;
        RECT 262.235 37.595 262.405 37.765 ;
        RECT 360.795 37.405 360.965 37.575 ;
        RECT 361.655 37.405 361.825 37.575 ;
        RECT 362.685 37.405 362.855 37.575 ;
        RECT 363.545 37.405 363.715 37.575 ;
        RECT 7.435 33.675 7.605 33.845 ;
        RECT 8.295 33.675 8.465 33.845 ;
        RECT 9.325 33.675 9.495 33.845 ;
        RECT 10.185 33.675 10.355 33.845 ;
        RECT 108.745 33.485 108.915 33.655 ;
        RECT 109.605 33.485 109.775 33.655 ;
        RECT 110.635 33.485 110.805 33.655 ;
        RECT 111.495 33.485 111.665 33.655 ;
        RECT 243.965 33.615 244.135 33.785 ;
        RECT 244.825 33.615 244.995 33.785 ;
        RECT 245.855 33.615 246.025 33.785 ;
        RECT 246.715 33.615 246.885 33.785 ;
        RECT 345.275 33.425 345.445 33.595 ;
        RECT 346.135 33.425 346.305 33.595 ;
        RECT 347.165 33.425 347.335 33.595 ;
        RECT 348.025 33.425 348.195 33.595 ;
        RECT 40.535 32.105 40.705 32.275 ;
        RECT 41.395 32.105 41.565 32.275 ;
        RECT 42.425 32.105 42.595 32.275 ;
        RECT 43.285 32.105 43.455 32.275 ;
        RECT 141.845 31.915 142.015 32.085 ;
        RECT 142.705 31.915 142.875 32.085 ;
        RECT 143.735 31.915 143.905 32.085 ;
        RECT 144.595 31.915 144.765 32.085 ;
        RECT 277.065 32.045 277.235 32.215 ;
        RECT 277.925 32.045 278.095 32.215 ;
        RECT 278.955 32.045 279.125 32.215 ;
        RECT 279.815 32.045 279.985 32.215 ;
        RECT 378.375 31.855 378.545 32.025 ;
        RECT 379.235 31.855 379.405 32.025 ;
        RECT 380.265 31.855 380.435 32.025 ;
        RECT 381.125 31.855 381.295 32.025 ;
        RECT 7.105 25.655 7.275 25.825 ;
        RECT 7.965 25.655 8.135 25.825 ;
        RECT 8.995 25.655 9.165 25.825 ;
        RECT 9.855 25.655 10.025 25.825 ;
        RECT 108.415 25.465 108.585 25.635 ;
        RECT 109.275 25.465 109.445 25.635 ;
        RECT 110.305 25.465 110.475 25.635 ;
        RECT 111.165 25.465 111.335 25.635 ;
        RECT 243.635 25.595 243.805 25.765 ;
        RECT 244.495 25.595 244.665 25.765 ;
        RECT 245.525 25.595 245.695 25.765 ;
        RECT 246.385 25.595 246.555 25.765 ;
        RECT 344.945 25.405 345.115 25.575 ;
        RECT 345.805 25.405 345.975 25.575 ;
        RECT 346.835 25.405 347.005 25.575 ;
        RECT 347.695 25.405 347.865 25.575 ;
        RECT 22.785 23.235 22.955 23.405 ;
        RECT 23.645 23.235 23.815 23.405 ;
        RECT 24.675 23.235 24.845 23.405 ;
        RECT 25.535 23.235 25.705 23.405 ;
        RECT 124.095 23.045 124.265 23.215 ;
        RECT 124.955 23.045 125.125 23.215 ;
        RECT 125.985 23.045 126.155 23.215 ;
        RECT 126.845 23.045 127.015 23.215 ;
        RECT 259.315 23.175 259.485 23.345 ;
        RECT 260.175 23.175 260.345 23.345 ;
        RECT 261.205 23.175 261.375 23.345 ;
        RECT 262.065 23.175 262.235 23.345 ;
        RECT 360.625 22.985 360.795 23.155 ;
        RECT 361.485 22.985 361.655 23.155 ;
        RECT 362.515 22.985 362.685 23.155 ;
        RECT 363.375 22.985 363.545 23.155 ;
        RECT 7.265 19.255 7.435 19.425 ;
        RECT 8.125 19.255 8.295 19.425 ;
        RECT 9.155 19.255 9.325 19.425 ;
        RECT 10.015 19.255 10.185 19.425 ;
        RECT 108.575 19.065 108.745 19.235 ;
        RECT 109.435 19.065 109.605 19.235 ;
        RECT 110.465 19.065 110.635 19.235 ;
        RECT 111.325 19.065 111.495 19.235 ;
        RECT 243.795 19.195 243.965 19.365 ;
        RECT 244.655 19.195 244.825 19.365 ;
        RECT 245.685 19.195 245.855 19.365 ;
        RECT 246.545 19.195 246.715 19.365 ;
        RECT 345.105 19.005 345.275 19.175 ;
        RECT 345.965 19.005 346.135 19.175 ;
        RECT 346.995 19.005 347.165 19.175 ;
        RECT 347.855 19.005 348.025 19.175 ;
      LAYER met1 ;
        RECT 7.950 250.620 11.280 250.990 ;
        RECT 7.950 250.610 11.580 250.620 ;
        RECT 7.950 250.450 11.640 250.610 ;
        RECT 7.940 250.170 11.640 250.450 ;
        RECT 109.260 250.430 112.590 250.800 ;
        RECT 244.480 250.560 247.810 250.930 ;
        RECT 244.480 250.550 248.110 250.560 ;
        RECT 109.260 250.420 112.890 250.430 ;
        RECT 109.260 250.260 112.950 250.420 ;
        RECT 244.480 250.390 248.170 250.550 ;
        RECT 7.940 250.140 11.230 250.170 ;
        RECT 109.250 249.980 112.950 250.260 ;
        RECT 244.470 250.110 248.170 250.390 ;
        RECT 345.790 250.370 349.120 250.740 ;
        RECT 345.790 250.360 349.420 250.370 ;
        RECT 345.790 250.200 349.480 250.360 ;
        RECT 244.470 250.080 247.760 250.110 ;
        RECT 109.250 249.950 112.540 249.980 ;
        RECT 345.780 249.920 349.480 250.200 ;
        RECT 345.780 249.890 349.070 249.920 ;
        RECT 23.630 248.200 26.930 248.570 ;
        RECT 23.630 248.030 27.490 248.200 ;
        RECT 23.620 247.730 27.490 248.030 ;
        RECT 124.940 248.010 128.240 248.380 ;
        RECT 260.160 248.140 263.460 248.510 ;
        RECT 124.940 247.840 128.800 248.010 ;
        RECT 260.160 247.970 264.020 248.140 ;
        RECT 23.620 247.720 26.910 247.730 ;
        RECT 124.930 247.540 128.800 247.840 ;
        RECT 260.150 247.670 264.020 247.970 ;
        RECT 361.470 247.950 364.770 248.320 ;
        RECT 361.470 247.780 365.330 247.950 ;
        RECT 260.150 247.660 263.440 247.670 ;
        RECT 124.930 247.530 128.220 247.540 ;
        RECT 361.460 247.480 365.330 247.780 ;
        RECT 361.460 247.470 364.750 247.480 ;
        RECT 8.110 244.220 11.410 244.590 ;
        RECT 8.110 244.050 11.830 244.220 ;
        RECT 8.100 243.750 11.830 244.050 ;
        RECT 109.420 244.030 112.720 244.400 ;
        RECT 244.640 244.160 247.940 244.530 ;
        RECT 109.420 243.860 113.140 244.030 ;
        RECT 244.640 243.990 248.360 244.160 ;
        RECT 8.100 243.740 11.390 243.750 ;
        RECT 109.410 243.560 113.140 243.860 ;
        RECT 244.630 243.690 248.360 243.990 ;
        RECT 345.950 243.970 349.250 244.340 ;
        RECT 345.950 243.800 349.670 243.970 ;
        RECT 244.630 243.680 247.920 243.690 ;
        RECT 109.410 243.550 112.700 243.560 ;
        RECT 345.940 243.500 349.670 243.800 ;
        RECT 345.940 243.490 349.230 243.500 ;
        RECT 41.210 242.580 44.510 243.020 ;
        RECT 41.210 242.480 45.010 242.580 ;
        RECT 41.200 242.170 45.010 242.480 ;
        RECT 142.520 242.390 145.820 242.830 ;
        RECT 277.740 242.520 281.040 242.960 ;
        RECT 277.740 242.420 281.540 242.520 ;
        RECT 142.520 242.290 146.320 242.390 ;
        RECT 142.510 241.980 146.320 242.290 ;
        RECT 277.730 242.110 281.540 242.420 ;
        RECT 379.050 242.330 382.350 242.770 ;
        RECT 379.050 242.230 382.850 242.330 ;
        RECT 379.040 241.920 382.850 242.230 ;
        RECT 7.780 236.200 11.110 236.570 ;
        RECT 7.780 236.190 11.410 236.200 ;
        RECT 7.780 236.030 11.470 236.190 ;
        RECT 7.770 235.750 11.470 236.030 ;
        RECT 109.090 236.010 112.420 236.380 ;
        RECT 244.310 236.140 247.640 236.510 ;
        RECT 244.310 236.130 247.940 236.140 ;
        RECT 109.090 236.000 112.720 236.010 ;
        RECT 109.090 235.840 112.780 236.000 ;
        RECT 244.310 235.970 248.000 236.130 ;
        RECT 7.770 235.720 11.060 235.750 ;
        RECT 109.080 235.560 112.780 235.840 ;
        RECT 244.300 235.690 248.000 235.970 ;
        RECT 345.620 235.950 348.950 236.320 ;
        RECT 345.620 235.940 349.250 235.950 ;
        RECT 345.620 235.780 349.310 235.940 ;
        RECT 244.300 235.660 247.590 235.690 ;
        RECT 109.080 235.530 112.370 235.560 ;
        RECT 345.610 235.500 349.310 235.780 ;
        RECT 345.610 235.470 348.900 235.500 ;
        RECT 23.460 233.780 26.760 234.150 ;
        RECT 23.460 233.610 27.320 233.780 ;
        RECT 23.450 233.310 27.320 233.610 ;
        RECT 124.770 233.590 128.070 233.960 ;
        RECT 259.990 233.720 263.290 234.090 ;
        RECT 124.770 233.420 128.630 233.590 ;
        RECT 259.990 233.550 263.850 233.720 ;
        RECT 23.450 233.300 26.740 233.310 ;
        RECT 124.760 233.120 128.630 233.420 ;
        RECT 259.980 233.250 263.850 233.550 ;
        RECT 361.300 233.530 364.600 233.900 ;
        RECT 361.300 233.360 365.160 233.530 ;
        RECT 259.980 233.240 263.270 233.250 ;
        RECT 124.760 233.110 128.050 233.120 ;
        RECT 361.290 233.060 365.160 233.360 ;
        RECT 361.290 233.050 364.580 233.060 ;
        RECT 7.940 229.800 11.240 230.170 ;
        RECT 7.940 229.630 11.660 229.800 ;
        RECT 7.930 229.330 11.660 229.630 ;
        RECT 109.250 229.610 112.550 229.980 ;
        RECT 244.470 229.740 247.770 230.110 ;
        RECT 109.250 229.440 112.970 229.610 ;
        RECT 244.470 229.570 248.190 229.740 ;
        RECT 7.930 229.320 11.220 229.330 ;
        RECT 109.240 229.140 112.970 229.440 ;
        RECT 244.460 229.270 248.190 229.570 ;
        RECT 345.780 229.550 349.080 229.920 ;
        RECT 345.780 229.380 349.500 229.550 ;
        RECT 244.460 229.260 247.750 229.270 ;
        RECT 109.240 229.130 112.530 229.140 ;
        RECT 345.770 229.080 349.500 229.380 ;
        RECT 345.770 229.070 349.060 229.080 ;
        RECT 58.740 226.550 62.040 227.000 ;
        RECT 58.740 226.460 62.480 226.550 ;
        RECT 58.730 226.160 62.480 226.460 ;
        RECT 160.050 226.360 163.350 226.810 ;
        RECT 295.270 226.490 298.570 226.940 ;
        RECT 295.270 226.400 299.010 226.490 ;
        RECT 160.050 226.270 163.790 226.360 ;
        RECT 58.730 226.150 62.020 226.160 ;
        RECT 160.040 225.970 163.790 226.270 ;
        RECT 295.260 226.100 299.010 226.400 ;
        RECT 396.580 226.300 399.880 226.750 ;
        RECT 396.580 226.210 400.320 226.300 ;
        RECT 295.260 226.090 298.550 226.100 ;
        RECT 160.040 225.960 163.330 225.970 ;
        RECT 396.570 225.910 400.320 226.210 ;
        RECT 396.570 225.900 399.860 225.910 ;
        RECT 7.920 220.550 11.250 220.920 ;
        RECT 7.920 220.540 11.550 220.550 ;
        RECT 7.920 220.380 11.610 220.540 ;
        RECT 7.910 220.100 11.610 220.380 ;
        RECT 109.230 220.360 112.560 220.730 ;
        RECT 244.450 220.490 247.780 220.860 ;
        RECT 244.450 220.480 248.080 220.490 ;
        RECT 109.230 220.350 112.860 220.360 ;
        RECT 109.230 220.190 112.920 220.350 ;
        RECT 244.450 220.320 248.140 220.480 ;
        RECT 7.910 220.070 11.200 220.100 ;
        RECT 109.220 219.910 112.920 220.190 ;
        RECT 244.440 220.040 248.140 220.320 ;
        RECT 345.760 220.300 349.090 220.670 ;
        RECT 345.760 220.290 349.390 220.300 ;
        RECT 345.760 220.130 349.450 220.290 ;
        RECT 244.440 220.010 247.730 220.040 ;
        RECT 109.220 219.880 112.510 219.910 ;
        RECT 345.750 219.850 349.450 220.130 ;
        RECT 345.750 219.820 349.040 219.850 ;
        RECT 23.600 218.130 26.900 218.500 ;
        RECT 23.600 217.960 27.460 218.130 ;
        RECT 23.590 217.660 27.460 217.960 ;
        RECT 124.910 217.940 128.210 218.310 ;
        RECT 260.130 218.070 263.430 218.440 ;
        RECT 124.910 217.770 128.770 217.940 ;
        RECT 260.130 217.900 263.990 218.070 ;
        RECT 23.590 217.650 26.880 217.660 ;
        RECT 124.900 217.470 128.770 217.770 ;
        RECT 260.120 217.600 263.990 217.900 ;
        RECT 361.440 217.880 364.740 218.250 ;
        RECT 361.440 217.710 365.300 217.880 ;
        RECT 260.120 217.590 263.410 217.600 ;
        RECT 124.900 217.460 128.190 217.470 ;
        RECT 361.430 217.410 365.300 217.710 ;
        RECT 361.430 217.400 364.720 217.410 ;
        RECT 8.080 214.150 11.380 214.520 ;
        RECT 8.080 213.980 11.800 214.150 ;
        RECT 8.070 213.680 11.800 213.980 ;
        RECT 109.390 213.960 112.690 214.330 ;
        RECT 244.610 214.090 247.910 214.460 ;
        RECT 109.390 213.790 113.110 213.960 ;
        RECT 244.610 213.920 248.330 214.090 ;
        RECT 8.070 213.670 11.360 213.680 ;
        RECT 109.380 213.490 113.110 213.790 ;
        RECT 244.600 213.620 248.330 213.920 ;
        RECT 345.920 213.900 349.220 214.270 ;
        RECT 345.920 213.730 349.640 213.900 ;
        RECT 244.600 213.610 247.890 213.620 ;
        RECT 109.380 213.480 112.670 213.490 ;
        RECT 345.910 213.430 349.640 213.730 ;
        RECT 345.910 213.420 349.200 213.430 ;
        RECT 41.180 212.510 44.480 212.950 ;
        RECT 41.180 212.410 44.980 212.510 ;
        RECT 41.170 212.100 44.980 212.410 ;
        RECT 142.490 212.320 145.790 212.760 ;
        RECT 277.710 212.450 281.010 212.890 ;
        RECT 277.710 212.350 281.510 212.450 ;
        RECT 142.490 212.220 146.290 212.320 ;
        RECT 142.480 211.910 146.290 212.220 ;
        RECT 277.700 212.040 281.510 212.350 ;
        RECT 379.020 212.260 382.320 212.700 ;
        RECT 379.020 212.160 382.820 212.260 ;
        RECT 379.010 211.850 382.820 212.160 ;
        RECT 7.750 206.130 11.080 206.500 ;
        RECT 7.750 206.120 11.380 206.130 ;
        RECT 7.750 205.960 11.440 206.120 ;
        RECT 7.740 205.680 11.440 205.960 ;
        RECT 109.060 205.940 112.390 206.310 ;
        RECT 244.280 206.070 247.610 206.440 ;
        RECT 244.280 206.060 247.910 206.070 ;
        RECT 109.060 205.930 112.690 205.940 ;
        RECT 109.060 205.770 112.750 205.930 ;
        RECT 244.280 205.900 247.970 206.060 ;
        RECT 7.740 205.650 11.030 205.680 ;
        RECT 109.050 205.490 112.750 205.770 ;
        RECT 244.270 205.620 247.970 205.900 ;
        RECT 345.590 205.880 348.920 206.250 ;
        RECT 345.590 205.870 349.220 205.880 ;
        RECT 345.590 205.710 349.280 205.870 ;
        RECT 244.270 205.590 247.560 205.620 ;
        RECT 109.050 205.460 112.340 205.490 ;
        RECT 345.580 205.430 349.280 205.710 ;
        RECT 345.580 205.400 348.870 205.430 ;
        RECT 23.430 203.710 26.730 204.080 ;
        RECT 23.430 203.540 27.290 203.710 ;
        RECT 23.420 203.240 27.290 203.540 ;
        RECT 124.740 203.520 128.040 203.890 ;
        RECT 259.960 203.650 263.260 204.020 ;
        RECT 124.740 203.350 128.600 203.520 ;
        RECT 259.960 203.480 263.820 203.650 ;
        RECT 23.420 203.230 26.710 203.240 ;
        RECT 124.730 203.050 128.600 203.350 ;
        RECT 259.950 203.180 263.820 203.480 ;
        RECT 361.270 203.460 364.570 203.830 ;
        RECT 361.270 203.290 365.130 203.460 ;
        RECT 259.950 203.170 263.240 203.180 ;
        RECT 124.730 203.040 128.020 203.050 ;
        RECT 361.260 202.990 365.130 203.290 ;
        RECT 361.260 202.980 364.550 202.990 ;
        RECT 72.940 200.360 76.240 200.710 ;
        RECT 72.940 200.170 76.810 200.360 ;
        RECT 7.910 199.730 11.210 200.100 ;
        RECT 72.930 199.880 76.810 200.170 ;
        RECT 174.250 200.170 177.550 200.520 ;
        RECT 309.470 200.300 312.770 200.650 ;
        RECT 174.250 199.980 178.120 200.170 ;
        RECT 309.470 200.110 313.340 200.300 ;
        RECT 72.930 199.860 76.220 199.880 ;
        RECT 7.910 199.560 11.630 199.730 ;
        RECT 7.900 199.260 11.630 199.560 ;
        RECT 109.220 199.540 112.520 199.910 ;
        RECT 174.240 199.690 178.120 199.980 ;
        RECT 174.240 199.670 177.530 199.690 ;
        RECT 244.440 199.670 247.740 200.040 ;
        RECT 309.460 199.820 313.340 200.110 ;
        RECT 410.780 200.110 414.080 200.460 ;
        RECT 410.780 199.920 414.650 200.110 ;
        RECT 309.460 199.800 312.750 199.820 ;
        RECT 109.220 199.370 112.940 199.540 ;
        RECT 244.440 199.500 248.160 199.670 ;
        RECT 7.900 199.250 11.190 199.260 ;
        RECT 109.210 199.070 112.940 199.370 ;
        RECT 244.430 199.200 248.160 199.500 ;
        RECT 345.750 199.480 349.050 199.850 ;
        RECT 410.770 199.630 414.650 199.920 ;
        RECT 410.770 199.610 414.060 199.630 ;
        RECT 345.750 199.310 349.470 199.480 ;
        RECT 244.430 199.190 247.720 199.200 ;
        RECT 109.210 199.060 112.500 199.070 ;
        RECT 345.740 199.010 349.470 199.310 ;
        RECT 345.740 199.000 349.030 199.010 ;
        RECT 7.600 190.700 10.930 191.070 ;
        RECT 7.600 190.690 11.230 190.700 ;
        RECT 7.600 190.530 11.290 190.690 ;
        RECT 7.590 190.250 11.290 190.530 ;
        RECT 108.910 190.510 112.240 190.880 ;
        RECT 244.130 190.640 247.460 191.010 ;
        RECT 244.130 190.630 247.760 190.640 ;
        RECT 108.910 190.500 112.540 190.510 ;
        RECT 108.910 190.340 112.600 190.500 ;
        RECT 244.130 190.470 247.820 190.630 ;
        RECT 7.590 190.220 10.880 190.250 ;
        RECT 108.900 190.060 112.600 190.340 ;
        RECT 244.120 190.190 247.820 190.470 ;
        RECT 345.440 190.450 348.770 190.820 ;
        RECT 345.440 190.440 349.070 190.450 ;
        RECT 345.440 190.280 349.130 190.440 ;
        RECT 244.120 190.160 247.410 190.190 ;
        RECT 108.900 190.030 112.190 190.060 ;
        RECT 345.430 190.000 349.130 190.280 ;
        RECT 345.430 189.970 348.720 190.000 ;
        RECT 23.280 188.280 26.580 188.650 ;
        RECT 23.280 188.110 27.140 188.280 ;
        RECT 23.270 187.810 27.140 188.110 ;
        RECT 124.590 188.090 127.890 188.460 ;
        RECT 259.810 188.220 263.110 188.590 ;
        RECT 124.590 187.920 128.450 188.090 ;
        RECT 259.810 188.050 263.670 188.220 ;
        RECT 23.270 187.800 26.560 187.810 ;
        RECT 124.580 187.620 128.450 187.920 ;
        RECT 259.800 187.750 263.670 188.050 ;
        RECT 361.120 188.030 364.420 188.400 ;
        RECT 361.120 187.860 364.980 188.030 ;
        RECT 259.800 187.740 263.090 187.750 ;
        RECT 124.580 187.610 127.870 187.620 ;
        RECT 361.110 187.560 364.980 187.860 ;
        RECT 361.110 187.550 364.400 187.560 ;
        RECT 7.760 184.300 11.060 184.670 ;
        RECT 7.760 184.130 11.480 184.300 ;
        RECT 7.750 183.830 11.480 184.130 ;
        RECT 109.070 184.110 112.370 184.480 ;
        RECT 244.290 184.240 247.590 184.610 ;
        RECT 109.070 183.940 112.790 184.110 ;
        RECT 244.290 184.070 248.010 184.240 ;
        RECT 7.750 183.820 11.040 183.830 ;
        RECT 109.060 183.640 112.790 183.940 ;
        RECT 244.280 183.770 248.010 184.070 ;
        RECT 345.600 184.050 348.900 184.420 ;
        RECT 345.600 183.880 349.320 184.050 ;
        RECT 244.280 183.760 247.570 183.770 ;
        RECT 109.060 183.630 112.350 183.640 ;
        RECT 345.590 183.580 349.320 183.880 ;
        RECT 345.590 183.570 348.880 183.580 ;
        RECT 40.860 182.660 44.160 183.100 ;
        RECT 40.860 182.560 44.660 182.660 ;
        RECT 40.850 182.250 44.660 182.560 ;
        RECT 142.170 182.470 145.470 182.910 ;
        RECT 277.390 182.600 280.690 183.040 ;
        RECT 277.390 182.500 281.190 182.600 ;
        RECT 142.170 182.370 145.970 182.470 ;
        RECT 142.160 182.060 145.970 182.370 ;
        RECT 277.380 182.190 281.190 182.500 ;
        RECT 378.700 182.410 382.000 182.850 ;
        RECT 378.700 182.310 382.500 182.410 ;
        RECT 378.690 182.000 382.500 182.310 ;
        RECT 7.430 176.280 10.760 176.650 ;
        RECT 7.430 176.270 11.060 176.280 ;
        RECT 7.430 176.110 11.120 176.270 ;
        RECT 7.420 175.830 11.120 176.110 ;
        RECT 108.740 176.090 112.070 176.460 ;
        RECT 243.960 176.220 247.290 176.590 ;
        RECT 243.960 176.210 247.590 176.220 ;
        RECT 108.740 176.080 112.370 176.090 ;
        RECT 108.740 175.920 112.430 176.080 ;
        RECT 243.960 176.050 247.650 176.210 ;
        RECT 7.420 175.800 10.710 175.830 ;
        RECT 108.730 175.640 112.430 175.920 ;
        RECT 243.950 175.770 247.650 176.050 ;
        RECT 345.270 176.030 348.600 176.400 ;
        RECT 345.270 176.020 348.900 176.030 ;
        RECT 345.270 175.860 348.960 176.020 ;
        RECT 243.950 175.740 247.240 175.770 ;
        RECT 108.730 175.610 112.020 175.640 ;
        RECT 345.260 175.580 348.960 175.860 ;
        RECT 345.260 175.550 348.550 175.580 ;
        RECT 23.110 173.860 26.410 174.230 ;
        RECT 23.110 173.690 26.970 173.860 ;
        RECT 23.100 173.390 26.970 173.690 ;
        RECT 124.420 173.670 127.720 174.040 ;
        RECT 259.640 173.800 262.940 174.170 ;
        RECT 124.420 173.500 128.280 173.670 ;
        RECT 259.640 173.630 263.500 173.800 ;
        RECT 23.100 173.380 26.390 173.390 ;
        RECT 124.410 173.200 128.280 173.500 ;
        RECT 259.630 173.330 263.500 173.630 ;
        RECT 360.950 173.610 364.250 173.980 ;
        RECT 360.950 173.440 364.810 173.610 ;
        RECT 259.630 173.320 262.920 173.330 ;
        RECT 124.410 173.190 127.700 173.200 ;
        RECT 360.940 173.140 364.810 173.440 ;
        RECT 360.940 173.130 364.230 173.140 ;
        RECT 7.590 169.880 10.890 170.250 ;
        RECT 7.590 169.710 11.310 169.880 ;
        RECT 7.580 169.410 11.310 169.710 ;
        RECT 108.900 169.690 112.200 170.060 ;
        RECT 244.120 169.820 247.420 170.190 ;
        RECT 108.900 169.520 112.620 169.690 ;
        RECT 244.120 169.650 247.840 169.820 ;
        RECT 7.580 169.400 10.870 169.410 ;
        RECT 108.890 169.220 112.620 169.520 ;
        RECT 244.110 169.350 247.840 169.650 ;
        RECT 345.430 169.630 348.730 170.000 ;
        RECT 345.430 169.460 349.150 169.630 ;
        RECT 244.110 169.340 247.400 169.350 ;
        RECT 108.890 169.210 112.180 169.220 ;
        RECT 345.420 169.160 349.150 169.460 ;
        RECT 345.420 169.150 348.710 169.160 ;
        RECT 58.390 166.630 61.690 167.080 ;
        RECT 58.390 166.540 62.130 166.630 ;
        RECT 58.380 166.240 62.130 166.540 ;
        RECT 159.700 166.440 163.000 166.890 ;
        RECT 294.920 166.570 298.220 167.020 ;
        RECT 294.920 166.480 298.660 166.570 ;
        RECT 159.700 166.350 163.440 166.440 ;
        RECT 58.380 166.230 61.670 166.240 ;
        RECT 159.690 166.050 163.440 166.350 ;
        RECT 294.910 166.180 298.660 166.480 ;
        RECT 396.230 166.380 399.530 166.830 ;
        RECT 396.230 166.290 399.970 166.380 ;
        RECT 294.910 166.170 298.200 166.180 ;
        RECT 159.690 166.040 162.980 166.050 ;
        RECT 396.220 165.990 399.970 166.290 ;
        RECT 396.220 165.980 399.510 165.990 ;
        RECT 7.570 160.630 10.900 161.000 ;
        RECT 7.570 160.620 11.200 160.630 ;
        RECT 7.570 160.460 11.260 160.620 ;
        RECT 7.560 160.180 11.260 160.460 ;
        RECT 108.880 160.440 112.210 160.810 ;
        RECT 244.100 160.570 247.430 160.940 ;
        RECT 244.100 160.560 247.730 160.570 ;
        RECT 108.880 160.430 112.510 160.440 ;
        RECT 108.880 160.270 112.570 160.430 ;
        RECT 244.100 160.400 247.790 160.560 ;
        RECT 7.560 160.150 10.850 160.180 ;
        RECT 108.870 159.990 112.570 160.270 ;
        RECT 244.090 160.120 247.790 160.400 ;
        RECT 345.410 160.380 348.740 160.750 ;
        RECT 345.410 160.370 349.040 160.380 ;
        RECT 345.410 160.210 349.100 160.370 ;
        RECT 244.090 160.090 247.380 160.120 ;
        RECT 108.870 159.960 112.160 159.990 ;
        RECT 345.400 159.930 349.100 160.210 ;
        RECT 345.400 159.900 348.690 159.930 ;
        RECT 23.250 158.210 26.550 158.580 ;
        RECT 23.250 158.040 27.110 158.210 ;
        RECT 23.240 157.740 27.110 158.040 ;
        RECT 124.560 158.020 127.860 158.390 ;
        RECT 259.780 158.150 263.080 158.520 ;
        RECT 124.560 157.850 128.420 158.020 ;
        RECT 259.780 157.980 263.640 158.150 ;
        RECT 23.240 157.730 26.530 157.740 ;
        RECT 124.550 157.550 128.420 157.850 ;
        RECT 259.770 157.680 263.640 157.980 ;
        RECT 361.090 157.960 364.390 158.330 ;
        RECT 361.090 157.790 364.950 157.960 ;
        RECT 259.770 157.670 263.060 157.680 ;
        RECT 124.550 157.540 127.840 157.550 ;
        RECT 361.080 157.490 364.950 157.790 ;
        RECT 361.080 157.480 364.370 157.490 ;
        RECT 7.730 154.230 11.030 154.600 ;
        RECT 7.730 154.060 11.450 154.230 ;
        RECT 7.720 153.760 11.450 154.060 ;
        RECT 109.040 154.040 112.340 154.410 ;
        RECT 244.260 154.170 247.560 154.540 ;
        RECT 109.040 153.870 112.760 154.040 ;
        RECT 244.260 154.000 247.980 154.170 ;
        RECT 7.720 153.750 11.010 153.760 ;
        RECT 109.030 153.570 112.760 153.870 ;
        RECT 244.250 153.700 247.980 154.000 ;
        RECT 345.570 153.980 348.870 154.350 ;
        RECT 345.570 153.810 349.290 153.980 ;
        RECT 244.250 153.690 247.540 153.700 ;
        RECT 109.030 153.560 112.320 153.570 ;
        RECT 345.560 153.510 349.290 153.810 ;
        RECT 345.560 153.500 348.850 153.510 ;
        RECT 40.830 152.590 44.130 153.030 ;
        RECT 40.830 152.490 44.630 152.590 ;
        RECT 40.820 152.180 44.630 152.490 ;
        RECT 142.140 152.400 145.440 152.840 ;
        RECT 277.360 152.530 280.660 152.970 ;
        RECT 277.360 152.430 281.160 152.530 ;
        RECT 142.140 152.300 145.940 152.400 ;
        RECT 142.130 151.990 145.940 152.300 ;
        RECT 277.350 152.120 281.160 152.430 ;
        RECT 378.670 152.340 381.970 152.780 ;
        RECT 378.670 152.240 382.470 152.340 ;
        RECT 378.660 151.930 382.470 152.240 ;
        RECT 7.400 146.210 10.730 146.580 ;
        RECT 7.400 146.200 11.030 146.210 ;
        RECT 7.400 146.040 11.090 146.200 ;
        RECT 7.390 145.760 11.090 146.040 ;
        RECT 108.710 146.020 112.040 146.390 ;
        RECT 243.930 146.150 247.260 146.520 ;
        RECT 243.930 146.140 247.560 146.150 ;
        RECT 108.710 146.010 112.340 146.020 ;
        RECT 108.710 145.850 112.400 146.010 ;
        RECT 243.930 145.980 247.620 146.140 ;
        RECT 7.390 145.730 10.680 145.760 ;
        RECT 108.700 145.570 112.400 145.850 ;
        RECT 243.920 145.700 247.620 145.980 ;
        RECT 345.240 145.960 348.570 146.330 ;
        RECT 345.240 145.950 348.870 145.960 ;
        RECT 345.240 145.790 348.930 145.950 ;
        RECT 243.920 145.670 247.210 145.700 ;
        RECT 108.700 145.540 111.990 145.570 ;
        RECT 345.230 145.510 348.930 145.790 ;
        RECT 345.230 145.480 348.520 145.510 ;
        RECT 23.080 143.790 26.380 144.160 ;
        RECT 23.080 143.620 26.940 143.790 ;
        RECT 23.070 143.320 26.940 143.620 ;
        RECT 124.390 143.600 127.690 143.970 ;
        RECT 259.610 143.730 262.910 144.100 ;
        RECT 124.390 143.430 128.250 143.600 ;
        RECT 259.610 143.560 263.470 143.730 ;
        RECT 23.070 143.310 26.360 143.320 ;
        RECT 124.380 143.130 128.250 143.430 ;
        RECT 259.600 143.260 263.470 143.560 ;
        RECT 360.920 143.540 364.220 143.910 ;
        RECT 360.920 143.370 364.780 143.540 ;
        RECT 259.600 143.250 262.890 143.260 ;
        RECT 124.380 143.120 127.670 143.130 ;
        RECT 360.910 143.070 364.780 143.370 ;
        RECT 360.910 143.060 364.200 143.070 ;
        RECT 7.560 139.810 10.860 140.180 ;
        RECT 7.560 139.640 11.280 139.810 ;
        RECT 7.550 139.340 11.280 139.640 ;
        RECT 108.870 139.620 112.170 139.990 ;
        RECT 244.090 139.750 247.390 140.120 ;
        RECT 108.870 139.450 112.590 139.620 ;
        RECT 7.550 139.330 10.840 139.340 ;
        RECT 108.860 139.150 112.590 139.450 ;
        RECT 216.860 139.240 220.160 139.710 ;
        RECT 244.090 139.580 247.810 139.750 ;
        RECT 244.080 139.280 247.810 139.580 ;
        RECT 345.400 139.560 348.700 139.930 ;
        RECT 345.400 139.390 349.120 139.560 ;
        RECT 244.080 139.270 247.370 139.280 ;
        RECT 216.860 139.170 220.670 139.240 ;
        RECT 108.860 139.140 112.150 139.150 ;
        RECT 216.850 138.860 220.670 139.170 ;
        RECT 345.390 139.090 349.120 139.390 ;
        RECT 453.390 139.180 456.690 139.650 ;
        RECT 453.390 139.110 457.200 139.180 ;
        RECT 345.390 139.080 348.680 139.090 ;
        RECT 453.380 138.800 457.200 139.110 ;
        RECT 89.270 137.130 92.570 137.570 ;
        RECT 89.270 137.030 93.070 137.130 ;
        RECT 89.260 136.730 93.070 137.030 ;
        RECT 190.580 136.940 193.880 137.380 ;
        RECT 325.800 137.070 329.100 137.510 ;
        RECT 325.800 136.970 329.600 137.070 ;
        RECT 190.580 136.840 194.380 136.940 ;
        RECT 89.260 136.720 92.550 136.730 ;
        RECT 190.570 136.540 194.380 136.840 ;
        RECT 325.790 136.670 329.600 136.970 ;
        RECT 427.110 136.880 430.410 137.320 ;
        RECT 427.110 136.780 430.910 136.880 ;
        RECT 325.790 136.660 329.080 136.670 ;
        RECT 190.570 136.530 193.860 136.540 ;
        RECT 427.100 136.480 430.910 136.780 ;
        RECT 470.690 136.830 473.990 137.300 ;
        RECT 470.690 136.760 474.400 136.830 ;
        RECT 427.100 136.470 430.390 136.480 ;
        RECT 470.680 136.450 474.400 136.760 ;
        RECT 7.450 130.380 10.780 130.750 ;
        RECT 7.450 130.370 11.080 130.380 ;
        RECT 7.450 130.210 11.140 130.370 ;
        RECT 7.440 129.930 11.140 130.210 ;
        RECT 108.760 130.190 112.090 130.560 ;
        RECT 243.980 130.320 247.310 130.690 ;
        RECT 243.980 130.310 247.610 130.320 ;
        RECT 108.760 130.180 112.390 130.190 ;
        RECT 108.760 130.020 112.450 130.180 ;
        RECT 243.980 130.150 247.670 130.310 ;
        RECT 7.440 129.900 10.730 129.930 ;
        RECT 108.750 129.740 112.450 130.020 ;
        RECT 243.970 129.870 247.670 130.150 ;
        RECT 345.290 130.130 348.620 130.500 ;
        RECT 345.290 130.120 348.920 130.130 ;
        RECT 345.290 129.960 348.980 130.120 ;
        RECT 243.970 129.840 247.260 129.870 ;
        RECT 108.750 129.710 112.040 129.740 ;
        RECT 345.280 129.680 348.980 129.960 ;
        RECT 345.280 129.650 348.570 129.680 ;
        RECT 23.130 127.960 26.430 128.330 ;
        RECT 23.130 127.790 26.990 127.960 ;
        RECT 23.120 127.490 26.990 127.790 ;
        RECT 124.440 127.770 127.740 128.140 ;
        RECT 259.660 127.900 262.960 128.270 ;
        RECT 124.440 127.600 128.300 127.770 ;
        RECT 259.660 127.730 263.520 127.900 ;
        RECT 23.120 127.480 26.410 127.490 ;
        RECT 124.430 127.300 128.300 127.600 ;
        RECT 259.650 127.430 263.520 127.730 ;
        RECT 360.970 127.710 364.270 128.080 ;
        RECT 360.970 127.540 364.830 127.710 ;
        RECT 259.650 127.420 262.940 127.430 ;
        RECT 124.430 127.290 127.720 127.300 ;
        RECT 360.960 127.240 364.830 127.540 ;
        RECT 360.960 127.230 364.250 127.240 ;
        RECT 7.610 123.980 10.910 124.350 ;
        RECT 7.610 123.810 11.330 123.980 ;
        RECT 7.600 123.510 11.330 123.810 ;
        RECT 108.920 123.790 112.220 124.160 ;
        RECT 244.140 123.920 247.440 124.290 ;
        RECT 108.920 123.620 112.640 123.790 ;
        RECT 244.140 123.750 247.860 123.920 ;
        RECT 7.600 123.500 10.890 123.510 ;
        RECT 108.910 123.320 112.640 123.620 ;
        RECT 244.130 123.450 247.860 123.750 ;
        RECT 345.450 123.730 348.750 124.100 ;
        RECT 345.450 123.560 349.170 123.730 ;
        RECT 244.130 123.440 247.420 123.450 ;
        RECT 108.910 123.310 112.200 123.320 ;
        RECT 345.440 123.260 349.170 123.560 ;
        RECT 345.440 123.250 348.730 123.260 ;
        RECT 40.710 122.340 44.010 122.780 ;
        RECT 40.710 122.240 44.510 122.340 ;
        RECT 40.700 121.930 44.510 122.240 ;
        RECT 142.020 122.150 145.320 122.590 ;
        RECT 277.240 122.280 280.540 122.720 ;
        RECT 277.240 122.180 281.040 122.280 ;
        RECT 142.020 122.050 145.820 122.150 ;
        RECT 142.010 121.740 145.820 122.050 ;
        RECT 277.230 121.870 281.040 122.180 ;
        RECT 378.550 122.090 381.850 122.530 ;
        RECT 378.550 121.990 382.350 122.090 ;
        RECT 378.540 121.680 382.350 121.990 ;
        RECT 7.280 115.960 10.610 116.330 ;
        RECT 7.280 115.950 10.910 115.960 ;
        RECT 7.280 115.790 10.970 115.950 ;
        RECT 7.270 115.510 10.970 115.790 ;
        RECT 108.590 115.770 111.920 116.140 ;
        RECT 243.810 115.900 247.140 116.270 ;
        RECT 243.810 115.890 247.440 115.900 ;
        RECT 108.590 115.760 112.220 115.770 ;
        RECT 108.590 115.600 112.280 115.760 ;
        RECT 243.810 115.730 247.500 115.890 ;
        RECT 7.270 115.480 10.560 115.510 ;
        RECT 108.580 115.320 112.280 115.600 ;
        RECT 243.800 115.450 247.500 115.730 ;
        RECT 345.120 115.710 348.450 116.080 ;
        RECT 345.120 115.700 348.750 115.710 ;
        RECT 345.120 115.540 348.810 115.700 ;
        RECT 243.800 115.420 247.090 115.450 ;
        RECT 108.580 115.290 111.870 115.320 ;
        RECT 345.110 115.260 348.810 115.540 ;
        RECT 345.110 115.230 348.400 115.260 ;
        RECT 22.960 113.540 26.260 113.910 ;
        RECT 22.960 113.370 26.820 113.540 ;
        RECT 22.950 113.070 26.820 113.370 ;
        RECT 124.270 113.350 127.570 113.720 ;
        RECT 259.490 113.480 262.790 113.850 ;
        RECT 124.270 113.180 128.130 113.350 ;
        RECT 259.490 113.310 263.350 113.480 ;
        RECT 22.950 113.060 26.240 113.070 ;
        RECT 124.260 112.880 128.130 113.180 ;
        RECT 259.480 113.010 263.350 113.310 ;
        RECT 360.800 113.290 364.100 113.660 ;
        RECT 360.800 113.120 364.660 113.290 ;
        RECT 259.480 113.000 262.770 113.010 ;
        RECT 124.260 112.870 127.550 112.880 ;
        RECT 360.790 112.820 364.660 113.120 ;
        RECT 360.790 112.810 364.080 112.820 ;
        RECT 7.440 109.560 10.740 109.930 ;
        RECT 7.440 109.390 11.160 109.560 ;
        RECT 7.430 109.090 11.160 109.390 ;
        RECT 108.750 109.370 112.050 109.740 ;
        RECT 243.970 109.500 247.270 109.870 ;
        RECT 108.750 109.200 112.470 109.370 ;
        RECT 243.970 109.330 247.690 109.500 ;
        RECT 7.430 109.080 10.720 109.090 ;
        RECT 108.740 108.900 112.470 109.200 ;
        RECT 243.960 109.030 247.690 109.330 ;
        RECT 345.280 109.310 348.580 109.680 ;
        RECT 345.280 109.140 349.000 109.310 ;
        RECT 243.960 109.020 247.250 109.030 ;
        RECT 108.740 108.890 112.030 108.900 ;
        RECT 345.270 108.840 349.000 109.140 ;
        RECT 345.270 108.830 348.560 108.840 ;
        RECT 58.240 106.310 61.540 106.760 ;
        RECT 58.240 106.220 61.980 106.310 ;
        RECT 58.230 105.920 61.980 106.220 ;
        RECT 159.550 106.120 162.850 106.570 ;
        RECT 294.770 106.250 298.070 106.700 ;
        RECT 294.770 106.160 298.510 106.250 ;
        RECT 159.550 106.030 163.290 106.120 ;
        RECT 58.230 105.910 61.520 105.920 ;
        RECT 159.540 105.730 163.290 106.030 ;
        RECT 294.760 105.860 298.510 106.160 ;
        RECT 396.080 106.060 399.380 106.510 ;
        RECT 396.080 105.970 399.820 106.060 ;
        RECT 294.760 105.850 298.050 105.860 ;
        RECT 159.540 105.720 162.830 105.730 ;
        RECT 396.070 105.670 399.820 105.970 ;
        RECT 396.070 105.660 399.360 105.670 ;
        RECT 7.420 100.310 10.750 100.680 ;
        RECT 7.420 100.300 11.050 100.310 ;
        RECT 7.420 100.140 11.110 100.300 ;
        RECT 7.410 99.860 11.110 100.140 ;
        RECT 108.730 100.120 112.060 100.490 ;
        RECT 243.950 100.250 247.280 100.620 ;
        RECT 243.950 100.240 247.580 100.250 ;
        RECT 108.730 100.110 112.360 100.120 ;
        RECT 108.730 99.950 112.420 100.110 ;
        RECT 243.950 100.080 247.640 100.240 ;
        RECT 7.410 99.830 10.700 99.860 ;
        RECT 108.720 99.670 112.420 99.950 ;
        RECT 243.940 99.800 247.640 100.080 ;
        RECT 345.260 100.060 348.590 100.430 ;
        RECT 345.260 100.050 348.890 100.060 ;
        RECT 345.260 99.890 348.950 100.050 ;
        RECT 243.940 99.770 247.230 99.800 ;
        RECT 108.720 99.640 112.010 99.670 ;
        RECT 345.250 99.610 348.950 99.890 ;
        RECT 345.250 99.580 348.540 99.610 ;
        RECT 23.100 97.890 26.400 98.260 ;
        RECT 23.100 97.720 26.960 97.890 ;
        RECT 23.090 97.420 26.960 97.720 ;
        RECT 124.410 97.700 127.710 98.070 ;
        RECT 259.630 97.830 262.930 98.200 ;
        RECT 124.410 97.530 128.270 97.700 ;
        RECT 259.630 97.660 263.490 97.830 ;
        RECT 23.090 97.410 26.380 97.420 ;
        RECT 124.400 97.230 128.270 97.530 ;
        RECT 259.620 97.360 263.490 97.660 ;
        RECT 360.940 97.640 364.240 98.010 ;
        RECT 360.940 97.470 364.800 97.640 ;
        RECT 259.620 97.350 262.910 97.360 ;
        RECT 124.400 97.220 127.690 97.230 ;
        RECT 360.930 97.170 364.800 97.470 ;
        RECT 360.930 97.160 364.220 97.170 ;
        RECT 7.580 93.910 10.880 94.280 ;
        RECT 7.580 93.740 11.300 93.910 ;
        RECT 7.570 93.440 11.300 93.740 ;
        RECT 108.890 93.720 112.190 94.090 ;
        RECT 244.110 93.850 247.410 94.220 ;
        RECT 108.890 93.550 112.610 93.720 ;
        RECT 244.110 93.680 247.830 93.850 ;
        RECT 7.570 93.430 10.860 93.440 ;
        RECT 108.880 93.250 112.610 93.550 ;
        RECT 244.100 93.380 247.830 93.680 ;
        RECT 345.420 93.660 348.720 94.030 ;
        RECT 345.420 93.490 349.140 93.660 ;
        RECT 244.100 93.370 247.390 93.380 ;
        RECT 108.880 93.240 112.170 93.250 ;
        RECT 345.410 93.190 349.140 93.490 ;
        RECT 345.410 93.180 348.700 93.190 ;
        RECT 40.680 92.270 43.980 92.710 ;
        RECT 40.680 92.170 44.480 92.270 ;
        RECT 40.670 91.860 44.480 92.170 ;
        RECT 141.990 92.080 145.290 92.520 ;
        RECT 277.210 92.210 280.510 92.650 ;
        RECT 277.210 92.110 281.010 92.210 ;
        RECT 141.990 91.980 145.790 92.080 ;
        RECT 141.980 91.670 145.790 91.980 ;
        RECT 277.200 91.800 281.010 92.110 ;
        RECT 378.520 92.020 381.820 92.460 ;
        RECT 378.520 91.920 382.320 92.020 ;
        RECT 378.510 91.610 382.320 91.920 ;
        RECT 7.250 85.890 10.580 86.260 ;
        RECT 7.250 85.880 10.880 85.890 ;
        RECT 7.250 85.720 10.940 85.880 ;
        RECT 7.240 85.440 10.940 85.720 ;
        RECT 108.560 85.700 111.890 86.070 ;
        RECT 243.780 85.830 247.110 86.200 ;
        RECT 243.780 85.820 247.410 85.830 ;
        RECT 108.560 85.690 112.190 85.700 ;
        RECT 108.560 85.530 112.250 85.690 ;
        RECT 243.780 85.660 247.470 85.820 ;
        RECT 7.240 85.410 10.530 85.440 ;
        RECT 108.550 85.250 112.250 85.530 ;
        RECT 243.770 85.380 247.470 85.660 ;
        RECT 345.090 85.640 348.420 86.010 ;
        RECT 345.090 85.630 348.720 85.640 ;
        RECT 345.090 85.470 348.780 85.630 ;
        RECT 243.770 85.350 247.060 85.380 ;
        RECT 108.550 85.220 111.840 85.250 ;
        RECT 345.080 85.190 348.780 85.470 ;
        RECT 345.080 85.160 348.370 85.190 ;
        RECT 22.930 83.470 26.230 83.840 ;
        RECT 22.930 83.300 26.790 83.470 ;
        RECT 22.920 83.000 26.790 83.300 ;
        RECT 124.240 83.280 127.540 83.650 ;
        RECT 259.460 83.410 262.760 83.780 ;
        RECT 124.240 83.110 128.100 83.280 ;
        RECT 259.460 83.240 263.320 83.410 ;
        RECT 22.920 82.990 26.210 83.000 ;
        RECT 124.230 82.810 128.100 83.110 ;
        RECT 259.450 82.940 263.320 83.240 ;
        RECT 360.770 83.220 364.070 83.590 ;
        RECT 360.770 83.050 364.630 83.220 ;
        RECT 259.450 82.930 262.740 82.940 ;
        RECT 124.230 82.800 127.520 82.810 ;
        RECT 360.760 82.750 364.630 83.050 ;
        RECT 360.760 82.740 364.050 82.750 ;
        RECT 72.440 80.120 75.740 80.470 ;
        RECT 72.440 79.930 76.310 80.120 ;
        RECT 7.410 79.490 10.710 79.860 ;
        RECT 72.430 79.640 76.310 79.930 ;
        RECT 173.750 79.930 177.050 80.280 ;
        RECT 308.970 80.060 312.270 80.410 ;
        RECT 173.750 79.740 177.620 79.930 ;
        RECT 308.970 79.870 312.840 80.060 ;
        RECT 72.430 79.620 75.720 79.640 ;
        RECT 7.410 79.320 11.130 79.490 ;
        RECT 7.400 79.020 11.130 79.320 ;
        RECT 108.720 79.300 112.020 79.670 ;
        RECT 173.740 79.450 177.620 79.740 ;
        RECT 173.740 79.430 177.030 79.450 ;
        RECT 243.940 79.430 247.240 79.800 ;
        RECT 308.960 79.580 312.840 79.870 ;
        RECT 410.280 79.870 413.580 80.220 ;
        RECT 410.280 79.680 414.150 79.870 ;
        RECT 308.960 79.560 312.250 79.580 ;
        RECT 108.720 79.130 112.440 79.300 ;
        RECT 243.940 79.260 247.660 79.430 ;
        RECT 7.400 79.010 10.690 79.020 ;
        RECT 108.710 78.830 112.440 79.130 ;
        RECT 243.930 78.960 247.660 79.260 ;
        RECT 345.250 79.240 348.550 79.610 ;
        RECT 410.270 79.390 414.150 79.680 ;
        RECT 410.270 79.370 413.560 79.390 ;
        RECT 345.250 79.070 348.970 79.240 ;
        RECT 243.930 78.950 247.220 78.960 ;
        RECT 108.710 78.820 112.000 78.830 ;
        RECT 345.240 78.770 348.970 79.070 ;
        RECT 345.240 78.760 348.530 78.770 ;
        RECT 7.100 70.460 10.430 70.830 ;
        RECT 7.100 70.450 10.730 70.460 ;
        RECT 7.100 70.290 10.790 70.450 ;
        RECT 7.090 70.010 10.790 70.290 ;
        RECT 108.410 70.270 111.740 70.640 ;
        RECT 243.630 70.400 246.960 70.770 ;
        RECT 243.630 70.390 247.260 70.400 ;
        RECT 108.410 70.260 112.040 70.270 ;
        RECT 108.410 70.100 112.100 70.260 ;
        RECT 243.630 70.230 247.320 70.390 ;
        RECT 7.090 69.980 10.380 70.010 ;
        RECT 108.400 69.820 112.100 70.100 ;
        RECT 243.620 69.950 247.320 70.230 ;
        RECT 344.940 70.210 348.270 70.580 ;
        RECT 344.940 70.200 348.570 70.210 ;
        RECT 344.940 70.040 348.630 70.200 ;
        RECT 243.620 69.920 246.910 69.950 ;
        RECT 108.400 69.790 111.690 69.820 ;
        RECT 344.930 69.760 348.630 70.040 ;
        RECT 344.930 69.730 348.220 69.760 ;
        RECT 22.780 68.040 26.080 68.410 ;
        RECT 22.780 67.870 26.640 68.040 ;
        RECT 22.770 67.570 26.640 67.870 ;
        RECT 124.090 67.850 127.390 68.220 ;
        RECT 259.310 67.980 262.610 68.350 ;
        RECT 124.090 67.680 127.950 67.850 ;
        RECT 259.310 67.810 263.170 67.980 ;
        RECT 22.770 67.560 26.060 67.570 ;
        RECT 124.080 67.380 127.950 67.680 ;
        RECT 259.300 67.510 263.170 67.810 ;
        RECT 360.620 67.790 363.920 68.160 ;
        RECT 360.620 67.620 364.480 67.790 ;
        RECT 259.300 67.500 262.590 67.510 ;
        RECT 124.080 67.370 127.370 67.380 ;
        RECT 360.610 67.320 364.480 67.620 ;
        RECT 360.610 67.310 363.900 67.320 ;
        RECT 7.260 64.060 10.560 64.430 ;
        RECT 7.260 63.890 10.980 64.060 ;
        RECT 7.250 63.590 10.980 63.890 ;
        RECT 108.570 63.870 111.870 64.240 ;
        RECT 243.790 64.000 247.090 64.370 ;
        RECT 108.570 63.700 112.290 63.870 ;
        RECT 243.790 63.830 247.510 64.000 ;
        RECT 7.250 63.580 10.540 63.590 ;
        RECT 108.560 63.400 112.290 63.700 ;
        RECT 243.780 63.530 247.510 63.830 ;
        RECT 345.100 63.810 348.400 64.180 ;
        RECT 345.100 63.640 348.820 63.810 ;
        RECT 243.780 63.520 247.070 63.530 ;
        RECT 108.560 63.390 111.850 63.400 ;
        RECT 345.090 63.340 348.820 63.640 ;
        RECT 345.090 63.330 348.380 63.340 ;
        RECT 40.360 62.420 43.660 62.860 ;
        RECT 40.360 62.320 44.160 62.420 ;
        RECT 40.350 62.010 44.160 62.320 ;
        RECT 141.670 62.230 144.970 62.670 ;
        RECT 276.890 62.360 280.190 62.800 ;
        RECT 276.890 62.260 280.690 62.360 ;
        RECT 141.670 62.130 145.470 62.230 ;
        RECT 141.660 61.820 145.470 62.130 ;
        RECT 276.880 61.950 280.690 62.260 ;
        RECT 378.200 62.170 381.500 62.610 ;
        RECT 378.200 62.070 382.000 62.170 ;
        RECT 378.190 61.760 382.000 62.070 ;
        RECT 6.930 56.040 10.260 56.410 ;
        RECT 6.930 56.030 10.560 56.040 ;
        RECT 6.930 55.870 10.620 56.030 ;
        RECT 6.920 55.590 10.620 55.870 ;
        RECT 108.240 55.850 111.570 56.220 ;
        RECT 243.460 55.980 246.790 56.350 ;
        RECT 243.460 55.970 247.090 55.980 ;
        RECT 108.240 55.840 111.870 55.850 ;
        RECT 108.240 55.680 111.930 55.840 ;
        RECT 243.460 55.810 247.150 55.970 ;
        RECT 6.920 55.560 10.210 55.590 ;
        RECT 108.230 55.400 111.930 55.680 ;
        RECT 243.450 55.530 247.150 55.810 ;
        RECT 344.770 55.790 348.100 56.160 ;
        RECT 344.770 55.780 348.400 55.790 ;
        RECT 344.770 55.620 348.460 55.780 ;
        RECT 243.450 55.500 246.740 55.530 ;
        RECT 108.230 55.370 111.520 55.400 ;
        RECT 344.760 55.340 348.460 55.620 ;
        RECT 344.760 55.310 348.050 55.340 ;
        RECT 22.610 53.620 25.910 53.990 ;
        RECT 22.610 53.450 26.470 53.620 ;
        RECT 22.600 53.150 26.470 53.450 ;
        RECT 123.920 53.430 127.220 53.800 ;
        RECT 259.140 53.560 262.440 53.930 ;
        RECT 123.920 53.260 127.780 53.430 ;
        RECT 259.140 53.390 263.000 53.560 ;
        RECT 22.600 53.140 25.890 53.150 ;
        RECT 123.910 52.960 127.780 53.260 ;
        RECT 259.130 53.090 263.000 53.390 ;
        RECT 360.450 53.370 363.750 53.740 ;
        RECT 360.450 53.200 364.310 53.370 ;
        RECT 259.130 53.080 262.420 53.090 ;
        RECT 123.910 52.950 127.200 52.960 ;
        RECT 360.440 52.900 364.310 53.200 ;
        RECT 360.440 52.890 363.730 52.900 ;
        RECT 7.090 49.640 10.390 50.010 ;
        RECT 7.090 49.470 10.810 49.640 ;
        RECT 7.080 49.170 10.810 49.470 ;
        RECT 108.400 49.450 111.700 49.820 ;
        RECT 243.620 49.580 246.920 49.950 ;
        RECT 108.400 49.280 112.120 49.450 ;
        RECT 243.620 49.410 247.340 49.580 ;
        RECT 7.080 49.160 10.370 49.170 ;
        RECT 108.390 48.980 112.120 49.280 ;
        RECT 243.610 49.110 247.340 49.410 ;
        RECT 344.930 49.390 348.230 49.760 ;
        RECT 344.930 49.220 348.650 49.390 ;
        RECT 243.610 49.100 246.900 49.110 ;
        RECT 108.390 48.970 111.680 48.980 ;
        RECT 344.920 48.920 348.650 49.220 ;
        RECT 344.920 48.910 348.210 48.920 ;
        RECT 57.890 46.390 61.190 46.840 ;
        RECT 57.890 46.300 61.630 46.390 ;
        RECT 57.880 46.000 61.630 46.300 ;
        RECT 159.200 46.200 162.500 46.650 ;
        RECT 294.420 46.330 297.720 46.780 ;
        RECT 294.420 46.240 298.160 46.330 ;
        RECT 159.200 46.110 162.940 46.200 ;
        RECT 57.880 45.990 61.170 46.000 ;
        RECT 159.190 45.810 162.940 46.110 ;
        RECT 294.410 45.940 298.160 46.240 ;
        RECT 395.730 46.140 399.030 46.590 ;
        RECT 395.730 46.050 399.470 46.140 ;
        RECT 294.410 45.930 297.700 45.940 ;
        RECT 159.190 45.800 162.480 45.810 ;
        RECT 395.720 45.750 399.470 46.050 ;
        RECT 395.720 45.740 399.010 45.750 ;
        RECT 7.070 40.390 10.400 40.760 ;
        RECT 7.070 40.380 10.700 40.390 ;
        RECT 7.070 40.220 10.760 40.380 ;
        RECT 7.060 39.940 10.760 40.220 ;
        RECT 108.380 40.200 111.710 40.570 ;
        RECT 243.600 40.330 246.930 40.700 ;
        RECT 243.600 40.320 247.230 40.330 ;
        RECT 108.380 40.190 112.010 40.200 ;
        RECT 108.380 40.030 112.070 40.190 ;
        RECT 243.600 40.160 247.290 40.320 ;
        RECT 7.060 39.910 10.350 39.940 ;
        RECT 108.370 39.750 112.070 40.030 ;
        RECT 243.590 39.880 247.290 40.160 ;
        RECT 344.910 40.140 348.240 40.510 ;
        RECT 344.910 40.130 348.540 40.140 ;
        RECT 344.910 39.970 348.600 40.130 ;
        RECT 243.590 39.850 246.880 39.880 ;
        RECT 108.370 39.720 111.660 39.750 ;
        RECT 344.900 39.690 348.600 39.970 ;
        RECT 344.900 39.660 348.190 39.690 ;
        RECT 22.750 37.970 26.050 38.340 ;
        RECT 22.750 37.800 26.610 37.970 ;
        RECT 22.740 37.500 26.610 37.800 ;
        RECT 124.060 37.780 127.360 38.150 ;
        RECT 259.280 37.910 262.580 38.280 ;
        RECT 124.060 37.610 127.920 37.780 ;
        RECT 259.280 37.740 263.140 37.910 ;
        RECT 22.740 37.490 26.030 37.500 ;
        RECT 124.050 37.310 127.920 37.610 ;
        RECT 259.270 37.440 263.140 37.740 ;
        RECT 360.590 37.720 363.890 38.090 ;
        RECT 360.590 37.550 364.450 37.720 ;
        RECT 259.270 37.430 262.560 37.440 ;
        RECT 124.050 37.300 127.340 37.310 ;
        RECT 360.580 37.250 364.450 37.550 ;
        RECT 360.580 37.240 363.870 37.250 ;
        RECT 7.230 33.990 10.530 34.360 ;
        RECT 7.230 33.820 10.950 33.990 ;
        RECT 7.220 33.520 10.950 33.820 ;
        RECT 108.540 33.800 111.840 34.170 ;
        RECT 243.760 33.930 247.060 34.300 ;
        RECT 108.540 33.630 112.260 33.800 ;
        RECT 243.760 33.760 247.480 33.930 ;
        RECT 7.220 33.510 10.510 33.520 ;
        RECT 108.530 33.330 112.260 33.630 ;
        RECT 243.750 33.460 247.480 33.760 ;
        RECT 345.070 33.740 348.370 34.110 ;
        RECT 345.070 33.570 348.790 33.740 ;
        RECT 243.750 33.450 247.040 33.460 ;
        RECT 108.530 33.320 111.820 33.330 ;
        RECT 345.060 33.270 348.790 33.570 ;
        RECT 345.060 33.260 348.350 33.270 ;
        RECT 40.330 32.350 43.630 32.790 ;
        RECT 40.330 32.250 44.130 32.350 ;
        RECT 40.320 31.940 44.130 32.250 ;
        RECT 141.640 32.160 144.940 32.600 ;
        RECT 276.860 32.290 280.160 32.730 ;
        RECT 276.860 32.190 280.660 32.290 ;
        RECT 141.640 32.060 145.440 32.160 ;
        RECT 141.630 31.750 145.440 32.060 ;
        RECT 276.850 31.880 280.660 32.190 ;
        RECT 378.170 32.100 381.470 32.540 ;
        RECT 378.170 32.000 381.970 32.100 ;
        RECT 378.160 31.690 381.970 32.000 ;
        RECT 6.900 25.970 10.230 26.340 ;
        RECT 6.900 25.960 10.530 25.970 ;
        RECT 6.900 25.800 10.590 25.960 ;
        RECT 6.890 25.520 10.590 25.800 ;
        RECT 108.210 25.780 111.540 26.150 ;
        RECT 243.430 25.910 246.760 26.280 ;
        RECT 243.430 25.900 247.060 25.910 ;
        RECT 108.210 25.770 111.840 25.780 ;
        RECT 108.210 25.610 111.900 25.770 ;
        RECT 243.430 25.740 247.120 25.900 ;
        RECT 6.890 25.490 10.180 25.520 ;
        RECT 108.200 25.330 111.900 25.610 ;
        RECT 243.420 25.460 247.120 25.740 ;
        RECT 344.740 25.720 348.070 26.090 ;
        RECT 344.740 25.710 348.370 25.720 ;
        RECT 344.740 25.550 348.430 25.710 ;
        RECT 243.420 25.430 246.710 25.460 ;
        RECT 108.200 25.300 111.490 25.330 ;
        RECT 344.730 25.270 348.430 25.550 ;
        RECT 344.730 25.240 348.020 25.270 ;
        RECT 22.580 23.550 25.880 23.920 ;
        RECT 22.580 23.380 26.440 23.550 ;
        RECT 22.570 23.080 26.440 23.380 ;
        RECT 123.890 23.360 127.190 23.730 ;
        RECT 259.110 23.490 262.410 23.860 ;
        RECT 123.890 23.190 127.750 23.360 ;
        RECT 259.110 23.320 262.970 23.490 ;
        RECT 22.570 23.070 25.860 23.080 ;
        RECT 123.880 22.890 127.750 23.190 ;
        RECT 259.100 23.020 262.970 23.320 ;
        RECT 360.420 23.300 363.720 23.670 ;
        RECT 360.420 23.130 364.280 23.300 ;
        RECT 259.100 23.010 262.390 23.020 ;
        RECT 123.880 22.880 127.170 22.890 ;
        RECT 360.410 22.830 364.280 23.130 ;
        RECT 360.410 22.820 363.700 22.830 ;
        RECT 7.060 19.570 10.360 19.940 ;
        RECT 7.060 19.400 10.780 19.570 ;
        RECT 7.050 19.100 10.780 19.400 ;
        RECT 108.370 19.380 111.670 19.750 ;
        RECT 243.590 19.510 246.890 19.880 ;
        RECT 108.370 19.210 112.090 19.380 ;
        RECT 243.590 19.340 247.310 19.510 ;
        RECT 7.050 19.090 10.340 19.100 ;
        RECT 108.360 18.910 112.090 19.210 ;
        RECT 243.580 19.040 247.310 19.340 ;
        RECT 344.900 19.320 348.200 19.690 ;
        RECT 344.900 19.150 348.620 19.320 ;
        RECT 243.580 19.030 246.870 19.040 ;
        RECT 108.360 18.900 111.650 18.910 ;
        RECT 344.890 18.850 348.620 19.150 ;
        RECT 344.890 18.840 348.180 18.850 ;
      LAYER via ;
        RECT 11.320 250.260 11.580 250.520 ;
        RECT 112.630 250.070 112.890 250.330 ;
        RECT 247.850 250.200 248.110 250.460 ;
        RECT 349.160 250.010 349.420 250.270 ;
        RECT 27.115 247.830 27.375 248.090 ;
        RECT 128.425 247.640 128.685 247.900 ;
        RECT 263.645 247.770 263.905 248.030 ;
        RECT 364.955 247.580 365.215 247.840 ;
        RECT 11.495 243.845 11.755 244.105 ;
        RECT 112.805 243.655 113.065 243.915 ;
        RECT 248.025 243.785 248.285 244.045 ;
        RECT 349.335 243.595 349.595 243.855 ;
        RECT 44.645 242.230 44.905 242.490 ;
        RECT 145.955 242.040 146.215 242.300 ;
        RECT 281.175 242.170 281.435 242.430 ;
        RECT 382.485 241.980 382.745 242.240 ;
        RECT 11.150 235.840 11.410 236.100 ;
        RECT 112.460 235.650 112.720 235.910 ;
        RECT 247.680 235.780 247.940 236.040 ;
        RECT 348.990 235.590 349.250 235.850 ;
        RECT 26.945 233.410 27.205 233.670 ;
        RECT 128.255 233.220 128.515 233.480 ;
        RECT 263.475 233.350 263.735 233.610 ;
        RECT 364.785 233.160 365.045 233.420 ;
        RECT 11.325 229.425 11.585 229.685 ;
        RECT 112.635 229.235 112.895 229.495 ;
        RECT 247.855 229.365 248.115 229.625 ;
        RECT 349.165 229.175 349.425 229.435 ;
        RECT 62.145 226.215 62.405 226.475 ;
        RECT 163.455 226.025 163.715 226.285 ;
        RECT 298.675 226.155 298.935 226.415 ;
        RECT 399.985 225.965 400.245 226.225 ;
        RECT 11.290 220.190 11.550 220.450 ;
        RECT 112.600 220.000 112.860 220.260 ;
        RECT 247.820 220.130 248.080 220.390 ;
        RECT 349.130 219.940 349.390 220.200 ;
        RECT 27.085 217.760 27.345 218.020 ;
        RECT 128.395 217.570 128.655 217.830 ;
        RECT 263.615 217.700 263.875 217.960 ;
        RECT 364.925 217.510 365.185 217.770 ;
        RECT 11.465 213.775 11.725 214.035 ;
        RECT 112.775 213.585 113.035 213.845 ;
        RECT 247.995 213.715 248.255 213.975 ;
        RECT 349.305 213.525 349.565 213.785 ;
        RECT 44.615 212.160 44.875 212.420 ;
        RECT 145.925 211.970 146.185 212.230 ;
        RECT 281.145 212.100 281.405 212.360 ;
        RECT 382.455 211.910 382.715 212.170 ;
        RECT 11.120 205.770 11.380 206.030 ;
        RECT 112.430 205.580 112.690 205.840 ;
        RECT 247.650 205.710 247.910 205.970 ;
        RECT 348.960 205.520 349.220 205.780 ;
        RECT 26.915 203.340 27.175 203.600 ;
        RECT 128.225 203.150 128.485 203.410 ;
        RECT 263.445 203.280 263.705 203.540 ;
        RECT 364.755 203.090 365.015 203.350 ;
        RECT 76.445 199.970 76.705 200.230 ;
        RECT 11.295 199.355 11.555 199.615 ;
        RECT 177.755 199.780 178.015 200.040 ;
        RECT 312.975 199.910 313.235 200.170 ;
        RECT 112.605 199.165 112.865 199.425 ;
        RECT 247.825 199.295 248.085 199.555 ;
        RECT 414.285 199.720 414.545 199.980 ;
        RECT 349.135 199.105 349.395 199.365 ;
        RECT 10.970 190.340 11.230 190.600 ;
        RECT 112.280 190.150 112.540 190.410 ;
        RECT 247.500 190.280 247.760 190.540 ;
        RECT 348.810 190.090 349.070 190.350 ;
        RECT 26.765 187.910 27.025 188.170 ;
        RECT 128.075 187.720 128.335 187.980 ;
        RECT 263.295 187.850 263.555 188.110 ;
        RECT 364.605 187.660 364.865 187.920 ;
        RECT 11.145 183.925 11.405 184.185 ;
        RECT 112.455 183.735 112.715 183.995 ;
        RECT 247.675 183.865 247.935 184.125 ;
        RECT 348.985 183.675 349.245 183.935 ;
        RECT 44.295 182.310 44.555 182.570 ;
        RECT 145.605 182.120 145.865 182.380 ;
        RECT 280.825 182.250 281.085 182.510 ;
        RECT 382.135 182.060 382.395 182.320 ;
        RECT 10.800 175.920 11.060 176.180 ;
        RECT 112.110 175.730 112.370 175.990 ;
        RECT 247.330 175.860 247.590 176.120 ;
        RECT 348.640 175.670 348.900 175.930 ;
        RECT 26.595 173.490 26.855 173.750 ;
        RECT 127.905 173.300 128.165 173.560 ;
        RECT 263.125 173.430 263.385 173.690 ;
        RECT 364.435 173.240 364.695 173.500 ;
        RECT 10.975 169.505 11.235 169.765 ;
        RECT 112.285 169.315 112.545 169.575 ;
        RECT 247.505 169.445 247.765 169.705 ;
        RECT 348.815 169.255 349.075 169.515 ;
        RECT 61.795 166.295 62.055 166.555 ;
        RECT 163.105 166.105 163.365 166.365 ;
        RECT 298.325 166.235 298.585 166.495 ;
        RECT 399.635 166.045 399.895 166.305 ;
        RECT 10.940 160.270 11.200 160.530 ;
        RECT 112.250 160.080 112.510 160.340 ;
        RECT 247.470 160.210 247.730 160.470 ;
        RECT 348.780 160.020 349.040 160.280 ;
        RECT 26.735 157.840 26.995 158.100 ;
        RECT 128.045 157.650 128.305 157.910 ;
        RECT 263.265 157.780 263.525 158.040 ;
        RECT 364.575 157.590 364.835 157.850 ;
        RECT 11.115 153.855 11.375 154.115 ;
        RECT 112.425 153.665 112.685 153.925 ;
        RECT 247.645 153.795 247.905 154.055 ;
        RECT 348.955 153.605 349.215 153.865 ;
        RECT 44.265 152.240 44.525 152.500 ;
        RECT 145.575 152.050 145.835 152.310 ;
        RECT 280.795 152.180 281.055 152.440 ;
        RECT 382.105 151.990 382.365 152.250 ;
        RECT 10.770 145.850 11.030 146.110 ;
        RECT 112.080 145.660 112.340 145.920 ;
        RECT 247.300 145.790 247.560 146.050 ;
        RECT 348.610 145.600 348.870 145.860 ;
        RECT 26.565 143.420 26.825 143.680 ;
        RECT 127.875 143.230 128.135 143.490 ;
        RECT 263.095 143.360 263.355 143.620 ;
        RECT 364.405 143.170 364.665 143.430 ;
        RECT 10.945 139.435 11.205 139.695 ;
        RECT 112.255 139.245 112.515 139.505 ;
        RECT 247.475 139.375 247.735 139.635 ;
        RECT 220.315 138.910 220.575 139.170 ;
        RECT 348.785 139.185 349.045 139.445 ;
        RECT 456.845 138.850 457.105 139.110 ;
        RECT 92.690 136.805 92.950 137.065 ;
        RECT 194.000 136.615 194.260 136.875 ;
        RECT 329.220 136.745 329.480 137.005 ;
        RECT 430.530 136.555 430.790 136.815 ;
        RECT 474.125 136.510 474.385 136.770 ;
        RECT 10.820 130.020 11.080 130.280 ;
        RECT 112.130 129.830 112.390 130.090 ;
        RECT 247.350 129.960 247.610 130.220 ;
        RECT 348.660 129.770 348.920 130.030 ;
        RECT 26.615 127.590 26.875 127.850 ;
        RECT 127.925 127.400 128.185 127.660 ;
        RECT 263.145 127.530 263.405 127.790 ;
        RECT 364.455 127.340 364.715 127.600 ;
        RECT 10.995 123.605 11.255 123.865 ;
        RECT 112.305 123.415 112.565 123.675 ;
        RECT 247.525 123.545 247.785 123.805 ;
        RECT 348.835 123.355 349.095 123.615 ;
        RECT 44.145 121.990 44.405 122.250 ;
        RECT 145.455 121.800 145.715 122.060 ;
        RECT 280.675 121.930 280.935 122.190 ;
        RECT 381.985 121.740 382.245 122.000 ;
        RECT 10.650 115.600 10.910 115.860 ;
        RECT 111.960 115.410 112.220 115.670 ;
        RECT 247.180 115.540 247.440 115.800 ;
        RECT 348.490 115.350 348.750 115.610 ;
        RECT 26.445 113.170 26.705 113.430 ;
        RECT 127.755 112.980 128.015 113.240 ;
        RECT 262.975 113.110 263.235 113.370 ;
        RECT 364.285 112.920 364.545 113.180 ;
        RECT 10.825 109.185 11.085 109.445 ;
        RECT 112.135 108.995 112.395 109.255 ;
        RECT 247.355 109.125 247.615 109.385 ;
        RECT 348.665 108.935 348.925 109.195 ;
        RECT 61.645 105.975 61.905 106.235 ;
        RECT 162.955 105.785 163.215 106.045 ;
        RECT 298.175 105.915 298.435 106.175 ;
        RECT 399.485 105.725 399.745 105.985 ;
        RECT 10.790 99.950 11.050 100.210 ;
        RECT 112.100 99.760 112.360 100.020 ;
        RECT 247.320 99.890 247.580 100.150 ;
        RECT 348.630 99.700 348.890 99.960 ;
        RECT 26.585 97.520 26.845 97.780 ;
        RECT 127.895 97.330 128.155 97.590 ;
        RECT 263.115 97.460 263.375 97.720 ;
        RECT 364.425 97.270 364.685 97.530 ;
        RECT 10.965 93.535 11.225 93.795 ;
        RECT 112.275 93.345 112.535 93.605 ;
        RECT 247.495 93.475 247.755 93.735 ;
        RECT 348.805 93.285 349.065 93.545 ;
        RECT 44.115 91.920 44.375 92.180 ;
        RECT 145.425 91.730 145.685 91.990 ;
        RECT 280.645 91.860 280.905 92.120 ;
        RECT 381.955 91.670 382.215 91.930 ;
        RECT 10.620 85.530 10.880 85.790 ;
        RECT 111.930 85.340 112.190 85.600 ;
        RECT 247.150 85.470 247.410 85.730 ;
        RECT 348.460 85.280 348.720 85.540 ;
        RECT 26.415 83.100 26.675 83.360 ;
        RECT 127.725 82.910 127.985 83.170 ;
        RECT 262.945 83.040 263.205 83.300 ;
        RECT 364.255 82.850 364.515 83.110 ;
        RECT 75.945 79.730 76.205 79.990 ;
        RECT 10.795 79.115 11.055 79.375 ;
        RECT 177.255 79.540 177.515 79.800 ;
        RECT 312.475 79.670 312.735 79.930 ;
        RECT 112.105 78.925 112.365 79.185 ;
        RECT 247.325 79.055 247.585 79.315 ;
        RECT 413.785 79.480 414.045 79.740 ;
        RECT 348.635 78.865 348.895 79.125 ;
        RECT 10.470 70.100 10.730 70.360 ;
        RECT 111.780 69.910 112.040 70.170 ;
        RECT 247.000 70.040 247.260 70.300 ;
        RECT 348.310 69.850 348.570 70.110 ;
        RECT 26.265 67.670 26.525 67.930 ;
        RECT 127.575 67.480 127.835 67.740 ;
        RECT 262.795 67.610 263.055 67.870 ;
        RECT 364.105 67.420 364.365 67.680 ;
        RECT 10.645 63.685 10.905 63.945 ;
        RECT 111.955 63.495 112.215 63.755 ;
        RECT 247.175 63.625 247.435 63.885 ;
        RECT 348.485 63.435 348.745 63.695 ;
        RECT 43.795 62.070 44.055 62.330 ;
        RECT 145.105 61.880 145.365 62.140 ;
        RECT 280.325 62.010 280.585 62.270 ;
        RECT 381.635 61.820 381.895 62.080 ;
        RECT 10.300 55.680 10.560 55.940 ;
        RECT 111.610 55.490 111.870 55.750 ;
        RECT 246.830 55.620 247.090 55.880 ;
        RECT 348.140 55.430 348.400 55.690 ;
        RECT 26.095 53.250 26.355 53.510 ;
        RECT 127.405 53.060 127.665 53.320 ;
        RECT 262.625 53.190 262.885 53.450 ;
        RECT 363.935 53.000 364.195 53.260 ;
        RECT 10.475 49.265 10.735 49.525 ;
        RECT 111.785 49.075 112.045 49.335 ;
        RECT 247.005 49.205 247.265 49.465 ;
        RECT 348.315 49.015 348.575 49.275 ;
        RECT 61.295 46.055 61.555 46.315 ;
        RECT 162.605 45.865 162.865 46.125 ;
        RECT 297.825 45.995 298.085 46.255 ;
        RECT 399.135 45.805 399.395 46.065 ;
        RECT 10.440 40.030 10.700 40.290 ;
        RECT 111.750 39.840 112.010 40.100 ;
        RECT 246.970 39.970 247.230 40.230 ;
        RECT 348.280 39.780 348.540 40.040 ;
        RECT 26.235 37.600 26.495 37.860 ;
        RECT 127.545 37.410 127.805 37.670 ;
        RECT 262.765 37.540 263.025 37.800 ;
        RECT 364.075 37.350 364.335 37.610 ;
        RECT 10.615 33.615 10.875 33.875 ;
        RECT 111.925 33.425 112.185 33.685 ;
        RECT 247.145 33.555 247.405 33.815 ;
        RECT 348.455 33.365 348.715 33.625 ;
        RECT 43.765 32.000 44.025 32.260 ;
        RECT 145.075 31.810 145.335 32.070 ;
        RECT 280.295 31.940 280.555 32.200 ;
        RECT 381.605 31.750 381.865 32.010 ;
        RECT 10.270 25.610 10.530 25.870 ;
        RECT 111.580 25.420 111.840 25.680 ;
        RECT 246.800 25.550 247.060 25.810 ;
        RECT 348.110 25.360 348.370 25.620 ;
        RECT 26.065 23.180 26.325 23.440 ;
        RECT 127.375 22.990 127.635 23.250 ;
        RECT 262.595 23.120 262.855 23.380 ;
        RECT 363.905 22.930 364.165 23.190 ;
        RECT 10.445 19.195 10.705 19.455 ;
        RECT 111.755 19.005 112.015 19.265 ;
        RECT 246.975 19.135 247.235 19.395 ;
        RECT 348.285 18.945 348.545 19.205 ;
      LAYER met2 ;
        RECT 11.280 250.640 11.700 251.160 ;
        RECT 11.280 250.160 11.640 250.640 ;
        RECT 112.590 250.450 113.010 250.970 ;
        RECT 247.810 250.580 248.230 251.100 ;
        RECT 112.590 249.970 112.950 250.450 ;
        RECT 247.810 250.100 248.170 250.580 ;
        RECT 349.120 250.390 349.540 250.910 ;
        RECT 349.120 249.910 349.480 250.390 ;
        RECT 27.000 247.730 27.500 248.750 ;
        RECT 128.310 247.540 128.810 248.560 ;
        RECT 263.530 247.670 264.030 248.690 ;
        RECT 364.840 247.480 365.340 248.500 ;
        RECT 11.450 243.750 11.830 244.660 ;
        RECT 112.760 243.560 113.140 244.470 ;
        RECT 247.980 243.690 248.360 244.600 ;
        RECT 349.290 243.500 349.670 244.410 ;
        RECT 44.570 242.170 45.020 243.030 ;
        RECT 145.880 241.980 146.330 242.840 ;
        RECT 281.100 242.110 281.550 242.970 ;
        RECT 382.410 241.920 382.860 242.780 ;
        RECT 11.110 236.220 11.530 236.740 ;
        RECT 11.110 235.740 11.470 236.220 ;
        RECT 112.420 236.030 112.840 236.550 ;
        RECT 247.640 236.160 248.060 236.680 ;
        RECT 112.420 235.550 112.780 236.030 ;
        RECT 247.640 235.680 248.000 236.160 ;
        RECT 348.950 235.970 349.370 236.490 ;
        RECT 348.950 235.490 349.310 235.970 ;
        RECT 26.830 233.310 27.330 234.330 ;
        RECT 128.140 233.120 128.640 234.140 ;
        RECT 263.360 233.250 263.860 234.270 ;
        RECT 364.670 233.060 365.170 234.080 ;
        RECT 11.280 229.330 11.660 230.240 ;
        RECT 112.590 229.140 112.970 230.050 ;
        RECT 247.810 229.270 248.190 230.180 ;
        RECT 349.120 229.080 349.500 229.990 ;
        RECT 62.090 226.170 62.470 227.030 ;
        RECT 163.400 225.980 163.780 226.840 ;
        RECT 298.620 226.110 299.000 226.970 ;
        RECT 399.930 225.920 400.310 226.780 ;
        RECT 11.250 220.570 11.670 221.090 ;
        RECT 11.250 220.090 11.610 220.570 ;
        RECT 112.560 220.380 112.980 220.900 ;
        RECT 247.780 220.510 248.200 221.030 ;
        RECT 112.560 219.900 112.920 220.380 ;
        RECT 247.780 220.030 248.140 220.510 ;
        RECT 349.090 220.320 349.510 220.840 ;
        RECT 349.090 219.840 349.450 220.320 ;
        RECT 26.970 217.660 27.470 218.680 ;
        RECT 128.280 217.470 128.780 218.490 ;
        RECT 263.500 217.600 264.000 218.620 ;
        RECT 364.810 217.410 365.310 218.430 ;
        RECT 11.420 213.680 11.800 214.590 ;
        RECT 112.730 213.490 113.110 214.400 ;
        RECT 247.950 213.620 248.330 214.530 ;
        RECT 349.260 213.430 349.640 214.340 ;
        RECT 44.540 212.100 44.990 212.960 ;
        RECT 145.850 211.910 146.300 212.770 ;
        RECT 281.070 212.040 281.520 212.900 ;
        RECT 382.380 211.850 382.830 212.710 ;
        RECT 11.080 206.150 11.500 206.670 ;
        RECT 11.080 205.670 11.440 206.150 ;
        RECT 112.390 205.960 112.810 206.480 ;
        RECT 247.610 206.090 248.030 206.610 ;
        RECT 112.390 205.480 112.750 205.960 ;
        RECT 247.610 205.610 247.970 206.090 ;
        RECT 348.920 205.900 349.340 206.420 ;
        RECT 348.920 205.420 349.280 205.900 ;
        RECT 26.800 203.240 27.300 204.260 ;
        RECT 128.110 203.050 128.610 204.070 ;
        RECT 263.330 203.180 263.830 204.200 ;
        RECT 364.640 202.990 365.140 204.010 ;
        RECT 76.330 200.850 76.830 200.930 ;
        RECT 76.320 200.370 76.830 200.850 ;
        RECT 312.860 200.790 313.360 200.870 ;
        RECT 177.640 200.660 178.140 200.740 ;
        RECT 11.250 199.260 11.630 200.170 ;
        RECT 76.320 199.890 76.820 200.370 ;
        RECT 177.630 200.180 178.140 200.660 ;
        RECT 312.850 200.310 313.360 200.790 ;
        RECT 414.170 200.600 414.670 200.680 ;
        RECT 112.560 199.070 112.940 199.980 ;
        RECT 177.630 199.700 178.130 200.180 ;
        RECT 247.780 199.200 248.160 200.110 ;
        RECT 312.850 199.830 313.350 200.310 ;
        RECT 414.160 200.120 414.670 200.600 ;
        RECT 349.090 199.010 349.470 199.920 ;
        RECT 414.160 199.640 414.660 200.120 ;
        RECT 10.930 190.720 11.350 191.240 ;
        RECT 10.930 190.240 11.290 190.720 ;
        RECT 112.240 190.530 112.660 191.050 ;
        RECT 247.460 190.660 247.880 191.180 ;
        RECT 112.240 190.050 112.600 190.530 ;
        RECT 247.460 190.180 247.820 190.660 ;
        RECT 348.770 190.470 349.190 190.990 ;
        RECT 348.770 189.990 349.130 190.470 ;
        RECT 26.650 187.810 27.150 188.830 ;
        RECT 127.960 187.620 128.460 188.640 ;
        RECT 263.180 187.750 263.680 188.770 ;
        RECT 364.490 187.560 364.990 188.580 ;
        RECT 11.100 183.830 11.480 184.740 ;
        RECT 112.410 183.640 112.790 184.550 ;
        RECT 247.630 183.770 248.010 184.680 ;
        RECT 348.940 183.580 349.320 184.490 ;
        RECT 44.220 182.250 44.670 183.110 ;
        RECT 145.530 182.060 145.980 182.920 ;
        RECT 280.750 182.190 281.200 183.050 ;
        RECT 382.060 182.000 382.510 182.860 ;
        RECT 10.760 176.300 11.180 176.820 ;
        RECT 10.760 175.820 11.120 176.300 ;
        RECT 112.070 176.110 112.490 176.630 ;
        RECT 247.290 176.240 247.710 176.760 ;
        RECT 112.070 175.630 112.430 176.110 ;
        RECT 247.290 175.760 247.650 176.240 ;
        RECT 348.600 176.050 349.020 176.570 ;
        RECT 348.600 175.570 348.960 176.050 ;
        RECT 26.480 173.390 26.980 174.410 ;
        RECT 127.790 173.200 128.290 174.220 ;
        RECT 263.010 173.330 263.510 174.350 ;
        RECT 364.320 173.140 364.820 174.160 ;
        RECT 10.930 169.410 11.310 170.320 ;
        RECT 112.240 169.220 112.620 170.130 ;
        RECT 247.460 169.350 247.840 170.260 ;
        RECT 348.770 169.160 349.150 170.070 ;
        RECT 61.740 166.250 62.120 167.110 ;
        RECT 163.050 166.060 163.430 166.920 ;
        RECT 298.270 166.190 298.650 167.050 ;
        RECT 399.580 166.000 399.960 166.860 ;
        RECT 10.900 160.650 11.320 161.170 ;
        RECT 10.900 160.170 11.260 160.650 ;
        RECT 112.210 160.460 112.630 160.980 ;
        RECT 247.430 160.590 247.850 161.110 ;
        RECT 112.210 159.980 112.570 160.460 ;
        RECT 247.430 160.110 247.790 160.590 ;
        RECT 348.740 160.400 349.160 160.920 ;
        RECT 348.740 159.920 349.100 160.400 ;
        RECT 26.620 157.740 27.120 158.760 ;
        RECT 127.930 157.550 128.430 158.570 ;
        RECT 263.150 157.680 263.650 158.700 ;
        RECT 364.460 157.490 364.960 158.510 ;
        RECT 11.070 153.760 11.450 154.670 ;
        RECT 112.380 153.570 112.760 154.480 ;
        RECT 247.600 153.700 247.980 154.610 ;
        RECT 348.910 153.510 349.290 154.420 ;
        RECT 44.190 152.180 44.640 153.040 ;
        RECT 145.500 151.990 145.950 152.850 ;
        RECT 280.720 152.120 281.170 152.980 ;
        RECT 382.030 151.930 382.480 152.790 ;
        RECT 10.730 146.230 11.150 146.750 ;
        RECT 10.730 145.750 11.090 146.230 ;
        RECT 112.040 146.040 112.460 146.560 ;
        RECT 247.260 146.170 247.680 146.690 ;
        RECT 112.040 145.560 112.400 146.040 ;
        RECT 247.260 145.690 247.620 146.170 ;
        RECT 348.570 145.980 348.990 146.500 ;
        RECT 348.570 145.500 348.930 145.980 ;
        RECT 26.450 143.320 26.950 144.340 ;
        RECT 127.760 143.130 128.260 144.150 ;
        RECT 262.980 143.260 263.480 144.280 ;
        RECT 364.290 143.070 364.790 144.090 ;
        RECT 10.900 139.340 11.280 140.250 ;
        RECT 112.210 139.150 112.590 140.060 ;
        RECT 220.220 138.860 220.690 139.690 ;
        RECT 247.430 139.280 247.810 140.190 ;
        RECT 348.740 139.090 349.120 140.000 ;
        RECT 456.750 138.800 457.220 139.630 ;
        RECT 92.620 137.440 93.080 137.630 ;
        RECT 92.630 136.730 93.080 137.440 ;
        RECT 193.930 137.250 194.390 137.440 ;
        RECT 329.150 137.380 329.610 137.570 ;
        RECT 193.940 136.540 194.390 137.250 ;
        RECT 329.160 136.670 329.610 137.380 ;
        RECT 430.460 137.190 430.920 137.380 ;
        RECT 430.470 136.480 430.920 137.190 ;
        RECT 474.050 136.460 474.400 137.230 ;
        RECT 10.780 130.400 11.200 130.920 ;
        RECT 10.780 129.920 11.140 130.400 ;
        RECT 112.090 130.210 112.510 130.730 ;
        RECT 247.310 130.340 247.730 130.860 ;
        RECT 112.090 129.730 112.450 130.210 ;
        RECT 247.310 129.860 247.670 130.340 ;
        RECT 348.620 130.150 349.040 130.670 ;
        RECT 348.620 129.670 348.980 130.150 ;
        RECT 26.500 127.490 27.000 128.510 ;
        RECT 127.810 127.300 128.310 128.320 ;
        RECT 263.030 127.430 263.530 128.450 ;
        RECT 364.340 127.240 364.840 128.260 ;
        RECT 10.950 123.510 11.330 124.420 ;
        RECT 112.260 123.320 112.640 124.230 ;
        RECT 247.480 123.450 247.860 124.360 ;
        RECT 348.790 123.260 349.170 124.170 ;
        RECT 44.070 121.930 44.520 122.790 ;
        RECT 145.380 121.740 145.830 122.600 ;
        RECT 280.600 121.870 281.050 122.730 ;
        RECT 381.910 121.680 382.360 122.540 ;
        RECT 10.610 115.980 11.030 116.500 ;
        RECT 10.610 115.500 10.970 115.980 ;
        RECT 111.920 115.790 112.340 116.310 ;
        RECT 247.140 115.920 247.560 116.440 ;
        RECT 111.920 115.310 112.280 115.790 ;
        RECT 247.140 115.440 247.500 115.920 ;
        RECT 348.450 115.730 348.870 116.250 ;
        RECT 348.450 115.250 348.810 115.730 ;
        RECT 26.330 113.070 26.830 114.090 ;
        RECT 127.640 112.880 128.140 113.900 ;
        RECT 262.860 113.010 263.360 114.030 ;
        RECT 364.170 112.820 364.670 113.840 ;
        RECT 10.780 109.090 11.160 110.000 ;
        RECT 112.090 108.900 112.470 109.810 ;
        RECT 247.310 109.030 247.690 109.940 ;
        RECT 348.620 108.840 349.000 109.750 ;
        RECT 61.590 105.930 61.970 106.790 ;
        RECT 162.900 105.740 163.280 106.600 ;
        RECT 298.120 105.870 298.500 106.730 ;
        RECT 399.430 105.680 399.810 106.540 ;
        RECT 10.750 100.330 11.170 100.850 ;
        RECT 10.750 99.850 11.110 100.330 ;
        RECT 112.060 100.140 112.480 100.660 ;
        RECT 247.280 100.270 247.700 100.790 ;
        RECT 112.060 99.660 112.420 100.140 ;
        RECT 247.280 99.790 247.640 100.270 ;
        RECT 348.590 100.080 349.010 100.600 ;
        RECT 348.590 99.600 348.950 100.080 ;
        RECT 26.470 97.420 26.970 98.440 ;
        RECT 127.780 97.230 128.280 98.250 ;
        RECT 263.000 97.360 263.500 98.380 ;
        RECT 364.310 97.170 364.810 98.190 ;
        RECT 10.920 93.440 11.300 94.350 ;
        RECT 112.230 93.250 112.610 94.160 ;
        RECT 247.450 93.380 247.830 94.290 ;
        RECT 348.760 93.190 349.140 94.100 ;
        RECT 44.040 91.860 44.490 92.720 ;
        RECT 145.350 91.670 145.800 92.530 ;
        RECT 280.570 91.800 281.020 92.660 ;
        RECT 381.880 91.610 382.330 92.470 ;
        RECT 10.580 85.910 11.000 86.430 ;
        RECT 10.580 85.430 10.940 85.910 ;
        RECT 111.890 85.720 112.310 86.240 ;
        RECT 247.110 85.850 247.530 86.370 ;
        RECT 111.890 85.240 112.250 85.720 ;
        RECT 247.110 85.370 247.470 85.850 ;
        RECT 348.420 85.660 348.840 86.180 ;
        RECT 348.420 85.180 348.780 85.660 ;
        RECT 26.300 83.000 26.800 84.020 ;
        RECT 127.610 82.810 128.110 83.830 ;
        RECT 262.830 82.940 263.330 83.960 ;
        RECT 364.140 82.750 364.640 83.770 ;
        RECT 75.830 80.610 76.330 80.690 ;
        RECT 75.820 80.130 76.330 80.610 ;
        RECT 312.360 80.550 312.860 80.630 ;
        RECT 177.140 80.420 177.640 80.500 ;
        RECT 10.750 79.020 11.130 79.930 ;
        RECT 75.820 79.650 76.320 80.130 ;
        RECT 177.130 79.940 177.640 80.420 ;
        RECT 312.350 80.070 312.860 80.550 ;
        RECT 413.670 80.360 414.170 80.440 ;
        RECT 112.060 78.830 112.440 79.740 ;
        RECT 177.130 79.460 177.630 79.940 ;
        RECT 247.280 78.960 247.660 79.870 ;
        RECT 312.350 79.590 312.850 80.070 ;
        RECT 413.660 79.880 414.170 80.360 ;
        RECT 348.590 78.770 348.970 79.680 ;
        RECT 413.660 79.400 414.160 79.880 ;
        RECT 10.430 70.480 10.850 71.000 ;
        RECT 10.430 70.000 10.790 70.480 ;
        RECT 111.740 70.290 112.160 70.810 ;
        RECT 246.960 70.420 247.380 70.940 ;
        RECT 111.740 69.810 112.100 70.290 ;
        RECT 246.960 69.940 247.320 70.420 ;
        RECT 348.270 70.230 348.690 70.750 ;
        RECT 348.270 69.750 348.630 70.230 ;
        RECT 26.150 67.570 26.650 68.590 ;
        RECT 127.460 67.380 127.960 68.400 ;
        RECT 262.680 67.510 263.180 68.530 ;
        RECT 363.990 67.320 364.490 68.340 ;
        RECT 10.600 63.590 10.980 64.500 ;
        RECT 111.910 63.400 112.290 64.310 ;
        RECT 247.130 63.530 247.510 64.440 ;
        RECT 348.440 63.340 348.820 64.250 ;
        RECT 43.720 62.010 44.170 62.870 ;
        RECT 145.030 61.820 145.480 62.680 ;
        RECT 280.250 61.950 280.700 62.810 ;
        RECT 381.560 61.760 382.010 62.620 ;
        RECT 10.260 56.060 10.680 56.580 ;
        RECT 10.260 55.580 10.620 56.060 ;
        RECT 111.570 55.870 111.990 56.390 ;
        RECT 246.790 56.000 247.210 56.520 ;
        RECT 111.570 55.390 111.930 55.870 ;
        RECT 246.790 55.520 247.150 56.000 ;
        RECT 348.100 55.810 348.520 56.330 ;
        RECT 348.100 55.330 348.460 55.810 ;
        RECT 25.980 53.150 26.480 54.170 ;
        RECT 127.290 52.960 127.790 53.980 ;
        RECT 262.510 53.090 263.010 54.110 ;
        RECT 363.820 52.900 364.320 53.920 ;
        RECT 10.430 49.170 10.810 50.080 ;
        RECT 111.740 48.980 112.120 49.890 ;
        RECT 246.960 49.110 247.340 50.020 ;
        RECT 348.270 48.920 348.650 49.830 ;
        RECT 61.240 46.010 61.620 46.870 ;
        RECT 162.550 45.820 162.930 46.680 ;
        RECT 297.770 45.950 298.150 46.810 ;
        RECT 399.080 45.760 399.460 46.620 ;
        RECT 10.400 40.410 10.820 40.930 ;
        RECT 10.400 39.930 10.760 40.410 ;
        RECT 111.710 40.220 112.130 40.740 ;
        RECT 246.930 40.350 247.350 40.870 ;
        RECT 111.710 39.740 112.070 40.220 ;
        RECT 246.930 39.870 247.290 40.350 ;
        RECT 348.240 40.160 348.660 40.680 ;
        RECT 348.240 39.680 348.600 40.160 ;
        RECT 26.120 37.500 26.620 38.520 ;
        RECT 127.430 37.310 127.930 38.330 ;
        RECT 262.650 37.440 263.150 38.460 ;
        RECT 363.960 37.250 364.460 38.270 ;
        RECT 10.570 33.520 10.950 34.430 ;
        RECT 111.880 33.330 112.260 34.240 ;
        RECT 247.100 33.460 247.480 34.370 ;
        RECT 348.410 33.270 348.790 34.180 ;
        RECT 43.690 31.940 44.140 32.800 ;
        RECT 145.000 31.750 145.450 32.610 ;
        RECT 280.220 31.880 280.670 32.740 ;
        RECT 381.530 31.690 381.980 32.550 ;
        RECT 10.230 25.990 10.650 26.510 ;
        RECT 10.230 25.510 10.590 25.990 ;
        RECT 111.540 25.800 111.960 26.320 ;
        RECT 246.760 25.930 247.180 26.450 ;
        RECT 111.540 25.320 111.900 25.800 ;
        RECT 246.760 25.450 247.120 25.930 ;
        RECT 348.070 25.740 348.490 26.260 ;
        RECT 348.070 25.260 348.430 25.740 ;
        RECT 25.950 23.080 26.450 24.100 ;
        RECT 127.260 22.890 127.760 23.910 ;
        RECT 262.480 23.020 262.980 24.040 ;
        RECT 363.790 22.830 364.290 23.850 ;
        RECT 10.400 19.100 10.780 20.010 ;
        RECT 111.710 18.910 112.090 19.820 ;
        RECT 246.930 19.040 247.310 19.950 ;
        RECT 348.240 18.850 348.620 19.760 ;
      LAYER via2 ;
        RECT 11.345 250.720 11.625 251.000 ;
        RECT 112.655 250.530 112.935 250.810 ;
        RECT 247.875 250.660 248.155 250.940 ;
        RECT 349.185 250.470 349.465 250.750 ;
        RECT 27.110 248.315 27.390 248.595 ;
        RECT 128.420 248.125 128.700 248.405 ;
        RECT 263.640 248.255 263.920 248.535 ;
        RECT 364.950 248.065 365.230 248.345 ;
        RECT 11.495 244.295 11.775 244.575 ;
        RECT 112.805 244.105 113.085 244.385 ;
        RECT 248.025 244.235 248.305 244.515 ;
        RECT 349.335 244.045 349.615 244.325 ;
        RECT 44.645 242.655 44.925 242.935 ;
        RECT 145.955 242.465 146.235 242.745 ;
        RECT 281.175 242.595 281.455 242.875 ;
        RECT 382.485 242.405 382.765 242.685 ;
        RECT 11.175 236.300 11.455 236.580 ;
        RECT 112.485 236.110 112.765 236.390 ;
        RECT 247.705 236.240 247.985 236.520 ;
        RECT 349.015 236.050 349.295 236.330 ;
        RECT 26.940 233.895 27.220 234.175 ;
        RECT 128.250 233.705 128.530 233.985 ;
        RECT 263.470 233.835 263.750 234.115 ;
        RECT 364.780 233.645 365.060 233.925 ;
        RECT 11.325 229.875 11.605 230.155 ;
        RECT 112.635 229.685 112.915 229.965 ;
        RECT 247.855 229.815 248.135 230.095 ;
        RECT 349.165 229.625 349.445 229.905 ;
        RECT 62.150 226.675 62.430 226.955 ;
        RECT 163.460 226.485 163.740 226.765 ;
        RECT 298.680 226.615 298.960 226.895 ;
        RECT 399.990 226.425 400.270 226.705 ;
        RECT 11.315 220.650 11.595 220.930 ;
        RECT 112.625 220.460 112.905 220.740 ;
        RECT 247.845 220.590 248.125 220.870 ;
        RECT 349.155 220.400 349.435 220.680 ;
        RECT 27.080 218.245 27.360 218.525 ;
        RECT 128.390 218.055 128.670 218.335 ;
        RECT 263.610 218.185 263.890 218.465 ;
        RECT 364.920 217.995 365.200 218.275 ;
        RECT 11.465 214.225 11.745 214.505 ;
        RECT 112.775 214.035 113.055 214.315 ;
        RECT 247.995 214.165 248.275 214.445 ;
        RECT 349.305 213.975 349.585 214.255 ;
        RECT 44.615 212.585 44.895 212.865 ;
        RECT 145.925 212.395 146.205 212.675 ;
        RECT 281.145 212.525 281.425 212.805 ;
        RECT 382.455 212.335 382.735 212.615 ;
        RECT 11.145 206.230 11.425 206.510 ;
        RECT 112.455 206.040 112.735 206.320 ;
        RECT 247.675 206.170 247.955 206.450 ;
        RECT 348.985 205.980 349.265 206.260 ;
        RECT 26.910 203.825 27.190 204.105 ;
        RECT 128.220 203.635 128.500 203.915 ;
        RECT 263.440 203.765 263.720 204.045 ;
        RECT 364.750 203.575 365.030 203.855 ;
        RECT 76.445 200.550 76.725 200.830 ;
        RECT 11.295 199.805 11.575 200.085 ;
        RECT 177.755 200.360 178.035 200.640 ;
        RECT 312.975 200.490 313.255 200.770 ;
        RECT 112.605 199.615 112.885 199.895 ;
        RECT 247.825 199.745 248.105 200.025 ;
        RECT 414.285 200.300 414.565 200.580 ;
        RECT 349.135 199.555 349.415 199.835 ;
        RECT 10.995 190.800 11.275 191.080 ;
        RECT 112.305 190.610 112.585 190.890 ;
        RECT 247.525 190.740 247.805 191.020 ;
        RECT 348.835 190.550 349.115 190.830 ;
        RECT 26.760 188.395 27.040 188.675 ;
        RECT 128.070 188.205 128.350 188.485 ;
        RECT 263.290 188.335 263.570 188.615 ;
        RECT 364.600 188.145 364.880 188.425 ;
        RECT 11.145 184.375 11.425 184.655 ;
        RECT 112.455 184.185 112.735 184.465 ;
        RECT 247.675 184.315 247.955 184.595 ;
        RECT 348.985 184.125 349.265 184.405 ;
        RECT 44.295 182.735 44.575 183.015 ;
        RECT 145.605 182.545 145.885 182.825 ;
        RECT 280.825 182.675 281.105 182.955 ;
        RECT 382.135 182.485 382.415 182.765 ;
        RECT 10.825 176.380 11.105 176.660 ;
        RECT 112.135 176.190 112.415 176.470 ;
        RECT 247.355 176.320 247.635 176.600 ;
        RECT 348.665 176.130 348.945 176.410 ;
        RECT 26.590 173.975 26.870 174.255 ;
        RECT 127.900 173.785 128.180 174.065 ;
        RECT 263.120 173.915 263.400 174.195 ;
        RECT 364.430 173.725 364.710 174.005 ;
        RECT 10.975 169.955 11.255 170.235 ;
        RECT 112.285 169.765 112.565 170.045 ;
        RECT 247.505 169.895 247.785 170.175 ;
        RECT 348.815 169.705 349.095 169.985 ;
        RECT 61.800 166.755 62.080 167.035 ;
        RECT 163.110 166.565 163.390 166.845 ;
        RECT 298.330 166.695 298.610 166.975 ;
        RECT 399.640 166.505 399.920 166.785 ;
        RECT 10.965 160.730 11.245 161.010 ;
        RECT 112.275 160.540 112.555 160.820 ;
        RECT 247.495 160.670 247.775 160.950 ;
        RECT 348.805 160.480 349.085 160.760 ;
        RECT 26.730 158.325 27.010 158.605 ;
        RECT 128.040 158.135 128.320 158.415 ;
        RECT 263.260 158.265 263.540 158.545 ;
        RECT 364.570 158.075 364.850 158.355 ;
        RECT 11.115 154.305 11.395 154.585 ;
        RECT 112.425 154.115 112.705 154.395 ;
        RECT 247.645 154.245 247.925 154.525 ;
        RECT 348.955 154.055 349.235 154.335 ;
        RECT 44.265 152.665 44.545 152.945 ;
        RECT 145.575 152.475 145.855 152.755 ;
        RECT 280.795 152.605 281.075 152.885 ;
        RECT 382.105 152.415 382.385 152.695 ;
        RECT 10.795 146.310 11.075 146.590 ;
        RECT 112.105 146.120 112.385 146.400 ;
        RECT 247.325 146.250 247.605 146.530 ;
        RECT 348.635 146.060 348.915 146.340 ;
        RECT 26.560 143.905 26.840 144.185 ;
        RECT 127.870 143.715 128.150 143.995 ;
        RECT 263.090 143.845 263.370 144.125 ;
        RECT 364.400 143.655 364.680 143.935 ;
        RECT 10.945 139.885 11.225 140.165 ;
        RECT 112.255 139.695 112.535 139.975 ;
        RECT 247.475 139.825 247.755 140.105 ;
        RECT 220.305 139.320 220.585 139.600 ;
        RECT 348.785 139.635 349.065 139.915 ;
        RECT 456.835 139.260 457.115 139.540 ;
        RECT 92.730 137.205 93.010 137.485 ;
        RECT 194.040 137.015 194.320 137.295 ;
        RECT 329.260 137.145 329.540 137.425 ;
        RECT 430.570 136.955 430.850 137.235 ;
        RECT 474.080 136.900 474.360 137.180 ;
        RECT 10.845 130.480 11.125 130.760 ;
        RECT 112.155 130.290 112.435 130.570 ;
        RECT 247.375 130.420 247.655 130.700 ;
        RECT 348.685 130.230 348.965 130.510 ;
        RECT 26.610 128.075 26.890 128.355 ;
        RECT 127.920 127.885 128.200 128.165 ;
        RECT 263.140 128.015 263.420 128.295 ;
        RECT 364.450 127.825 364.730 128.105 ;
        RECT 10.995 124.055 11.275 124.335 ;
        RECT 112.305 123.865 112.585 124.145 ;
        RECT 247.525 123.995 247.805 124.275 ;
        RECT 348.835 123.805 349.115 124.085 ;
        RECT 44.145 122.415 44.425 122.695 ;
        RECT 145.455 122.225 145.735 122.505 ;
        RECT 280.675 122.355 280.955 122.635 ;
        RECT 381.985 122.165 382.265 122.445 ;
        RECT 10.675 116.060 10.955 116.340 ;
        RECT 111.985 115.870 112.265 116.150 ;
        RECT 247.205 116.000 247.485 116.280 ;
        RECT 348.515 115.810 348.795 116.090 ;
        RECT 26.440 113.655 26.720 113.935 ;
        RECT 127.750 113.465 128.030 113.745 ;
        RECT 262.970 113.595 263.250 113.875 ;
        RECT 364.280 113.405 364.560 113.685 ;
        RECT 10.825 109.635 11.105 109.915 ;
        RECT 112.135 109.445 112.415 109.725 ;
        RECT 247.355 109.575 247.635 109.855 ;
        RECT 348.665 109.385 348.945 109.665 ;
        RECT 61.650 106.435 61.930 106.715 ;
        RECT 162.960 106.245 163.240 106.525 ;
        RECT 298.180 106.375 298.460 106.655 ;
        RECT 399.490 106.185 399.770 106.465 ;
        RECT 10.815 100.410 11.095 100.690 ;
        RECT 112.125 100.220 112.405 100.500 ;
        RECT 247.345 100.350 247.625 100.630 ;
        RECT 348.655 100.160 348.935 100.440 ;
        RECT 26.580 98.005 26.860 98.285 ;
        RECT 127.890 97.815 128.170 98.095 ;
        RECT 263.110 97.945 263.390 98.225 ;
        RECT 364.420 97.755 364.700 98.035 ;
        RECT 10.965 93.985 11.245 94.265 ;
        RECT 112.275 93.795 112.555 94.075 ;
        RECT 247.495 93.925 247.775 94.205 ;
        RECT 348.805 93.735 349.085 94.015 ;
        RECT 44.115 92.345 44.395 92.625 ;
        RECT 145.425 92.155 145.705 92.435 ;
        RECT 280.645 92.285 280.925 92.565 ;
        RECT 381.955 92.095 382.235 92.375 ;
        RECT 10.645 85.990 10.925 86.270 ;
        RECT 111.955 85.800 112.235 86.080 ;
        RECT 247.175 85.930 247.455 86.210 ;
        RECT 348.485 85.740 348.765 86.020 ;
        RECT 26.410 83.585 26.690 83.865 ;
        RECT 127.720 83.395 128.000 83.675 ;
        RECT 262.940 83.525 263.220 83.805 ;
        RECT 364.250 83.335 364.530 83.615 ;
        RECT 75.945 80.310 76.225 80.590 ;
        RECT 10.795 79.565 11.075 79.845 ;
        RECT 177.255 80.120 177.535 80.400 ;
        RECT 312.475 80.250 312.755 80.530 ;
        RECT 112.105 79.375 112.385 79.655 ;
        RECT 247.325 79.505 247.605 79.785 ;
        RECT 413.785 80.060 414.065 80.340 ;
        RECT 348.635 79.315 348.915 79.595 ;
        RECT 10.495 70.560 10.775 70.840 ;
        RECT 111.805 70.370 112.085 70.650 ;
        RECT 247.025 70.500 247.305 70.780 ;
        RECT 348.335 70.310 348.615 70.590 ;
        RECT 26.260 68.155 26.540 68.435 ;
        RECT 127.570 67.965 127.850 68.245 ;
        RECT 262.790 68.095 263.070 68.375 ;
        RECT 364.100 67.905 364.380 68.185 ;
        RECT 10.645 64.135 10.925 64.415 ;
        RECT 111.955 63.945 112.235 64.225 ;
        RECT 247.175 64.075 247.455 64.355 ;
        RECT 348.485 63.885 348.765 64.165 ;
        RECT 43.795 62.495 44.075 62.775 ;
        RECT 145.105 62.305 145.385 62.585 ;
        RECT 280.325 62.435 280.605 62.715 ;
        RECT 381.635 62.245 381.915 62.525 ;
        RECT 10.325 56.140 10.605 56.420 ;
        RECT 111.635 55.950 111.915 56.230 ;
        RECT 246.855 56.080 247.135 56.360 ;
        RECT 348.165 55.890 348.445 56.170 ;
        RECT 26.090 53.735 26.370 54.015 ;
        RECT 127.400 53.545 127.680 53.825 ;
        RECT 262.620 53.675 262.900 53.955 ;
        RECT 363.930 53.485 364.210 53.765 ;
        RECT 10.475 49.715 10.755 49.995 ;
        RECT 111.785 49.525 112.065 49.805 ;
        RECT 247.005 49.655 247.285 49.935 ;
        RECT 348.315 49.465 348.595 49.745 ;
        RECT 61.300 46.515 61.580 46.795 ;
        RECT 162.610 46.325 162.890 46.605 ;
        RECT 297.830 46.455 298.110 46.735 ;
        RECT 399.140 46.265 399.420 46.545 ;
        RECT 10.465 40.490 10.745 40.770 ;
        RECT 111.775 40.300 112.055 40.580 ;
        RECT 246.995 40.430 247.275 40.710 ;
        RECT 348.305 40.240 348.585 40.520 ;
        RECT 26.230 38.085 26.510 38.365 ;
        RECT 127.540 37.895 127.820 38.175 ;
        RECT 262.760 38.025 263.040 38.305 ;
        RECT 364.070 37.835 364.350 38.115 ;
        RECT 10.615 34.065 10.895 34.345 ;
        RECT 111.925 33.875 112.205 34.155 ;
        RECT 247.145 34.005 247.425 34.285 ;
        RECT 348.455 33.815 348.735 34.095 ;
        RECT 43.765 32.425 44.045 32.705 ;
        RECT 145.075 32.235 145.355 32.515 ;
        RECT 280.295 32.365 280.575 32.645 ;
        RECT 381.605 32.175 381.885 32.455 ;
        RECT 10.295 26.070 10.575 26.350 ;
        RECT 111.605 25.880 111.885 26.160 ;
        RECT 246.825 26.010 247.105 26.290 ;
        RECT 348.135 25.820 348.415 26.100 ;
        RECT 26.060 23.665 26.340 23.945 ;
        RECT 127.370 23.475 127.650 23.755 ;
        RECT 262.590 23.605 262.870 23.885 ;
        RECT 363.900 23.415 364.180 23.695 ;
        RECT 10.445 19.645 10.725 19.925 ;
        RECT 111.755 19.455 112.035 19.735 ;
        RECT 246.975 19.585 247.255 19.865 ;
        RECT 348.285 19.395 348.565 19.675 ;
      LAYER met3 ;
        RECT 11.270 251.570 11.810 252.120 ;
        RECT 11.280 251.160 11.680 251.570 ;
        RECT 112.580 251.380 113.120 251.930 ;
        RECT 247.800 251.510 248.340 252.060 ;
        RECT 11.280 250.640 11.700 251.160 ;
        RECT 112.590 250.970 112.990 251.380 ;
        RECT 247.810 251.100 248.210 251.510 ;
        RECT 349.110 251.320 349.650 251.870 ;
        RECT 11.280 250.620 11.640 250.640 ;
        RECT 112.590 250.450 113.010 250.970 ;
        RECT 247.810 250.580 248.230 251.100 ;
        RECT 349.120 250.910 349.520 251.320 ;
        RECT 247.810 250.560 248.170 250.580 ;
        RECT 112.590 250.430 112.950 250.450 ;
        RECT 349.120 250.390 349.540 250.910 ;
        RECT 349.120 250.370 349.480 250.390 ;
        RECT 27.000 249.280 27.510 249.770 ;
        RECT 27.000 248.200 27.500 249.280 ;
        RECT 128.310 249.090 128.820 249.580 ;
        RECT 263.530 249.220 264.040 249.710 ;
        RECT 128.310 248.010 128.810 249.090 ;
        RECT 263.530 248.140 264.030 249.220 ;
        RECT 364.840 249.030 365.350 249.520 ;
        RECT 364.840 247.950 365.340 249.030 ;
        RECT 11.450 245.080 11.900 245.510 ;
        RECT 11.450 244.220 11.890 245.080 ;
        RECT 112.760 244.890 113.210 245.320 ;
        RECT 247.980 245.020 248.430 245.450 ;
        RECT 112.760 244.030 113.200 244.890 ;
        RECT 247.980 244.160 248.420 245.020 ;
        RECT 349.290 244.830 349.740 245.260 ;
        RECT 349.290 243.970 349.730 244.830 ;
        RECT 44.570 242.590 45.020 243.760 ;
        RECT 145.880 242.400 146.330 243.570 ;
        RECT 281.100 242.530 281.550 243.700 ;
        RECT 382.410 242.340 382.860 243.510 ;
        RECT 11.100 237.150 11.640 237.700 ;
        RECT 11.110 236.740 11.510 237.150 ;
        RECT 112.410 236.960 112.950 237.510 ;
        RECT 247.630 237.090 248.170 237.640 ;
        RECT 11.110 236.220 11.530 236.740 ;
        RECT 112.420 236.550 112.820 236.960 ;
        RECT 247.640 236.680 248.040 237.090 ;
        RECT 348.940 236.900 349.480 237.450 ;
        RECT 11.110 236.200 11.470 236.220 ;
        RECT 112.420 236.030 112.840 236.550 ;
        RECT 247.640 236.160 248.060 236.680 ;
        RECT 348.950 236.490 349.350 236.900 ;
        RECT 247.640 236.140 248.000 236.160 ;
        RECT 112.420 236.010 112.780 236.030 ;
        RECT 348.950 235.970 349.370 236.490 ;
        RECT 348.950 235.950 349.310 235.970 ;
        RECT 26.830 234.860 27.340 235.350 ;
        RECT 26.830 233.780 27.330 234.860 ;
        RECT 128.140 234.670 128.650 235.160 ;
        RECT 263.360 234.800 263.870 235.290 ;
        RECT 128.140 233.590 128.640 234.670 ;
        RECT 263.360 233.720 263.860 234.800 ;
        RECT 364.670 234.610 365.180 235.100 ;
        RECT 364.670 233.530 365.170 234.610 ;
        RECT 11.280 230.660 11.730 231.090 ;
        RECT 11.280 229.800 11.720 230.660 ;
        RECT 112.590 230.470 113.040 230.900 ;
        RECT 247.810 230.600 248.260 231.030 ;
        RECT 112.590 229.610 113.030 230.470 ;
        RECT 247.810 229.740 248.250 230.600 ;
        RECT 349.120 230.410 349.570 230.840 ;
        RECT 349.120 229.550 349.560 230.410 ;
        RECT 62.100 227.380 62.480 227.720 ;
        RECT 62.090 226.620 62.480 227.380 ;
        RECT 163.410 227.190 163.790 227.530 ;
        RECT 298.630 227.320 299.010 227.660 ;
        RECT 163.400 226.430 163.790 227.190 ;
        RECT 298.620 226.560 299.010 227.320 ;
        RECT 399.940 227.130 400.320 227.470 ;
        RECT 399.930 226.370 400.320 227.130 ;
        RECT 11.240 221.500 11.780 222.050 ;
        RECT 11.250 221.090 11.650 221.500 ;
        RECT 112.550 221.310 113.090 221.860 ;
        RECT 247.770 221.440 248.310 221.990 ;
        RECT 11.250 220.570 11.670 221.090 ;
        RECT 112.560 220.900 112.960 221.310 ;
        RECT 247.780 221.030 248.180 221.440 ;
        RECT 349.080 221.250 349.620 221.800 ;
        RECT 11.250 220.550 11.610 220.570 ;
        RECT 112.560 220.380 112.980 220.900 ;
        RECT 247.780 220.510 248.200 221.030 ;
        RECT 349.090 220.840 349.490 221.250 ;
        RECT 247.780 220.490 248.140 220.510 ;
        RECT 112.560 220.360 112.920 220.380 ;
        RECT 349.090 220.320 349.510 220.840 ;
        RECT 349.090 220.300 349.450 220.320 ;
        RECT 26.970 219.210 27.480 219.700 ;
        RECT 26.970 218.130 27.470 219.210 ;
        RECT 128.280 219.020 128.790 219.510 ;
        RECT 263.500 219.150 264.010 219.640 ;
        RECT 128.280 217.940 128.780 219.020 ;
        RECT 263.500 218.070 264.000 219.150 ;
        RECT 364.810 218.960 365.320 219.450 ;
        RECT 364.810 217.880 365.310 218.960 ;
        RECT 11.420 215.010 11.870 215.440 ;
        RECT 11.420 214.150 11.860 215.010 ;
        RECT 112.730 214.820 113.180 215.250 ;
        RECT 247.950 214.950 248.400 215.380 ;
        RECT 112.730 213.960 113.170 214.820 ;
        RECT 247.950 214.090 248.390 214.950 ;
        RECT 349.260 214.760 349.710 215.190 ;
        RECT 349.260 213.900 349.700 214.760 ;
        RECT 44.540 212.520 44.990 213.690 ;
        RECT 145.850 212.330 146.300 213.500 ;
        RECT 281.070 212.460 281.520 213.630 ;
        RECT 382.380 212.270 382.830 213.440 ;
        RECT 11.070 207.080 11.610 207.630 ;
        RECT 11.080 206.670 11.480 207.080 ;
        RECT 112.380 206.890 112.920 207.440 ;
        RECT 247.600 207.020 248.140 207.570 ;
        RECT 11.080 206.150 11.500 206.670 ;
        RECT 112.390 206.480 112.790 206.890 ;
        RECT 247.610 206.610 248.010 207.020 ;
        RECT 348.910 206.830 349.450 207.380 ;
        RECT 11.080 206.130 11.440 206.150 ;
        RECT 112.390 205.960 112.810 206.480 ;
        RECT 247.610 206.090 248.030 206.610 ;
        RECT 348.920 206.420 349.320 206.830 ;
        RECT 247.610 206.070 247.970 206.090 ;
        RECT 112.390 205.940 112.750 205.960 ;
        RECT 348.920 205.900 349.340 206.420 ;
        RECT 348.920 205.880 349.280 205.900 ;
        RECT 26.800 204.790 27.310 205.280 ;
        RECT 26.800 203.710 27.300 204.790 ;
        RECT 128.110 204.600 128.620 205.090 ;
        RECT 263.330 204.730 263.840 205.220 ;
        RECT 128.110 203.520 128.610 204.600 ;
        RECT 263.330 203.650 263.830 204.730 ;
        RECT 364.640 204.540 365.150 205.030 ;
        RECT 364.640 203.460 365.140 204.540 ;
        RECT 11.250 200.590 11.700 201.020 ;
        RECT 76.310 200.980 76.900 201.580 ;
        RECT 11.250 199.730 11.690 200.590 ;
        RECT 76.330 200.450 76.810 200.980 ;
        RECT 112.560 200.400 113.010 200.830 ;
        RECT 177.620 200.790 178.210 201.390 ;
        RECT 112.560 199.540 113.000 200.400 ;
        RECT 177.640 200.260 178.120 200.790 ;
        RECT 247.780 200.530 248.230 200.960 ;
        RECT 312.840 200.920 313.430 201.520 ;
        RECT 247.780 199.670 248.220 200.530 ;
        RECT 312.860 200.390 313.340 200.920 ;
        RECT 349.090 200.340 349.540 200.770 ;
        RECT 414.150 200.730 414.740 201.330 ;
        RECT 349.090 199.480 349.530 200.340 ;
        RECT 414.170 200.200 414.650 200.730 ;
        RECT 10.920 191.650 11.460 192.200 ;
        RECT 10.930 191.240 11.330 191.650 ;
        RECT 112.230 191.460 112.770 192.010 ;
        RECT 247.450 191.590 247.990 192.140 ;
        RECT 10.930 190.720 11.350 191.240 ;
        RECT 112.240 191.050 112.640 191.460 ;
        RECT 247.460 191.180 247.860 191.590 ;
        RECT 348.760 191.400 349.300 191.950 ;
        RECT 10.930 190.700 11.290 190.720 ;
        RECT 112.240 190.530 112.660 191.050 ;
        RECT 247.460 190.660 247.880 191.180 ;
        RECT 348.770 190.990 349.170 191.400 ;
        RECT 247.460 190.640 247.820 190.660 ;
        RECT 112.240 190.510 112.600 190.530 ;
        RECT 348.770 190.470 349.190 190.990 ;
        RECT 348.770 190.450 349.130 190.470 ;
        RECT 26.650 189.360 27.160 189.850 ;
        RECT 26.650 188.280 27.150 189.360 ;
        RECT 127.960 189.170 128.470 189.660 ;
        RECT 263.180 189.300 263.690 189.790 ;
        RECT 127.960 188.090 128.460 189.170 ;
        RECT 263.180 188.220 263.680 189.300 ;
        RECT 364.490 189.110 365.000 189.600 ;
        RECT 364.490 188.030 364.990 189.110 ;
        RECT 11.100 185.160 11.550 185.590 ;
        RECT 11.100 184.300 11.540 185.160 ;
        RECT 112.410 184.970 112.860 185.400 ;
        RECT 247.630 185.100 248.080 185.530 ;
        RECT 112.410 184.110 112.850 184.970 ;
        RECT 247.630 184.240 248.070 185.100 ;
        RECT 348.940 184.910 349.390 185.340 ;
        RECT 348.940 184.050 349.380 184.910 ;
        RECT 44.220 182.670 44.670 183.840 ;
        RECT 145.530 182.480 145.980 183.650 ;
        RECT 280.750 182.610 281.200 183.780 ;
        RECT 382.060 182.420 382.510 183.590 ;
        RECT 10.750 177.230 11.290 177.780 ;
        RECT 10.760 176.820 11.160 177.230 ;
        RECT 112.060 177.040 112.600 177.590 ;
        RECT 247.280 177.170 247.820 177.720 ;
        RECT 10.760 176.300 11.180 176.820 ;
        RECT 112.070 176.630 112.470 177.040 ;
        RECT 247.290 176.760 247.690 177.170 ;
        RECT 348.590 176.980 349.130 177.530 ;
        RECT 10.760 176.280 11.120 176.300 ;
        RECT 112.070 176.110 112.490 176.630 ;
        RECT 247.290 176.240 247.710 176.760 ;
        RECT 348.600 176.570 349.000 176.980 ;
        RECT 247.290 176.220 247.650 176.240 ;
        RECT 112.070 176.090 112.430 176.110 ;
        RECT 348.600 176.050 349.020 176.570 ;
        RECT 348.600 176.030 348.960 176.050 ;
        RECT 26.480 174.940 26.990 175.430 ;
        RECT 26.480 173.860 26.980 174.940 ;
        RECT 127.790 174.750 128.300 175.240 ;
        RECT 263.010 174.880 263.520 175.370 ;
        RECT 127.790 173.670 128.290 174.750 ;
        RECT 263.010 173.800 263.510 174.880 ;
        RECT 364.320 174.690 364.830 175.180 ;
        RECT 364.320 173.610 364.820 174.690 ;
        RECT 10.930 170.740 11.380 171.170 ;
        RECT 10.930 169.880 11.370 170.740 ;
        RECT 112.240 170.550 112.690 170.980 ;
        RECT 247.460 170.680 247.910 171.110 ;
        RECT 112.240 169.690 112.680 170.550 ;
        RECT 247.460 169.820 247.900 170.680 ;
        RECT 348.770 170.490 349.220 170.920 ;
        RECT 348.770 169.630 349.210 170.490 ;
        RECT 61.750 167.460 62.130 167.800 ;
        RECT 61.740 166.700 62.130 167.460 ;
        RECT 163.060 167.270 163.440 167.610 ;
        RECT 298.280 167.400 298.660 167.740 ;
        RECT 163.050 166.510 163.440 167.270 ;
        RECT 298.270 166.640 298.660 167.400 ;
        RECT 399.590 167.210 399.970 167.550 ;
        RECT 399.580 166.450 399.970 167.210 ;
        RECT 10.890 161.580 11.430 162.130 ;
        RECT 10.900 161.170 11.300 161.580 ;
        RECT 112.200 161.390 112.740 161.940 ;
        RECT 247.420 161.520 247.960 162.070 ;
        RECT 10.900 160.650 11.320 161.170 ;
        RECT 112.210 160.980 112.610 161.390 ;
        RECT 247.430 161.110 247.830 161.520 ;
        RECT 348.730 161.330 349.270 161.880 ;
        RECT 10.900 160.630 11.260 160.650 ;
        RECT 112.210 160.460 112.630 160.980 ;
        RECT 247.430 160.590 247.850 161.110 ;
        RECT 348.740 160.920 349.140 161.330 ;
        RECT 247.430 160.570 247.790 160.590 ;
        RECT 112.210 160.440 112.570 160.460 ;
        RECT 348.740 160.400 349.160 160.920 ;
        RECT 348.740 160.380 349.100 160.400 ;
        RECT 26.620 159.290 27.130 159.780 ;
        RECT 26.620 158.210 27.120 159.290 ;
        RECT 127.930 159.100 128.440 159.590 ;
        RECT 263.150 159.230 263.660 159.720 ;
        RECT 127.930 158.020 128.430 159.100 ;
        RECT 263.150 158.150 263.650 159.230 ;
        RECT 364.460 159.040 364.970 159.530 ;
        RECT 364.460 157.960 364.960 159.040 ;
        RECT 11.070 155.090 11.520 155.520 ;
        RECT 11.070 154.230 11.510 155.090 ;
        RECT 112.380 154.900 112.830 155.330 ;
        RECT 247.600 155.030 248.050 155.460 ;
        RECT 112.380 154.040 112.820 154.900 ;
        RECT 247.600 154.170 248.040 155.030 ;
        RECT 348.910 154.840 349.360 155.270 ;
        RECT 348.910 153.980 349.350 154.840 ;
        RECT 44.190 152.600 44.640 153.770 ;
        RECT 145.500 152.410 145.950 153.580 ;
        RECT 280.720 152.540 281.170 153.710 ;
        RECT 382.030 152.350 382.480 153.520 ;
        RECT 10.720 147.160 11.260 147.710 ;
        RECT 10.730 146.750 11.130 147.160 ;
        RECT 112.030 146.970 112.570 147.520 ;
        RECT 247.250 147.100 247.790 147.650 ;
        RECT 10.730 146.230 11.150 146.750 ;
        RECT 112.040 146.560 112.440 146.970 ;
        RECT 247.260 146.690 247.660 147.100 ;
        RECT 348.560 146.910 349.100 147.460 ;
        RECT 10.730 146.210 11.090 146.230 ;
        RECT 112.040 146.040 112.460 146.560 ;
        RECT 247.260 146.170 247.680 146.690 ;
        RECT 348.570 146.500 348.970 146.910 ;
        RECT 247.260 146.150 247.620 146.170 ;
        RECT 112.040 146.020 112.400 146.040 ;
        RECT 348.570 145.980 348.990 146.500 ;
        RECT 348.570 145.960 348.930 145.980 ;
        RECT 26.450 144.870 26.960 145.360 ;
        RECT 26.450 143.790 26.950 144.870 ;
        RECT 127.760 144.680 128.270 145.170 ;
        RECT 262.980 144.810 263.490 145.300 ;
        RECT 127.760 143.600 128.260 144.680 ;
        RECT 262.980 143.730 263.480 144.810 ;
        RECT 364.290 144.620 364.800 145.110 ;
        RECT 364.290 143.540 364.790 144.620 ;
        RECT 10.900 140.670 11.350 141.100 ;
        RECT 10.900 139.810 11.340 140.670 ;
        RECT 112.210 140.480 112.660 140.910 ;
        RECT 247.430 140.610 247.880 141.040 ;
        RECT 112.210 139.620 112.650 140.480 ;
        RECT 220.210 139.270 220.710 140.150 ;
        RECT 247.430 139.750 247.870 140.610 ;
        RECT 348.740 140.420 349.190 140.850 ;
        RECT 348.740 139.560 349.180 140.420 ;
        RECT 456.740 139.210 457.240 140.090 ;
        RECT 92.630 137.150 93.080 138.240 ;
        RECT 193.940 136.960 194.390 138.050 ;
        RECT 329.160 137.090 329.610 138.180 ;
        RECT 430.470 136.900 430.920 137.990 ;
        RECT 474.050 137.280 474.450 137.690 ;
        RECT 474.050 136.860 474.400 137.280 ;
        RECT 10.770 131.330 11.310 131.880 ;
        RECT 10.780 130.920 11.180 131.330 ;
        RECT 112.080 131.140 112.620 131.690 ;
        RECT 247.300 131.270 247.840 131.820 ;
        RECT 10.780 130.400 11.200 130.920 ;
        RECT 112.090 130.730 112.490 131.140 ;
        RECT 247.310 130.860 247.710 131.270 ;
        RECT 348.610 131.080 349.150 131.630 ;
        RECT 10.780 130.380 11.140 130.400 ;
        RECT 112.090 130.210 112.510 130.730 ;
        RECT 247.310 130.340 247.730 130.860 ;
        RECT 348.620 130.670 349.020 131.080 ;
        RECT 247.310 130.320 247.670 130.340 ;
        RECT 112.090 130.190 112.450 130.210 ;
        RECT 348.620 130.150 349.040 130.670 ;
        RECT 348.620 130.130 348.980 130.150 ;
        RECT 26.500 129.040 27.010 129.530 ;
        RECT 26.500 127.960 27.000 129.040 ;
        RECT 127.810 128.850 128.320 129.340 ;
        RECT 263.030 128.980 263.540 129.470 ;
        RECT 127.810 127.770 128.310 128.850 ;
        RECT 263.030 127.900 263.530 128.980 ;
        RECT 364.340 128.790 364.850 129.280 ;
        RECT 364.340 127.710 364.840 128.790 ;
        RECT 10.950 124.840 11.400 125.270 ;
        RECT 10.950 123.980 11.390 124.840 ;
        RECT 112.260 124.650 112.710 125.080 ;
        RECT 247.480 124.780 247.930 125.210 ;
        RECT 112.260 123.790 112.700 124.650 ;
        RECT 247.480 123.920 247.920 124.780 ;
        RECT 348.790 124.590 349.240 125.020 ;
        RECT 348.790 123.730 349.230 124.590 ;
        RECT 44.070 122.350 44.520 123.520 ;
        RECT 145.380 122.160 145.830 123.330 ;
        RECT 280.600 122.290 281.050 123.460 ;
        RECT 381.910 122.100 382.360 123.270 ;
        RECT 10.600 116.910 11.140 117.460 ;
        RECT 10.610 116.500 11.010 116.910 ;
        RECT 111.910 116.720 112.450 117.270 ;
        RECT 247.130 116.850 247.670 117.400 ;
        RECT 10.610 115.980 11.030 116.500 ;
        RECT 111.920 116.310 112.320 116.720 ;
        RECT 247.140 116.440 247.540 116.850 ;
        RECT 348.440 116.660 348.980 117.210 ;
        RECT 10.610 115.960 10.970 115.980 ;
        RECT 111.920 115.790 112.340 116.310 ;
        RECT 247.140 115.920 247.560 116.440 ;
        RECT 348.450 116.250 348.850 116.660 ;
        RECT 247.140 115.900 247.500 115.920 ;
        RECT 111.920 115.770 112.280 115.790 ;
        RECT 348.450 115.730 348.870 116.250 ;
        RECT 348.450 115.710 348.810 115.730 ;
        RECT 26.330 114.620 26.840 115.110 ;
        RECT 26.330 113.540 26.830 114.620 ;
        RECT 127.640 114.430 128.150 114.920 ;
        RECT 262.860 114.560 263.370 115.050 ;
        RECT 127.640 113.350 128.140 114.430 ;
        RECT 262.860 113.480 263.360 114.560 ;
        RECT 364.170 114.370 364.680 114.860 ;
        RECT 364.170 113.290 364.670 114.370 ;
        RECT 10.780 110.420 11.230 110.850 ;
        RECT 10.780 109.560 11.220 110.420 ;
        RECT 112.090 110.230 112.540 110.660 ;
        RECT 247.310 110.360 247.760 110.790 ;
        RECT 112.090 109.370 112.530 110.230 ;
        RECT 247.310 109.500 247.750 110.360 ;
        RECT 348.620 110.170 349.070 110.600 ;
        RECT 348.620 109.310 349.060 110.170 ;
        RECT 61.600 107.140 61.980 107.480 ;
        RECT 61.590 106.380 61.980 107.140 ;
        RECT 162.910 106.950 163.290 107.290 ;
        RECT 298.130 107.080 298.510 107.420 ;
        RECT 162.900 106.190 163.290 106.950 ;
        RECT 298.120 106.320 298.510 107.080 ;
        RECT 399.440 106.890 399.820 107.230 ;
        RECT 399.430 106.130 399.820 106.890 ;
        RECT 10.740 101.260 11.280 101.810 ;
        RECT 10.750 100.850 11.150 101.260 ;
        RECT 112.050 101.070 112.590 101.620 ;
        RECT 247.270 101.200 247.810 101.750 ;
        RECT 10.750 100.330 11.170 100.850 ;
        RECT 112.060 100.660 112.460 101.070 ;
        RECT 247.280 100.790 247.680 101.200 ;
        RECT 348.580 101.010 349.120 101.560 ;
        RECT 10.750 100.310 11.110 100.330 ;
        RECT 112.060 100.140 112.480 100.660 ;
        RECT 247.280 100.270 247.700 100.790 ;
        RECT 348.590 100.600 348.990 101.010 ;
        RECT 247.280 100.250 247.640 100.270 ;
        RECT 112.060 100.120 112.420 100.140 ;
        RECT 348.590 100.080 349.010 100.600 ;
        RECT 348.590 100.060 348.950 100.080 ;
        RECT 26.470 98.970 26.980 99.460 ;
        RECT 26.470 97.890 26.970 98.970 ;
        RECT 127.780 98.780 128.290 99.270 ;
        RECT 263.000 98.910 263.510 99.400 ;
        RECT 127.780 97.700 128.280 98.780 ;
        RECT 263.000 97.830 263.500 98.910 ;
        RECT 364.310 98.720 364.820 99.210 ;
        RECT 364.310 97.640 364.810 98.720 ;
        RECT 10.920 94.770 11.370 95.200 ;
        RECT 10.920 93.910 11.360 94.770 ;
        RECT 112.230 94.580 112.680 95.010 ;
        RECT 247.450 94.710 247.900 95.140 ;
        RECT 112.230 93.720 112.670 94.580 ;
        RECT 247.450 93.850 247.890 94.710 ;
        RECT 348.760 94.520 349.210 94.950 ;
        RECT 348.760 93.660 349.200 94.520 ;
        RECT 44.040 92.280 44.490 93.450 ;
        RECT 145.350 92.090 145.800 93.260 ;
        RECT 280.570 92.220 281.020 93.390 ;
        RECT 381.880 92.030 382.330 93.200 ;
        RECT 10.570 86.840 11.110 87.390 ;
        RECT 10.580 86.430 10.980 86.840 ;
        RECT 111.880 86.650 112.420 87.200 ;
        RECT 247.100 86.780 247.640 87.330 ;
        RECT 10.580 85.910 11.000 86.430 ;
        RECT 111.890 86.240 112.290 86.650 ;
        RECT 247.110 86.370 247.510 86.780 ;
        RECT 348.410 86.590 348.950 87.140 ;
        RECT 10.580 85.890 10.940 85.910 ;
        RECT 111.890 85.720 112.310 86.240 ;
        RECT 247.110 85.850 247.530 86.370 ;
        RECT 348.420 86.180 348.820 86.590 ;
        RECT 247.110 85.830 247.470 85.850 ;
        RECT 111.890 85.700 112.250 85.720 ;
        RECT 348.420 85.660 348.840 86.180 ;
        RECT 348.420 85.640 348.780 85.660 ;
        RECT 26.300 84.550 26.810 85.040 ;
        RECT 26.300 83.470 26.800 84.550 ;
        RECT 127.610 84.360 128.120 84.850 ;
        RECT 262.830 84.490 263.340 84.980 ;
        RECT 127.610 83.280 128.110 84.360 ;
        RECT 262.830 83.410 263.330 84.490 ;
        RECT 364.140 84.300 364.650 84.790 ;
        RECT 364.140 83.220 364.640 84.300 ;
        RECT 10.750 80.350 11.200 80.780 ;
        RECT 75.810 80.740 76.400 81.340 ;
        RECT 10.750 79.490 11.190 80.350 ;
        RECT 75.830 80.210 76.310 80.740 ;
        RECT 112.060 80.160 112.510 80.590 ;
        RECT 177.120 80.550 177.710 81.150 ;
        RECT 112.060 79.300 112.500 80.160 ;
        RECT 177.140 80.020 177.620 80.550 ;
        RECT 247.280 80.290 247.730 80.720 ;
        RECT 312.340 80.680 312.930 81.280 ;
        RECT 247.280 79.430 247.720 80.290 ;
        RECT 312.360 80.150 312.840 80.680 ;
        RECT 348.590 80.100 349.040 80.530 ;
        RECT 413.650 80.490 414.240 81.090 ;
        RECT 348.590 79.240 349.030 80.100 ;
        RECT 413.670 79.960 414.150 80.490 ;
        RECT 10.420 71.410 10.960 71.960 ;
        RECT 10.430 71.000 10.830 71.410 ;
        RECT 111.730 71.220 112.270 71.770 ;
        RECT 246.950 71.350 247.490 71.900 ;
        RECT 10.430 70.480 10.850 71.000 ;
        RECT 111.740 70.810 112.140 71.220 ;
        RECT 246.960 70.940 247.360 71.350 ;
        RECT 348.260 71.160 348.800 71.710 ;
        RECT 10.430 70.460 10.790 70.480 ;
        RECT 111.740 70.290 112.160 70.810 ;
        RECT 246.960 70.420 247.380 70.940 ;
        RECT 348.270 70.750 348.670 71.160 ;
        RECT 246.960 70.400 247.320 70.420 ;
        RECT 111.740 70.270 112.100 70.290 ;
        RECT 348.270 70.230 348.690 70.750 ;
        RECT 348.270 70.210 348.630 70.230 ;
        RECT 26.150 69.120 26.660 69.610 ;
        RECT 26.150 68.040 26.650 69.120 ;
        RECT 127.460 68.930 127.970 69.420 ;
        RECT 262.680 69.060 263.190 69.550 ;
        RECT 127.460 67.850 127.960 68.930 ;
        RECT 262.680 67.980 263.180 69.060 ;
        RECT 363.990 68.870 364.500 69.360 ;
        RECT 363.990 67.790 364.490 68.870 ;
        RECT 10.600 64.920 11.050 65.350 ;
        RECT 10.600 64.060 11.040 64.920 ;
        RECT 111.910 64.730 112.360 65.160 ;
        RECT 247.130 64.860 247.580 65.290 ;
        RECT 111.910 63.870 112.350 64.730 ;
        RECT 247.130 64.000 247.570 64.860 ;
        RECT 348.440 64.670 348.890 65.100 ;
        RECT 348.440 63.810 348.880 64.670 ;
        RECT 43.720 62.430 44.170 63.600 ;
        RECT 145.030 62.240 145.480 63.410 ;
        RECT 280.250 62.370 280.700 63.540 ;
        RECT 381.560 62.180 382.010 63.350 ;
        RECT 10.250 56.990 10.790 57.540 ;
        RECT 10.260 56.580 10.660 56.990 ;
        RECT 111.560 56.800 112.100 57.350 ;
        RECT 246.780 56.930 247.320 57.480 ;
        RECT 10.260 56.060 10.680 56.580 ;
        RECT 111.570 56.390 111.970 56.800 ;
        RECT 246.790 56.520 247.190 56.930 ;
        RECT 348.090 56.740 348.630 57.290 ;
        RECT 10.260 56.040 10.620 56.060 ;
        RECT 111.570 55.870 111.990 56.390 ;
        RECT 246.790 56.000 247.210 56.520 ;
        RECT 348.100 56.330 348.500 56.740 ;
        RECT 246.790 55.980 247.150 56.000 ;
        RECT 111.570 55.850 111.930 55.870 ;
        RECT 348.100 55.810 348.520 56.330 ;
        RECT 348.100 55.790 348.460 55.810 ;
        RECT 25.980 54.700 26.490 55.190 ;
        RECT 25.980 53.620 26.480 54.700 ;
        RECT 127.290 54.510 127.800 55.000 ;
        RECT 262.510 54.640 263.020 55.130 ;
        RECT 127.290 53.430 127.790 54.510 ;
        RECT 262.510 53.560 263.010 54.640 ;
        RECT 363.820 54.450 364.330 54.940 ;
        RECT 363.820 53.370 364.320 54.450 ;
        RECT 10.430 50.500 10.880 50.930 ;
        RECT 10.430 49.640 10.870 50.500 ;
        RECT 111.740 50.310 112.190 50.740 ;
        RECT 246.960 50.440 247.410 50.870 ;
        RECT 111.740 49.450 112.180 50.310 ;
        RECT 246.960 49.580 247.400 50.440 ;
        RECT 348.270 50.250 348.720 50.680 ;
        RECT 348.270 49.390 348.710 50.250 ;
        RECT 61.250 47.220 61.630 47.560 ;
        RECT 61.240 46.460 61.630 47.220 ;
        RECT 162.560 47.030 162.940 47.370 ;
        RECT 297.780 47.160 298.160 47.500 ;
        RECT 162.550 46.270 162.940 47.030 ;
        RECT 297.770 46.400 298.160 47.160 ;
        RECT 399.090 46.970 399.470 47.310 ;
        RECT 399.080 46.210 399.470 46.970 ;
        RECT 10.390 41.340 10.930 41.890 ;
        RECT 10.400 40.930 10.800 41.340 ;
        RECT 111.700 41.150 112.240 41.700 ;
        RECT 246.920 41.280 247.460 41.830 ;
        RECT 10.400 40.410 10.820 40.930 ;
        RECT 111.710 40.740 112.110 41.150 ;
        RECT 246.930 40.870 247.330 41.280 ;
        RECT 348.230 41.090 348.770 41.640 ;
        RECT 10.400 40.390 10.760 40.410 ;
        RECT 111.710 40.220 112.130 40.740 ;
        RECT 246.930 40.350 247.350 40.870 ;
        RECT 348.240 40.680 348.640 41.090 ;
        RECT 246.930 40.330 247.290 40.350 ;
        RECT 111.710 40.200 112.070 40.220 ;
        RECT 348.240 40.160 348.660 40.680 ;
        RECT 348.240 40.140 348.600 40.160 ;
        RECT 26.120 39.050 26.630 39.540 ;
        RECT 26.120 37.970 26.620 39.050 ;
        RECT 127.430 38.860 127.940 39.350 ;
        RECT 262.650 38.990 263.160 39.480 ;
        RECT 127.430 37.780 127.930 38.860 ;
        RECT 262.650 37.910 263.150 38.990 ;
        RECT 363.960 38.800 364.470 39.290 ;
        RECT 363.960 37.720 364.460 38.800 ;
        RECT 10.570 34.850 11.020 35.280 ;
        RECT 10.570 33.990 11.010 34.850 ;
        RECT 111.880 34.660 112.330 35.090 ;
        RECT 247.100 34.790 247.550 35.220 ;
        RECT 111.880 33.800 112.320 34.660 ;
        RECT 247.100 33.930 247.540 34.790 ;
        RECT 348.410 34.600 348.860 35.030 ;
        RECT 348.410 33.740 348.850 34.600 ;
        RECT 43.690 32.360 44.140 33.530 ;
        RECT 145.000 32.170 145.450 33.340 ;
        RECT 280.220 32.300 280.670 33.470 ;
        RECT 381.530 32.110 381.980 33.280 ;
        RECT 10.220 26.920 10.760 27.470 ;
        RECT 10.230 26.510 10.630 26.920 ;
        RECT 111.530 26.730 112.070 27.280 ;
        RECT 246.750 26.860 247.290 27.410 ;
        RECT 10.230 25.990 10.650 26.510 ;
        RECT 111.540 26.320 111.940 26.730 ;
        RECT 246.760 26.450 247.160 26.860 ;
        RECT 348.060 26.670 348.600 27.220 ;
        RECT 10.230 25.970 10.590 25.990 ;
        RECT 111.540 25.800 111.960 26.320 ;
        RECT 246.760 25.930 247.180 26.450 ;
        RECT 348.070 26.260 348.470 26.670 ;
        RECT 246.760 25.910 247.120 25.930 ;
        RECT 111.540 25.780 111.900 25.800 ;
        RECT 348.070 25.740 348.490 26.260 ;
        RECT 348.070 25.720 348.430 25.740 ;
        RECT 25.950 24.630 26.460 25.120 ;
        RECT 25.950 23.550 26.450 24.630 ;
        RECT 127.260 24.440 127.770 24.930 ;
        RECT 262.480 24.570 262.990 25.060 ;
        RECT 127.260 23.360 127.760 24.440 ;
        RECT 262.480 23.490 262.980 24.570 ;
        RECT 363.790 24.380 364.300 24.870 ;
        RECT 363.790 23.300 364.290 24.380 ;
        RECT 10.400 20.430 10.850 20.860 ;
        RECT 10.400 19.570 10.840 20.430 ;
        RECT 111.710 20.240 112.160 20.670 ;
        RECT 246.930 20.370 247.380 20.800 ;
        RECT 111.710 19.380 112.150 20.240 ;
        RECT 246.930 19.510 247.370 20.370 ;
        RECT 348.240 20.180 348.690 20.610 ;
        RECT 348.240 19.320 348.680 20.180 ;
      LAYER via3 ;
        RECT 11.350 251.680 11.670 252.000 ;
        RECT 112.660 251.490 112.980 251.810 ;
        RECT 247.880 251.620 248.200 251.940 ;
        RECT 349.190 251.430 349.510 251.750 ;
        RECT 27.090 249.370 27.410 249.690 ;
        RECT 128.400 249.180 128.720 249.500 ;
        RECT 263.620 249.310 263.940 249.630 ;
        RECT 364.930 249.120 365.250 249.440 ;
        RECT 11.510 245.115 11.830 245.435 ;
        RECT 112.820 244.925 113.140 245.245 ;
        RECT 248.040 245.055 248.360 245.375 ;
        RECT 349.350 244.865 349.670 245.185 ;
        RECT 44.640 243.365 44.960 243.685 ;
        RECT 145.950 243.175 146.270 243.495 ;
        RECT 281.170 243.305 281.490 243.625 ;
        RECT 382.480 243.115 382.800 243.435 ;
        RECT 11.180 237.260 11.500 237.580 ;
        RECT 112.490 237.070 112.810 237.390 ;
        RECT 247.710 237.200 248.030 237.520 ;
        RECT 349.020 237.010 349.340 237.330 ;
        RECT 26.920 234.950 27.240 235.270 ;
        RECT 128.230 234.760 128.550 235.080 ;
        RECT 263.450 234.890 263.770 235.210 ;
        RECT 364.760 234.700 365.080 235.020 ;
        RECT 11.340 230.695 11.660 231.015 ;
        RECT 112.650 230.505 112.970 230.825 ;
        RECT 247.870 230.635 248.190 230.955 ;
        RECT 349.180 230.445 349.500 230.765 ;
        RECT 62.150 227.330 62.470 227.650 ;
        RECT 163.460 227.140 163.780 227.460 ;
        RECT 298.680 227.270 299.000 227.590 ;
        RECT 399.990 227.080 400.310 227.400 ;
        RECT 11.320 221.610 11.640 221.930 ;
        RECT 112.630 221.420 112.950 221.740 ;
        RECT 247.850 221.550 248.170 221.870 ;
        RECT 349.160 221.360 349.480 221.680 ;
        RECT 27.060 219.300 27.380 219.620 ;
        RECT 128.370 219.110 128.690 219.430 ;
        RECT 263.590 219.240 263.910 219.560 ;
        RECT 364.900 219.050 365.220 219.370 ;
        RECT 11.480 215.045 11.800 215.365 ;
        RECT 112.790 214.855 113.110 215.175 ;
        RECT 248.010 214.985 248.330 215.305 ;
        RECT 349.320 214.795 349.640 215.115 ;
        RECT 44.610 213.295 44.930 213.615 ;
        RECT 145.920 213.105 146.240 213.425 ;
        RECT 281.140 213.235 281.460 213.555 ;
        RECT 382.450 213.045 382.770 213.365 ;
        RECT 11.150 207.190 11.470 207.510 ;
        RECT 112.460 207.000 112.780 207.320 ;
        RECT 247.680 207.130 248.000 207.450 ;
        RECT 348.990 206.940 349.310 207.260 ;
        RECT 26.890 204.880 27.210 205.200 ;
        RECT 128.200 204.690 128.520 205.010 ;
        RECT 263.420 204.820 263.740 205.140 ;
        RECT 364.730 204.630 365.050 204.950 ;
        RECT 76.460 201.090 76.780 201.410 ;
        RECT 11.310 200.625 11.630 200.945 ;
        RECT 177.770 200.900 178.090 201.220 ;
        RECT 312.990 201.030 313.310 201.350 ;
        RECT 112.620 200.435 112.940 200.755 ;
        RECT 247.840 200.565 248.160 200.885 ;
        RECT 414.300 200.840 414.620 201.160 ;
        RECT 349.150 200.375 349.470 200.695 ;
        RECT 11.000 191.760 11.320 192.080 ;
        RECT 112.310 191.570 112.630 191.890 ;
        RECT 247.530 191.700 247.850 192.020 ;
        RECT 348.840 191.510 349.160 191.830 ;
        RECT 26.740 189.450 27.060 189.770 ;
        RECT 128.050 189.260 128.370 189.580 ;
        RECT 263.270 189.390 263.590 189.710 ;
        RECT 364.580 189.200 364.900 189.520 ;
        RECT 11.160 185.195 11.480 185.515 ;
        RECT 112.470 185.005 112.790 185.325 ;
        RECT 247.690 185.135 248.010 185.455 ;
        RECT 349.000 184.945 349.320 185.265 ;
        RECT 44.290 183.445 44.610 183.765 ;
        RECT 145.600 183.255 145.920 183.575 ;
        RECT 280.820 183.385 281.140 183.705 ;
        RECT 382.130 183.195 382.450 183.515 ;
        RECT 10.830 177.340 11.150 177.660 ;
        RECT 112.140 177.150 112.460 177.470 ;
        RECT 247.360 177.280 247.680 177.600 ;
        RECT 348.670 177.090 348.990 177.410 ;
        RECT 26.570 175.030 26.890 175.350 ;
        RECT 127.880 174.840 128.200 175.160 ;
        RECT 263.100 174.970 263.420 175.290 ;
        RECT 364.410 174.780 364.730 175.100 ;
        RECT 10.990 170.775 11.310 171.095 ;
        RECT 112.300 170.585 112.620 170.905 ;
        RECT 247.520 170.715 247.840 171.035 ;
        RECT 348.830 170.525 349.150 170.845 ;
        RECT 61.800 167.410 62.120 167.730 ;
        RECT 163.110 167.220 163.430 167.540 ;
        RECT 298.330 167.350 298.650 167.670 ;
        RECT 399.640 167.160 399.960 167.480 ;
        RECT 10.970 161.690 11.290 162.010 ;
        RECT 112.280 161.500 112.600 161.820 ;
        RECT 247.500 161.630 247.820 161.950 ;
        RECT 348.810 161.440 349.130 161.760 ;
        RECT 26.710 159.380 27.030 159.700 ;
        RECT 128.020 159.190 128.340 159.510 ;
        RECT 263.240 159.320 263.560 159.640 ;
        RECT 364.550 159.130 364.870 159.450 ;
        RECT 11.130 155.125 11.450 155.445 ;
        RECT 112.440 154.935 112.760 155.255 ;
        RECT 247.660 155.065 247.980 155.385 ;
        RECT 348.970 154.875 349.290 155.195 ;
        RECT 44.260 153.375 44.580 153.695 ;
        RECT 145.570 153.185 145.890 153.505 ;
        RECT 280.790 153.315 281.110 153.635 ;
        RECT 382.100 153.125 382.420 153.445 ;
        RECT 10.800 147.270 11.120 147.590 ;
        RECT 112.110 147.080 112.430 147.400 ;
        RECT 247.330 147.210 247.650 147.530 ;
        RECT 348.640 147.020 348.960 147.340 ;
        RECT 26.540 144.960 26.860 145.280 ;
        RECT 127.850 144.770 128.170 145.090 ;
        RECT 263.070 144.900 263.390 145.220 ;
        RECT 364.380 144.710 364.700 145.030 ;
        RECT 10.960 140.705 11.280 141.025 ;
        RECT 112.270 140.515 112.590 140.835 ;
        RECT 247.490 140.645 247.810 140.965 ;
        RECT 220.315 139.790 220.635 140.110 ;
        RECT 348.800 140.455 349.120 140.775 ;
        RECT 456.845 139.730 457.165 140.050 ;
        RECT 92.705 137.820 93.025 138.140 ;
        RECT 194.015 137.630 194.335 137.950 ;
        RECT 329.235 137.760 329.555 138.080 ;
        RECT 430.545 137.570 430.865 137.890 ;
        RECT 474.100 137.330 474.420 137.650 ;
        RECT 10.850 131.440 11.170 131.760 ;
        RECT 112.160 131.250 112.480 131.570 ;
        RECT 247.380 131.380 247.700 131.700 ;
        RECT 348.690 131.190 349.010 131.510 ;
        RECT 26.590 129.130 26.910 129.450 ;
        RECT 127.900 128.940 128.220 129.260 ;
        RECT 263.120 129.070 263.440 129.390 ;
        RECT 364.430 128.880 364.750 129.200 ;
        RECT 11.010 124.875 11.330 125.195 ;
        RECT 112.320 124.685 112.640 125.005 ;
        RECT 247.540 124.815 247.860 125.135 ;
        RECT 348.850 124.625 349.170 124.945 ;
        RECT 44.140 123.125 44.460 123.445 ;
        RECT 145.450 122.935 145.770 123.255 ;
        RECT 280.670 123.065 280.990 123.385 ;
        RECT 381.980 122.875 382.300 123.195 ;
        RECT 10.680 117.020 11.000 117.340 ;
        RECT 111.990 116.830 112.310 117.150 ;
        RECT 247.210 116.960 247.530 117.280 ;
        RECT 348.520 116.770 348.840 117.090 ;
        RECT 26.420 114.710 26.740 115.030 ;
        RECT 127.730 114.520 128.050 114.840 ;
        RECT 262.950 114.650 263.270 114.970 ;
        RECT 364.260 114.460 364.580 114.780 ;
        RECT 10.840 110.455 11.160 110.775 ;
        RECT 112.150 110.265 112.470 110.585 ;
        RECT 247.370 110.395 247.690 110.715 ;
        RECT 348.680 110.205 349.000 110.525 ;
        RECT 61.650 107.090 61.970 107.410 ;
        RECT 162.960 106.900 163.280 107.220 ;
        RECT 298.180 107.030 298.500 107.350 ;
        RECT 399.490 106.840 399.810 107.160 ;
        RECT 10.820 101.370 11.140 101.690 ;
        RECT 112.130 101.180 112.450 101.500 ;
        RECT 247.350 101.310 247.670 101.630 ;
        RECT 348.660 101.120 348.980 101.440 ;
        RECT 26.560 99.060 26.880 99.380 ;
        RECT 127.870 98.870 128.190 99.190 ;
        RECT 263.090 99.000 263.410 99.320 ;
        RECT 364.400 98.810 364.720 99.130 ;
        RECT 10.980 94.805 11.300 95.125 ;
        RECT 112.290 94.615 112.610 94.935 ;
        RECT 247.510 94.745 247.830 95.065 ;
        RECT 348.820 94.555 349.140 94.875 ;
        RECT 44.110 93.055 44.430 93.375 ;
        RECT 145.420 92.865 145.740 93.185 ;
        RECT 280.640 92.995 280.960 93.315 ;
        RECT 381.950 92.805 382.270 93.125 ;
        RECT 10.650 86.950 10.970 87.270 ;
        RECT 111.960 86.760 112.280 87.080 ;
        RECT 247.180 86.890 247.500 87.210 ;
        RECT 348.490 86.700 348.810 87.020 ;
        RECT 26.390 84.640 26.710 84.960 ;
        RECT 127.700 84.450 128.020 84.770 ;
        RECT 262.920 84.580 263.240 84.900 ;
        RECT 364.230 84.390 364.550 84.710 ;
        RECT 75.960 80.850 76.280 81.170 ;
        RECT 10.810 80.385 11.130 80.705 ;
        RECT 177.270 80.660 177.590 80.980 ;
        RECT 312.490 80.790 312.810 81.110 ;
        RECT 112.120 80.195 112.440 80.515 ;
        RECT 247.340 80.325 247.660 80.645 ;
        RECT 413.800 80.600 414.120 80.920 ;
        RECT 348.650 80.135 348.970 80.455 ;
        RECT 10.500 71.520 10.820 71.840 ;
        RECT 111.810 71.330 112.130 71.650 ;
        RECT 247.030 71.460 247.350 71.780 ;
        RECT 348.340 71.270 348.660 71.590 ;
        RECT 26.240 69.210 26.560 69.530 ;
        RECT 127.550 69.020 127.870 69.340 ;
        RECT 262.770 69.150 263.090 69.470 ;
        RECT 364.080 68.960 364.400 69.280 ;
        RECT 10.660 64.955 10.980 65.275 ;
        RECT 111.970 64.765 112.290 65.085 ;
        RECT 247.190 64.895 247.510 65.215 ;
        RECT 348.500 64.705 348.820 65.025 ;
        RECT 43.790 63.205 44.110 63.525 ;
        RECT 145.100 63.015 145.420 63.335 ;
        RECT 280.320 63.145 280.640 63.465 ;
        RECT 381.630 62.955 381.950 63.275 ;
        RECT 10.330 57.100 10.650 57.420 ;
        RECT 111.640 56.910 111.960 57.230 ;
        RECT 246.860 57.040 247.180 57.360 ;
        RECT 348.170 56.850 348.490 57.170 ;
        RECT 26.070 54.790 26.390 55.110 ;
        RECT 127.380 54.600 127.700 54.920 ;
        RECT 262.600 54.730 262.920 55.050 ;
        RECT 363.910 54.540 364.230 54.860 ;
        RECT 10.490 50.535 10.810 50.855 ;
        RECT 111.800 50.345 112.120 50.665 ;
        RECT 247.020 50.475 247.340 50.795 ;
        RECT 348.330 50.285 348.650 50.605 ;
        RECT 61.300 47.170 61.620 47.490 ;
        RECT 162.610 46.980 162.930 47.300 ;
        RECT 297.830 47.110 298.150 47.430 ;
        RECT 399.140 46.920 399.460 47.240 ;
        RECT 10.470 41.450 10.790 41.770 ;
        RECT 111.780 41.260 112.100 41.580 ;
        RECT 247.000 41.390 247.320 41.710 ;
        RECT 348.310 41.200 348.630 41.520 ;
        RECT 26.210 39.140 26.530 39.460 ;
        RECT 127.520 38.950 127.840 39.270 ;
        RECT 262.740 39.080 263.060 39.400 ;
        RECT 364.050 38.890 364.370 39.210 ;
        RECT 10.630 34.885 10.950 35.205 ;
        RECT 111.940 34.695 112.260 35.015 ;
        RECT 247.160 34.825 247.480 35.145 ;
        RECT 348.470 34.635 348.790 34.955 ;
        RECT 43.760 33.135 44.080 33.455 ;
        RECT 145.070 32.945 145.390 33.265 ;
        RECT 280.290 33.075 280.610 33.395 ;
        RECT 381.600 32.885 381.920 33.205 ;
        RECT 10.300 27.030 10.620 27.350 ;
        RECT 111.610 26.840 111.930 27.160 ;
        RECT 246.830 26.970 247.150 27.290 ;
        RECT 348.140 26.780 348.460 27.100 ;
        RECT 26.040 24.720 26.360 25.040 ;
        RECT 127.350 24.530 127.670 24.850 ;
        RECT 262.570 24.660 262.890 24.980 ;
        RECT 363.880 24.470 364.200 24.790 ;
        RECT 10.460 20.465 10.780 20.785 ;
        RECT 111.770 20.275 112.090 20.595 ;
        RECT 246.990 20.405 247.310 20.725 ;
        RECT 348.300 20.215 348.620 20.535 ;
      LAYER met4 ;
        RECT 14.180 252.130 19.500 276.245 ;
        RECT 118.810 257.480 248.820 257.500 ;
        RECT 113.760 257.170 248.820 257.480 ;
        RECT 113.760 257.160 119.040 257.170 ;
        RECT 113.820 253.510 114.240 257.160 ;
        RECT 39.990 253.490 40.470 253.510 ;
        RECT 113.560 253.490 114.240 253.510 ;
        RECT 39.990 253.110 114.240 253.490 ;
        RECT 39.990 253.080 114.210 253.110 ;
        RECT 14.110 252.120 23.380 252.130 ;
        RECT 25.610 252.120 27.520 252.140 ;
        RECT 11.280 251.600 27.520 252.120 ;
        RECT 11.280 251.590 25.690 251.600 ;
        RECT 11.280 251.580 14.120 251.590 ;
        RECT 23.330 251.580 25.690 251.590 ;
        RECT 11.890 245.500 12.440 251.580 ;
        RECT 27.000 250.120 27.490 251.600 ;
        RECT 36.990 250.170 37.500 250.300 ;
        RECT 39.990 250.170 40.470 253.080 ;
        RECT 113.560 253.070 114.210 253.080 ;
        RECT 113.830 251.930 114.210 253.070 ;
        RECT 248.460 252.060 248.810 257.170 ;
        RECT 276.520 253.430 277.000 253.450 ;
        RECT 350.090 253.430 350.740 253.450 ;
        RECT 276.520 253.020 350.740 253.430 ;
        RECT 250.640 252.060 259.910 252.070 ;
        RECT 262.140 252.060 264.050 252.080 ;
        RECT 115.420 251.930 124.690 251.940 ;
        RECT 126.920 251.930 128.830 251.950 ;
        RECT 112.590 251.410 128.830 251.930 ;
        RECT 247.810 251.540 264.050 252.060 ;
        RECT 247.810 251.530 262.220 251.540 ;
        RECT 247.810 251.520 250.650 251.530 ;
        RECT 259.860 251.520 262.220 251.530 ;
        RECT 112.590 251.400 127.000 251.410 ;
        RECT 112.590 251.390 115.430 251.400 ;
        RECT 124.640 251.390 127.000 251.400 ;
        RECT 41.720 250.170 45.050 250.190 ;
        RECT 34.820 250.140 45.050 250.170 ;
        RECT 34.260 250.130 45.050 250.140 ;
        RECT 32.550 250.120 45.050 250.130 ;
        RECT 27.000 249.770 45.050 250.120 ;
        RECT 27.000 249.760 34.330 249.770 ;
        RECT 27.000 249.750 32.620 249.760 ;
        RECT 27.000 249.280 27.510 249.750 ;
        RECT 34.820 249.730 45.050 249.770 ;
        RECT 11.450 245.100 12.440 245.500 ;
        RECT 11.450 245.080 12.030 245.100 ;
        RECT 36.990 238.250 37.500 249.730 ;
        RECT 39.990 249.710 40.470 249.730 ;
        RECT 41.720 249.690 45.050 249.730 ;
        RECT 44.580 243.940 45.020 249.690 ;
        RECT 113.200 245.310 113.750 251.390 ;
        RECT 128.310 249.930 128.800 251.410 ;
        RECT 138.300 249.980 138.810 250.110 ;
        RECT 143.030 249.980 146.360 250.000 ;
        RECT 136.130 249.950 146.360 249.980 ;
        RECT 135.570 249.940 146.360 249.950 ;
        RECT 133.860 249.930 146.360 249.940 ;
        RECT 128.310 249.580 146.360 249.930 ;
        RECT 128.310 249.570 135.640 249.580 ;
        RECT 128.310 249.560 133.930 249.570 ;
        RECT 128.310 249.090 128.820 249.560 ;
        RECT 136.130 249.540 146.360 249.580 ;
        RECT 112.760 244.910 113.750 245.310 ;
        RECT 112.760 244.890 113.340 244.910 ;
        RECT 44.570 243.320 45.020 243.940 ;
        RECT 36.990 237.940 37.480 238.250 ;
        RECT 30.310 237.740 37.480 237.940 ;
        RECT 138.300 238.060 138.810 249.540 ;
        RECT 143.030 249.500 146.360 249.540 ;
        RECT 145.890 243.750 146.330 249.500 ;
        RECT 248.420 245.440 248.970 251.520 ;
        RECT 263.530 250.060 264.020 251.540 ;
        RECT 273.520 250.110 274.030 250.240 ;
        RECT 276.520 250.110 277.000 253.020 ;
        RECT 350.090 253.010 350.740 253.020 ;
        RECT 350.360 251.870 350.740 253.010 ;
        RECT 351.950 251.870 361.220 251.880 ;
        RECT 363.450 251.870 365.360 251.890 ;
        RECT 349.120 251.350 365.360 251.870 ;
        RECT 349.120 251.340 363.530 251.350 ;
        RECT 349.120 251.330 351.960 251.340 ;
        RECT 361.170 251.330 363.530 251.340 ;
        RECT 278.250 250.110 281.580 250.130 ;
        RECT 271.350 250.080 281.580 250.110 ;
        RECT 270.790 250.070 281.580 250.080 ;
        RECT 269.080 250.060 281.580 250.070 ;
        RECT 263.530 249.710 281.580 250.060 ;
        RECT 263.530 249.700 270.860 249.710 ;
        RECT 263.530 249.690 269.150 249.700 ;
        RECT 263.530 249.220 264.040 249.690 ;
        RECT 271.350 249.670 281.580 249.710 ;
        RECT 247.980 245.040 248.970 245.440 ;
        RECT 247.980 245.020 248.560 245.040 ;
        RECT 145.880 243.130 146.330 243.750 ;
        RECT 273.520 238.190 274.030 249.670 ;
        RECT 276.520 249.650 277.000 249.670 ;
        RECT 278.250 249.630 281.580 249.670 ;
        RECT 281.110 243.880 281.550 249.630 ;
        RECT 349.730 245.250 350.280 251.330 ;
        RECT 364.840 249.870 365.330 251.350 ;
        RECT 374.830 249.920 375.340 250.050 ;
        RECT 379.560 249.920 382.890 249.940 ;
        RECT 372.660 249.890 382.890 249.920 ;
        RECT 372.100 249.880 382.890 249.890 ;
        RECT 370.390 249.870 382.890 249.880 ;
        RECT 364.840 249.520 382.890 249.870 ;
        RECT 364.840 249.510 372.170 249.520 ;
        RECT 364.840 249.500 370.460 249.510 ;
        RECT 364.840 249.030 365.350 249.500 ;
        RECT 372.660 249.480 382.890 249.520 ;
        RECT 349.290 244.850 350.280 245.250 ;
        RECT 349.290 244.830 349.870 244.850 ;
        RECT 281.100 243.260 281.550 243.880 ;
        RECT 138.300 237.750 138.790 238.060 ;
        RECT 273.520 237.880 274.010 238.190 ;
        RECT 26.770 237.720 37.480 237.740 ;
        RECT 13.940 237.700 23.210 237.710 ;
        RECT 25.440 237.700 37.480 237.720 ;
        RECT 11.110 237.180 37.480 237.700 ;
        RECT 131.620 237.550 138.790 237.750 ;
        RECT 266.840 237.680 274.010 237.880 ;
        RECT 374.830 238.000 375.340 249.480 ;
        RECT 379.560 249.440 382.890 249.480 ;
        RECT 382.420 243.690 382.860 249.440 ;
        RECT 382.410 243.070 382.860 243.690 ;
        RECT 374.830 237.690 375.320 238.000 ;
        RECT 263.300 237.660 274.010 237.680 ;
        RECT 250.470 237.640 259.740 237.650 ;
        RECT 261.970 237.640 274.010 237.660 ;
        RECT 128.080 237.530 138.790 237.550 ;
        RECT 115.250 237.510 124.520 237.520 ;
        RECT 126.750 237.510 138.790 237.530 ;
        RECT 11.110 237.170 25.520 237.180 ;
        RECT 11.110 237.160 13.950 237.170 ;
        RECT 23.160 237.160 25.520 237.170 ;
        RECT 26.770 237.160 37.480 237.180 ;
        RECT 11.720 231.080 12.270 237.160 ;
        RECT 26.770 237.140 30.590 237.160 ;
        RECT 26.830 235.350 27.320 237.140 ;
        RECT 26.830 234.860 27.340 235.350 ;
        RECT 11.280 230.680 12.270 231.080 ;
        RECT 11.280 230.660 11.860 230.680 ;
        RECT 37.060 228.330 37.450 237.160 ;
        RECT 112.420 236.990 138.790 237.510 ;
        RECT 247.640 237.120 274.010 237.640 ;
        RECT 368.150 237.490 375.320 237.690 ;
        RECT 364.610 237.470 375.320 237.490 ;
        RECT 351.780 237.450 361.050 237.460 ;
        RECT 363.280 237.450 375.320 237.470 ;
        RECT 247.640 237.110 262.050 237.120 ;
        RECT 247.640 237.100 250.480 237.110 ;
        RECT 259.690 237.100 262.050 237.110 ;
        RECT 263.300 237.100 274.010 237.120 ;
        RECT 112.420 236.980 126.830 236.990 ;
        RECT 112.420 236.970 115.260 236.980 ;
        RECT 124.470 236.970 126.830 236.980 ;
        RECT 128.080 236.970 138.790 236.990 ;
        RECT 113.030 230.890 113.580 236.970 ;
        RECT 128.080 236.950 131.900 236.970 ;
        RECT 128.140 235.160 128.630 236.950 ;
        RECT 128.140 234.670 128.650 235.160 ;
        RECT 112.590 230.490 113.580 230.890 ;
        RECT 112.590 230.470 113.170 230.490 ;
        RECT 53.490 228.330 53.930 228.340 ;
        RECT 36.950 227.940 62.480 228.330 ;
        RECT 138.370 228.140 138.760 236.970 ;
        RECT 248.250 231.020 248.800 237.100 ;
        RECT 263.300 237.080 267.120 237.100 ;
        RECT 263.360 235.290 263.850 237.080 ;
        RECT 263.360 234.800 263.870 235.290 ;
        RECT 247.810 230.620 248.800 231.020 ;
        RECT 247.810 230.600 248.390 230.620 ;
        RECT 273.590 228.270 273.980 237.100 ;
        RECT 348.950 236.930 375.320 237.450 ;
        RECT 348.950 236.920 363.360 236.930 ;
        RECT 348.950 236.910 351.790 236.920 ;
        RECT 361.000 236.910 363.360 236.920 ;
        RECT 364.610 236.910 375.320 236.930 ;
        RECT 349.560 230.830 350.110 236.910 ;
        RECT 364.610 236.890 368.430 236.910 ;
        RECT 364.670 235.100 365.160 236.890 ;
        RECT 364.670 234.610 365.180 235.100 ;
        RECT 349.120 230.430 350.110 230.830 ;
        RECT 349.120 230.410 349.700 230.430 ;
        RECT 290.020 228.270 290.460 228.280 ;
        RECT 154.800 228.140 155.240 228.150 ;
        RECT 14.080 222.050 23.350 222.060 ;
        RECT 25.580 222.050 27.490 222.070 ;
        RECT 11.250 221.530 27.490 222.050 ;
        RECT 11.250 221.520 25.660 221.530 ;
        RECT 11.250 221.510 14.090 221.520 ;
        RECT 23.300 221.510 25.660 221.520 ;
        RECT 11.860 215.430 12.410 221.510 ;
        RECT 26.970 220.050 27.460 221.530 ;
        RECT 37.060 220.230 37.450 227.940 ;
        RECT 36.960 220.100 37.470 220.230 ;
        RECT 41.690 220.100 45.020 220.120 ;
        RECT 34.790 220.070 45.020 220.100 ;
        RECT 34.230 220.060 45.020 220.070 ;
        RECT 32.520 220.050 45.020 220.060 ;
        RECT 26.970 219.700 45.020 220.050 ;
        RECT 26.970 219.690 34.300 219.700 ;
        RECT 26.970 219.680 32.590 219.690 ;
        RECT 26.970 219.210 27.480 219.680 ;
        RECT 34.790 219.660 45.020 219.700 ;
        RECT 11.420 215.030 12.410 215.430 ;
        RECT 11.420 215.010 12.000 215.030 ;
        RECT 36.960 208.180 37.470 219.660 ;
        RECT 41.690 219.620 45.020 219.660 ;
        RECT 44.550 213.870 44.990 219.620 ;
        RECT 44.540 213.250 44.990 213.870 ;
        RECT 53.490 209.890 53.930 227.940 ;
        RECT 62.100 227.270 62.480 227.940 ;
        RECT 138.260 227.750 163.790 228.140 ;
        RECT 273.480 227.880 299.010 228.270 ;
        RECT 374.900 228.080 375.290 236.910 ;
        RECT 391.330 228.080 391.770 228.090 ;
        RECT 115.390 221.860 124.660 221.870 ;
        RECT 126.890 221.860 128.800 221.880 ;
        RECT 112.560 221.340 128.800 221.860 ;
        RECT 112.560 221.330 126.970 221.340 ;
        RECT 112.560 221.320 115.400 221.330 ;
        RECT 124.610 221.320 126.970 221.330 ;
        RECT 113.170 215.240 113.720 221.320 ;
        RECT 128.280 219.860 128.770 221.340 ;
        RECT 138.370 220.040 138.760 227.750 ;
        RECT 138.270 219.910 138.780 220.040 ;
        RECT 143.000 219.910 146.330 219.930 ;
        RECT 136.100 219.880 146.330 219.910 ;
        RECT 135.540 219.870 146.330 219.880 ;
        RECT 133.830 219.860 146.330 219.870 ;
        RECT 128.280 219.510 146.330 219.860 ;
        RECT 128.280 219.500 135.610 219.510 ;
        RECT 128.280 219.490 133.900 219.500 ;
        RECT 128.280 219.020 128.790 219.490 ;
        RECT 136.100 219.470 146.330 219.510 ;
        RECT 112.730 214.840 113.720 215.240 ;
        RECT 112.730 214.820 113.310 214.840 ;
        RECT 36.960 207.870 37.450 208.180 ;
        RECT 30.280 207.670 37.450 207.870 ;
        RECT 26.740 207.650 37.450 207.670 ;
        RECT 13.910 207.630 23.180 207.640 ;
        RECT 25.410 207.630 37.450 207.650 ;
        RECT 11.080 207.110 37.450 207.630 ;
        RECT 11.080 207.100 25.490 207.110 ;
        RECT 11.080 207.090 13.920 207.100 ;
        RECT 23.130 207.090 25.490 207.100 ;
        RECT 26.740 207.090 37.450 207.110 ;
        RECT 11.690 201.010 12.240 207.090 ;
        RECT 26.740 207.070 30.560 207.090 ;
        RECT 26.800 205.280 27.290 207.070 ;
        RECT 26.800 204.790 27.310 205.280 ;
        RECT 53.490 202.400 53.940 209.890 ;
        RECT 138.270 207.990 138.780 219.470 ;
        RECT 143.000 219.430 146.330 219.470 ;
        RECT 145.860 213.680 146.300 219.430 ;
        RECT 145.850 213.060 146.300 213.680 ;
        RECT 154.800 209.700 155.240 227.750 ;
        RECT 163.410 227.080 163.790 227.750 ;
        RECT 250.610 221.990 259.880 222.000 ;
        RECT 262.110 221.990 264.020 222.010 ;
        RECT 247.780 221.470 264.020 221.990 ;
        RECT 247.780 221.460 262.190 221.470 ;
        RECT 247.780 221.450 250.620 221.460 ;
        RECT 259.830 221.450 262.190 221.460 ;
        RECT 248.390 215.370 248.940 221.450 ;
        RECT 263.500 219.990 263.990 221.470 ;
        RECT 273.590 220.170 273.980 227.880 ;
        RECT 273.490 220.040 274.000 220.170 ;
        RECT 278.220 220.040 281.550 220.060 ;
        RECT 271.320 220.010 281.550 220.040 ;
        RECT 270.760 220.000 281.550 220.010 ;
        RECT 269.050 219.990 281.550 220.000 ;
        RECT 263.500 219.640 281.550 219.990 ;
        RECT 263.500 219.630 270.830 219.640 ;
        RECT 263.500 219.620 269.120 219.630 ;
        RECT 263.500 219.150 264.010 219.620 ;
        RECT 271.320 219.600 281.550 219.640 ;
        RECT 247.950 214.970 248.940 215.370 ;
        RECT 247.950 214.950 248.530 214.970 ;
        RECT 138.270 207.680 138.760 207.990 ;
        RECT 131.590 207.480 138.760 207.680 ;
        RECT 128.050 207.460 138.760 207.480 ;
        RECT 115.220 207.440 124.490 207.450 ;
        RECT 126.720 207.440 138.760 207.460 ;
        RECT 112.390 206.920 138.760 207.440 ;
        RECT 112.390 206.910 126.800 206.920 ;
        RECT 112.390 206.900 115.230 206.910 ;
        RECT 124.440 206.900 126.800 206.910 ;
        RECT 128.050 206.900 138.760 206.920 ;
        RECT 76.310 202.400 76.890 202.420 ;
        RECT 53.470 201.840 76.890 202.400 ;
        RECT 11.250 200.610 12.240 201.010 ;
        RECT 11.250 200.590 11.830 200.610 ;
        RECT 13.760 192.200 23.030 192.210 ;
        RECT 25.260 192.200 27.170 192.220 ;
        RECT 10.930 191.680 27.170 192.200 ;
        RECT 10.930 191.670 25.340 191.680 ;
        RECT 10.930 191.660 13.770 191.670 ;
        RECT 22.980 191.660 25.340 191.670 ;
        RECT 11.540 185.580 12.090 191.660 ;
        RECT 26.650 190.200 27.140 191.680 ;
        RECT 36.640 190.250 37.150 190.380 ;
        RECT 41.370 190.250 44.700 190.270 ;
        RECT 34.470 190.220 44.700 190.250 ;
        RECT 33.910 190.210 44.700 190.220 ;
        RECT 32.200 190.200 44.700 190.210 ;
        RECT 26.650 189.850 44.700 190.200 ;
        RECT 26.650 189.840 33.980 189.850 ;
        RECT 26.650 189.830 32.270 189.840 ;
        RECT 26.650 189.360 27.160 189.830 ;
        RECT 34.470 189.810 44.700 189.850 ;
        RECT 11.100 185.180 12.090 185.580 ;
        RECT 11.100 185.160 11.680 185.180 ;
        RECT 36.640 178.330 37.150 189.810 ;
        RECT 41.370 189.770 44.700 189.810 ;
        RECT 44.230 184.020 44.670 189.770 ;
        RECT 44.220 183.400 44.670 184.020 ;
        RECT 36.640 178.020 37.130 178.330 ;
        RECT 29.960 177.820 37.130 178.020 ;
        RECT 26.420 177.800 37.130 177.820 ;
        RECT 13.590 177.780 22.860 177.790 ;
        RECT 25.090 177.780 37.130 177.800 ;
        RECT 10.760 177.260 37.130 177.780 ;
        RECT 10.760 177.250 25.170 177.260 ;
        RECT 10.760 177.240 13.600 177.250 ;
        RECT 22.810 177.240 25.170 177.250 ;
        RECT 26.420 177.240 37.130 177.260 ;
        RECT 11.370 171.160 11.920 177.240 ;
        RECT 26.420 177.220 30.240 177.240 ;
        RECT 26.480 175.430 26.970 177.220 ;
        RECT 26.480 174.940 26.990 175.430 ;
        RECT 10.930 170.760 11.920 171.160 ;
        RECT 10.930 170.740 11.510 170.760 ;
        RECT 36.710 168.410 37.100 177.240 ;
        RECT 53.490 168.410 53.940 201.840 ;
        RECT 76.310 200.980 76.890 201.840 ;
        RECT 113.000 200.820 113.550 206.900 ;
        RECT 128.050 206.880 131.870 206.900 ;
        RECT 128.110 205.090 128.600 206.880 ;
        RECT 128.110 204.600 128.620 205.090 ;
        RECT 154.800 202.210 155.250 209.700 ;
        RECT 273.490 208.120 274.000 219.600 ;
        RECT 278.220 219.560 281.550 219.600 ;
        RECT 281.080 213.810 281.520 219.560 ;
        RECT 281.070 213.190 281.520 213.810 ;
        RECT 290.020 209.830 290.460 227.880 ;
        RECT 298.630 227.210 299.010 227.880 ;
        RECT 374.790 227.690 400.320 228.080 ;
        RECT 351.920 221.800 361.190 221.810 ;
        RECT 363.420 221.800 365.330 221.820 ;
        RECT 349.090 221.280 365.330 221.800 ;
        RECT 349.090 221.270 363.500 221.280 ;
        RECT 349.090 221.260 351.930 221.270 ;
        RECT 361.140 221.260 363.500 221.270 ;
        RECT 349.700 215.180 350.250 221.260 ;
        RECT 364.810 219.800 365.300 221.280 ;
        RECT 374.900 219.980 375.290 227.690 ;
        RECT 374.800 219.850 375.310 219.980 ;
        RECT 379.530 219.850 382.860 219.870 ;
        RECT 372.630 219.820 382.860 219.850 ;
        RECT 372.070 219.810 382.860 219.820 ;
        RECT 370.360 219.800 382.860 219.810 ;
        RECT 364.810 219.450 382.860 219.800 ;
        RECT 364.810 219.440 372.140 219.450 ;
        RECT 364.810 219.430 370.430 219.440 ;
        RECT 364.810 218.960 365.320 219.430 ;
        RECT 372.630 219.410 382.860 219.450 ;
        RECT 349.260 214.780 350.250 215.180 ;
        RECT 349.260 214.760 349.840 214.780 ;
        RECT 273.490 207.810 273.980 208.120 ;
        RECT 266.810 207.610 273.980 207.810 ;
        RECT 263.270 207.590 273.980 207.610 ;
        RECT 250.440 207.570 259.710 207.580 ;
        RECT 261.940 207.570 273.980 207.590 ;
        RECT 247.610 207.050 273.980 207.570 ;
        RECT 247.610 207.040 262.020 207.050 ;
        RECT 247.610 207.030 250.450 207.040 ;
        RECT 259.660 207.030 262.020 207.040 ;
        RECT 263.270 207.030 273.980 207.050 ;
        RECT 177.620 202.210 178.200 202.230 ;
        RECT 154.780 201.650 178.200 202.210 ;
        RECT 112.560 200.420 113.550 200.820 ;
        RECT 112.560 200.400 113.140 200.420 ;
        RECT 115.070 192.010 124.340 192.020 ;
        RECT 126.570 192.010 128.480 192.030 ;
        RECT 112.240 191.490 128.480 192.010 ;
        RECT 112.240 191.480 126.650 191.490 ;
        RECT 112.240 191.470 115.080 191.480 ;
        RECT 124.290 191.470 126.650 191.480 ;
        RECT 112.850 185.390 113.400 191.470 ;
        RECT 127.960 190.010 128.450 191.490 ;
        RECT 137.950 190.060 138.460 190.190 ;
        RECT 142.680 190.060 146.010 190.080 ;
        RECT 135.780 190.030 146.010 190.060 ;
        RECT 135.220 190.020 146.010 190.030 ;
        RECT 133.510 190.010 146.010 190.020 ;
        RECT 127.960 189.660 146.010 190.010 ;
        RECT 127.960 189.650 135.290 189.660 ;
        RECT 127.960 189.640 133.580 189.650 ;
        RECT 127.960 189.170 128.470 189.640 ;
        RECT 135.780 189.620 146.010 189.660 ;
        RECT 112.410 184.990 113.400 185.390 ;
        RECT 112.410 184.970 112.990 184.990 ;
        RECT 137.950 178.140 138.460 189.620 ;
        RECT 142.680 189.580 146.010 189.620 ;
        RECT 145.540 183.830 145.980 189.580 ;
        RECT 145.530 183.210 145.980 183.830 ;
        RECT 137.950 177.830 138.440 178.140 ;
        RECT 131.270 177.630 138.440 177.830 ;
        RECT 127.730 177.610 138.440 177.630 ;
        RECT 114.900 177.590 124.170 177.600 ;
        RECT 126.400 177.590 138.440 177.610 ;
        RECT 112.070 177.070 138.440 177.590 ;
        RECT 112.070 177.060 126.480 177.070 ;
        RECT 112.070 177.050 114.910 177.060 ;
        RECT 124.120 177.050 126.480 177.060 ;
        RECT 127.730 177.050 138.440 177.070 ;
        RECT 112.680 170.970 113.230 177.050 ;
        RECT 127.730 177.030 131.550 177.050 ;
        RECT 127.790 175.240 128.280 177.030 ;
        RECT 127.790 174.750 128.300 175.240 ;
        RECT 112.240 170.570 113.230 170.970 ;
        RECT 112.240 170.550 112.820 170.570 ;
        RECT 89.680 168.540 93.040 168.550 ;
        RECT 85.430 168.530 93.040 168.540 ;
        RECT 81.930 168.510 93.040 168.530 ;
        RECT 78.090 168.500 93.040 168.510 ;
        RECT 69.820 168.460 93.040 168.500 ;
        RECT 65.730 168.430 93.040 168.460 ;
        RECT 61.690 168.410 93.040 168.430 ;
        RECT 36.600 168.190 93.040 168.410 ;
        RECT 138.020 168.220 138.410 177.050 ;
        RECT 154.800 168.220 155.250 201.650 ;
        RECT 177.620 200.790 178.200 201.650 ;
        RECT 248.220 200.950 248.770 207.030 ;
        RECT 263.270 207.010 267.090 207.030 ;
        RECT 263.330 205.220 263.820 207.010 ;
        RECT 263.330 204.730 263.840 205.220 ;
        RECT 290.020 202.340 290.470 209.830 ;
        RECT 374.800 207.930 375.310 219.410 ;
        RECT 379.530 219.370 382.860 219.410 ;
        RECT 382.390 213.620 382.830 219.370 ;
        RECT 382.380 213.000 382.830 213.620 ;
        RECT 391.330 209.640 391.770 227.690 ;
        RECT 399.940 227.020 400.320 227.690 ;
        RECT 374.800 207.620 375.290 207.930 ;
        RECT 368.120 207.420 375.290 207.620 ;
        RECT 364.580 207.400 375.290 207.420 ;
        RECT 351.750 207.380 361.020 207.390 ;
        RECT 363.250 207.380 375.290 207.400 ;
        RECT 348.920 206.860 375.290 207.380 ;
        RECT 348.920 206.850 363.330 206.860 ;
        RECT 348.920 206.840 351.760 206.850 ;
        RECT 360.970 206.840 363.330 206.850 ;
        RECT 364.580 206.840 375.290 206.860 ;
        RECT 312.840 202.340 313.420 202.360 ;
        RECT 290.000 201.780 313.420 202.340 ;
        RECT 247.780 200.550 248.770 200.950 ;
        RECT 247.780 200.530 248.360 200.550 ;
        RECT 250.290 192.140 259.560 192.150 ;
        RECT 261.790 192.140 263.700 192.160 ;
        RECT 247.460 191.620 263.700 192.140 ;
        RECT 247.460 191.610 261.870 191.620 ;
        RECT 247.460 191.600 250.300 191.610 ;
        RECT 259.510 191.600 261.870 191.610 ;
        RECT 248.070 185.520 248.620 191.600 ;
        RECT 263.180 190.140 263.670 191.620 ;
        RECT 273.170 190.190 273.680 190.320 ;
        RECT 277.900 190.190 281.230 190.210 ;
        RECT 271.000 190.160 281.230 190.190 ;
        RECT 270.440 190.150 281.230 190.160 ;
        RECT 268.730 190.140 281.230 190.150 ;
        RECT 263.180 189.790 281.230 190.140 ;
        RECT 263.180 189.780 270.510 189.790 ;
        RECT 263.180 189.770 268.800 189.780 ;
        RECT 263.180 189.300 263.690 189.770 ;
        RECT 271.000 189.750 281.230 189.790 ;
        RECT 247.630 185.120 248.620 185.520 ;
        RECT 247.630 185.100 248.210 185.120 ;
        RECT 273.170 178.270 273.680 189.750 ;
        RECT 277.900 189.710 281.230 189.750 ;
        RECT 280.760 183.960 281.200 189.710 ;
        RECT 280.750 183.340 281.200 183.960 ;
        RECT 273.170 177.960 273.660 178.270 ;
        RECT 266.490 177.760 273.660 177.960 ;
        RECT 262.950 177.740 273.660 177.760 ;
        RECT 250.120 177.720 259.390 177.730 ;
        RECT 261.620 177.720 273.660 177.740 ;
        RECT 247.290 177.200 273.660 177.720 ;
        RECT 247.290 177.190 261.700 177.200 ;
        RECT 247.290 177.180 250.130 177.190 ;
        RECT 259.340 177.180 261.700 177.190 ;
        RECT 262.950 177.180 273.660 177.200 ;
        RECT 247.900 171.100 248.450 177.180 ;
        RECT 262.950 177.160 266.770 177.180 ;
        RECT 263.010 175.370 263.500 177.160 ;
        RECT 263.010 174.880 263.520 175.370 ;
        RECT 247.460 170.700 248.450 171.100 ;
        RECT 247.460 170.680 248.040 170.700 ;
        RECT 190.990 168.350 194.350 168.360 ;
        RECT 273.240 168.350 273.630 177.180 ;
        RECT 290.020 168.350 290.470 201.780 ;
        RECT 312.840 200.920 313.420 201.780 ;
        RECT 349.530 200.760 350.080 206.840 ;
        RECT 364.580 206.820 368.400 206.840 ;
        RECT 364.640 205.030 365.130 206.820 ;
        RECT 364.640 204.540 365.150 205.030 ;
        RECT 391.330 202.150 391.780 209.640 ;
        RECT 414.150 202.150 414.730 202.170 ;
        RECT 391.310 201.590 414.730 202.150 ;
        RECT 349.090 200.360 350.080 200.760 ;
        RECT 349.090 200.340 349.670 200.360 ;
        RECT 351.600 191.950 360.870 191.960 ;
        RECT 363.100 191.950 365.010 191.970 ;
        RECT 348.770 191.430 365.010 191.950 ;
        RECT 348.770 191.420 363.180 191.430 ;
        RECT 348.770 191.410 351.610 191.420 ;
        RECT 360.820 191.410 363.180 191.420 ;
        RECT 349.380 185.330 349.930 191.410 ;
        RECT 364.490 189.950 364.980 191.430 ;
        RECT 374.480 190.000 374.990 190.130 ;
        RECT 379.210 190.000 382.540 190.020 ;
        RECT 372.310 189.970 382.540 190.000 ;
        RECT 371.750 189.960 382.540 189.970 ;
        RECT 370.040 189.950 382.540 189.960 ;
        RECT 364.490 189.600 382.540 189.950 ;
        RECT 364.490 189.590 371.820 189.600 ;
        RECT 364.490 189.580 370.110 189.590 ;
        RECT 364.490 189.110 365.000 189.580 ;
        RECT 372.310 189.560 382.540 189.600 ;
        RECT 348.940 184.930 349.930 185.330 ;
        RECT 348.940 184.910 349.520 184.930 ;
        RECT 374.480 178.080 374.990 189.560 ;
        RECT 379.210 189.520 382.540 189.560 ;
        RECT 382.070 183.770 382.510 189.520 ;
        RECT 382.060 183.150 382.510 183.770 ;
        RECT 374.480 177.770 374.970 178.080 ;
        RECT 367.800 177.570 374.970 177.770 ;
        RECT 364.260 177.550 374.970 177.570 ;
        RECT 351.430 177.530 360.700 177.540 ;
        RECT 362.930 177.530 374.970 177.550 ;
        RECT 348.600 177.010 374.970 177.530 ;
        RECT 348.600 177.000 363.010 177.010 ;
        RECT 348.600 176.990 351.440 177.000 ;
        RECT 360.650 176.990 363.010 177.000 ;
        RECT 364.260 176.990 374.970 177.010 ;
        RECT 349.210 170.910 349.760 176.990 ;
        RECT 364.260 176.970 368.080 176.990 ;
        RECT 364.320 175.180 364.810 176.970 ;
        RECT 364.320 174.690 364.830 175.180 ;
        RECT 348.770 170.510 349.760 170.910 ;
        RECT 348.770 170.490 349.350 170.510 ;
        RECT 326.210 168.480 329.570 168.490 ;
        RECT 321.960 168.470 329.570 168.480 ;
        RECT 318.460 168.450 329.570 168.470 ;
        RECT 314.620 168.440 329.570 168.450 ;
        RECT 306.350 168.400 329.570 168.440 ;
        RECT 302.260 168.370 329.570 168.400 ;
        RECT 298.220 168.350 329.570 168.370 ;
        RECT 186.740 168.340 194.350 168.350 ;
        RECT 183.240 168.320 194.350 168.340 ;
        RECT 179.400 168.310 194.350 168.320 ;
        RECT 171.130 168.270 194.350 168.310 ;
        RECT 167.040 168.240 194.350 168.270 ;
        RECT 163.000 168.220 194.350 168.240 ;
        RECT 36.600 168.180 86.380 168.190 ;
        RECT 36.600 168.160 82.540 168.180 ;
        RECT 36.600 168.150 78.340 168.160 ;
        RECT 36.600 168.110 70.180 168.150 ;
        RECT 36.600 168.080 66.140 168.110 ;
        RECT 36.600 168.020 62.130 168.080 ;
        RECT 13.730 162.130 23.000 162.140 ;
        RECT 25.230 162.130 27.140 162.150 ;
        RECT 10.900 161.610 27.140 162.130 ;
        RECT 10.900 161.600 25.310 161.610 ;
        RECT 10.900 161.590 13.740 161.600 ;
        RECT 22.950 161.590 25.310 161.600 ;
        RECT 11.510 155.510 12.060 161.590 ;
        RECT 26.620 160.130 27.110 161.610 ;
        RECT 36.710 160.310 37.100 168.020 ;
        RECT 53.490 167.780 53.940 168.020 ;
        RECT 61.750 167.350 62.130 168.020 ;
        RECT 36.610 160.180 37.120 160.310 ;
        RECT 41.340 160.180 44.670 160.200 ;
        RECT 34.440 160.150 44.670 160.180 ;
        RECT 33.880 160.140 44.670 160.150 ;
        RECT 32.170 160.130 44.670 160.140 ;
        RECT 26.620 159.780 44.670 160.130 ;
        RECT 26.620 159.770 33.950 159.780 ;
        RECT 26.620 159.760 32.240 159.770 ;
        RECT 26.620 159.290 27.130 159.760 ;
        RECT 34.440 159.740 44.670 159.780 ;
        RECT 11.070 155.110 12.060 155.510 ;
        RECT 11.070 155.090 11.650 155.110 ;
        RECT 36.610 148.260 37.120 159.740 ;
        RECT 41.340 159.700 44.670 159.740 ;
        RECT 44.200 153.950 44.640 159.700 ;
        RECT 44.190 153.330 44.640 153.950 ;
        RECT 92.630 150.270 93.040 168.190 ;
        RECT 137.910 168.000 194.350 168.220 ;
        RECT 137.910 167.990 187.690 168.000 ;
        RECT 137.910 167.970 183.850 167.990 ;
        RECT 137.910 167.960 179.650 167.970 ;
        RECT 137.910 167.920 171.490 167.960 ;
        RECT 137.910 167.890 167.450 167.920 ;
        RECT 137.910 167.830 163.440 167.890 ;
        RECT 115.040 161.940 124.310 161.950 ;
        RECT 126.540 161.940 128.450 161.960 ;
        RECT 112.210 161.420 128.450 161.940 ;
        RECT 112.210 161.410 126.620 161.420 ;
        RECT 112.210 161.400 115.050 161.410 ;
        RECT 124.260 161.400 126.620 161.410 ;
        RECT 112.820 155.320 113.370 161.400 ;
        RECT 127.930 159.940 128.420 161.420 ;
        RECT 138.020 160.120 138.410 167.830 ;
        RECT 154.800 167.590 155.250 167.830 ;
        RECT 163.060 167.160 163.440 167.830 ;
        RECT 137.920 159.990 138.430 160.120 ;
        RECT 142.650 159.990 145.980 160.010 ;
        RECT 135.750 159.960 145.980 159.990 ;
        RECT 135.190 159.950 145.980 159.960 ;
        RECT 133.480 159.940 145.980 159.950 ;
        RECT 127.930 159.590 145.980 159.940 ;
        RECT 127.930 159.580 135.260 159.590 ;
        RECT 127.930 159.570 133.550 159.580 ;
        RECT 127.930 159.100 128.440 159.570 ;
        RECT 135.750 159.550 145.980 159.590 ;
        RECT 112.380 154.920 113.370 155.320 ;
        RECT 112.380 154.900 112.960 154.920 ;
        RECT 92.630 149.920 93.060 150.270 ;
        RECT 36.610 147.950 37.100 148.260 ;
        RECT 29.930 147.750 37.100 147.950 ;
        RECT 26.390 147.730 37.100 147.750 ;
        RECT 13.560 147.710 22.830 147.720 ;
        RECT 25.060 147.710 37.100 147.730 ;
        RECT 10.730 147.190 37.100 147.710 ;
        RECT 10.730 147.180 25.140 147.190 ;
        RECT 10.730 147.170 13.570 147.180 ;
        RECT 22.780 147.170 25.140 147.180 ;
        RECT 26.390 147.170 37.100 147.190 ;
        RECT 11.340 141.090 11.890 147.170 ;
        RECT 26.390 147.150 30.210 147.170 ;
        RECT 26.450 145.360 26.940 147.150 ;
        RECT 92.630 145.630 93.100 149.920 ;
        RECT 137.920 148.070 138.430 159.550 ;
        RECT 142.650 159.510 145.980 159.550 ;
        RECT 145.510 153.760 145.950 159.510 ;
        RECT 145.500 153.140 145.950 153.760 ;
        RECT 193.940 150.080 194.350 168.000 ;
        RECT 273.130 168.130 329.570 168.350 ;
        RECT 374.550 168.160 374.940 176.990 ;
        RECT 391.330 168.160 391.780 201.590 ;
        RECT 414.150 200.730 414.730 201.590 ;
        RECT 427.520 168.290 430.880 168.300 ;
        RECT 423.270 168.280 430.880 168.290 ;
        RECT 419.770 168.260 430.880 168.280 ;
        RECT 415.930 168.250 430.880 168.260 ;
        RECT 407.660 168.210 430.880 168.250 ;
        RECT 403.570 168.180 430.880 168.210 ;
        RECT 399.530 168.160 430.880 168.180 ;
        RECT 273.130 168.120 322.910 168.130 ;
        RECT 273.130 168.100 319.070 168.120 ;
        RECT 273.130 168.090 314.870 168.100 ;
        RECT 273.130 168.050 306.710 168.090 ;
        RECT 273.130 168.020 302.670 168.050 ;
        RECT 273.130 167.960 298.660 168.020 ;
        RECT 250.260 162.070 259.530 162.080 ;
        RECT 261.760 162.070 263.670 162.090 ;
        RECT 247.430 161.550 263.670 162.070 ;
        RECT 247.430 161.540 261.840 161.550 ;
        RECT 247.430 161.530 250.270 161.540 ;
        RECT 259.480 161.530 261.840 161.540 ;
        RECT 248.040 155.450 248.590 161.530 ;
        RECT 263.150 160.070 263.640 161.550 ;
        RECT 273.240 160.250 273.630 167.960 ;
        RECT 290.020 167.720 290.470 167.960 ;
        RECT 298.280 167.290 298.660 167.960 ;
        RECT 273.140 160.120 273.650 160.250 ;
        RECT 277.870 160.120 281.200 160.140 ;
        RECT 270.970 160.090 281.200 160.120 ;
        RECT 270.410 160.080 281.200 160.090 ;
        RECT 268.700 160.070 281.200 160.080 ;
        RECT 263.150 159.720 281.200 160.070 ;
        RECT 263.150 159.710 270.480 159.720 ;
        RECT 263.150 159.700 268.770 159.710 ;
        RECT 263.150 159.230 263.660 159.700 ;
        RECT 270.970 159.680 281.200 159.720 ;
        RECT 247.600 155.050 248.590 155.450 ;
        RECT 247.600 155.030 248.180 155.050 ;
        RECT 193.940 149.730 194.370 150.080 ;
        RECT 137.920 147.760 138.410 148.070 ;
        RECT 131.240 147.560 138.410 147.760 ;
        RECT 127.700 147.540 138.410 147.560 ;
        RECT 114.870 147.520 124.140 147.530 ;
        RECT 126.370 147.520 138.410 147.540 ;
        RECT 112.040 147.000 138.410 147.520 ;
        RECT 112.040 146.990 126.450 147.000 ;
        RECT 112.040 146.980 114.880 146.990 ;
        RECT 124.090 146.980 126.450 146.990 ;
        RECT 127.700 146.980 138.410 147.000 ;
        RECT 26.450 144.870 26.960 145.360 ;
        RECT 92.640 143.710 93.100 145.630 ;
        RECT 92.340 143.680 93.100 143.710 ;
        RECT 75.820 143.420 93.100 143.680 ;
        RECT 10.900 140.690 11.890 141.090 ;
        RECT 75.780 143.280 93.100 143.420 ;
        RECT 10.900 140.670 11.480 140.690 ;
        RECT 13.610 131.880 22.880 131.890 ;
        RECT 25.110 131.880 27.020 131.900 ;
        RECT 10.780 131.360 27.020 131.880 ;
        RECT 10.780 131.350 25.190 131.360 ;
        RECT 10.780 131.340 13.620 131.350 ;
        RECT 22.830 131.340 25.190 131.350 ;
        RECT 11.390 125.260 11.940 131.340 ;
        RECT 26.500 129.880 26.990 131.360 ;
        RECT 36.490 129.930 37.000 130.060 ;
        RECT 41.220 129.930 44.550 129.950 ;
        RECT 34.320 129.900 44.550 129.930 ;
        RECT 33.760 129.890 44.550 129.900 ;
        RECT 32.050 129.880 44.550 129.890 ;
        RECT 26.500 129.530 44.550 129.880 ;
        RECT 26.500 129.520 33.830 129.530 ;
        RECT 26.500 129.510 32.120 129.520 ;
        RECT 26.500 129.040 27.010 129.510 ;
        RECT 34.320 129.490 44.550 129.530 ;
        RECT 10.950 124.860 11.940 125.260 ;
        RECT 10.950 124.840 11.530 124.860 ;
        RECT 36.490 118.010 37.000 129.490 ;
        RECT 41.220 129.450 44.550 129.490 ;
        RECT 44.080 123.700 44.520 129.450 ;
        RECT 44.070 123.080 44.520 123.700 ;
        RECT 36.490 117.700 36.980 118.010 ;
        RECT 29.810 117.500 36.980 117.700 ;
        RECT 26.270 117.480 36.980 117.500 ;
        RECT 13.440 117.460 22.710 117.470 ;
        RECT 24.940 117.460 36.980 117.480 ;
        RECT 10.610 116.940 36.980 117.460 ;
        RECT 10.610 116.930 25.020 116.940 ;
        RECT 10.610 116.920 13.450 116.930 ;
        RECT 22.660 116.920 25.020 116.930 ;
        RECT 26.270 116.920 36.980 116.940 ;
        RECT 11.220 110.840 11.770 116.920 ;
        RECT 26.270 116.900 30.090 116.920 ;
        RECT 26.330 115.110 26.820 116.900 ;
        RECT 26.330 114.620 26.840 115.110 ;
        RECT 10.780 110.440 11.770 110.840 ;
        RECT 10.780 110.420 11.360 110.440 ;
        RECT 36.560 108.090 36.950 116.920 ;
        RECT 52.990 108.090 53.430 108.100 ;
        RECT 36.450 107.700 61.980 108.090 ;
        RECT 13.580 101.810 22.850 101.820 ;
        RECT 25.080 101.810 26.990 101.830 ;
        RECT 10.750 101.290 26.990 101.810 ;
        RECT 10.750 101.280 25.160 101.290 ;
        RECT 10.750 101.270 13.590 101.280 ;
        RECT 22.800 101.270 25.160 101.280 ;
        RECT 11.360 95.190 11.910 101.270 ;
        RECT 26.470 99.810 26.960 101.290 ;
        RECT 36.560 99.990 36.950 107.700 ;
        RECT 36.460 99.860 36.970 99.990 ;
        RECT 41.190 99.860 44.520 99.880 ;
        RECT 34.290 99.830 44.520 99.860 ;
        RECT 33.730 99.820 44.520 99.830 ;
        RECT 32.020 99.810 44.520 99.820 ;
        RECT 26.470 99.460 44.520 99.810 ;
        RECT 26.470 99.450 33.800 99.460 ;
        RECT 26.470 99.440 32.090 99.450 ;
        RECT 26.470 98.970 26.980 99.440 ;
        RECT 34.290 99.420 44.520 99.460 ;
        RECT 10.920 94.790 11.910 95.190 ;
        RECT 10.920 94.770 11.500 94.790 ;
        RECT 36.460 87.940 36.970 99.420 ;
        RECT 41.190 99.380 44.520 99.420 ;
        RECT 44.050 93.630 44.490 99.380 ;
        RECT 44.040 93.010 44.490 93.630 ;
        RECT 52.990 89.650 53.430 107.700 ;
        RECT 61.600 107.030 61.980 107.700 ;
        RECT 36.460 87.630 36.950 87.940 ;
        RECT 29.780 87.430 36.950 87.630 ;
        RECT 26.240 87.410 36.950 87.430 ;
        RECT 13.410 87.390 22.680 87.400 ;
        RECT 24.910 87.390 36.950 87.410 ;
        RECT 10.580 86.870 36.950 87.390 ;
        RECT 10.580 86.860 24.990 86.870 ;
        RECT 10.580 86.850 13.420 86.860 ;
        RECT 22.630 86.850 24.990 86.860 ;
        RECT 26.240 86.850 36.950 86.870 ;
        RECT 11.190 80.770 11.740 86.850 ;
        RECT 26.240 86.830 30.060 86.850 ;
        RECT 26.300 85.040 26.790 86.830 ;
        RECT 26.300 84.550 26.810 85.040 ;
        RECT 52.990 82.160 53.440 89.650 ;
        RECT 75.780 86.760 76.310 143.280 ;
        RECT 92.340 143.270 93.100 143.280 ;
        RECT 92.640 142.040 93.100 143.270 ;
        RECT 92.630 141.960 93.100 142.040 ;
        RECT 92.630 138.310 93.090 141.960 ;
        RECT 112.650 140.900 113.200 146.980 ;
        RECT 127.700 146.960 131.520 146.980 ;
        RECT 127.760 145.170 128.250 146.960 ;
        RECT 193.940 145.440 194.410 149.730 ;
        RECT 273.140 148.200 273.650 159.680 ;
        RECT 277.870 159.640 281.200 159.680 ;
        RECT 280.730 153.890 281.170 159.640 ;
        RECT 280.720 153.270 281.170 153.890 ;
        RECT 329.160 150.210 329.570 168.130 ;
        RECT 374.440 167.940 430.880 168.160 ;
        RECT 374.440 167.930 424.220 167.940 ;
        RECT 374.440 167.910 420.380 167.930 ;
        RECT 374.440 167.900 416.180 167.910 ;
        RECT 374.440 167.860 408.020 167.900 ;
        RECT 374.440 167.830 403.980 167.860 ;
        RECT 374.440 167.770 399.970 167.830 ;
        RECT 351.570 161.880 360.840 161.890 ;
        RECT 363.070 161.880 364.980 161.900 ;
        RECT 348.740 161.360 364.980 161.880 ;
        RECT 348.740 161.350 363.150 161.360 ;
        RECT 348.740 161.340 351.580 161.350 ;
        RECT 360.790 161.340 363.150 161.350 ;
        RECT 349.350 155.260 349.900 161.340 ;
        RECT 364.460 159.880 364.950 161.360 ;
        RECT 374.550 160.060 374.940 167.770 ;
        RECT 391.330 167.530 391.780 167.770 ;
        RECT 399.590 167.100 399.970 167.770 ;
        RECT 374.450 159.930 374.960 160.060 ;
        RECT 379.180 159.930 382.510 159.950 ;
        RECT 372.280 159.900 382.510 159.930 ;
        RECT 371.720 159.890 382.510 159.900 ;
        RECT 370.010 159.880 382.510 159.890 ;
        RECT 364.460 159.530 382.510 159.880 ;
        RECT 364.460 159.520 371.790 159.530 ;
        RECT 364.460 159.510 370.080 159.520 ;
        RECT 364.460 159.040 364.970 159.510 ;
        RECT 372.280 159.490 382.510 159.530 ;
        RECT 348.910 154.860 349.900 155.260 ;
        RECT 348.910 154.840 349.490 154.860 ;
        RECT 329.160 149.860 329.590 150.210 ;
        RECT 273.140 147.890 273.630 148.200 ;
        RECT 266.460 147.690 273.630 147.890 ;
        RECT 262.920 147.670 273.630 147.690 ;
        RECT 250.090 147.650 259.360 147.660 ;
        RECT 261.590 147.650 273.630 147.670 ;
        RECT 247.260 147.130 273.630 147.650 ;
        RECT 247.260 147.120 261.670 147.130 ;
        RECT 247.260 147.110 250.100 147.120 ;
        RECT 259.310 147.110 261.670 147.120 ;
        RECT 262.920 147.110 273.630 147.130 ;
        RECT 127.760 144.680 128.270 145.170 ;
        RECT 193.950 143.520 194.410 145.440 ;
        RECT 193.650 143.490 194.410 143.520 ;
        RECT 177.130 143.480 194.410 143.490 ;
        RECT 177.130 143.470 214.450 143.480 ;
        RECT 220.200 143.470 220.680 143.480 ;
        RECT 177.130 143.230 220.680 143.470 ;
        RECT 112.210 140.500 113.200 140.900 ;
        RECT 177.090 143.130 220.680 143.230 ;
        RECT 177.090 143.100 214.450 143.130 ;
        RECT 177.090 143.090 194.410 143.100 ;
        RECT 112.210 140.480 112.790 140.500 ;
        RECT 92.630 137.740 93.080 138.310 ;
        RECT 114.920 131.690 124.190 131.700 ;
        RECT 126.420 131.690 128.330 131.710 ;
        RECT 112.090 131.170 128.330 131.690 ;
        RECT 112.090 131.160 126.500 131.170 ;
        RECT 112.090 131.150 114.930 131.160 ;
        RECT 124.140 131.150 126.500 131.160 ;
        RECT 112.700 125.070 113.250 131.150 ;
        RECT 127.810 129.690 128.300 131.170 ;
        RECT 137.800 129.740 138.310 129.870 ;
        RECT 142.530 129.740 145.860 129.760 ;
        RECT 135.630 129.710 145.860 129.740 ;
        RECT 135.070 129.700 145.860 129.710 ;
        RECT 133.360 129.690 145.860 129.700 ;
        RECT 127.810 129.340 145.860 129.690 ;
        RECT 127.810 129.330 135.140 129.340 ;
        RECT 127.810 129.320 133.430 129.330 ;
        RECT 127.810 128.850 128.320 129.320 ;
        RECT 135.630 129.300 145.860 129.340 ;
        RECT 112.260 124.670 113.250 125.070 ;
        RECT 112.260 124.650 112.840 124.670 ;
        RECT 137.800 117.820 138.310 129.300 ;
        RECT 142.530 129.260 145.860 129.300 ;
        RECT 145.390 123.510 145.830 129.260 ;
        RECT 145.380 122.890 145.830 123.510 ;
        RECT 137.800 117.510 138.290 117.820 ;
        RECT 131.120 117.310 138.290 117.510 ;
        RECT 127.580 117.290 138.290 117.310 ;
        RECT 114.750 117.270 124.020 117.280 ;
        RECT 126.250 117.270 138.290 117.290 ;
        RECT 111.920 116.750 138.290 117.270 ;
        RECT 111.920 116.740 126.330 116.750 ;
        RECT 111.920 116.730 114.760 116.740 ;
        RECT 123.970 116.730 126.330 116.740 ;
        RECT 127.580 116.730 138.290 116.750 ;
        RECT 112.530 110.650 113.080 116.730 ;
        RECT 127.580 116.710 131.400 116.730 ;
        RECT 127.640 114.920 128.130 116.710 ;
        RECT 127.640 114.430 128.150 114.920 ;
        RECT 112.090 110.250 113.080 110.650 ;
        RECT 112.090 110.230 112.670 110.250 ;
        RECT 137.870 107.900 138.260 116.730 ;
        RECT 154.300 107.900 154.740 107.910 ;
        RECT 137.760 107.510 163.290 107.900 ;
        RECT 114.890 101.620 124.160 101.630 ;
        RECT 126.390 101.620 128.300 101.640 ;
        RECT 112.060 101.100 128.300 101.620 ;
        RECT 112.060 101.090 126.470 101.100 ;
        RECT 112.060 101.080 114.900 101.090 ;
        RECT 124.110 101.080 126.470 101.090 ;
        RECT 112.670 95.000 113.220 101.080 ;
        RECT 127.780 99.620 128.270 101.100 ;
        RECT 137.870 99.800 138.260 107.510 ;
        RECT 137.770 99.670 138.280 99.800 ;
        RECT 142.500 99.670 145.830 99.690 ;
        RECT 135.600 99.640 145.830 99.670 ;
        RECT 135.040 99.630 145.830 99.640 ;
        RECT 133.330 99.620 145.830 99.630 ;
        RECT 127.780 99.270 145.830 99.620 ;
        RECT 127.780 99.260 135.110 99.270 ;
        RECT 127.780 99.250 133.400 99.260 ;
        RECT 127.780 98.780 128.290 99.250 ;
        RECT 135.600 99.230 145.830 99.270 ;
        RECT 112.230 94.600 113.220 95.000 ;
        RECT 112.230 94.580 112.810 94.600 ;
        RECT 137.770 87.750 138.280 99.230 ;
        RECT 142.500 99.190 145.830 99.230 ;
        RECT 145.360 93.440 145.800 99.190 ;
        RECT 145.350 92.820 145.800 93.440 ;
        RECT 154.300 89.460 154.740 107.510 ;
        RECT 162.910 106.840 163.290 107.510 ;
        RECT 137.770 87.440 138.260 87.750 ;
        RECT 131.090 87.240 138.260 87.440 ;
        RECT 127.550 87.220 138.260 87.240 ;
        RECT 114.720 87.200 123.990 87.210 ;
        RECT 126.220 87.200 138.260 87.220 ;
        RECT 75.780 86.410 76.400 86.760 ;
        RECT 111.890 86.680 138.260 87.200 ;
        RECT 111.890 86.670 126.300 86.680 ;
        RECT 111.890 86.660 114.730 86.670 ;
        RECT 123.940 86.660 126.300 86.670 ;
        RECT 127.550 86.660 138.260 86.680 ;
        RECT 75.820 82.180 76.400 86.410 ;
        RECT 75.810 82.160 76.400 82.180 ;
        RECT 52.970 81.630 76.400 82.160 ;
        RECT 52.970 81.600 76.390 81.630 ;
        RECT 10.750 80.370 11.740 80.770 ;
        RECT 10.750 80.350 11.330 80.370 ;
        RECT 13.260 71.960 22.530 71.970 ;
        RECT 24.760 71.960 26.670 71.980 ;
        RECT 10.430 71.440 26.670 71.960 ;
        RECT 10.430 71.430 24.840 71.440 ;
        RECT 10.430 71.420 13.270 71.430 ;
        RECT 22.480 71.420 24.840 71.430 ;
        RECT 11.040 65.340 11.590 71.420 ;
        RECT 26.150 69.960 26.640 71.440 ;
        RECT 36.140 70.010 36.650 70.140 ;
        RECT 40.870 70.010 44.200 70.030 ;
        RECT 33.970 69.980 44.200 70.010 ;
        RECT 33.410 69.970 44.200 69.980 ;
        RECT 31.700 69.960 44.200 69.970 ;
        RECT 26.150 69.610 44.200 69.960 ;
        RECT 26.150 69.600 33.480 69.610 ;
        RECT 26.150 69.590 31.770 69.600 ;
        RECT 26.150 69.120 26.660 69.590 ;
        RECT 33.970 69.570 44.200 69.610 ;
        RECT 10.600 64.940 11.590 65.340 ;
        RECT 10.600 64.920 11.180 64.940 ;
        RECT 36.140 58.090 36.650 69.570 ;
        RECT 40.870 69.530 44.200 69.570 ;
        RECT 43.730 63.780 44.170 69.530 ;
        RECT 43.720 63.160 44.170 63.780 ;
        RECT 36.140 57.780 36.630 58.090 ;
        RECT 29.460 57.580 36.630 57.780 ;
        RECT 25.920 57.560 36.630 57.580 ;
        RECT 13.090 57.540 22.360 57.550 ;
        RECT 24.590 57.540 36.630 57.560 ;
        RECT 10.260 57.020 36.630 57.540 ;
        RECT 10.260 57.010 24.670 57.020 ;
        RECT 10.260 57.000 13.100 57.010 ;
        RECT 22.310 57.000 24.670 57.010 ;
        RECT 25.920 57.000 36.630 57.020 ;
        RECT 10.870 50.920 11.420 57.000 ;
        RECT 25.920 56.980 29.740 57.000 ;
        RECT 25.980 55.190 26.470 56.980 ;
        RECT 25.980 54.700 26.490 55.190 ;
        RECT 10.430 50.520 11.420 50.920 ;
        RECT 10.430 50.500 11.010 50.520 ;
        RECT 36.210 48.170 36.600 57.000 ;
        RECT 52.990 48.170 53.440 81.600 ;
        RECT 75.810 80.740 76.390 81.600 ;
        RECT 112.500 80.580 113.050 86.660 ;
        RECT 127.550 86.640 131.370 86.660 ;
        RECT 127.610 84.850 128.100 86.640 ;
        RECT 127.610 84.360 128.120 84.850 ;
        RECT 154.300 81.970 154.750 89.460 ;
        RECT 177.090 86.570 177.620 143.090 ;
        RECT 193.650 143.080 194.410 143.090 ;
        RECT 193.950 141.850 194.410 143.080 ;
        RECT 193.940 141.770 194.410 141.850 ;
        RECT 193.940 138.120 194.400 141.770 ;
        RECT 220.200 140.410 220.680 143.130 ;
        RECT 247.870 141.030 248.420 147.110 ;
        RECT 262.920 147.090 266.740 147.110 ;
        RECT 262.980 145.300 263.470 147.090 ;
        RECT 329.160 145.570 329.630 149.860 ;
        RECT 374.450 148.010 374.960 159.490 ;
        RECT 379.180 159.450 382.510 159.490 ;
        RECT 382.040 153.700 382.480 159.450 ;
        RECT 382.030 153.080 382.480 153.700 ;
        RECT 430.470 150.020 430.880 167.940 ;
        RECT 430.470 149.670 430.900 150.020 ;
        RECT 374.450 147.700 374.940 148.010 ;
        RECT 367.770 147.500 374.940 147.700 ;
        RECT 364.230 147.480 374.940 147.500 ;
        RECT 351.400 147.460 360.670 147.470 ;
        RECT 362.900 147.460 374.940 147.480 ;
        RECT 348.570 146.940 374.940 147.460 ;
        RECT 348.570 146.930 362.980 146.940 ;
        RECT 348.570 146.920 351.410 146.930 ;
        RECT 360.620 146.920 362.980 146.930 ;
        RECT 364.230 146.920 374.940 146.940 ;
        RECT 262.980 144.810 263.490 145.300 ;
        RECT 329.170 143.650 329.630 145.570 ;
        RECT 328.870 143.620 329.630 143.650 ;
        RECT 312.350 143.360 329.630 143.620 ;
        RECT 247.430 140.630 248.420 141.030 ;
        RECT 312.310 143.220 329.630 143.360 ;
        RECT 247.430 140.610 248.010 140.630 ;
        RECT 220.200 140.340 220.710 140.410 ;
        RECT 220.210 139.750 220.710 140.340 ;
        RECT 193.940 137.550 194.390 138.120 ;
        RECT 250.140 131.820 259.410 131.830 ;
        RECT 261.640 131.820 263.550 131.840 ;
        RECT 247.310 131.300 263.550 131.820 ;
        RECT 247.310 131.290 261.720 131.300 ;
        RECT 247.310 131.280 250.150 131.290 ;
        RECT 259.360 131.280 261.720 131.290 ;
        RECT 247.920 125.200 248.470 131.280 ;
        RECT 263.030 129.820 263.520 131.300 ;
        RECT 273.020 129.870 273.530 130.000 ;
        RECT 277.750 129.870 281.080 129.890 ;
        RECT 270.850 129.840 281.080 129.870 ;
        RECT 270.290 129.830 281.080 129.840 ;
        RECT 268.580 129.820 281.080 129.830 ;
        RECT 263.030 129.470 281.080 129.820 ;
        RECT 263.030 129.460 270.360 129.470 ;
        RECT 263.030 129.450 268.650 129.460 ;
        RECT 263.030 128.980 263.540 129.450 ;
        RECT 270.850 129.430 281.080 129.470 ;
        RECT 247.480 124.800 248.470 125.200 ;
        RECT 247.480 124.780 248.060 124.800 ;
        RECT 273.020 117.950 273.530 129.430 ;
        RECT 277.750 129.390 281.080 129.430 ;
        RECT 280.610 123.640 281.050 129.390 ;
        RECT 280.600 123.020 281.050 123.640 ;
        RECT 273.020 117.640 273.510 117.950 ;
        RECT 266.340 117.440 273.510 117.640 ;
        RECT 262.800 117.420 273.510 117.440 ;
        RECT 249.970 117.400 259.240 117.410 ;
        RECT 261.470 117.400 273.510 117.420 ;
        RECT 247.140 116.880 273.510 117.400 ;
        RECT 247.140 116.870 261.550 116.880 ;
        RECT 247.140 116.860 249.980 116.870 ;
        RECT 259.190 116.860 261.550 116.870 ;
        RECT 262.800 116.860 273.510 116.880 ;
        RECT 247.750 110.780 248.300 116.860 ;
        RECT 262.800 116.840 266.620 116.860 ;
        RECT 262.860 115.050 263.350 116.840 ;
        RECT 262.860 114.560 263.370 115.050 ;
        RECT 247.310 110.380 248.300 110.780 ;
        RECT 247.310 110.360 247.890 110.380 ;
        RECT 273.090 108.030 273.480 116.860 ;
        RECT 289.520 108.030 289.960 108.040 ;
        RECT 272.980 107.640 298.510 108.030 ;
        RECT 250.110 101.750 259.380 101.760 ;
        RECT 261.610 101.750 263.520 101.770 ;
        RECT 247.280 101.230 263.520 101.750 ;
        RECT 247.280 101.220 261.690 101.230 ;
        RECT 247.280 101.210 250.120 101.220 ;
        RECT 259.330 101.210 261.690 101.220 ;
        RECT 247.890 95.130 248.440 101.210 ;
        RECT 263.000 99.750 263.490 101.230 ;
        RECT 273.090 99.930 273.480 107.640 ;
        RECT 272.990 99.800 273.500 99.930 ;
        RECT 277.720 99.800 281.050 99.820 ;
        RECT 270.820 99.770 281.050 99.800 ;
        RECT 270.260 99.760 281.050 99.770 ;
        RECT 268.550 99.750 281.050 99.760 ;
        RECT 263.000 99.400 281.050 99.750 ;
        RECT 263.000 99.390 270.330 99.400 ;
        RECT 263.000 99.380 268.620 99.390 ;
        RECT 263.000 98.910 263.510 99.380 ;
        RECT 270.820 99.360 281.050 99.400 ;
        RECT 247.450 94.730 248.440 95.130 ;
        RECT 247.450 94.710 248.030 94.730 ;
        RECT 272.990 87.880 273.500 99.360 ;
        RECT 277.720 99.320 281.050 99.360 ;
        RECT 280.580 93.570 281.020 99.320 ;
        RECT 280.570 92.950 281.020 93.570 ;
        RECT 289.520 89.590 289.960 107.640 ;
        RECT 298.130 106.970 298.510 107.640 ;
        RECT 272.990 87.570 273.480 87.880 ;
        RECT 266.310 87.370 273.480 87.570 ;
        RECT 262.770 87.350 273.480 87.370 ;
        RECT 249.940 87.330 259.210 87.340 ;
        RECT 261.440 87.330 273.480 87.350 ;
        RECT 247.110 86.810 273.480 87.330 ;
        RECT 247.110 86.800 261.520 86.810 ;
        RECT 247.110 86.790 249.950 86.800 ;
        RECT 259.160 86.790 261.520 86.800 ;
        RECT 262.770 86.790 273.480 86.810 ;
        RECT 177.090 86.220 177.710 86.570 ;
        RECT 177.130 81.990 177.710 86.220 ;
        RECT 177.120 81.970 177.710 81.990 ;
        RECT 154.280 81.440 177.710 81.970 ;
        RECT 154.280 81.410 177.700 81.440 ;
        RECT 112.060 80.180 113.050 80.580 ;
        RECT 112.060 80.160 112.640 80.180 ;
        RECT 114.570 71.770 123.840 71.780 ;
        RECT 126.070 71.770 127.980 71.790 ;
        RECT 111.740 71.250 127.980 71.770 ;
        RECT 111.740 71.240 126.150 71.250 ;
        RECT 111.740 71.230 114.580 71.240 ;
        RECT 123.790 71.230 126.150 71.240 ;
        RECT 112.350 65.150 112.900 71.230 ;
        RECT 127.460 69.770 127.950 71.250 ;
        RECT 137.450 69.820 137.960 69.950 ;
        RECT 142.180 69.820 145.510 69.840 ;
        RECT 135.280 69.790 145.510 69.820 ;
        RECT 134.720 69.780 145.510 69.790 ;
        RECT 133.010 69.770 145.510 69.780 ;
        RECT 127.460 69.420 145.510 69.770 ;
        RECT 127.460 69.410 134.790 69.420 ;
        RECT 127.460 69.400 133.080 69.410 ;
        RECT 127.460 68.930 127.970 69.400 ;
        RECT 135.280 69.380 145.510 69.420 ;
        RECT 111.910 64.750 112.900 65.150 ;
        RECT 111.910 64.730 112.490 64.750 ;
        RECT 137.450 57.900 137.960 69.380 ;
        RECT 142.180 69.340 145.510 69.380 ;
        RECT 145.040 63.590 145.480 69.340 ;
        RECT 145.030 62.970 145.480 63.590 ;
        RECT 137.450 57.590 137.940 57.900 ;
        RECT 130.770 57.390 137.940 57.590 ;
        RECT 127.230 57.370 137.940 57.390 ;
        RECT 114.400 57.350 123.670 57.360 ;
        RECT 125.900 57.350 137.940 57.370 ;
        RECT 111.570 56.830 137.940 57.350 ;
        RECT 111.570 56.820 125.980 56.830 ;
        RECT 111.570 56.810 114.410 56.820 ;
        RECT 123.620 56.810 125.980 56.820 ;
        RECT 127.230 56.810 137.940 56.830 ;
        RECT 112.180 50.730 112.730 56.810 ;
        RECT 127.230 56.790 131.050 56.810 ;
        RECT 127.290 55.000 127.780 56.790 ;
        RECT 127.290 54.510 127.800 55.000 ;
        RECT 111.740 50.330 112.730 50.730 ;
        RECT 111.740 50.310 112.320 50.330 ;
        RECT 36.100 47.780 61.630 48.170 ;
        RECT 137.520 47.980 137.910 56.810 ;
        RECT 154.300 47.980 154.750 81.410 ;
        RECT 177.120 80.550 177.700 81.410 ;
        RECT 247.720 80.710 248.270 86.790 ;
        RECT 262.770 86.770 266.590 86.790 ;
        RECT 262.830 84.980 263.320 86.770 ;
        RECT 262.830 84.490 263.340 84.980 ;
        RECT 289.520 82.100 289.970 89.590 ;
        RECT 312.310 86.700 312.840 143.220 ;
        RECT 328.870 143.210 329.630 143.220 ;
        RECT 329.170 141.980 329.630 143.210 ;
        RECT 329.160 141.900 329.630 141.980 ;
        RECT 329.160 138.250 329.620 141.900 ;
        RECT 349.180 140.840 349.730 146.920 ;
        RECT 364.230 146.900 368.050 146.920 ;
        RECT 364.290 145.110 364.780 146.900 ;
        RECT 430.470 145.380 430.940 149.670 ;
        RECT 364.290 144.620 364.800 145.110 ;
        RECT 430.480 143.460 430.940 145.380 ;
        RECT 430.180 143.430 430.940 143.460 ;
        RECT 413.660 143.420 430.940 143.430 ;
        RECT 413.660 143.410 450.980 143.420 ;
        RECT 456.730 143.410 457.210 143.420 ;
        RECT 413.660 143.170 457.210 143.410 ;
        RECT 348.740 140.440 349.730 140.840 ;
        RECT 413.620 143.070 457.210 143.170 ;
        RECT 413.620 143.040 450.980 143.070 ;
        RECT 413.620 143.030 430.940 143.040 ;
        RECT 348.740 140.420 349.320 140.440 ;
        RECT 329.160 137.680 329.610 138.250 ;
        RECT 351.450 131.630 360.720 131.640 ;
        RECT 362.950 131.630 364.860 131.650 ;
        RECT 348.620 131.110 364.860 131.630 ;
        RECT 348.620 131.100 363.030 131.110 ;
        RECT 348.620 131.090 351.460 131.100 ;
        RECT 360.670 131.090 363.030 131.100 ;
        RECT 349.230 125.010 349.780 131.090 ;
        RECT 364.340 129.630 364.830 131.110 ;
        RECT 374.330 129.680 374.840 129.810 ;
        RECT 379.060 129.680 382.390 129.700 ;
        RECT 372.160 129.650 382.390 129.680 ;
        RECT 371.600 129.640 382.390 129.650 ;
        RECT 369.890 129.630 382.390 129.640 ;
        RECT 364.340 129.280 382.390 129.630 ;
        RECT 364.340 129.270 371.670 129.280 ;
        RECT 364.340 129.260 369.960 129.270 ;
        RECT 364.340 128.790 364.850 129.260 ;
        RECT 372.160 129.240 382.390 129.280 ;
        RECT 348.790 124.610 349.780 125.010 ;
        RECT 348.790 124.590 349.370 124.610 ;
        RECT 374.330 117.760 374.840 129.240 ;
        RECT 379.060 129.200 382.390 129.240 ;
        RECT 381.920 123.450 382.360 129.200 ;
        RECT 381.910 122.830 382.360 123.450 ;
        RECT 374.330 117.450 374.820 117.760 ;
        RECT 367.650 117.250 374.820 117.450 ;
        RECT 364.110 117.230 374.820 117.250 ;
        RECT 351.280 117.210 360.550 117.220 ;
        RECT 362.780 117.210 374.820 117.230 ;
        RECT 348.450 116.690 374.820 117.210 ;
        RECT 348.450 116.680 362.860 116.690 ;
        RECT 348.450 116.670 351.290 116.680 ;
        RECT 360.500 116.670 362.860 116.680 ;
        RECT 364.110 116.670 374.820 116.690 ;
        RECT 349.060 110.590 349.610 116.670 ;
        RECT 364.110 116.650 367.930 116.670 ;
        RECT 364.170 114.860 364.660 116.650 ;
        RECT 364.170 114.370 364.680 114.860 ;
        RECT 348.620 110.190 349.610 110.590 ;
        RECT 348.620 110.170 349.200 110.190 ;
        RECT 374.400 107.840 374.790 116.670 ;
        RECT 390.830 107.840 391.270 107.850 ;
        RECT 374.290 107.450 399.820 107.840 ;
        RECT 351.420 101.560 360.690 101.570 ;
        RECT 362.920 101.560 364.830 101.580 ;
        RECT 348.590 101.040 364.830 101.560 ;
        RECT 348.590 101.030 363.000 101.040 ;
        RECT 348.590 101.020 351.430 101.030 ;
        RECT 360.640 101.020 363.000 101.030 ;
        RECT 349.200 94.940 349.750 101.020 ;
        RECT 364.310 99.560 364.800 101.040 ;
        RECT 374.400 99.740 374.790 107.450 ;
        RECT 374.300 99.610 374.810 99.740 ;
        RECT 379.030 99.610 382.360 99.630 ;
        RECT 372.130 99.580 382.360 99.610 ;
        RECT 371.570 99.570 382.360 99.580 ;
        RECT 369.860 99.560 382.360 99.570 ;
        RECT 364.310 99.210 382.360 99.560 ;
        RECT 364.310 99.200 371.640 99.210 ;
        RECT 364.310 99.190 369.930 99.200 ;
        RECT 364.310 98.720 364.820 99.190 ;
        RECT 372.130 99.170 382.360 99.210 ;
        RECT 348.760 94.540 349.750 94.940 ;
        RECT 348.760 94.520 349.340 94.540 ;
        RECT 374.300 87.690 374.810 99.170 ;
        RECT 379.030 99.130 382.360 99.170 ;
        RECT 381.890 93.380 382.330 99.130 ;
        RECT 381.880 92.760 382.330 93.380 ;
        RECT 390.830 89.400 391.270 107.450 ;
        RECT 399.440 106.780 399.820 107.450 ;
        RECT 374.300 87.380 374.790 87.690 ;
        RECT 367.620 87.180 374.790 87.380 ;
        RECT 364.080 87.160 374.790 87.180 ;
        RECT 351.250 87.140 360.520 87.150 ;
        RECT 362.750 87.140 374.790 87.160 ;
        RECT 312.310 86.350 312.930 86.700 ;
        RECT 348.420 86.620 374.790 87.140 ;
        RECT 348.420 86.610 362.830 86.620 ;
        RECT 348.420 86.600 351.260 86.610 ;
        RECT 360.470 86.600 362.830 86.610 ;
        RECT 364.080 86.600 374.790 86.620 ;
        RECT 312.350 82.120 312.930 86.350 ;
        RECT 312.340 82.100 312.930 82.120 ;
        RECT 289.500 81.570 312.930 82.100 ;
        RECT 289.500 81.540 312.920 81.570 ;
        RECT 247.280 80.310 248.270 80.710 ;
        RECT 247.280 80.290 247.860 80.310 ;
        RECT 249.790 71.900 259.060 71.910 ;
        RECT 261.290 71.900 263.200 71.920 ;
        RECT 246.960 71.380 263.200 71.900 ;
        RECT 246.960 71.370 261.370 71.380 ;
        RECT 246.960 71.360 249.800 71.370 ;
        RECT 259.010 71.360 261.370 71.370 ;
        RECT 247.570 65.280 248.120 71.360 ;
        RECT 262.680 69.900 263.170 71.380 ;
        RECT 272.670 69.950 273.180 70.080 ;
        RECT 277.400 69.950 280.730 69.970 ;
        RECT 270.500 69.920 280.730 69.950 ;
        RECT 269.940 69.910 280.730 69.920 ;
        RECT 268.230 69.900 280.730 69.910 ;
        RECT 262.680 69.550 280.730 69.900 ;
        RECT 262.680 69.540 270.010 69.550 ;
        RECT 262.680 69.530 268.300 69.540 ;
        RECT 262.680 69.060 263.190 69.530 ;
        RECT 270.500 69.510 280.730 69.550 ;
        RECT 247.130 64.880 248.120 65.280 ;
        RECT 247.130 64.860 247.710 64.880 ;
        RECT 272.670 58.030 273.180 69.510 ;
        RECT 277.400 69.470 280.730 69.510 ;
        RECT 280.260 63.720 280.700 69.470 ;
        RECT 280.250 63.100 280.700 63.720 ;
        RECT 272.670 57.720 273.160 58.030 ;
        RECT 265.990 57.520 273.160 57.720 ;
        RECT 262.450 57.500 273.160 57.520 ;
        RECT 249.620 57.480 258.890 57.490 ;
        RECT 261.120 57.480 273.160 57.500 ;
        RECT 246.790 56.960 273.160 57.480 ;
        RECT 246.790 56.950 261.200 56.960 ;
        RECT 246.790 56.940 249.630 56.950 ;
        RECT 258.840 56.940 261.200 56.950 ;
        RECT 262.450 56.940 273.160 56.960 ;
        RECT 247.400 50.860 247.950 56.940 ;
        RECT 262.450 56.920 266.270 56.940 ;
        RECT 262.510 55.130 263.000 56.920 ;
        RECT 262.510 54.640 263.020 55.130 ;
        RECT 246.960 50.460 247.950 50.860 ;
        RECT 246.960 50.440 247.540 50.460 ;
        RECT 272.740 48.110 273.130 56.940 ;
        RECT 289.520 48.110 289.970 81.540 ;
        RECT 312.340 80.680 312.920 81.540 ;
        RECT 349.030 80.520 349.580 86.600 ;
        RECT 364.080 86.580 367.900 86.600 ;
        RECT 364.140 84.790 364.630 86.580 ;
        RECT 364.140 84.300 364.650 84.790 ;
        RECT 390.830 81.910 391.280 89.400 ;
        RECT 413.620 86.510 414.150 143.030 ;
        RECT 430.180 143.020 430.940 143.030 ;
        RECT 430.480 141.790 430.940 143.020 ;
        RECT 430.470 141.710 430.940 141.790 ;
        RECT 430.470 138.060 430.930 141.710 ;
        RECT 456.730 140.700 457.210 143.070 ;
        RECT 456.670 140.350 474.450 140.700 ;
        RECT 456.730 140.280 457.240 140.350 ;
        RECT 456.740 139.690 457.240 140.280 ;
        RECT 430.470 137.490 430.920 138.060 ;
        RECT 474.080 137.950 474.450 140.350 ;
        RECT 474.050 137.920 474.450 137.950 ;
        RECT 474.050 137.300 474.440 137.920 ;
        RECT 413.620 86.160 414.240 86.510 ;
        RECT 413.660 81.930 414.240 86.160 ;
        RECT 413.650 81.910 414.240 81.930 ;
        RECT 390.810 81.380 414.240 81.910 ;
        RECT 390.810 81.350 414.230 81.380 ;
        RECT 348.590 80.120 349.580 80.520 ;
        RECT 348.590 80.100 349.170 80.120 ;
        RECT 351.100 71.710 360.370 71.720 ;
        RECT 362.600 71.710 364.510 71.730 ;
        RECT 348.270 71.190 364.510 71.710 ;
        RECT 348.270 71.180 362.680 71.190 ;
        RECT 348.270 71.170 351.110 71.180 ;
        RECT 360.320 71.170 362.680 71.180 ;
        RECT 348.880 65.090 349.430 71.170 ;
        RECT 363.990 69.710 364.480 71.190 ;
        RECT 373.980 69.760 374.490 69.890 ;
        RECT 378.710 69.760 382.040 69.780 ;
        RECT 371.810 69.730 382.040 69.760 ;
        RECT 371.250 69.720 382.040 69.730 ;
        RECT 369.540 69.710 382.040 69.720 ;
        RECT 363.990 69.360 382.040 69.710 ;
        RECT 363.990 69.350 371.320 69.360 ;
        RECT 363.990 69.340 369.610 69.350 ;
        RECT 363.990 68.870 364.500 69.340 ;
        RECT 371.810 69.320 382.040 69.360 ;
        RECT 348.440 64.690 349.430 65.090 ;
        RECT 348.440 64.670 349.020 64.690 ;
        RECT 373.980 57.840 374.490 69.320 ;
        RECT 378.710 69.280 382.040 69.320 ;
        RECT 381.570 63.530 382.010 69.280 ;
        RECT 381.560 62.910 382.010 63.530 ;
        RECT 373.980 57.530 374.470 57.840 ;
        RECT 367.300 57.330 374.470 57.530 ;
        RECT 363.760 57.310 374.470 57.330 ;
        RECT 350.930 57.290 360.200 57.300 ;
        RECT 362.430 57.290 374.470 57.310 ;
        RECT 348.100 56.770 374.470 57.290 ;
        RECT 348.100 56.760 362.510 56.770 ;
        RECT 348.100 56.750 350.940 56.760 ;
        RECT 360.150 56.750 362.510 56.760 ;
        RECT 363.760 56.750 374.470 56.770 ;
        RECT 348.710 50.670 349.260 56.750 ;
        RECT 363.760 56.730 367.580 56.750 ;
        RECT 363.820 54.940 364.310 56.730 ;
        RECT 363.820 54.450 364.330 54.940 ;
        RECT 348.270 50.270 349.260 50.670 ;
        RECT 348.270 50.250 348.850 50.270 ;
        RECT 13.230 41.890 22.500 41.900 ;
        RECT 24.730 41.890 26.640 41.910 ;
        RECT 10.400 41.370 26.640 41.890 ;
        RECT 10.400 41.360 24.810 41.370 ;
        RECT 10.400 41.350 13.240 41.360 ;
        RECT 22.450 41.350 24.810 41.360 ;
        RECT 11.010 35.270 11.560 41.350 ;
        RECT 26.120 39.890 26.610 41.370 ;
        RECT 36.210 40.070 36.600 47.780 ;
        RECT 52.990 47.540 53.440 47.780 ;
        RECT 61.250 47.110 61.630 47.780 ;
        RECT 137.410 47.590 162.940 47.980 ;
        RECT 272.630 47.720 298.160 48.110 ;
        RECT 374.050 47.920 374.440 56.750 ;
        RECT 390.830 47.920 391.280 81.350 ;
        RECT 413.650 80.490 414.230 81.350 ;
        RECT 114.540 41.700 123.810 41.710 ;
        RECT 126.040 41.700 127.950 41.720 ;
        RECT 111.710 41.180 127.950 41.700 ;
        RECT 111.710 41.170 126.120 41.180 ;
        RECT 111.710 41.160 114.550 41.170 ;
        RECT 123.760 41.160 126.120 41.170 ;
        RECT 36.110 39.940 36.620 40.070 ;
        RECT 40.840 39.940 44.170 39.960 ;
        RECT 33.940 39.910 44.170 39.940 ;
        RECT 33.380 39.900 44.170 39.910 ;
        RECT 31.670 39.890 44.170 39.900 ;
        RECT 26.120 39.540 44.170 39.890 ;
        RECT 26.120 39.530 33.450 39.540 ;
        RECT 26.120 39.520 31.740 39.530 ;
        RECT 26.120 39.050 26.630 39.520 ;
        RECT 33.940 39.500 44.170 39.540 ;
        RECT 10.570 34.870 11.560 35.270 ;
        RECT 10.570 34.850 11.150 34.870 ;
        RECT 36.110 28.020 36.620 39.500 ;
        RECT 40.840 39.460 44.170 39.500 ;
        RECT 43.700 33.710 44.140 39.460 ;
        RECT 112.320 35.080 112.870 41.160 ;
        RECT 127.430 39.700 127.920 41.180 ;
        RECT 137.520 39.880 137.910 47.590 ;
        RECT 154.300 47.350 154.750 47.590 ;
        RECT 162.560 46.920 162.940 47.590 ;
        RECT 249.760 41.830 259.030 41.840 ;
        RECT 261.260 41.830 263.170 41.850 ;
        RECT 246.930 41.310 263.170 41.830 ;
        RECT 246.930 41.300 261.340 41.310 ;
        RECT 246.930 41.290 249.770 41.300 ;
        RECT 258.980 41.290 261.340 41.300 ;
        RECT 137.420 39.750 137.930 39.880 ;
        RECT 142.150 39.750 145.480 39.770 ;
        RECT 135.250 39.720 145.480 39.750 ;
        RECT 134.690 39.710 145.480 39.720 ;
        RECT 132.980 39.700 145.480 39.710 ;
        RECT 127.430 39.350 145.480 39.700 ;
        RECT 127.430 39.340 134.760 39.350 ;
        RECT 127.430 39.330 133.050 39.340 ;
        RECT 127.430 38.860 127.940 39.330 ;
        RECT 135.250 39.310 145.480 39.350 ;
        RECT 111.880 34.680 112.870 35.080 ;
        RECT 111.880 34.660 112.460 34.680 ;
        RECT 43.690 33.090 44.140 33.710 ;
        RECT 36.110 27.710 36.600 28.020 ;
        RECT 29.430 27.510 36.600 27.710 ;
        RECT 137.420 27.830 137.930 39.310 ;
        RECT 142.150 39.270 145.480 39.310 ;
        RECT 145.010 33.520 145.450 39.270 ;
        RECT 247.540 35.210 248.090 41.290 ;
        RECT 262.650 39.830 263.140 41.310 ;
        RECT 272.740 40.010 273.130 47.720 ;
        RECT 289.520 47.480 289.970 47.720 ;
        RECT 297.780 47.050 298.160 47.720 ;
        RECT 373.940 47.530 399.470 47.920 ;
        RECT 351.070 41.640 360.340 41.650 ;
        RECT 362.570 41.640 364.480 41.660 ;
        RECT 348.240 41.120 364.480 41.640 ;
        RECT 348.240 41.110 362.650 41.120 ;
        RECT 348.240 41.100 351.080 41.110 ;
        RECT 360.290 41.100 362.650 41.110 ;
        RECT 272.640 39.880 273.150 40.010 ;
        RECT 277.370 39.880 280.700 39.900 ;
        RECT 270.470 39.850 280.700 39.880 ;
        RECT 269.910 39.840 280.700 39.850 ;
        RECT 268.200 39.830 280.700 39.840 ;
        RECT 262.650 39.480 280.700 39.830 ;
        RECT 262.650 39.470 269.980 39.480 ;
        RECT 262.650 39.460 268.270 39.470 ;
        RECT 262.650 38.990 263.160 39.460 ;
        RECT 270.470 39.440 280.700 39.480 ;
        RECT 247.100 34.810 248.090 35.210 ;
        RECT 247.100 34.790 247.680 34.810 ;
        RECT 145.000 32.900 145.450 33.520 ;
        RECT 272.640 27.960 273.150 39.440 ;
        RECT 277.370 39.400 280.700 39.440 ;
        RECT 280.230 33.650 280.670 39.400 ;
        RECT 348.850 35.020 349.400 41.100 ;
        RECT 363.960 39.640 364.450 41.120 ;
        RECT 374.050 39.820 374.440 47.530 ;
        RECT 390.830 47.290 391.280 47.530 ;
        RECT 399.090 46.860 399.470 47.530 ;
        RECT 373.950 39.690 374.460 39.820 ;
        RECT 378.680 39.690 382.010 39.710 ;
        RECT 371.780 39.660 382.010 39.690 ;
        RECT 371.220 39.650 382.010 39.660 ;
        RECT 369.510 39.640 382.010 39.650 ;
        RECT 363.960 39.290 382.010 39.640 ;
        RECT 363.960 39.280 371.290 39.290 ;
        RECT 363.960 39.270 369.580 39.280 ;
        RECT 363.960 38.800 364.470 39.270 ;
        RECT 371.780 39.250 382.010 39.290 ;
        RECT 348.410 34.620 349.400 35.020 ;
        RECT 348.410 34.600 348.990 34.620 ;
        RECT 280.220 33.030 280.670 33.650 ;
        RECT 137.420 27.520 137.910 27.830 ;
        RECT 272.640 27.650 273.130 27.960 ;
        RECT 25.890 27.490 36.600 27.510 ;
        RECT 13.060 27.470 22.330 27.480 ;
        RECT 24.560 27.470 36.600 27.490 ;
        RECT 10.230 26.950 36.600 27.470 ;
        RECT 130.740 27.320 137.910 27.520 ;
        RECT 265.960 27.450 273.130 27.650 ;
        RECT 373.950 27.770 374.460 39.250 ;
        RECT 378.680 39.210 382.010 39.250 ;
        RECT 381.540 33.460 381.980 39.210 ;
        RECT 381.530 32.840 381.980 33.460 ;
        RECT 373.950 27.460 374.440 27.770 ;
        RECT 262.420 27.430 273.130 27.450 ;
        RECT 249.590 27.410 258.860 27.420 ;
        RECT 261.090 27.410 273.130 27.430 ;
        RECT 127.200 27.300 137.910 27.320 ;
        RECT 114.370 27.280 123.640 27.290 ;
        RECT 125.870 27.280 137.910 27.300 ;
        RECT 10.230 26.940 24.640 26.950 ;
        RECT 10.230 26.930 13.070 26.940 ;
        RECT 22.280 26.930 24.640 26.940 ;
        RECT 25.890 26.930 36.600 26.950 ;
        RECT 10.840 20.850 11.390 26.930 ;
        RECT 25.890 26.910 29.710 26.930 ;
        RECT 25.950 25.120 26.440 26.910 ;
        RECT 111.540 26.760 137.910 27.280 ;
        RECT 246.760 26.890 273.130 27.410 ;
        RECT 367.270 27.260 374.440 27.460 ;
        RECT 363.730 27.240 374.440 27.260 ;
        RECT 350.900 27.220 360.170 27.230 ;
        RECT 362.400 27.220 374.440 27.240 ;
        RECT 246.760 26.880 261.170 26.890 ;
        RECT 246.760 26.870 249.600 26.880 ;
        RECT 258.810 26.870 261.170 26.880 ;
        RECT 262.420 26.870 273.130 26.890 ;
        RECT 111.540 26.750 125.950 26.760 ;
        RECT 111.540 26.740 114.380 26.750 ;
        RECT 123.590 26.740 125.950 26.750 ;
        RECT 127.200 26.740 137.910 26.760 ;
        RECT 25.950 24.630 26.460 25.120 ;
        RECT 10.400 20.450 11.390 20.850 ;
        RECT 112.150 20.660 112.700 26.740 ;
        RECT 127.200 26.720 131.020 26.740 ;
        RECT 127.260 24.930 127.750 26.720 ;
        RECT 127.260 24.440 127.770 24.930 ;
        RECT 247.370 20.790 247.920 26.870 ;
        RECT 262.420 26.850 266.240 26.870 ;
        RECT 262.480 25.060 262.970 26.850 ;
        RECT 348.070 26.700 374.440 27.220 ;
        RECT 348.070 26.690 362.480 26.700 ;
        RECT 348.070 26.680 350.910 26.690 ;
        RECT 360.120 26.680 362.480 26.690 ;
        RECT 363.730 26.680 374.440 26.700 ;
        RECT 262.480 24.570 262.990 25.060 ;
        RECT 10.400 20.430 10.980 20.450 ;
        RECT 111.710 20.260 112.700 20.660 ;
        RECT 246.930 20.390 247.920 20.790 ;
        RECT 348.680 20.600 349.230 26.680 ;
        RECT 363.730 26.660 367.550 26.680 ;
        RECT 363.790 24.870 364.280 26.660 ;
        RECT 363.790 24.380 364.300 24.870 ;
        RECT 246.930 20.370 247.510 20.390 ;
        RECT 111.710 20.240 112.290 20.260 ;
        RECT 348.240 20.200 349.230 20.600 ;
        RECT 348.240 20.180 348.820 20.200 ;
    END
  END vdd
  PIN gnd
    ANTENNADIFFAREA 525.044983 ;
    PORT
      LAYER pwell ;
        RECT 8.030 246.920 9.320 247.880 ;
        RECT 9.920 246.920 11.210 247.880 ;
        RECT 7.920 246.070 9.470 246.920 ;
        RECT 9.810 246.070 11.360 246.920 ;
        RECT 109.340 246.730 110.630 247.690 ;
        RECT 111.230 246.730 112.520 247.690 ;
        RECT 244.560 246.860 245.850 247.820 ;
        RECT 246.450 246.860 247.740 247.820 ;
        RECT 109.230 245.880 110.780 246.730 ;
        RECT 111.120 245.880 112.670 246.730 ;
        RECT 244.450 246.010 246.000 246.860 ;
        RECT 246.340 246.010 247.890 246.860 ;
        RECT 345.870 246.670 347.160 247.630 ;
        RECT 347.760 246.670 349.050 247.630 ;
        RECT 345.760 245.820 347.310 246.670 ;
        RECT 347.650 245.820 349.200 246.670 ;
        RECT 23.710 244.500 25.000 245.460 ;
        RECT 25.600 244.500 26.890 245.460 ;
        RECT 23.600 243.650 25.150 244.500 ;
        RECT 25.490 243.650 27.040 244.500 ;
        RECT 125.020 244.310 126.310 245.270 ;
        RECT 126.910 244.310 128.200 245.270 ;
        RECT 260.240 244.440 261.530 245.400 ;
        RECT 262.130 244.440 263.420 245.400 ;
        RECT 124.910 243.460 126.460 244.310 ;
        RECT 126.800 243.460 128.350 244.310 ;
        RECT 260.130 243.590 261.680 244.440 ;
        RECT 262.020 243.590 263.570 244.440 ;
        RECT 361.550 244.250 362.840 245.210 ;
        RECT 363.440 244.250 364.730 245.210 ;
        RECT 361.440 243.400 362.990 244.250 ;
        RECT 363.330 243.400 364.880 244.250 ;
        RECT 8.190 240.520 9.480 241.480 ;
        RECT 10.080 240.520 11.370 241.480 ;
        RECT 8.080 239.670 9.630 240.520 ;
        RECT 9.970 239.670 11.520 240.520 ;
        RECT 109.500 240.330 110.790 241.290 ;
        RECT 111.390 240.330 112.680 241.290 ;
        RECT 244.720 240.460 246.010 241.420 ;
        RECT 246.610 240.460 247.900 241.420 ;
        RECT 41.290 238.950 42.580 239.910 ;
        RECT 43.180 238.950 44.470 239.910 ;
        RECT 109.390 239.480 110.940 240.330 ;
        RECT 111.280 239.480 112.830 240.330 ;
        RECT 41.180 238.100 42.730 238.950 ;
        RECT 43.070 238.100 44.620 238.950 ;
        RECT 142.600 238.760 143.890 239.720 ;
        RECT 144.490 238.760 145.780 239.720 ;
        RECT 244.610 239.610 246.160 240.460 ;
        RECT 246.500 239.610 248.050 240.460 ;
        RECT 346.030 240.270 347.320 241.230 ;
        RECT 347.920 240.270 349.210 241.230 ;
        RECT 277.820 238.890 279.110 239.850 ;
        RECT 279.710 238.890 281.000 239.850 ;
        RECT 345.920 239.420 347.470 240.270 ;
        RECT 347.810 239.420 349.360 240.270 ;
        RECT 142.490 237.910 144.040 238.760 ;
        RECT 144.380 237.910 145.930 238.760 ;
        RECT 277.710 238.040 279.260 238.890 ;
        RECT 279.600 238.040 281.150 238.890 ;
        RECT 379.130 238.700 380.420 239.660 ;
        RECT 381.020 238.700 382.310 239.660 ;
        RECT 379.020 237.850 380.570 238.700 ;
        RECT 380.910 237.850 382.460 238.700 ;
        RECT 7.860 232.500 9.150 233.460 ;
        RECT 9.750 232.500 11.040 233.460 ;
        RECT 7.750 231.650 9.300 232.500 ;
        RECT 9.640 231.650 11.190 232.500 ;
        RECT 109.170 232.310 110.460 233.270 ;
        RECT 111.060 232.310 112.350 233.270 ;
        RECT 244.390 232.440 245.680 233.400 ;
        RECT 246.280 232.440 247.570 233.400 ;
        RECT 109.060 231.460 110.610 232.310 ;
        RECT 110.950 231.460 112.500 232.310 ;
        RECT 244.280 231.590 245.830 232.440 ;
        RECT 246.170 231.590 247.720 232.440 ;
        RECT 345.700 232.250 346.990 233.210 ;
        RECT 347.590 232.250 348.880 233.210 ;
        RECT 345.590 231.400 347.140 232.250 ;
        RECT 347.480 231.400 349.030 232.250 ;
        RECT 23.540 230.080 24.830 231.040 ;
        RECT 25.430 230.080 26.720 231.040 ;
        RECT 23.430 229.230 24.980 230.080 ;
        RECT 25.320 229.230 26.870 230.080 ;
        RECT 124.850 229.890 126.140 230.850 ;
        RECT 126.740 229.890 128.030 230.850 ;
        RECT 260.070 230.020 261.360 230.980 ;
        RECT 261.960 230.020 263.250 230.980 ;
        RECT 124.740 229.040 126.290 229.890 ;
        RECT 126.630 229.040 128.180 229.890 ;
        RECT 259.960 229.170 261.510 230.020 ;
        RECT 261.850 229.170 263.400 230.020 ;
        RECT 361.380 229.830 362.670 230.790 ;
        RECT 363.270 229.830 364.560 230.790 ;
        RECT 361.270 228.980 362.820 229.830 ;
        RECT 363.160 228.980 364.710 229.830 ;
        RECT 8.020 226.100 9.310 227.060 ;
        RECT 9.910 226.100 11.200 227.060 ;
        RECT 7.910 225.250 9.460 226.100 ;
        RECT 9.800 225.250 11.350 226.100 ;
        RECT 109.330 225.910 110.620 226.870 ;
        RECT 111.220 225.910 112.510 226.870 ;
        RECT 244.550 226.040 245.840 227.000 ;
        RECT 246.440 226.040 247.730 227.000 ;
        RECT 109.220 225.060 110.770 225.910 ;
        RECT 111.110 225.060 112.660 225.910 ;
        RECT 244.440 225.190 245.990 226.040 ;
        RECT 246.330 225.190 247.880 226.040 ;
        RECT 345.860 225.850 347.150 226.810 ;
        RECT 347.750 225.850 349.040 226.810 ;
        RECT 345.750 225.000 347.300 225.850 ;
        RECT 347.640 225.000 349.190 225.850 ;
        RECT 58.820 222.930 60.110 223.890 ;
        RECT 60.710 222.930 62.000 223.890 ;
        RECT 58.710 222.080 60.260 222.930 ;
        RECT 60.600 222.080 62.150 222.930 ;
        RECT 160.130 222.740 161.420 223.700 ;
        RECT 162.020 222.740 163.310 223.700 ;
        RECT 295.350 222.870 296.640 223.830 ;
        RECT 297.240 222.870 298.530 223.830 ;
        RECT 160.020 221.890 161.570 222.740 ;
        RECT 161.910 221.890 163.460 222.740 ;
        RECT 295.240 222.020 296.790 222.870 ;
        RECT 297.130 222.020 298.680 222.870 ;
        RECT 396.660 222.680 397.950 223.640 ;
        RECT 398.550 222.680 399.840 223.640 ;
        RECT 396.550 221.830 398.100 222.680 ;
        RECT 398.440 221.830 399.990 222.680 ;
        RECT 8.000 216.850 9.290 217.810 ;
        RECT 9.890 216.850 11.180 217.810 ;
        RECT 7.890 216.000 9.440 216.850 ;
        RECT 9.780 216.000 11.330 216.850 ;
        RECT 109.310 216.660 110.600 217.620 ;
        RECT 111.200 216.660 112.490 217.620 ;
        RECT 244.530 216.790 245.820 217.750 ;
        RECT 246.420 216.790 247.710 217.750 ;
        RECT 109.200 215.810 110.750 216.660 ;
        RECT 111.090 215.810 112.640 216.660 ;
        RECT 244.420 215.940 245.970 216.790 ;
        RECT 246.310 215.940 247.860 216.790 ;
        RECT 345.840 216.600 347.130 217.560 ;
        RECT 347.730 216.600 349.020 217.560 ;
        RECT 345.730 215.750 347.280 216.600 ;
        RECT 347.620 215.750 349.170 216.600 ;
        RECT 23.680 214.430 24.970 215.390 ;
        RECT 25.570 214.430 26.860 215.390 ;
        RECT 23.570 213.580 25.120 214.430 ;
        RECT 25.460 213.580 27.010 214.430 ;
        RECT 124.990 214.240 126.280 215.200 ;
        RECT 126.880 214.240 128.170 215.200 ;
        RECT 260.210 214.370 261.500 215.330 ;
        RECT 262.100 214.370 263.390 215.330 ;
        RECT 124.880 213.390 126.430 214.240 ;
        RECT 126.770 213.390 128.320 214.240 ;
        RECT 260.100 213.520 261.650 214.370 ;
        RECT 261.990 213.520 263.540 214.370 ;
        RECT 361.520 214.180 362.810 215.140 ;
        RECT 363.410 214.180 364.700 215.140 ;
        RECT 361.410 213.330 362.960 214.180 ;
        RECT 363.300 213.330 364.850 214.180 ;
        RECT 8.160 210.450 9.450 211.410 ;
        RECT 10.050 210.450 11.340 211.410 ;
        RECT 8.050 209.600 9.600 210.450 ;
        RECT 9.940 209.600 11.490 210.450 ;
        RECT 109.470 210.260 110.760 211.220 ;
        RECT 111.360 210.260 112.650 211.220 ;
        RECT 244.690 210.390 245.980 211.350 ;
        RECT 246.580 210.390 247.870 211.350 ;
        RECT 41.260 208.880 42.550 209.840 ;
        RECT 43.150 208.880 44.440 209.840 ;
        RECT 109.360 209.410 110.910 210.260 ;
        RECT 111.250 209.410 112.800 210.260 ;
        RECT 41.150 208.030 42.700 208.880 ;
        RECT 43.040 208.030 44.590 208.880 ;
        RECT 142.570 208.690 143.860 209.650 ;
        RECT 144.460 208.690 145.750 209.650 ;
        RECT 244.580 209.540 246.130 210.390 ;
        RECT 246.470 209.540 248.020 210.390 ;
        RECT 346.000 210.200 347.290 211.160 ;
        RECT 347.890 210.200 349.180 211.160 ;
        RECT 277.790 208.820 279.080 209.780 ;
        RECT 279.680 208.820 280.970 209.780 ;
        RECT 345.890 209.350 347.440 210.200 ;
        RECT 347.780 209.350 349.330 210.200 ;
        RECT 142.460 207.840 144.010 208.690 ;
        RECT 144.350 207.840 145.900 208.690 ;
        RECT 277.680 207.970 279.230 208.820 ;
        RECT 279.570 207.970 281.120 208.820 ;
        RECT 379.100 208.630 380.390 209.590 ;
        RECT 380.990 208.630 382.280 209.590 ;
        RECT 378.990 207.780 380.540 208.630 ;
        RECT 380.880 207.780 382.430 208.630 ;
        RECT 7.830 202.430 9.120 203.390 ;
        RECT 9.720 202.430 11.010 203.390 ;
        RECT 7.720 201.580 9.270 202.430 ;
        RECT 9.610 201.580 11.160 202.430 ;
        RECT 109.140 202.240 110.430 203.200 ;
        RECT 111.030 202.240 112.320 203.200 ;
        RECT 244.360 202.370 245.650 203.330 ;
        RECT 246.250 202.370 247.540 203.330 ;
        RECT 109.030 201.390 110.580 202.240 ;
        RECT 110.920 201.390 112.470 202.240 ;
        RECT 244.250 201.520 245.800 202.370 ;
        RECT 246.140 201.520 247.690 202.370 ;
        RECT 345.670 202.180 346.960 203.140 ;
        RECT 347.560 202.180 348.850 203.140 ;
        RECT 345.560 201.330 347.110 202.180 ;
        RECT 347.450 201.330 349.000 202.180 ;
        RECT 23.510 200.010 24.800 200.970 ;
        RECT 25.400 200.010 26.690 200.970 ;
        RECT 23.400 199.160 24.950 200.010 ;
        RECT 25.290 199.160 26.840 200.010 ;
        RECT 124.820 199.820 126.110 200.780 ;
        RECT 126.710 199.820 128.000 200.780 ;
        RECT 260.040 199.950 261.330 200.910 ;
        RECT 261.930 199.950 263.220 200.910 ;
        RECT 124.710 198.970 126.260 199.820 ;
        RECT 126.600 198.970 128.150 199.820 ;
        RECT 259.930 199.100 261.480 199.950 ;
        RECT 261.820 199.100 263.370 199.950 ;
        RECT 361.350 199.760 362.640 200.720 ;
        RECT 363.240 199.760 364.530 200.720 ;
        RECT 361.240 198.910 362.790 199.760 ;
        RECT 363.130 198.910 364.680 199.760 ;
        RECT 7.990 196.030 9.280 196.990 ;
        RECT 9.880 196.030 11.170 196.990 ;
        RECT 73.020 196.640 74.310 197.600 ;
        RECT 74.910 196.640 76.200 197.600 ;
        RECT 7.880 195.180 9.430 196.030 ;
        RECT 9.770 195.180 11.320 196.030 ;
        RECT 72.910 195.790 74.460 196.640 ;
        RECT 74.800 195.790 76.350 196.640 ;
        RECT 109.300 195.840 110.590 196.800 ;
        RECT 111.190 195.840 112.480 196.800 ;
        RECT 174.330 196.450 175.620 197.410 ;
        RECT 176.220 196.450 177.510 197.410 ;
        RECT 109.190 194.990 110.740 195.840 ;
        RECT 111.080 194.990 112.630 195.840 ;
        RECT 174.220 195.600 175.770 196.450 ;
        RECT 176.110 195.600 177.660 196.450 ;
        RECT 244.520 195.970 245.810 196.930 ;
        RECT 246.410 195.970 247.700 196.930 ;
        RECT 309.550 196.580 310.840 197.540 ;
        RECT 311.440 196.580 312.730 197.540 ;
        RECT 244.410 195.120 245.960 195.970 ;
        RECT 246.300 195.120 247.850 195.970 ;
        RECT 309.440 195.730 310.990 196.580 ;
        RECT 311.330 195.730 312.880 196.580 ;
        RECT 345.830 195.780 347.120 196.740 ;
        RECT 347.720 195.780 349.010 196.740 ;
        RECT 410.860 196.390 412.150 197.350 ;
        RECT 412.750 196.390 414.040 197.350 ;
        RECT 345.720 194.930 347.270 195.780 ;
        RECT 347.610 194.930 349.160 195.780 ;
        RECT 410.750 195.540 412.300 196.390 ;
        RECT 412.640 195.540 414.190 196.390 ;
        RECT 7.680 187.000 8.970 187.960 ;
        RECT 9.570 187.000 10.860 187.960 ;
        RECT 7.570 186.150 9.120 187.000 ;
        RECT 9.460 186.150 11.010 187.000 ;
        RECT 108.990 186.810 110.280 187.770 ;
        RECT 110.880 186.810 112.170 187.770 ;
        RECT 244.210 186.940 245.500 187.900 ;
        RECT 246.100 186.940 247.390 187.900 ;
        RECT 108.880 185.960 110.430 186.810 ;
        RECT 110.770 185.960 112.320 186.810 ;
        RECT 244.100 186.090 245.650 186.940 ;
        RECT 245.990 186.090 247.540 186.940 ;
        RECT 345.520 186.750 346.810 187.710 ;
        RECT 347.410 186.750 348.700 187.710 ;
        RECT 345.410 185.900 346.960 186.750 ;
        RECT 347.300 185.900 348.850 186.750 ;
        RECT 23.360 184.580 24.650 185.540 ;
        RECT 25.250 184.580 26.540 185.540 ;
        RECT 23.250 183.730 24.800 184.580 ;
        RECT 25.140 183.730 26.690 184.580 ;
        RECT 124.670 184.390 125.960 185.350 ;
        RECT 126.560 184.390 127.850 185.350 ;
        RECT 259.890 184.520 261.180 185.480 ;
        RECT 261.780 184.520 263.070 185.480 ;
        RECT 124.560 183.540 126.110 184.390 ;
        RECT 126.450 183.540 128.000 184.390 ;
        RECT 259.780 183.670 261.330 184.520 ;
        RECT 261.670 183.670 263.220 184.520 ;
        RECT 361.200 184.330 362.490 185.290 ;
        RECT 363.090 184.330 364.380 185.290 ;
        RECT 361.090 183.480 362.640 184.330 ;
        RECT 362.980 183.480 364.530 184.330 ;
        RECT 7.840 180.600 9.130 181.560 ;
        RECT 9.730 180.600 11.020 181.560 ;
        RECT 7.730 179.750 9.280 180.600 ;
        RECT 9.620 179.750 11.170 180.600 ;
        RECT 109.150 180.410 110.440 181.370 ;
        RECT 111.040 180.410 112.330 181.370 ;
        RECT 244.370 180.540 245.660 181.500 ;
        RECT 246.260 180.540 247.550 181.500 ;
        RECT 40.940 179.030 42.230 179.990 ;
        RECT 42.830 179.030 44.120 179.990 ;
        RECT 109.040 179.560 110.590 180.410 ;
        RECT 110.930 179.560 112.480 180.410 ;
        RECT 40.830 178.180 42.380 179.030 ;
        RECT 42.720 178.180 44.270 179.030 ;
        RECT 142.250 178.840 143.540 179.800 ;
        RECT 144.140 178.840 145.430 179.800 ;
        RECT 244.260 179.690 245.810 180.540 ;
        RECT 246.150 179.690 247.700 180.540 ;
        RECT 345.680 180.350 346.970 181.310 ;
        RECT 347.570 180.350 348.860 181.310 ;
        RECT 277.470 178.970 278.760 179.930 ;
        RECT 279.360 178.970 280.650 179.930 ;
        RECT 345.570 179.500 347.120 180.350 ;
        RECT 347.460 179.500 349.010 180.350 ;
        RECT 142.140 177.990 143.690 178.840 ;
        RECT 144.030 177.990 145.580 178.840 ;
        RECT 277.360 178.120 278.910 178.970 ;
        RECT 279.250 178.120 280.800 178.970 ;
        RECT 378.780 178.780 380.070 179.740 ;
        RECT 380.670 178.780 381.960 179.740 ;
        RECT 378.670 177.930 380.220 178.780 ;
        RECT 380.560 177.930 382.110 178.780 ;
        RECT 7.510 172.580 8.800 173.540 ;
        RECT 9.400 172.580 10.690 173.540 ;
        RECT 7.400 171.730 8.950 172.580 ;
        RECT 9.290 171.730 10.840 172.580 ;
        RECT 108.820 172.390 110.110 173.350 ;
        RECT 110.710 172.390 112.000 173.350 ;
        RECT 244.040 172.520 245.330 173.480 ;
        RECT 245.930 172.520 247.220 173.480 ;
        RECT 108.710 171.540 110.260 172.390 ;
        RECT 110.600 171.540 112.150 172.390 ;
        RECT 243.930 171.670 245.480 172.520 ;
        RECT 245.820 171.670 247.370 172.520 ;
        RECT 345.350 172.330 346.640 173.290 ;
        RECT 347.240 172.330 348.530 173.290 ;
        RECT 345.240 171.480 346.790 172.330 ;
        RECT 347.130 171.480 348.680 172.330 ;
        RECT 23.190 170.160 24.480 171.120 ;
        RECT 25.080 170.160 26.370 171.120 ;
        RECT 23.080 169.310 24.630 170.160 ;
        RECT 24.970 169.310 26.520 170.160 ;
        RECT 124.500 169.970 125.790 170.930 ;
        RECT 126.390 169.970 127.680 170.930 ;
        RECT 259.720 170.100 261.010 171.060 ;
        RECT 261.610 170.100 262.900 171.060 ;
        RECT 124.390 169.120 125.940 169.970 ;
        RECT 126.280 169.120 127.830 169.970 ;
        RECT 259.610 169.250 261.160 170.100 ;
        RECT 261.500 169.250 263.050 170.100 ;
        RECT 361.030 169.910 362.320 170.870 ;
        RECT 362.920 169.910 364.210 170.870 ;
        RECT 360.920 169.060 362.470 169.910 ;
        RECT 362.810 169.060 364.360 169.910 ;
        RECT 7.670 166.180 8.960 167.140 ;
        RECT 9.560 166.180 10.850 167.140 ;
        RECT 7.560 165.330 9.110 166.180 ;
        RECT 9.450 165.330 11.000 166.180 ;
        RECT 108.980 165.990 110.270 166.950 ;
        RECT 110.870 165.990 112.160 166.950 ;
        RECT 244.200 166.120 245.490 167.080 ;
        RECT 246.090 166.120 247.380 167.080 ;
        RECT 108.870 165.140 110.420 165.990 ;
        RECT 110.760 165.140 112.310 165.990 ;
        RECT 244.090 165.270 245.640 166.120 ;
        RECT 245.980 165.270 247.530 166.120 ;
        RECT 345.510 165.930 346.800 166.890 ;
        RECT 347.400 165.930 348.690 166.890 ;
        RECT 345.400 165.080 346.950 165.930 ;
        RECT 347.290 165.080 348.840 165.930 ;
        RECT 58.470 163.010 59.760 163.970 ;
        RECT 60.360 163.010 61.650 163.970 ;
        RECT 58.360 162.160 59.910 163.010 ;
        RECT 60.250 162.160 61.800 163.010 ;
        RECT 159.780 162.820 161.070 163.780 ;
        RECT 161.670 162.820 162.960 163.780 ;
        RECT 295.000 162.950 296.290 163.910 ;
        RECT 296.890 162.950 298.180 163.910 ;
        RECT 159.670 161.970 161.220 162.820 ;
        RECT 161.560 161.970 163.110 162.820 ;
        RECT 294.890 162.100 296.440 162.950 ;
        RECT 296.780 162.100 298.330 162.950 ;
        RECT 396.310 162.760 397.600 163.720 ;
        RECT 398.200 162.760 399.490 163.720 ;
        RECT 396.200 161.910 397.750 162.760 ;
        RECT 398.090 161.910 399.640 162.760 ;
        RECT 7.650 156.930 8.940 157.890 ;
        RECT 9.540 156.930 10.830 157.890 ;
        RECT 7.540 156.080 9.090 156.930 ;
        RECT 9.430 156.080 10.980 156.930 ;
        RECT 108.960 156.740 110.250 157.700 ;
        RECT 110.850 156.740 112.140 157.700 ;
        RECT 244.180 156.870 245.470 157.830 ;
        RECT 246.070 156.870 247.360 157.830 ;
        RECT 108.850 155.890 110.400 156.740 ;
        RECT 110.740 155.890 112.290 156.740 ;
        RECT 244.070 156.020 245.620 156.870 ;
        RECT 245.960 156.020 247.510 156.870 ;
        RECT 345.490 156.680 346.780 157.640 ;
        RECT 347.380 156.680 348.670 157.640 ;
        RECT 345.380 155.830 346.930 156.680 ;
        RECT 347.270 155.830 348.820 156.680 ;
        RECT 23.330 154.510 24.620 155.470 ;
        RECT 25.220 154.510 26.510 155.470 ;
        RECT 23.220 153.660 24.770 154.510 ;
        RECT 25.110 153.660 26.660 154.510 ;
        RECT 124.640 154.320 125.930 155.280 ;
        RECT 126.530 154.320 127.820 155.280 ;
        RECT 259.860 154.450 261.150 155.410 ;
        RECT 261.750 154.450 263.040 155.410 ;
        RECT 124.530 153.470 126.080 154.320 ;
        RECT 126.420 153.470 127.970 154.320 ;
        RECT 259.750 153.600 261.300 154.450 ;
        RECT 261.640 153.600 263.190 154.450 ;
        RECT 361.170 154.260 362.460 155.220 ;
        RECT 363.060 154.260 364.350 155.220 ;
        RECT 361.060 153.410 362.610 154.260 ;
        RECT 362.950 153.410 364.500 154.260 ;
        RECT 7.810 150.530 9.100 151.490 ;
        RECT 9.700 150.530 10.990 151.490 ;
        RECT 7.700 149.680 9.250 150.530 ;
        RECT 9.590 149.680 11.140 150.530 ;
        RECT 109.120 150.340 110.410 151.300 ;
        RECT 111.010 150.340 112.300 151.300 ;
        RECT 244.340 150.470 245.630 151.430 ;
        RECT 246.230 150.470 247.520 151.430 ;
        RECT 40.910 148.960 42.200 149.920 ;
        RECT 42.800 148.960 44.090 149.920 ;
        RECT 109.010 149.490 110.560 150.340 ;
        RECT 110.900 149.490 112.450 150.340 ;
        RECT 40.800 148.110 42.350 148.960 ;
        RECT 42.690 148.110 44.240 148.960 ;
        RECT 142.220 148.770 143.510 149.730 ;
        RECT 144.110 148.770 145.400 149.730 ;
        RECT 244.230 149.620 245.780 150.470 ;
        RECT 246.120 149.620 247.670 150.470 ;
        RECT 345.650 150.280 346.940 151.240 ;
        RECT 347.540 150.280 348.830 151.240 ;
        RECT 277.440 148.900 278.730 149.860 ;
        RECT 279.330 148.900 280.620 149.860 ;
        RECT 345.540 149.430 347.090 150.280 ;
        RECT 347.430 149.430 348.980 150.280 ;
        RECT 142.110 147.920 143.660 148.770 ;
        RECT 144.000 147.920 145.550 148.770 ;
        RECT 277.330 148.050 278.880 148.900 ;
        RECT 279.220 148.050 280.770 148.900 ;
        RECT 378.750 148.710 380.040 149.670 ;
        RECT 380.640 148.710 381.930 149.670 ;
        RECT 378.640 147.860 380.190 148.710 ;
        RECT 380.530 147.860 382.080 148.710 ;
        RECT 7.480 142.510 8.770 143.470 ;
        RECT 9.370 142.510 10.660 143.470 ;
        RECT 7.370 141.660 8.920 142.510 ;
        RECT 9.260 141.660 10.810 142.510 ;
        RECT 108.790 142.320 110.080 143.280 ;
        RECT 110.680 142.320 111.970 143.280 ;
        RECT 244.010 142.450 245.300 143.410 ;
        RECT 245.900 142.450 247.190 143.410 ;
        RECT 108.680 141.470 110.230 142.320 ;
        RECT 110.570 141.470 112.120 142.320 ;
        RECT 243.900 141.600 245.450 142.450 ;
        RECT 245.790 141.600 247.340 142.450 ;
        RECT 345.320 142.260 346.610 143.220 ;
        RECT 347.210 142.260 348.500 143.220 ;
        RECT 345.210 141.410 346.760 142.260 ;
        RECT 347.100 141.410 348.650 142.260 ;
        RECT 23.160 140.090 24.450 141.050 ;
        RECT 25.050 140.090 26.340 141.050 ;
        RECT 23.050 139.240 24.600 140.090 ;
        RECT 24.940 139.240 26.490 140.090 ;
        RECT 124.470 139.900 125.760 140.860 ;
        RECT 126.360 139.900 127.650 140.860 ;
        RECT 259.690 140.030 260.980 140.990 ;
        RECT 261.580 140.030 262.870 140.990 ;
        RECT 124.360 139.050 125.910 139.900 ;
        RECT 126.250 139.050 127.800 139.900 ;
        RECT 259.580 139.180 261.130 140.030 ;
        RECT 261.470 139.180 263.020 140.030 ;
        RECT 361.000 139.840 362.290 140.800 ;
        RECT 362.890 139.840 364.180 140.800 ;
        RECT 360.890 138.990 362.440 139.840 ;
        RECT 362.780 138.990 364.330 139.840 ;
        RECT 7.640 136.110 8.930 137.070 ;
        RECT 9.530 136.110 10.820 137.070 ;
        RECT 7.530 135.260 9.080 136.110 ;
        RECT 9.420 135.260 10.970 136.110 ;
        RECT 108.950 135.920 110.240 136.880 ;
        RECT 110.840 135.920 112.130 136.880 ;
        RECT 108.840 135.070 110.390 135.920 ;
        RECT 110.730 135.070 112.280 135.920 ;
        RECT 216.940 135.640 218.230 136.600 ;
        RECT 218.830 135.640 220.120 136.600 ;
        RECT 244.170 136.050 245.460 137.010 ;
        RECT 246.060 136.050 247.350 137.010 ;
        RECT 216.830 134.790 218.380 135.640 ;
        RECT 218.720 134.790 220.270 135.640 ;
        RECT 244.060 135.200 245.610 136.050 ;
        RECT 245.950 135.200 247.500 136.050 ;
        RECT 345.480 135.860 346.770 136.820 ;
        RECT 347.370 135.860 348.660 136.820 ;
        RECT 345.370 135.010 346.920 135.860 ;
        RECT 347.260 135.010 348.810 135.860 ;
        RECT 453.470 135.580 454.760 136.540 ;
        RECT 455.360 135.580 456.650 136.540 ;
        RECT 453.360 134.730 454.910 135.580 ;
        RECT 455.250 134.730 456.800 135.580 ;
        RECT 89.350 133.500 90.640 134.460 ;
        RECT 91.240 133.500 92.530 134.460 ;
        RECT 89.240 132.650 90.790 133.500 ;
        RECT 91.130 132.650 92.680 133.500 ;
        RECT 190.660 133.310 191.950 134.270 ;
        RECT 192.550 133.310 193.840 134.270 ;
        RECT 325.880 133.440 327.170 134.400 ;
        RECT 327.770 133.440 329.060 134.400 ;
        RECT 190.550 132.460 192.100 133.310 ;
        RECT 192.440 132.460 193.990 133.310 ;
        RECT 325.770 132.590 327.320 133.440 ;
        RECT 327.660 132.590 329.210 133.440 ;
        RECT 427.190 133.250 428.480 134.210 ;
        RECT 429.080 133.250 430.370 134.210 ;
        RECT 427.080 132.400 428.630 133.250 ;
        RECT 428.970 132.400 430.520 133.250 ;
        RECT 470.770 133.230 472.060 134.190 ;
        RECT 472.660 133.230 473.950 134.190 ;
        RECT 470.660 132.380 472.210 133.230 ;
        RECT 472.550 132.380 474.100 133.230 ;
        RECT 7.530 126.680 8.820 127.640 ;
        RECT 9.420 126.680 10.710 127.640 ;
        RECT 7.420 125.830 8.970 126.680 ;
        RECT 9.310 125.830 10.860 126.680 ;
        RECT 108.840 126.490 110.130 127.450 ;
        RECT 110.730 126.490 112.020 127.450 ;
        RECT 244.060 126.620 245.350 127.580 ;
        RECT 245.950 126.620 247.240 127.580 ;
        RECT 108.730 125.640 110.280 126.490 ;
        RECT 110.620 125.640 112.170 126.490 ;
        RECT 243.950 125.770 245.500 126.620 ;
        RECT 245.840 125.770 247.390 126.620 ;
        RECT 345.370 126.430 346.660 127.390 ;
        RECT 347.260 126.430 348.550 127.390 ;
        RECT 345.260 125.580 346.810 126.430 ;
        RECT 347.150 125.580 348.700 126.430 ;
        RECT 23.210 124.260 24.500 125.220 ;
        RECT 25.100 124.260 26.390 125.220 ;
        RECT 23.100 123.410 24.650 124.260 ;
        RECT 24.990 123.410 26.540 124.260 ;
        RECT 124.520 124.070 125.810 125.030 ;
        RECT 126.410 124.070 127.700 125.030 ;
        RECT 259.740 124.200 261.030 125.160 ;
        RECT 261.630 124.200 262.920 125.160 ;
        RECT 124.410 123.220 125.960 124.070 ;
        RECT 126.300 123.220 127.850 124.070 ;
        RECT 259.630 123.350 261.180 124.200 ;
        RECT 261.520 123.350 263.070 124.200 ;
        RECT 361.050 124.010 362.340 124.970 ;
        RECT 362.940 124.010 364.230 124.970 ;
        RECT 360.940 123.160 362.490 124.010 ;
        RECT 362.830 123.160 364.380 124.010 ;
        RECT 7.690 120.280 8.980 121.240 ;
        RECT 9.580 120.280 10.870 121.240 ;
        RECT 7.580 119.430 9.130 120.280 ;
        RECT 9.470 119.430 11.020 120.280 ;
        RECT 109.000 120.090 110.290 121.050 ;
        RECT 110.890 120.090 112.180 121.050 ;
        RECT 244.220 120.220 245.510 121.180 ;
        RECT 246.110 120.220 247.400 121.180 ;
        RECT 40.790 118.710 42.080 119.670 ;
        RECT 42.680 118.710 43.970 119.670 ;
        RECT 108.890 119.240 110.440 120.090 ;
        RECT 110.780 119.240 112.330 120.090 ;
        RECT 40.680 117.860 42.230 118.710 ;
        RECT 42.570 117.860 44.120 118.710 ;
        RECT 142.100 118.520 143.390 119.480 ;
        RECT 143.990 118.520 145.280 119.480 ;
        RECT 244.110 119.370 245.660 120.220 ;
        RECT 246.000 119.370 247.550 120.220 ;
        RECT 345.530 120.030 346.820 120.990 ;
        RECT 347.420 120.030 348.710 120.990 ;
        RECT 277.320 118.650 278.610 119.610 ;
        RECT 279.210 118.650 280.500 119.610 ;
        RECT 345.420 119.180 346.970 120.030 ;
        RECT 347.310 119.180 348.860 120.030 ;
        RECT 141.990 117.670 143.540 118.520 ;
        RECT 143.880 117.670 145.430 118.520 ;
        RECT 277.210 117.800 278.760 118.650 ;
        RECT 279.100 117.800 280.650 118.650 ;
        RECT 378.630 118.460 379.920 119.420 ;
        RECT 380.520 118.460 381.810 119.420 ;
        RECT 378.520 117.610 380.070 118.460 ;
        RECT 380.410 117.610 381.960 118.460 ;
        RECT 7.360 112.260 8.650 113.220 ;
        RECT 9.250 112.260 10.540 113.220 ;
        RECT 7.250 111.410 8.800 112.260 ;
        RECT 9.140 111.410 10.690 112.260 ;
        RECT 108.670 112.070 109.960 113.030 ;
        RECT 110.560 112.070 111.850 113.030 ;
        RECT 243.890 112.200 245.180 113.160 ;
        RECT 245.780 112.200 247.070 113.160 ;
        RECT 108.560 111.220 110.110 112.070 ;
        RECT 110.450 111.220 112.000 112.070 ;
        RECT 243.780 111.350 245.330 112.200 ;
        RECT 245.670 111.350 247.220 112.200 ;
        RECT 345.200 112.010 346.490 112.970 ;
        RECT 347.090 112.010 348.380 112.970 ;
        RECT 345.090 111.160 346.640 112.010 ;
        RECT 346.980 111.160 348.530 112.010 ;
        RECT 23.040 109.840 24.330 110.800 ;
        RECT 24.930 109.840 26.220 110.800 ;
        RECT 22.930 108.990 24.480 109.840 ;
        RECT 24.820 108.990 26.370 109.840 ;
        RECT 124.350 109.650 125.640 110.610 ;
        RECT 126.240 109.650 127.530 110.610 ;
        RECT 259.570 109.780 260.860 110.740 ;
        RECT 261.460 109.780 262.750 110.740 ;
        RECT 124.240 108.800 125.790 109.650 ;
        RECT 126.130 108.800 127.680 109.650 ;
        RECT 259.460 108.930 261.010 109.780 ;
        RECT 261.350 108.930 262.900 109.780 ;
        RECT 360.880 109.590 362.170 110.550 ;
        RECT 362.770 109.590 364.060 110.550 ;
        RECT 360.770 108.740 362.320 109.590 ;
        RECT 362.660 108.740 364.210 109.590 ;
        RECT 7.520 105.860 8.810 106.820 ;
        RECT 9.410 105.860 10.700 106.820 ;
        RECT 7.410 105.010 8.960 105.860 ;
        RECT 9.300 105.010 10.850 105.860 ;
        RECT 108.830 105.670 110.120 106.630 ;
        RECT 110.720 105.670 112.010 106.630 ;
        RECT 244.050 105.800 245.340 106.760 ;
        RECT 245.940 105.800 247.230 106.760 ;
        RECT 108.720 104.820 110.270 105.670 ;
        RECT 110.610 104.820 112.160 105.670 ;
        RECT 243.940 104.950 245.490 105.800 ;
        RECT 245.830 104.950 247.380 105.800 ;
        RECT 345.360 105.610 346.650 106.570 ;
        RECT 347.250 105.610 348.540 106.570 ;
        RECT 345.250 104.760 346.800 105.610 ;
        RECT 347.140 104.760 348.690 105.610 ;
        RECT 58.320 102.690 59.610 103.650 ;
        RECT 60.210 102.690 61.500 103.650 ;
        RECT 58.210 101.840 59.760 102.690 ;
        RECT 60.100 101.840 61.650 102.690 ;
        RECT 159.630 102.500 160.920 103.460 ;
        RECT 161.520 102.500 162.810 103.460 ;
        RECT 294.850 102.630 296.140 103.590 ;
        RECT 296.740 102.630 298.030 103.590 ;
        RECT 159.520 101.650 161.070 102.500 ;
        RECT 161.410 101.650 162.960 102.500 ;
        RECT 294.740 101.780 296.290 102.630 ;
        RECT 296.630 101.780 298.180 102.630 ;
        RECT 396.160 102.440 397.450 103.400 ;
        RECT 398.050 102.440 399.340 103.400 ;
        RECT 396.050 101.590 397.600 102.440 ;
        RECT 397.940 101.590 399.490 102.440 ;
        RECT 7.500 96.610 8.790 97.570 ;
        RECT 9.390 96.610 10.680 97.570 ;
        RECT 7.390 95.760 8.940 96.610 ;
        RECT 9.280 95.760 10.830 96.610 ;
        RECT 108.810 96.420 110.100 97.380 ;
        RECT 110.700 96.420 111.990 97.380 ;
        RECT 244.030 96.550 245.320 97.510 ;
        RECT 245.920 96.550 247.210 97.510 ;
        RECT 108.700 95.570 110.250 96.420 ;
        RECT 110.590 95.570 112.140 96.420 ;
        RECT 243.920 95.700 245.470 96.550 ;
        RECT 245.810 95.700 247.360 96.550 ;
        RECT 345.340 96.360 346.630 97.320 ;
        RECT 347.230 96.360 348.520 97.320 ;
        RECT 345.230 95.510 346.780 96.360 ;
        RECT 347.120 95.510 348.670 96.360 ;
        RECT 23.180 94.190 24.470 95.150 ;
        RECT 25.070 94.190 26.360 95.150 ;
        RECT 23.070 93.340 24.620 94.190 ;
        RECT 24.960 93.340 26.510 94.190 ;
        RECT 124.490 94.000 125.780 94.960 ;
        RECT 126.380 94.000 127.670 94.960 ;
        RECT 259.710 94.130 261.000 95.090 ;
        RECT 261.600 94.130 262.890 95.090 ;
        RECT 124.380 93.150 125.930 94.000 ;
        RECT 126.270 93.150 127.820 94.000 ;
        RECT 259.600 93.280 261.150 94.130 ;
        RECT 261.490 93.280 263.040 94.130 ;
        RECT 361.020 93.940 362.310 94.900 ;
        RECT 362.910 93.940 364.200 94.900 ;
        RECT 360.910 93.090 362.460 93.940 ;
        RECT 362.800 93.090 364.350 93.940 ;
        RECT 7.660 90.210 8.950 91.170 ;
        RECT 9.550 90.210 10.840 91.170 ;
        RECT 7.550 89.360 9.100 90.210 ;
        RECT 9.440 89.360 10.990 90.210 ;
        RECT 108.970 90.020 110.260 90.980 ;
        RECT 110.860 90.020 112.150 90.980 ;
        RECT 244.190 90.150 245.480 91.110 ;
        RECT 246.080 90.150 247.370 91.110 ;
        RECT 40.760 88.640 42.050 89.600 ;
        RECT 42.650 88.640 43.940 89.600 ;
        RECT 108.860 89.170 110.410 90.020 ;
        RECT 110.750 89.170 112.300 90.020 ;
        RECT 40.650 87.790 42.200 88.640 ;
        RECT 42.540 87.790 44.090 88.640 ;
        RECT 142.070 88.450 143.360 89.410 ;
        RECT 143.960 88.450 145.250 89.410 ;
        RECT 244.080 89.300 245.630 90.150 ;
        RECT 245.970 89.300 247.520 90.150 ;
        RECT 345.500 89.960 346.790 90.920 ;
        RECT 347.390 89.960 348.680 90.920 ;
        RECT 277.290 88.580 278.580 89.540 ;
        RECT 279.180 88.580 280.470 89.540 ;
        RECT 345.390 89.110 346.940 89.960 ;
        RECT 347.280 89.110 348.830 89.960 ;
        RECT 141.960 87.600 143.510 88.450 ;
        RECT 143.850 87.600 145.400 88.450 ;
        RECT 277.180 87.730 278.730 88.580 ;
        RECT 279.070 87.730 280.620 88.580 ;
        RECT 378.600 88.390 379.890 89.350 ;
        RECT 380.490 88.390 381.780 89.350 ;
        RECT 378.490 87.540 380.040 88.390 ;
        RECT 380.380 87.540 381.930 88.390 ;
        RECT 7.330 82.190 8.620 83.150 ;
        RECT 9.220 82.190 10.510 83.150 ;
        RECT 7.220 81.340 8.770 82.190 ;
        RECT 9.110 81.340 10.660 82.190 ;
        RECT 108.640 82.000 109.930 82.960 ;
        RECT 110.530 82.000 111.820 82.960 ;
        RECT 243.860 82.130 245.150 83.090 ;
        RECT 245.750 82.130 247.040 83.090 ;
        RECT 108.530 81.150 110.080 82.000 ;
        RECT 110.420 81.150 111.970 82.000 ;
        RECT 243.750 81.280 245.300 82.130 ;
        RECT 245.640 81.280 247.190 82.130 ;
        RECT 345.170 81.940 346.460 82.900 ;
        RECT 347.060 81.940 348.350 82.900 ;
        RECT 345.060 81.090 346.610 81.940 ;
        RECT 346.950 81.090 348.500 81.940 ;
        RECT 23.010 79.770 24.300 80.730 ;
        RECT 24.900 79.770 26.190 80.730 ;
        RECT 22.900 78.920 24.450 79.770 ;
        RECT 24.790 78.920 26.340 79.770 ;
        RECT 124.320 79.580 125.610 80.540 ;
        RECT 126.210 79.580 127.500 80.540 ;
        RECT 259.540 79.710 260.830 80.670 ;
        RECT 261.430 79.710 262.720 80.670 ;
        RECT 124.210 78.730 125.760 79.580 ;
        RECT 126.100 78.730 127.650 79.580 ;
        RECT 259.430 78.860 260.980 79.710 ;
        RECT 261.320 78.860 262.870 79.710 ;
        RECT 360.850 79.520 362.140 80.480 ;
        RECT 362.740 79.520 364.030 80.480 ;
        RECT 360.740 78.670 362.290 79.520 ;
        RECT 362.630 78.670 364.180 79.520 ;
        RECT 7.490 75.790 8.780 76.750 ;
        RECT 9.380 75.790 10.670 76.750 ;
        RECT 72.520 76.400 73.810 77.360 ;
        RECT 74.410 76.400 75.700 77.360 ;
        RECT 7.380 74.940 8.930 75.790 ;
        RECT 9.270 74.940 10.820 75.790 ;
        RECT 72.410 75.550 73.960 76.400 ;
        RECT 74.300 75.550 75.850 76.400 ;
        RECT 108.800 75.600 110.090 76.560 ;
        RECT 110.690 75.600 111.980 76.560 ;
        RECT 173.830 76.210 175.120 77.170 ;
        RECT 175.720 76.210 177.010 77.170 ;
        RECT 108.690 74.750 110.240 75.600 ;
        RECT 110.580 74.750 112.130 75.600 ;
        RECT 173.720 75.360 175.270 76.210 ;
        RECT 175.610 75.360 177.160 76.210 ;
        RECT 244.020 75.730 245.310 76.690 ;
        RECT 245.910 75.730 247.200 76.690 ;
        RECT 309.050 76.340 310.340 77.300 ;
        RECT 310.940 76.340 312.230 77.300 ;
        RECT 243.910 74.880 245.460 75.730 ;
        RECT 245.800 74.880 247.350 75.730 ;
        RECT 308.940 75.490 310.490 76.340 ;
        RECT 310.830 75.490 312.380 76.340 ;
        RECT 345.330 75.540 346.620 76.500 ;
        RECT 347.220 75.540 348.510 76.500 ;
        RECT 410.360 76.150 411.650 77.110 ;
        RECT 412.250 76.150 413.540 77.110 ;
        RECT 345.220 74.690 346.770 75.540 ;
        RECT 347.110 74.690 348.660 75.540 ;
        RECT 410.250 75.300 411.800 76.150 ;
        RECT 412.140 75.300 413.690 76.150 ;
        RECT 7.180 66.760 8.470 67.720 ;
        RECT 9.070 66.760 10.360 67.720 ;
        RECT 7.070 65.910 8.620 66.760 ;
        RECT 8.960 65.910 10.510 66.760 ;
        RECT 108.490 66.570 109.780 67.530 ;
        RECT 110.380 66.570 111.670 67.530 ;
        RECT 243.710 66.700 245.000 67.660 ;
        RECT 245.600 66.700 246.890 67.660 ;
        RECT 108.380 65.720 109.930 66.570 ;
        RECT 110.270 65.720 111.820 66.570 ;
        RECT 243.600 65.850 245.150 66.700 ;
        RECT 245.490 65.850 247.040 66.700 ;
        RECT 345.020 66.510 346.310 67.470 ;
        RECT 346.910 66.510 348.200 67.470 ;
        RECT 344.910 65.660 346.460 66.510 ;
        RECT 346.800 65.660 348.350 66.510 ;
        RECT 22.860 64.340 24.150 65.300 ;
        RECT 24.750 64.340 26.040 65.300 ;
        RECT 22.750 63.490 24.300 64.340 ;
        RECT 24.640 63.490 26.190 64.340 ;
        RECT 124.170 64.150 125.460 65.110 ;
        RECT 126.060 64.150 127.350 65.110 ;
        RECT 259.390 64.280 260.680 65.240 ;
        RECT 261.280 64.280 262.570 65.240 ;
        RECT 124.060 63.300 125.610 64.150 ;
        RECT 125.950 63.300 127.500 64.150 ;
        RECT 259.280 63.430 260.830 64.280 ;
        RECT 261.170 63.430 262.720 64.280 ;
        RECT 360.700 64.090 361.990 65.050 ;
        RECT 362.590 64.090 363.880 65.050 ;
        RECT 360.590 63.240 362.140 64.090 ;
        RECT 362.480 63.240 364.030 64.090 ;
        RECT 7.340 60.360 8.630 61.320 ;
        RECT 9.230 60.360 10.520 61.320 ;
        RECT 7.230 59.510 8.780 60.360 ;
        RECT 9.120 59.510 10.670 60.360 ;
        RECT 108.650 60.170 109.940 61.130 ;
        RECT 110.540 60.170 111.830 61.130 ;
        RECT 243.870 60.300 245.160 61.260 ;
        RECT 245.760 60.300 247.050 61.260 ;
        RECT 40.440 58.790 41.730 59.750 ;
        RECT 42.330 58.790 43.620 59.750 ;
        RECT 108.540 59.320 110.090 60.170 ;
        RECT 110.430 59.320 111.980 60.170 ;
        RECT 40.330 57.940 41.880 58.790 ;
        RECT 42.220 57.940 43.770 58.790 ;
        RECT 141.750 58.600 143.040 59.560 ;
        RECT 143.640 58.600 144.930 59.560 ;
        RECT 243.760 59.450 245.310 60.300 ;
        RECT 245.650 59.450 247.200 60.300 ;
        RECT 345.180 60.110 346.470 61.070 ;
        RECT 347.070 60.110 348.360 61.070 ;
        RECT 276.970 58.730 278.260 59.690 ;
        RECT 278.860 58.730 280.150 59.690 ;
        RECT 345.070 59.260 346.620 60.110 ;
        RECT 346.960 59.260 348.510 60.110 ;
        RECT 141.640 57.750 143.190 58.600 ;
        RECT 143.530 57.750 145.080 58.600 ;
        RECT 276.860 57.880 278.410 58.730 ;
        RECT 278.750 57.880 280.300 58.730 ;
        RECT 378.280 58.540 379.570 59.500 ;
        RECT 380.170 58.540 381.460 59.500 ;
        RECT 378.170 57.690 379.720 58.540 ;
        RECT 380.060 57.690 381.610 58.540 ;
        RECT 7.010 52.340 8.300 53.300 ;
        RECT 8.900 52.340 10.190 53.300 ;
        RECT 6.900 51.490 8.450 52.340 ;
        RECT 8.790 51.490 10.340 52.340 ;
        RECT 108.320 52.150 109.610 53.110 ;
        RECT 110.210 52.150 111.500 53.110 ;
        RECT 243.540 52.280 244.830 53.240 ;
        RECT 245.430 52.280 246.720 53.240 ;
        RECT 108.210 51.300 109.760 52.150 ;
        RECT 110.100 51.300 111.650 52.150 ;
        RECT 243.430 51.430 244.980 52.280 ;
        RECT 245.320 51.430 246.870 52.280 ;
        RECT 344.850 52.090 346.140 53.050 ;
        RECT 346.740 52.090 348.030 53.050 ;
        RECT 344.740 51.240 346.290 52.090 ;
        RECT 346.630 51.240 348.180 52.090 ;
        RECT 22.690 49.920 23.980 50.880 ;
        RECT 24.580 49.920 25.870 50.880 ;
        RECT 22.580 49.070 24.130 49.920 ;
        RECT 24.470 49.070 26.020 49.920 ;
        RECT 124.000 49.730 125.290 50.690 ;
        RECT 125.890 49.730 127.180 50.690 ;
        RECT 259.220 49.860 260.510 50.820 ;
        RECT 261.110 49.860 262.400 50.820 ;
        RECT 123.890 48.880 125.440 49.730 ;
        RECT 125.780 48.880 127.330 49.730 ;
        RECT 259.110 49.010 260.660 49.860 ;
        RECT 261.000 49.010 262.550 49.860 ;
        RECT 360.530 49.670 361.820 50.630 ;
        RECT 362.420 49.670 363.710 50.630 ;
        RECT 360.420 48.820 361.970 49.670 ;
        RECT 362.310 48.820 363.860 49.670 ;
        RECT 7.170 45.940 8.460 46.900 ;
        RECT 9.060 45.940 10.350 46.900 ;
        RECT 7.060 45.090 8.610 45.940 ;
        RECT 8.950 45.090 10.500 45.940 ;
        RECT 108.480 45.750 109.770 46.710 ;
        RECT 110.370 45.750 111.660 46.710 ;
        RECT 243.700 45.880 244.990 46.840 ;
        RECT 245.590 45.880 246.880 46.840 ;
        RECT 108.370 44.900 109.920 45.750 ;
        RECT 110.260 44.900 111.810 45.750 ;
        RECT 243.590 45.030 245.140 45.880 ;
        RECT 245.480 45.030 247.030 45.880 ;
        RECT 345.010 45.690 346.300 46.650 ;
        RECT 346.900 45.690 348.190 46.650 ;
        RECT 344.900 44.840 346.450 45.690 ;
        RECT 346.790 44.840 348.340 45.690 ;
        RECT 57.970 42.770 59.260 43.730 ;
        RECT 59.860 42.770 61.150 43.730 ;
        RECT 57.860 41.920 59.410 42.770 ;
        RECT 59.750 41.920 61.300 42.770 ;
        RECT 159.280 42.580 160.570 43.540 ;
        RECT 161.170 42.580 162.460 43.540 ;
        RECT 294.500 42.710 295.790 43.670 ;
        RECT 296.390 42.710 297.680 43.670 ;
        RECT 159.170 41.730 160.720 42.580 ;
        RECT 161.060 41.730 162.610 42.580 ;
        RECT 294.390 41.860 295.940 42.710 ;
        RECT 296.280 41.860 297.830 42.710 ;
        RECT 395.810 42.520 397.100 43.480 ;
        RECT 397.700 42.520 398.990 43.480 ;
        RECT 395.700 41.670 397.250 42.520 ;
        RECT 397.590 41.670 399.140 42.520 ;
        RECT 7.150 36.690 8.440 37.650 ;
        RECT 9.040 36.690 10.330 37.650 ;
        RECT 7.040 35.840 8.590 36.690 ;
        RECT 8.930 35.840 10.480 36.690 ;
        RECT 108.460 36.500 109.750 37.460 ;
        RECT 110.350 36.500 111.640 37.460 ;
        RECT 243.680 36.630 244.970 37.590 ;
        RECT 245.570 36.630 246.860 37.590 ;
        RECT 108.350 35.650 109.900 36.500 ;
        RECT 110.240 35.650 111.790 36.500 ;
        RECT 243.570 35.780 245.120 36.630 ;
        RECT 245.460 35.780 247.010 36.630 ;
        RECT 344.990 36.440 346.280 37.400 ;
        RECT 346.880 36.440 348.170 37.400 ;
        RECT 344.880 35.590 346.430 36.440 ;
        RECT 346.770 35.590 348.320 36.440 ;
        RECT 22.830 34.270 24.120 35.230 ;
        RECT 24.720 34.270 26.010 35.230 ;
        RECT 22.720 33.420 24.270 34.270 ;
        RECT 24.610 33.420 26.160 34.270 ;
        RECT 124.140 34.080 125.430 35.040 ;
        RECT 126.030 34.080 127.320 35.040 ;
        RECT 259.360 34.210 260.650 35.170 ;
        RECT 261.250 34.210 262.540 35.170 ;
        RECT 124.030 33.230 125.580 34.080 ;
        RECT 125.920 33.230 127.470 34.080 ;
        RECT 259.250 33.360 260.800 34.210 ;
        RECT 261.140 33.360 262.690 34.210 ;
        RECT 360.670 34.020 361.960 34.980 ;
        RECT 362.560 34.020 363.850 34.980 ;
        RECT 360.560 33.170 362.110 34.020 ;
        RECT 362.450 33.170 364.000 34.020 ;
        RECT 7.310 30.290 8.600 31.250 ;
        RECT 9.200 30.290 10.490 31.250 ;
        RECT 7.200 29.440 8.750 30.290 ;
        RECT 9.090 29.440 10.640 30.290 ;
        RECT 108.620 30.100 109.910 31.060 ;
        RECT 110.510 30.100 111.800 31.060 ;
        RECT 243.840 30.230 245.130 31.190 ;
        RECT 245.730 30.230 247.020 31.190 ;
        RECT 40.410 28.720 41.700 29.680 ;
        RECT 42.300 28.720 43.590 29.680 ;
        RECT 108.510 29.250 110.060 30.100 ;
        RECT 110.400 29.250 111.950 30.100 ;
        RECT 40.300 27.870 41.850 28.720 ;
        RECT 42.190 27.870 43.740 28.720 ;
        RECT 141.720 28.530 143.010 29.490 ;
        RECT 143.610 28.530 144.900 29.490 ;
        RECT 243.730 29.380 245.280 30.230 ;
        RECT 245.620 29.380 247.170 30.230 ;
        RECT 345.150 30.040 346.440 31.000 ;
        RECT 347.040 30.040 348.330 31.000 ;
        RECT 276.940 28.660 278.230 29.620 ;
        RECT 278.830 28.660 280.120 29.620 ;
        RECT 345.040 29.190 346.590 30.040 ;
        RECT 346.930 29.190 348.480 30.040 ;
        RECT 141.610 27.680 143.160 28.530 ;
        RECT 143.500 27.680 145.050 28.530 ;
        RECT 276.830 27.810 278.380 28.660 ;
        RECT 278.720 27.810 280.270 28.660 ;
        RECT 378.250 28.470 379.540 29.430 ;
        RECT 380.140 28.470 381.430 29.430 ;
        RECT 378.140 27.620 379.690 28.470 ;
        RECT 380.030 27.620 381.580 28.470 ;
        RECT 6.980 22.270 8.270 23.230 ;
        RECT 8.870 22.270 10.160 23.230 ;
        RECT 6.870 21.420 8.420 22.270 ;
        RECT 8.760 21.420 10.310 22.270 ;
        RECT 108.290 22.080 109.580 23.040 ;
        RECT 110.180 22.080 111.470 23.040 ;
        RECT 243.510 22.210 244.800 23.170 ;
        RECT 245.400 22.210 246.690 23.170 ;
        RECT 108.180 21.230 109.730 22.080 ;
        RECT 110.070 21.230 111.620 22.080 ;
        RECT 243.400 21.360 244.950 22.210 ;
        RECT 245.290 21.360 246.840 22.210 ;
        RECT 344.820 22.020 346.110 22.980 ;
        RECT 346.710 22.020 348.000 22.980 ;
        RECT 344.710 21.170 346.260 22.020 ;
        RECT 346.600 21.170 348.150 22.020 ;
        RECT 22.660 19.850 23.950 20.810 ;
        RECT 24.550 19.850 25.840 20.810 ;
        RECT 22.550 19.000 24.100 19.850 ;
        RECT 24.440 19.000 25.990 19.850 ;
        RECT 123.970 19.660 125.260 20.620 ;
        RECT 125.860 19.660 127.150 20.620 ;
        RECT 259.190 19.790 260.480 20.750 ;
        RECT 261.080 19.790 262.370 20.750 ;
        RECT 123.860 18.810 125.410 19.660 ;
        RECT 125.750 18.810 127.300 19.660 ;
        RECT 259.080 18.940 260.630 19.790 ;
        RECT 260.970 18.940 262.520 19.790 ;
        RECT 360.500 19.600 361.790 20.560 ;
        RECT 362.390 19.600 363.680 20.560 ;
        RECT 360.390 18.750 361.940 19.600 ;
        RECT 362.280 18.750 363.830 19.600 ;
        RECT 7.140 15.870 8.430 16.830 ;
        RECT 9.030 15.870 10.320 16.830 ;
        RECT 7.030 15.020 8.580 15.870 ;
        RECT 8.920 15.020 10.470 15.870 ;
        RECT 108.450 15.680 109.740 16.640 ;
        RECT 110.340 15.680 111.630 16.640 ;
        RECT 243.670 15.810 244.960 16.770 ;
        RECT 245.560 15.810 246.850 16.770 ;
        RECT 108.340 14.830 109.890 15.680 ;
        RECT 110.230 14.830 111.780 15.680 ;
        RECT 243.560 14.960 245.110 15.810 ;
        RECT 245.450 14.960 247.000 15.810 ;
        RECT 344.980 15.620 346.270 16.580 ;
        RECT 346.870 15.620 348.160 16.580 ;
        RECT 344.870 14.770 346.420 15.620 ;
        RECT 346.760 14.770 348.310 15.620 ;
      LAYER li1 ;
        RECT 8.150 246.800 8.450 247.750 ;
        RECT 10.040 246.800 10.340 247.750 ;
        RECT 8.050 246.200 11.240 246.800 ;
        RECT 109.460 246.610 109.760 247.560 ;
        RECT 111.350 246.610 111.650 247.560 ;
        RECT 244.680 246.740 244.980 247.690 ;
        RECT 246.570 246.740 246.870 247.690 ;
        RECT 109.360 246.010 112.550 246.610 ;
        RECT 244.580 246.140 247.770 246.740 ;
        RECT 345.990 246.550 346.290 247.500 ;
        RECT 347.880 246.550 348.180 247.500 ;
        RECT 345.890 245.950 349.080 246.550 ;
        RECT 23.830 244.380 24.130 245.330 ;
        RECT 25.720 244.380 26.020 245.330 ;
        RECT 23.730 243.780 26.920 244.380 ;
        RECT 125.140 244.190 125.440 245.140 ;
        RECT 127.030 244.190 127.330 245.140 ;
        RECT 260.360 244.320 260.660 245.270 ;
        RECT 262.250 244.320 262.550 245.270 ;
        RECT 125.040 243.590 128.230 244.190 ;
        RECT 260.260 243.720 263.450 244.320 ;
        RECT 361.670 244.130 361.970 245.080 ;
        RECT 363.560 244.130 363.860 245.080 ;
        RECT 361.570 243.530 364.760 244.130 ;
        RECT 8.310 240.400 8.610 241.350 ;
        RECT 10.200 240.400 10.500 241.350 ;
        RECT 8.210 239.800 11.400 240.400 ;
        RECT 109.620 240.210 109.920 241.160 ;
        RECT 111.510 240.210 111.810 241.160 ;
        RECT 244.840 240.340 245.140 241.290 ;
        RECT 246.730 240.340 247.030 241.290 ;
        RECT 41.410 238.830 41.710 239.780 ;
        RECT 43.300 238.830 43.600 239.780 ;
        RECT 109.520 239.610 112.710 240.210 ;
        RECT 244.740 239.740 247.930 240.340 ;
        RECT 346.150 240.150 346.450 241.100 ;
        RECT 348.040 240.150 348.340 241.100 ;
        RECT 41.310 238.230 44.500 238.830 ;
        RECT 142.720 238.640 143.020 239.590 ;
        RECT 144.610 238.640 144.910 239.590 ;
        RECT 277.940 238.770 278.240 239.720 ;
        RECT 279.830 238.770 280.130 239.720 ;
        RECT 346.050 239.550 349.240 240.150 ;
        RECT 142.620 238.040 145.810 238.640 ;
        RECT 277.840 238.170 281.030 238.770 ;
        RECT 379.250 238.580 379.550 239.530 ;
        RECT 381.140 238.580 381.440 239.530 ;
        RECT 379.150 237.980 382.340 238.580 ;
        RECT 7.980 232.380 8.280 233.330 ;
        RECT 9.870 232.380 10.170 233.330 ;
        RECT 7.880 231.780 11.070 232.380 ;
        RECT 109.290 232.190 109.590 233.140 ;
        RECT 111.180 232.190 111.480 233.140 ;
        RECT 244.510 232.320 244.810 233.270 ;
        RECT 246.400 232.320 246.700 233.270 ;
        RECT 109.190 231.590 112.380 232.190 ;
        RECT 244.410 231.720 247.600 232.320 ;
        RECT 345.820 232.130 346.120 233.080 ;
        RECT 347.710 232.130 348.010 233.080 ;
        RECT 345.720 231.530 348.910 232.130 ;
        RECT 23.660 229.960 23.960 230.910 ;
        RECT 25.550 229.960 25.850 230.910 ;
        RECT 23.560 229.360 26.750 229.960 ;
        RECT 124.970 229.770 125.270 230.720 ;
        RECT 126.860 229.770 127.160 230.720 ;
        RECT 260.190 229.900 260.490 230.850 ;
        RECT 262.080 229.900 262.380 230.850 ;
        RECT 124.870 229.170 128.060 229.770 ;
        RECT 260.090 229.300 263.280 229.900 ;
        RECT 361.500 229.710 361.800 230.660 ;
        RECT 363.390 229.710 363.690 230.660 ;
        RECT 361.400 229.110 364.590 229.710 ;
        RECT 8.140 225.980 8.440 226.930 ;
        RECT 10.030 225.980 10.330 226.930 ;
        RECT 8.040 225.380 11.230 225.980 ;
        RECT 109.450 225.790 109.750 226.740 ;
        RECT 111.340 225.790 111.640 226.740 ;
        RECT 244.670 225.920 244.970 226.870 ;
        RECT 246.560 225.920 246.860 226.870 ;
        RECT 109.350 225.190 112.540 225.790 ;
        RECT 244.570 225.320 247.760 225.920 ;
        RECT 345.980 225.730 346.280 226.680 ;
        RECT 347.870 225.730 348.170 226.680 ;
        RECT 345.880 225.130 349.070 225.730 ;
        RECT 58.940 222.810 59.240 223.760 ;
        RECT 60.830 222.810 61.130 223.760 ;
        RECT 58.840 222.210 62.030 222.810 ;
        RECT 160.250 222.620 160.550 223.570 ;
        RECT 162.140 222.620 162.440 223.570 ;
        RECT 295.470 222.750 295.770 223.700 ;
        RECT 297.360 222.750 297.660 223.700 ;
        RECT 160.150 222.020 163.340 222.620 ;
        RECT 295.370 222.150 298.560 222.750 ;
        RECT 396.780 222.560 397.080 223.510 ;
        RECT 398.670 222.560 398.970 223.510 ;
        RECT 396.680 221.960 399.870 222.560 ;
        RECT 8.120 216.730 8.420 217.680 ;
        RECT 10.010 216.730 10.310 217.680 ;
        RECT 8.020 216.130 11.210 216.730 ;
        RECT 109.430 216.540 109.730 217.490 ;
        RECT 111.320 216.540 111.620 217.490 ;
        RECT 244.650 216.670 244.950 217.620 ;
        RECT 246.540 216.670 246.840 217.620 ;
        RECT 109.330 215.940 112.520 216.540 ;
        RECT 244.550 216.070 247.740 216.670 ;
        RECT 345.960 216.480 346.260 217.430 ;
        RECT 347.850 216.480 348.150 217.430 ;
        RECT 345.860 215.880 349.050 216.480 ;
        RECT 23.800 214.310 24.100 215.260 ;
        RECT 25.690 214.310 25.990 215.260 ;
        RECT 23.700 213.710 26.890 214.310 ;
        RECT 125.110 214.120 125.410 215.070 ;
        RECT 127.000 214.120 127.300 215.070 ;
        RECT 260.330 214.250 260.630 215.200 ;
        RECT 262.220 214.250 262.520 215.200 ;
        RECT 125.010 213.520 128.200 214.120 ;
        RECT 260.230 213.650 263.420 214.250 ;
        RECT 361.640 214.060 361.940 215.010 ;
        RECT 363.530 214.060 363.830 215.010 ;
        RECT 361.540 213.460 364.730 214.060 ;
        RECT 8.280 210.330 8.580 211.280 ;
        RECT 10.170 210.330 10.470 211.280 ;
        RECT 8.180 209.730 11.370 210.330 ;
        RECT 109.590 210.140 109.890 211.090 ;
        RECT 111.480 210.140 111.780 211.090 ;
        RECT 244.810 210.270 245.110 211.220 ;
        RECT 246.700 210.270 247.000 211.220 ;
        RECT 41.380 208.760 41.680 209.710 ;
        RECT 43.270 208.760 43.570 209.710 ;
        RECT 109.490 209.540 112.680 210.140 ;
        RECT 244.710 209.670 247.900 210.270 ;
        RECT 346.120 210.080 346.420 211.030 ;
        RECT 348.010 210.080 348.310 211.030 ;
        RECT 41.280 208.160 44.470 208.760 ;
        RECT 142.690 208.570 142.990 209.520 ;
        RECT 144.580 208.570 144.880 209.520 ;
        RECT 277.910 208.700 278.210 209.650 ;
        RECT 279.800 208.700 280.100 209.650 ;
        RECT 346.020 209.480 349.210 210.080 ;
        RECT 142.590 207.970 145.780 208.570 ;
        RECT 277.810 208.100 281.000 208.700 ;
        RECT 379.220 208.510 379.520 209.460 ;
        RECT 381.110 208.510 381.410 209.460 ;
        RECT 379.120 207.910 382.310 208.510 ;
        RECT 7.950 202.310 8.250 203.260 ;
        RECT 9.840 202.310 10.140 203.260 ;
        RECT 7.850 201.710 11.040 202.310 ;
        RECT 109.260 202.120 109.560 203.070 ;
        RECT 111.150 202.120 111.450 203.070 ;
        RECT 244.480 202.250 244.780 203.200 ;
        RECT 246.370 202.250 246.670 203.200 ;
        RECT 109.160 201.520 112.350 202.120 ;
        RECT 244.380 201.650 247.570 202.250 ;
        RECT 345.790 202.060 346.090 203.010 ;
        RECT 347.680 202.060 347.980 203.010 ;
        RECT 345.690 201.460 348.880 202.060 ;
        RECT 23.630 199.890 23.930 200.840 ;
        RECT 25.520 199.890 25.820 200.840 ;
        RECT 23.530 199.290 26.720 199.890 ;
        RECT 124.940 199.700 125.240 200.650 ;
        RECT 126.830 199.700 127.130 200.650 ;
        RECT 260.160 199.830 260.460 200.780 ;
        RECT 262.050 199.830 262.350 200.780 ;
        RECT 124.840 199.100 128.030 199.700 ;
        RECT 260.060 199.230 263.250 199.830 ;
        RECT 361.470 199.640 361.770 200.590 ;
        RECT 363.360 199.640 363.660 200.590 ;
        RECT 361.370 199.040 364.560 199.640 ;
        RECT 8.110 195.910 8.410 196.860 ;
        RECT 10.000 195.910 10.300 196.860 ;
        RECT 73.140 196.520 73.440 197.470 ;
        RECT 75.030 196.520 75.330 197.470 ;
        RECT 73.040 195.920 76.230 196.520 ;
        RECT 8.010 195.310 11.200 195.910 ;
        RECT 109.420 195.720 109.720 196.670 ;
        RECT 111.310 195.720 111.610 196.670 ;
        RECT 174.450 196.330 174.750 197.280 ;
        RECT 176.340 196.330 176.640 197.280 ;
        RECT 174.350 195.730 177.540 196.330 ;
        RECT 244.640 195.850 244.940 196.800 ;
        RECT 246.530 195.850 246.830 196.800 ;
        RECT 309.670 196.460 309.970 197.410 ;
        RECT 311.560 196.460 311.860 197.410 ;
        RECT 309.570 195.860 312.760 196.460 ;
        RECT 109.320 195.120 112.510 195.720 ;
        RECT 244.540 195.250 247.730 195.850 ;
        RECT 345.950 195.660 346.250 196.610 ;
        RECT 347.840 195.660 348.140 196.610 ;
        RECT 410.980 196.270 411.280 197.220 ;
        RECT 412.870 196.270 413.170 197.220 ;
        RECT 410.880 195.670 414.070 196.270 ;
        RECT 345.850 195.060 349.040 195.660 ;
        RECT 7.800 186.880 8.100 187.830 ;
        RECT 9.690 186.880 9.990 187.830 ;
        RECT 7.700 186.280 10.890 186.880 ;
        RECT 109.110 186.690 109.410 187.640 ;
        RECT 111.000 186.690 111.300 187.640 ;
        RECT 244.330 186.820 244.630 187.770 ;
        RECT 246.220 186.820 246.520 187.770 ;
        RECT 109.010 186.090 112.200 186.690 ;
        RECT 244.230 186.220 247.420 186.820 ;
        RECT 345.640 186.630 345.940 187.580 ;
        RECT 347.530 186.630 347.830 187.580 ;
        RECT 345.540 186.030 348.730 186.630 ;
        RECT 23.480 184.460 23.780 185.410 ;
        RECT 25.370 184.460 25.670 185.410 ;
        RECT 23.380 183.860 26.570 184.460 ;
        RECT 124.790 184.270 125.090 185.220 ;
        RECT 126.680 184.270 126.980 185.220 ;
        RECT 260.010 184.400 260.310 185.350 ;
        RECT 261.900 184.400 262.200 185.350 ;
        RECT 124.690 183.670 127.880 184.270 ;
        RECT 259.910 183.800 263.100 184.400 ;
        RECT 361.320 184.210 361.620 185.160 ;
        RECT 363.210 184.210 363.510 185.160 ;
        RECT 361.220 183.610 364.410 184.210 ;
        RECT 7.960 180.480 8.260 181.430 ;
        RECT 9.850 180.480 10.150 181.430 ;
        RECT 7.860 179.880 11.050 180.480 ;
        RECT 109.270 180.290 109.570 181.240 ;
        RECT 111.160 180.290 111.460 181.240 ;
        RECT 244.490 180.420 244.790 181.370 ;
        RECT 246.380 180.420 246.680 181.370 ;
        RECT 41.060 178.910 41.360 179.860 ;
        RECT 42.950 178.910 43.250 179.860 ;
        RECT 109.170 179.690 112.360 180.290 ;
        RECT 244.390 179.820 247.580 180.420 ;
        RECT 345.800 180.230 346.100 181.180 ;
        RECT 347.690 180.230 347.990 181.180 ;
        RECT 40.960 178.310 44.150 178.910 ;
        RECT 142.370 178.720 142.670 179.670 ;
        RECT 144.260 178.720 144.560 179.670 ;
        RECT 277.590 178.850 277.890 179.800 ;
        RECT 279.480 178.850 279.780 179.800 ;
        RECT 345.700 179.630 348.890 180.230 ;
        RECT 142.270 178.120 145.460 178.720 ;
        RECT 277.490 178.250 280.680 178.850 ;
        RECT 378.900 178.660 379.200 179.610 ;
        RECT 380.790 178.660 381.090 179.610 ;
        RECT 378.800 178.060 381.990 178.660 ;
        RECT 7.630 172.460 7.930 173.410 ;
        RECT 9.520 172.460 9.820 173.410 ;
        RECT 7.530 171.860 10.720 172.460 ;
        RECT 108.940 172.270 109.240 173.220 ;
        RECT 110.830 172.270 111.130 173.220 ;
        RECT 244.160 172.400 244.460 173.350 ;
        RECT 246.050 172.400 246.350 173.350 ;
        RECT 108.840 171.670 112.030 172.270 ;
        RECT 244.060 171.800 247.250 172.400 ;
        RECT 345.470 172.210 345.770 173.160 ;
        RECT 347.360 172.210 347.660 173.160 ;
        RECT 345.370 171.610 348.560 172.210 ;
        RECT 23.310 170.040 23.610 170.990 ;
        RECT 25.200 170.040 25.500 170.990 ;
        RECT 23.210 169.440 26.400 170.040 ;
        RECT 124.620 169.850 124.920 170.800 ;
        RECT 126.510 169.850 126.810 170.800 ;
        RECT 259.840 169.980 260.140 170.930 ;
        RECT 261.730 169.980 262.030 170.930 ;
        RECT 124.520 169.250 127.710 169.850 ;
        RECT 259.740 169.380 262.930 169.980 ;
        RECT 361.150 169.790 361.450 170.740 ;
        RECT 363.040 169.790 363.340 170.740 ;
        RECT 361.050 169.190 364.240 169.790 ;
        RECT 7.790 166.060 8.090 167.010 ;
        RECT 9.680 166.060 9.980 167.010 ;
        RECT 7.690 165.460 10.880 166.060 ;
        RECT 109.100 165.870 109.400 166.820 ;
        RECT 110.990 165.870 111.290 166.820 ;
        RECT 244.320 166.000 244.620 166.950 ;
        RECT 246.210 166.000 246.510 166.950 ;
        RECT 109.000 165.270 112.190 165.870 ;
        RECT 244.220 165.400 247.410 166.000 ;
        RECT 345.630 165.810 345.930 166.760 ;
        RECT 347.520 165.810 347.820 166.760 ;
        RECT 345.530 165.210 348.720 165.810 ;
        RECT 58.590 162.890 58.890 163.840 ;
        RECT 60.480 162.890 60.780 163.840 ;
        RECT 58.490 162.290 61.680 162.890 ;
        RECT 159.900 162.700 160.200 163.650 ;
        RECT 161.790 162.700 162.090 163.650 ;
        RECT 295.120 162.830 295.420 163.780 ;
        RECT 297.010 162.830 297.310 163.780 ;
        RECT 159.800 162.100 162.990 162.700 ;
        RECT 295.020 162.230 298.210 162.830 ;
        RECT 396.430 162.640 396.730 163.590 ;
        RECT 398.320 162.640 398.620 163.590 ;
        RECT 396.330 162.040 399.520 162.640 ;
        RECT 7.770 156.810 8.070 157.760 ;
        RECT 9.660 156.810 9.960 157.760 ;
        RECT 7.670 156.210 10.860 156.810 ;
        RECT 109.080 156.620 109.380 157.570 ;
        RECT 110.970 156.620 111.270 157.570 ;
        RECT 244.300 156.750 244.600 157.700 ;
        RECT 246.190 156.750 246.490 157.700 ;
        RECT 108.980 156.020 112.170 156.620 ;
        RECT 244.200 156.150 247.390 156.750 ;
        RECT 345.610 156.560 345.910 157.510 ;
        RECT 347.500 156.560 347.800 157.510 ;
        RECT 345.510 155.960 348.700 156.560 ;
        RECT 23.450 154.390 23.750 155.340 ;
        RECT 25.340 154.390 25.640 155.340 ;
        RECT 23.350 153.790 26.540 154.390 ;
        RECT 124.760 154.200 125.060 155.150 ;
        RECT 126.650 154.200 126.950 155.150 ;
        RECT 259.980 154.330 260.280 155.280 ;
        RECT 261.870 154.330 262.170 155.280 ;
        RECT 124.660 153.600 127.850 154.200 ;
        RECT 259.880 153.730 263.070 154.330 ;
        RECT 361.290 154.140 361.590 155.090 ;
        RECT 363.180 154.140 363.480 155.090 ;
        RECT 361.190 153.540 364.380 154.140 ;
        RECT 7.930 150.410 8.230 151.360 ;
        RECT 9.820 150.410 10.120 151.360 ;
        RECT 7.830 149.810 11.020 150.410 ;
        RECT 109.240 150.220 109.540 151.170 ;
        RECT 111.130 150.220 111.430 151.170 ;
        RECT 244.460 150.350 244.760 151.300 ;
        RECT 246.350 150.350 246.650 151.300 ;
        RECT 41.030 148.840 41.330 149.790 ;
        RECT 42.920 148.840 43.220 149.790 ;
        RECT 109.140 149.620 112.330 150.220 ;
        RECT 244.360 149.750 247.550 150.350 ;
        RECT 345.770 150.160 346.070 151.110 ;
        RECT 347.660 150.160 347.960 151.110 ;
        RECT 40.930 148.240 44.120 148.840 ;
        RECT 142.340 148.650 142.640 149.600 ;
        RECT 144.230 148.650 144.530 149.600 ;
        RECT 277.560 148.780 277.860 149.730 ;
        RECT 279.450 148.780 279.750 149.730 ;
        RECT 345.670 149.560 348.860 150.160 ;
        RECT 142.240 148.050 145.430 148.650 ;
        RECT 277.460 148.180 280.650 148.780 ;
        RECT 378.870 148.590 379.170 149.540 ;
        RECT 380.760 148.590 381.060 149.540 ;
        RECT 378.770 147.990 381.960 148.590 ;
        RECT 7.600 142.390 7.900 143.340 ;
        RECT 9.490 142.390 9.790 143.340 ;
        RECT 7.500 141.790 10.690 142.390 ;
        RECT 108.910 142.200 109.210 143.150 ;
        RECT 110.800 142.200 111.100 143.150 ;
        RECT 244.130 142.330 244.430 143.280 ;
        RECT 246.020 142.330 246.320 143.280 ;
        RECT 108.810 141.600 112.000 142.200 ;
        RECT 244.030 141.730 247.220 142.330 ;
        RECT 345.440 142.140 345.740 143.090 ;
        RECT 347.330 142.140 347.630 143.090 ;
        RECT 345.340 141.540 348.530 142.140 ;
        RECT 23.280 139.970 23.580 140.920 ;
        RECT 25.170 139.970 25.470 140.920 ;
        RECT 23.180 139.370 26.370 139.970 ;
        RECT 124.590 139.780 124.890 140.730 ;
        RECT 126.480 139.780 126.780 140.730 ;
        RECT 259.810 139.910 260.110 140.860 ;
        RECT 261.700 139.910 262.000 140.860 ;
        RECT 124.490 139.180 127.680 139.780 ;
        RECT 259.710 139.310 262.900 139.910 ;
        RECT 361.120 139.720 361.420 140.670 ;
        RECT 363.010 139.720 363.310 140.670 ;
        RECT 361.020 139.120 364.210 139.720 ;
        RECT 7.760 135.990 8.060 136.940 ;
        RECT 9.650 135.990 9.950 136.940 ;
        RECT 7.660 135.390 10.850 135.990 ;
        RECT 109.070 135.800 109.370 136.750 ;
        RECT 110.960 135.800 111.260 136.750 ;
        RECT 108.970 135.200 112.160 135.800 ;
        RECT 217.060 135.520 217.360 136.470 ;
        RECT 218.950 135.520 219.250 136.470 ;
        RECT 244.290 135.930 244.590 136.880 ;
        RECT 246.180 135.930 246.480 136.880 ;
        RECT 216.960 134.920 220.150 135.520 ;
        RECT 244.190 135.330 247.380 135.930 ;
        RECT 345.600 135.740 345.900 136.690 ;
        RECT 347.490 135.740 347.790 136.690 ;
        RECT 345.500 135.140 348.690 135.740 ;
        RECT 453.590 135.460 453.890 136.410 ;
        RECT 455.480 135.460 455.780 136.410 ;
        RECT 453.490 134.860 456.680 135.460 ;
        RECT 89.470 133.380 89.770 134.330 ;
        RECT 91.360 133.380 91.660 134.330 ;
        RECT 89.370 132.780 92.560 133.380 ;
        RECT 190.780 133.190 191.080 134.140 ;
        RECT 192.670 133.190 192.970 134.140 ;
        RECT 326.000 133.320 326.300 134.270 ;
        RECT 327.890 133.320 328.190 134.270 ;
        RECT 190.680 132.590 193.870 133.190 ;
        RECT 325.900 132.720 329.090 133.320 ;
        RECT 427.310 133.130 427.610 134.080 ;
        RECT 429.200 133.130 429.500 134.080 ;
        RECT 427.210 132.530 430.400 133.130 ;
        RECT 470.890 133.110 471.190 134.060 ;
        RECT 472.780 133.110 473.080 134.060 ;
        RECT 470.790 132.510 473.980 133.110 ;
        RECT 7.650 126.560 7.950 127.510 ;
        RECT 9.540 126.560 9.840 127.510 ;
        RECT 7.550 125.960 10.740 126.560 ;
        RECT 108.960 126.370 109.260 127.320 ;
        RECT 110.850 126.370 111.150 127.320 ;
        RECT 244.180 126.500 244.480 127.450 ;
        RECT 246.070 126.500 246.370 127.450 ;
        RECT 108.860 125.770 112.050 126.370 ;
        RECT 244.080 125.900 247.270 126.500 ;
        RECT 345.490 126.310 345.790 127.260 ;
        RECT 347.380 126.310 347.680 127.260 ;
        RECT 345.390 125.710 348.580 126.310 ;
        RECT 23.330 124.140 23.630 125.090 ;
        RECT 25.220 124.140 25.520 125.090 ;
        RECT 23.230 123.540 26.420 124.140 ;
        RECT 124.640 123.950 124.940 124.900 ;
        RECT 126.530 123.950 126.830 124.900 ;
        RECT 259.860 124.080 260.160 125.030 ;
        RECT 261.750 124.080 262.050 125.030 ;
        RECT 124.540 123.350 127.730 123.950 ;
        RECT 259.760 123.480 262.950 124.080 ;
        RECT 361.170 123.890 361.470 124.840 ;
        RECT 363.060 123.890 363.360 124.840 ;
        RECT 361.070 123.290 364.260 123.890 ;
        RECT 7.810 120.160 8.110 121.110 ;
        RECT 9.700 120.160 10.000 121.110 ;
        RECT 7.710 119.560 10.900 120.160 ;
        RECT 109.120 119.970 109.420 120.920 ;
        RECT 111.010 119.970 111.310 120.920 ;
        RECT 244.340 120.100 244.640 121.050 ;
        RECT 246.230 120.100 246.530 121.050 ;
        RECT 40.910 118.590 41.210 119.540 ;
        RECT 42.800 118.590 43.100 119.540 ;
        RECT 109.020 119.370 112.210 119.970 ;
        RECT 244.240 119.500 247.430 120.100 ;
        RECT 345.650 119.910 345.950 120.860 ;
        RECT 347.540 119.910 347.840 120.860 ;
        RECT 40.810 117.990 44.000 118.590 ;
        RECT 142.220 118.400 142.520 119.350 ;
        RECT 144.110 118.400 144.410 119.350 ;
        RECT 277.440 118.530 277.740 119.480 ;
        RECT 279.330 118.530 279.630 119.480 ;
        RECT 345.550 119.310 348.740 119.910 ;
        RECT 142.120 117.800 145.310 118.400 ;
        RECT 277.340 117.930 280.530 118.530 ;
        RECT 378.750 118.340 379.050 119.290 ;
        RECT 380.640 118.340 380.940 119.290 ;
        RECT 378.650 117.740 381.840 118.340 ;
        RECT 7.480 112.140 7.780 113.090 ;
        RECT 9.370 112.140 9.670 113.090 ;
        RECT 7.380 111.540 10.570 112.140 ;
        RECT 108.790 111.950 109.090 112.900 ;
        RECT 110.680 111.950 110.980 112.900 ;
        RECT 244.010 112.080 244.310 113.030 ;
        RECT 245.900 112.080 246.200 113.030 ;
        RECT 108.690 111.350 111.880 111.950 ;
        RECT 243.910 111.480 247.100 112.080 ;
        RECT 345.320 111.890 345.620 112.840 ;
        RECT 347.210 111.890 347.510 112.840 ;
        RECT 345.220 111.290 348.410 111.890 ;
        RECT 23.160 109.720 23.460 110.670 ;
        RECT 25.050 109.720 25.350 110.670 ;
        RECT 23.060 109.120 26.250 109.720 ;
        RECT 124.470 109.530 124.770 110.480 ;
        RECT 126.360 109.530 126.660 110.480 ;
        RECT 259.690 109.660 259.990 110.610 ;
        RECT 261.580 109.660 261.880 110.610 ;
        RECT 124.370 108.930 127.560 109.530 ;
        RECT 259.590 109.060 262.780 109.660 ;
        RECT 361.000 109.470 361.300 110.420 ;
        RECT 362.890 109.470 363.190 110.420 ;
        RECT 360.900 108.870 364.090 109.470 ;
        RECT 7.640 105.740 7.940 106.690 ;
        RECT 9.530 105.740 9.830 106.690 ;
        RECT 7.540 105.140 10.730 105.740 ;
        RECT 108.950 105.550 109.250 106.500 ;
        RECT 110.840 105.550 111.140 106.500 ;
        RECT 244.170 105.680 244.470 106.630 ;
        RECT 246.060 105.680 246.360 106.630 ;
        RECT 108.850 104.950 112.040 105.550 ;
        RECT 244.070 105.080 247.260 105.680 ;
        RECT 345.480 105.490 345.780 106.440 ;
        RECT 347.370 105.490 347.670 106.440 ;
        RECT 345.380 104.890 348.570 105.490 ;
        RECT 58.440 102.570 58.740 103.520 ;
        RECT 60.330 102.570 60.630 103.520 ;
        RECT 58.340 101.970 61.530 102.570 ;
        RECT 159.750 102.380 160.050 103.330 ;
        RECT 161.640 102.380 161.940 103.330 ;
        RECT 294.970 102.510 295.270 103.460 ;
        RECT 296.860 102.510 297.160 103.460 ;
        RECT 159.650 101.780 162.840 102.380 ;
        RECT 294.870 101.910 298.060 102.510 ;
        RECT 396.280 102.320 396.580 103.270 ;
        RECT 398.170 102.320 398.470 103.270 ;
        RECT 396.180 101.720 399.370 102.320 ;
        RECT 7.620 96.490 7.920 97.440 ;
        RECT 9.510 96.490 9.810 97.440 ;
        RECT 7.520 95.890 10.710 96.490 ;
        RECT 108.930 96.300 109.230 97.250 ;
        RECT 110.820 96.300 111.120 97.250 ;
        RECT 244.150 96.430 244.450 97.380 ;
        RECT 246.040 96.430 246.340 97.380 ;
        RECT 108.830 95.700 112.020 96.300 ;
        RECT 244.050 95.830 247.240 96.430 ;
        RECT 345.460 96.240 345.760 97.190 ;
        RECT 347.350 96.240 347.650 97.190 ;
        RECT 345.360 95.640 348.550 96.240 ;
        RECT 23.300 94.070 23.600 95.020 ;
        RECT 25.190 94.070 25.490 95.020 ;
        RECT 23.200 93.470 26.390 94.070 ;
        RECT 124.610 93.880 124.910 94.830 ;
        RECT 126.500 93.880 126.800 94.830 ;
        RECT 259.830 94.010 260.130 94.960 ;
        RECT 261.720 94.010 262.020 94.960 ;
        RECT 124.510 93.280 127.700 93.880 ;
        RECT 259.730 93.410 262.920 94.010 ;
        RECT 361.140 93.820 361.440 94.770 ;
        RECT 363.030 93.820 363.330 94.770 ;
        RECT 361.040 93.220 364.230 93.820 ;
        RECT 7.780 90.090 8.080 91.040 ;
        RECT 9.670 90.090 9.970 91.040 ;
        RECT 7.680 89.490 10.870 90.090 ;
        RECT 109.090 89.900 109.390 90.850 ;
        RECT 110.980 89.900 111.280 90.850 ;
        RECT 244.310 90.030 244.610 90.980 ;
        RECT 246.200 90.030 246.500 90.980 ;
        RECT 40.880 88.520 41.180 89.470 ;
        RECT 42.770 88.520 43.070 89.470 ;
        RECT 108.990 89.300 112.180 89.900 ;
        RECT 244.210 89.430 247.400 90.030 ;
        RECT 345.620 89.840 345.920 90.790 ;
        RECT 347.510 89.840 347.810 90.790 ;
        RECT 40.780 87.920 43.970 88.520 ;
        RECT 142.190 88.330 142.490 89.280 ;
        RECT 144.080 88.330 144.380 89.280 ;
        RECT 277.410 88.460 277.710 89.410 ;
        RECT 279.300 88.460 279.600 89.410 ;
        RECT 345.520 89.240 348.710 89.840 ;
        RECT 142.090 87.730 145.280 88.330 ;
        RECT 277.310 87.860 280.500 88.460 ;
        RECT 378.720 88.270 379.020 89.220 ;
        RECT 380.610 88.270 380.910 89.220 ;
        RECT 378.620 87.670 381.810 88.270 ;
        RECT 7.450 82.070 7.750 83.020 ;
        RECT 9.340 82.070 9.640 83.020 ;
        RECT 7.350 81.470 10.540 82.070 ;
        RECT 108.760 81.880 109.060 82.830 ;
        RECT 110.650 81.880 110.950 82.830 ;
        RECT 243.980 82.010 244.280 82.960 ;
        RECT 245.870 82.010 246.170 82.960 ;
        RECT 108.660 81.280 111.850 81.880 ;
        RECT 243.880 81.410 247.070 82.010 ;
        RECT 345.290 81.820 345.590 82.770 ;
        RECT 347.180 81.820 347.480 82.770 ;
        RECT 345.190 81.220 348.380 81.820 ;
        RECT 23.130 79.650 23.430 80.600 ;
        RECT 25.020 79.650 25.320 80.600 ;
        RECT 23.030 79.050 26.220 79.650 ;
        RECT 124.440 79.460 124.740 80.410 ;
        RECT 126.330 79.460 126.630 80.410 ;
        RECT 259.660 79.590 259.960 80.540 ;
        RECT 261.550 79.590 261.850 80.540 ;
        RECT 124.340 78.860 127.530 79.460 ;
        RECT 259.560 78.990 262.750 79.590 ;
        RECT 360.970 79.400 361.270 80.350 ;
        RECT 362.860 79.400 363.160 80.350 ;
        RECT 360.870 78.800 364.060 79.400 ;
        RECT 7.610 75.670 7.910 76.620 ;
        RECT 9.500 75.670 9.800 76.620 ;
        RECT 72.640 76.280 72.940 77.230 ;
        RECT 74.530 76.280 74.830 77.230 ;
        RECT 72.540 75.680 75.730 76.280 ;
        RECT 7.510 75.070 10.700 75.670 ;
        RECT 108.920 75.480 109.220 76.430 ;
        RECT 110.810 75.480 111.110 76.430 ;
        RECT 173.950 76.090 174.250 77.040 ;
        RECT 175.840 76.090 176.140 77.040 ;
        RECT 173.850 75.490 177.040 76.090 ;
        RECT 244.140 75.610 244.440 76.560 ;
        RECT 246.030 75.610 246.330 76.560 ;
        RECT 309.170 76.220 309.470 77.170 ;
        RECT 311.060 76.220 311.360 77.170 ;
        RECT 309.070 75.620 312.260 76.220 ;
        RECT 108.820 74.880 112.010 75.480 ;
        RECT 244.040 75.010 247.230 75.610 ;
        RECT 345.450 75.420 345.750 76.370 ;
        RECT 347.340 75.420 347.640 76.370 ;
        RECT 410.480 76.030 410.780 76.980 ;
        RECT 412.370 76.030 412.670 76.980 ;
        RECT 410.380 75.430 413.570 76.030 ;
        RECT 345.350 74.820 348.540 75.420 ;
        RECT 7.300 66.640 7.600 67.590 ;
        RECT 9.190 66.640 9.490 67.590 ;
        RECT 7.200 66.040 10.390 66.640 ;
        RECT 108.610 66.450 108.910 67.400 ;
        RECT 110.500 66.450 110.800 67.400 ;
        RECT 243.830 66.580 244.130 67.530 ;
        RECT 245.720 66.580 246.020 67.530 ;
        RECT 108.510 65.850 111.700 66.450 ;
        RECT 243.730 65.980 246.920 66.580 ;
        RECT 345.140 66.390 345.440 67.340 ;
        RECT 347.030 66.390 347.330 67.340 ;
        RECT 345.040 65.790 348.230 66.390 ;
        RECT 22.980 64.220 23.280 65.170 ;
        RECT 24.870 64.220 25.170 65.170 ;
        RECT 22.880 63.620 26.070 64.220 ;
        RECT 124.290 64.030 124.590 64.980 ;
        RECT 126.180 64.030 126.480 64.980 ;
        RECT 259.510 64.160 259.810 65.110 ;
        RECT 261.400 64.160 261.700 65.110 ;
        RECT 124.190 63.430 127.380 64.030 ;
        RECT 259.410 63.560 262.600 64.160 ;
        RECT 360.820 63.970 361.120 64.920 ;
        RECT 362.710 63.970 363.010 64.920 ;
        RECT 360.720 63.370 363.910 63.970 ;
        RECT 7.460 60.240 7.760 61.190 ;
        RECT 9.350 60.240 9.650 61.190 ;
        RECT 7.360 59.640 10.550 60.240 ;
        RECT 108.770 60.050 109.070 61.000 ;
        RECT 110.660 60.050 110.960 61.000 ;
        RECT 243.990 60.180 244.290 61.130 ;
        RECT 245.880 60.180 246.180 61.130 ;
        RECT 40.560 58.670 40.860 59.620 ;
        RECT 42.450 58.670 42.750 59.620 ;
        RECT 108.670 59.450 111.860 60.050 ;
        RECT 243.890 59.580 247.080 60.180 ;
        RECT 345.300 59.990 345.600 60.940 ;
        RECT 347.190 59.990 347.490 60.940 ;
        RECT 40.460 58.070 43.650 58.670 ;
        RECT 141.870 58.480 142.170 59.430 ;
        RECT 143.760 58.480 144.060 59.430 ;
        RECT 277.090 58.610 277.390 59.560 ;
        RECT 278.980 58.610 279.280 59.560 ;
        RECT 345.200 59.390 348.390 59.990 ;
        RECT 141.770 57.880 144.960 58.480 ;
        RECT 276.990 58.010 280.180 58.610 ;
        RECT 378.400 58.420 378.700 59.370 ;
        RECT 380.290 58.420 380.590 59.370 ;
        RECT 378.300 57.820 381.490 58.420 ;
        RECT 7.130 52.220 7.430 53.170 ;
        RECT 9.020 52.220 9.320 53.170 ;
        RECT 7.030 51.620 10.220 52.220 ;
        RECT 108.440 52.030 108.740 52.980 ;
        RECT 110.330 52.030 110.630 52.980 ;
        RECT 243.660 52.160 243.960 53.110 ;
        RECT 245.550 52.160 245.850 53.110 ;
        RECT 108.340 51.430 111.530 52.030 ;
        RECT 243.560 51.560 246.750 52.160 ;
        RECT 344.970 51.970 345.270 52.920 ;
        RECT 346.860 51.970 347.160 52.920 ;
        RECT 344.870 51.370 348.060 51.970 ;
        RECT 22.810 49.800 23.110 50.750 ;
        RECT 24.700 49.800 25.000 50.750 ;
        RECT 22.710 49.200 25.900 49.800 ;
        RECT 124.120 49.610 124.420 50.560 ;
        RECT 126.010 49.610 126.310 50.560 ;
        RECT 259.340 49.740 259.640 50.690 ;
        RECT 261.230 49.740 261.530 50.690 ;
        RECT 124.020 49.010 127.210 49.610 ;
        RECT 259.240 49.140 262.430 49.740 ;
        RECT 360.650 49.550 360.950 50.500 ;
        RECT 362.540 49.550 362.840 50.500 ;
        RECT 360.550 48.950 363.740 49.550 ;
        RECT 7.290 45.820 7.590 46.770 ;
        RECT 9.180 45.820 9.480 46.770 ;
        RECT 7.190 45.220 10.380 45.820 ;
        RECT 108.600 45.630 108.900 46.580 ;
        RECT 110.490 45.630 110.790 46.580 ;
        RECT 243.820 45.760 244.120 46.710 ;
        RECT 245.710 45.760 246.010 46.710 ;
        RECT 108.500 45.030 111.690 45.630 ;
        RECT 243.720 45.160 246.910 45.760 ;
        RECT 345.130 45.570 345.430 46.520 ;
        RECT 347.020 45.570 347.320 46.520 ;
        RECT 345.030 44.970 348.220 45.570 ;
        RECT 58.090 42.650 58.390 43.600 ;
        RECT 59.980 42.650 60.280 43.600 ;
        RECT 57.990 42.050 61.180 42.650 ;
        RECT 159.400 42.460 159.700 43.410 ;
        RECT 161.290 42.460 161.590 43.410 ;
        RECT 294.620 42.590 294.920 43.540 ;
        RECT 296.510 42.590 296.810 43.540 ;
        RECT 159.300 41.860 162.490 42.460 ;
        RECT 294.520 41.990 297.710 42.590 ;
        RECT 395.930 42.400 396.230 43.350 ;
        RECT 397.820 42.400 398.120 43.350 ;
        RECT 395.830 41.800 399.020 42.400 ;
        RECT 7.270 36.570 7.570 37.520 ;
        RECT 9.160 36.570 9.460 37.520 ;
        RECT 7.170 35.970 10.360 36.570 ;
        RECT 108.580 36.380 108.880 37.330 ;
        RECT 110.470 36.380 110.770 37.330 ;
        RECT 243.800 36.510 244.100 37.460 ;
        RECT 245.690 36.510 245.990 37.460 ;
        RECT 108.480 35.780 111.670 36.380 ;
        RECT 243.700 35.910 246.890 36.510 ;
        RECT 345.110 36.320 345.410 37.270 ;
        RECT 347.000 36.320 347.300 37.270 ;
        RECT 345.010 35.720 348.200 36.320 ;
        RECT 22.950 34.150 23.250 35.100 ;
        RECT 24.840 34.150 25.140 35.100 ;
        RECT 22.850 33.550 26.040 34.150 ;
        RECT 124.260 33.960 124.560 34.910 ;
        RECT 126.150 33.960 126.450 34.910 ;
        RECT 259.480 34.090 259.780 35.040 ;
        RECT 261.370 34.090 261.670 35.040 ;
        RECT 124.160 33.360 127.350 33.960 ;
        RECT 259.380 33.490 262.570 34.090 ;
        RECT 360.790 33.900 361.090 34.850 ;
        RECT 362.680 33.900 362.980 34.850 ;
        RECT 360.690 33.300 363.880 33.900 ;
        RECT 7.430 30.170 7.730 31.120 ;
        RECT 9.320 30.170 9.620 31.120 ;
        RECT 7.330 29.570 10.520 30.170 ;
        RECT 108.740 29.980 109.040 30.930 ;
        RECT 110.630 29.980 110.930 30.930 ;
        RECT 243.960 30.110 244.260 31.060 ;
        RECT 245.850 30.110 246.150 31.060 ;
        RECT 40.530 28.600 40.830 29.550 ;
        RECT 42.420 28.600 42.720 29.550 ;
        RECT 108.640 29.380 111.830 29.980 ;
        RECT 243.860 29.510 247.050 30.110 ;
        RECT 345.270 29.920 345.570 30.870 ;
        RECT 347.160 29.920 347.460 30.870 ;
        RECT 40.430 28.000 43.620 28.600 ;
        RECT 141.840 28.410 142.140 29.360 ;
        RECT 143.730 28.410 144.030 29.360 ;
        RECT 277.060 28.540 277.360 29.490 ;
        RECT 278.950 28.540 279.250 29.490 ;
        RECT 345.170 29.320 348.360 29.920 ;
        RECT 141.740 27.810 144.930 28.410 ;
        RECT 276.960 27.940 280.150 28.540 ;
        RECT 378.370 28.350 378.670 29.300 ;
        RECT 380.260 28.350 380.560 29.300 ;
        RECT 378.270 27.750 381.460 28.350 ;
        RECT 7.100 22.150 7.400 23.100 ;
        RECT 8.990 22.150 9.290 23.100 ;
        RECT 7.000 21.550 10.190 22.150 ;
        RECT 108.410 21.960 108.710 22.910 ;
        RECT 110.300 21.960 110.600 22.910 ;
        RECT 243.630 22.090 243.930 23.040 ;
        RECT 245.520 22.090 245.820 23.040 ;
        RECT 108.310 21.360 111.500 21.960 ;
        RECT 243.530 21.490 246.720 22.090 ;
        RECT 344.940 21.900 345.240 22.850 ;
        RECT 346.830 21.900 347.130 22.850 ;
        RECT 344.840 21.300 348.030 21.900 ;
        RECT 22.780 19.730 23.080 20.680 ;
        RECT 24.670 19.730 24.970 20.680 ;
        RECT 22.680 19.130 25.870 19.730 ;
        RECT 124.090 19.540 124.390 20.490 ;
        RECT 125.980 19.540 126.280 20.490 ;
        RECT 259.310 19.670 259.610 20.620 ;
        RECT 261.200 19.670 261.500 20.620 ;
        RECT 123.990 18.940 127.180 19.540 ;
        RECT 259.210 19.070 262.400 19.670 ;
        RECT 360.620 19.480 360.920 20.430 ;
        RECT 362.510 19.480 362.810 20.430 ;
        RECT 360.520 18.880 363.710 19.480 ;
        RECT 7.260 15.750 7.560 16.700 ;
        RECT 9.150 15.750 9.450 16.700 ;
        RECT 7.160 15.150 10.350 15.750 ;
        RECT 108.570 15.560 108.870 16.510 ;
        RECT 110.460 15.560 110.760 16.510 ;
        RECT 243.790 15.690 244.090 16.640 ;
        RECT 245.680 15.690 245.980 16.640 ;
        RECT 108.470 14.960 111.660 15.560 ;
        RECT 243.690 15.090 246.880 15.690 ;
        RECT 345.100 15.500 345.400 16.450 ;
        RECT 346.990 15.500 347.290 16.450 ;
        RECT 345.000 14.900 348.190 15.500 ;
      LAYER mcon ;
        RECT 8.210 246.500 8.380 246.670 ;
        RECT 9.070 246.490 9.240 246.660 ;
        RECT 10.100 246.500 10.270 246.670 ;
        RECT 10.960 246.490 11.130 246.660 ;
        RECT 109.520 246.310 109.690 246.480 ;
        RECT 110.380 246.300 110.550 246.470 ;
        RECT 111.410 246.310 111.580 246.480 ;
        RECT 112.270 246.300 112.440 246.470 ;
        RECT 244.740 246.440 244.910 246.610 ;
        RECT 245.600 246.430 245.770 246.600 ;
        RECT 246.630 246.440 246.800 246.610 ;
        RECT 247.490 246.430 247.660 246.600 ;
        RECT 346.050 246.250 346.220 246.420 ;
        RECT 346.910 246.240 347.080 246.410 ;
        RECT 347.940 246.250 348.110 246.420 ;
        RECT 348.800 246.240 348.970 246.410 ;
        RECT 23.890 244.080 24.060 244.250 ;
        RECT 24.750 244.070 24.920 244.240 ;
        RECT 25.780 244.080 25.950 244.250 ;
        RECT 26.640 244.070 26.810 244.240 ;
        RECT 125.200 243.890 125.370 244.060 ;
        RECT 126.060 243.880 126.230 244.050 ;
        RECT 127.090 243.890 127.260 244.060 ;
        RECT 127.950 243.880 128.120 244.050 ;
        RECT 260.420 244.020 260.590 244.190 ;
        RECT 261.280 244.010 261.450 244.180 ;
        RECT 262.310 244.020 262.480 244.190 ;
        RECT 263.170 244.010 263.340 244.180 ;
        RECT 361.730 243.830 361.900 244.000 ;
        RECT 362.590 243.820 362.760 243.990 ;
        RECT 363.620 243.830 363.790 244.000 ;
        RECT 364.480 243.820 364.650 243.990 ;
        RECT 8.370 240.100 8.540 240.270 ;
        RECT 9.230 240.090 9.400 240.260 ;
        RECT 10.260 240.100 10.430 240.270 ;
        RECT 11.120 240.090 11.290 240.260 ;
        RECT 109.680 239.910 109.850 240.080 ;
        RECT 110.540 239.900 110.710 240.070 ;
        RECT 111.570 239.910 111.740 240.080 ;
        RECT 112.430 239.900 112.600 240.070 ;
        RECT 244.900 240.040 245.070 240.210 ;
        RECT 245.760 240.030 245.930 240.200 ;
        RECT 246.790 240.040 246.960 240.210 ;
        RECT 247.650 240.030 247.820 240.200 ;
        RECT 346.210 239.850 346.380 240.020 ;
        RECT 347.070 239.840 347.240 240.010 ;
        RECT 348.100 239.850 348.270 240.020 ;
        RECT 348.960 239.840 349.130 240.010 ;
        RECT 41.470 238.530 41.640 238.700 ;
        RECT 42.330 238.520 42.500 238.690 ;
        RECT 43.360 238.530 43.530 238.700 ;
        RECT 44.220 238.520 44.390 238.690 ;
        RECT 142.780 238.340 142.950 238.510 ;
        RECT 143.640 238.330 143.810 238.500 ;
        RECT 144.670 238.340 144.840 238.510 ;
        RECT 145.530 238.330 145.700 238.500 ;
        RECT 278.000 238.470 278.170 238.640 ;
        RECT 278.860 238.460 279.030 238.630 ;
        RECT 279.890 238.470 280.060 238.640 ;
        RECT 280.750 238.460 280.920 238.630 ;
        RECT 379.310 238.280 379.480 238.450 ;
        RECT 380.170 238.270 380.340 238.440 ;
        RECT 381.200 238.280 381.370 238.450 ;
        RECT 382.060 238.270 382.230 238.440 ;
        RECT 8.040 232.080 8.210 232.250 ;
        RECT 8.900 232.070 9.070 232.240 ;
        RECT 9.930 232.080 10.100 232.250 ;
        RECT 10.790 232.070 10.960 232.240 ;
        RECT 109.350 231.890 109.520 232.060 ;
        RECT 110.210 231.880 110.380 232.050 ;
        RECT 111.240 231.890 111.410 232.060 ;
        RECT 112.100 231.880 112.270 232.050 ;
        RECT 244.570 232.020 244.740 232.190 ;
        RECT 245.430 232.010 245.600 232.180 ;
        RECT 246.460 232.020 246.630 232.190 ;
        RECT 247.320 232.010 247.490 232.180 ;
        RECT 345.880 231.830 346.050 232.000 ;
        RECT 346.740 231.820 346.910 231.990 ;
        RECT 347.770 231.830 347.940 232.000 ;
        RECT 348.630 231.820 348.800 231.990 ;
        RECT 23.720 229.660 23.890 229.830 ;
        RECT 24.580 229.650 24.750 229.820 ;
        RECT 25.610 229.660 25.780 229.830 ;
        RECT 26.470 229.650 26.640 229.820 ;
        RECT 125.030 229.470 125.200 229.640 ;
        RECT 125.890 229.460 126.060 229.630 ;
        RECT 126.920 229.470 127.090 229.640 ;
        RECT 127.780 229.460 127.950 229.630 ;
        RECT 260.250 229.600 260.420 229.770 ;
        RECT 261.110 229.590 261.280 229.760 ;
        RECT 262.140 229.600 262.310 229.770 ;
        RECT 263.000 229.590 263.170 229.760 ;
        RECT 361.560 229.410 361.730 229.580 ;
        RECT 362.420 229.400 362.590 229.570 ;
        RECT 363.450 229.410 363.620 229.580 ;
        RECT 364.310 229.400 364.480 229.570 ;
        RECT 8.200 225.680 8.370 225.850 ;
        RECT 9.060 225.670 9.230 225.840 ;
        RECT 10.090 225.680 10.260 225.850 ;
        RECT 10.950 225.670 11.120 225.840 ;
        RECT 109.510 225.490 109.680 225.660 ;
        RECT 110.370 225.480 110.540 225.650 ;
        RECT 111.400 225.490 111.570 225.660 ;
        RECT 112.260 225.480 112.430 225.650 ;
        RECT 244.730 225.620 244.900 225.790 ;
        RECT 245.590 225.610 245.760 225.780 ;
        RECT 246.620 225.620 246.790 225.790 ;
        RECT 247.480 225.610 247.650 225.780 ;
        RECT 346.040 225.430 346.210 225.600 ;
        RECT 346.900 225.420 347.070 225.590 ;
        RECT 347.930 225.430 348.100 225.600 ;
        RECT 348.790 225.420 348.960 225.590 ;
        RECT 59.000 222.510 59.170 222.680 ;
        RECT 59.860 222.500 60.030 222.670 ;
        RECT 60.890 222.510 61.060 222.680 ;
        RECT 61.750 222.500 61.920 222.670 ;
        RECT 160.310 222.320 160.480 222.490 ;
        RECT 161.170 222.310 161.340 222.480 ;
        RECT 162.200 222.320 162.370 222.490 ;
        RECT 163.060 222.310 163.230 222.480 ;
        RECT 295.530 222.450 295.700 222.620 ;
        RECT 296.390 222.440 296.560 222.610 ;
        RECT 297.420 222.450 297.590 222.620 ;
        RECT 298.280 222.440 298.450 222.610 ;
        RECT 396.840 222.260 397.010 222.430 ;
        RECT 397.700 222.250 397.870 222.420 ;
        RECT 398.730 222.260 398.900 222.430 ;
        RECT 399.590 222.250 399.760 222.420 ;
        RECT 8.180 216.430 8.350 216.600 ;
        RECT 9.040 216.420 9.210 216.590 ;
        RECT 10.070 216.430 10.240 216.600 ;
        RECT 10.930 216.420 11.100 216.590 ;
        RECT 109.490 216.240 109.660 216.410 ;
        RECT 110.350 216.230 110.520 216.400 ;
        RECT 111.380 216.240 111.550 216.410 ;
        RECT 112.240 216.230 112.410 216.400 ;
        RECT 244.710 216.370 244.880 216.540 ;
        RECT 245.570 216.360 245.740 216.530 ;
        RECT 246.600 216.370 246.770 216.540 ;
        RECT 247.460 216.360 247.630 216.530 ;
        RECT 346.020 216.180 346.190 216.350 ;
        RECT 346.880 216.170 347.050 216.340 ;
        RECT 347.910 216.180 348.080 216.350 ;
        RECT 348.770 216.170 348.940 216.340 ;
        RECT 23.860 214.010 24.030 214.180 ;
        RECT 24.720 214.000 24.890 214.170 ;
        RECT 25.750 214.010 25.920 214.180 ;
        RECT 26.610 214.000 26.780 214.170 ;
        RECT 125.170 213.820 125.340 213.990 ;
        RECT 126.030 213.810 126.200 213.980 ;
        RECT 127.060 213.820 127.230 213.990 ;
        RECT 127.920 213.810 128.090 213.980 ;
        RECT 260.390 213.950 260.560 214.120 ;
        RECT 261.250 213.940 261.420 214.110 ;
        RECT 262.280 213.950 262.450 214.120 ;
        RECT 263.140 213.940 263.310 214.110 ;
        RECT 361.700 213.760 361.870 213.930 ;
        RECT 362.560 213.750 362.730 213.920 ;
        RECT 363.590 213.760 363.760 213.930 ;
        RECT 364.450 213.750 364.620 213.920 ;
        RECT 8.340 210.030 8.510 210.200 ;
        RECT 9.200 210.020 9.370 210.190 ;
        RECT 10.230 210.030 10.400 210.200 ;
        RECT 11.090 210.020 11.260 210.190 ;
        RECT 109.650 209.840 109.820 210.010 ;
        RECT 110.510 209.830 110.680 210.000 ;
        RECT 111.540 209.840 111.710 210.010 ;
        RECT 112.400 209.830 112.570 210.000 ;
        RECT 244.870 209.970 245.040 210.140 ;
        RECT 245.730 209.960 245.900 210.130 ;
        RECT 246.760 209.970 246.930 210.140 ;
        RECT 247.620 209.960 247.790 210.130 ;
        RECT 346.180 209.780 346.350 209.950 ;
        RECT 347.040 209.770 347.210 209.940 ;
        RECT 348.070 209.780 348.240 209.950 ;
        RECT 348.930 209.770 349.100 209.940 ;
        RECT 41.440 208.460 41.610 208.630 ;
        RECT 42.300 208.450 42.470 208.620 ;
        RECT 43.330 208.460 43.500 208.630 ;
        RECT 44.190 208.450 44.360 208.620 ;
        RECT 142.750 208.270 142.920 208.440 ;
        RECT 143.610 208.260 143.780 208.430 ;
        RECT 144.640 208.270 144.810 208.440 ;
        RECT 145.500 208.260 145.670 208.430 ;
        RECT 277.970 208.400 278.140 208.570 ;
        RECT 278.830 208.390 279.000 208.560 ;
        RECT 279.860 208.400 280.030 208.570 ;
        RECT 280.720 208.390 280.890 208.560 ;
        RECT 379.280 208.210 379.450 208.380 ;
        RECT 380.140 208.200 380.310 208.370 ;
        RECT 381.170 208.210 381.340 208.380 ;
        RECT 382.030 208.200 382.200 208.370 ;
        RECT 8.010 202.010 8.180 202.180 ;
        RECT 8.870 202.000 9.040 202.170 ;
        RECT 9.900 202.010 10.070 202.180 ;
        RECT 10.760 202.000 10.930 202.170 ;
        RECT 109.320 201.820 109.490 201.990 ;
        RECT 110.180 201.810 110.350 201.980 ;
        RECT 111.210 201.820 111.380 201.990 ;
        RECT 112.070 201.810 112.240 201.980 ;
        RECT 244.540 201.950 244.710 202.120 ;
        RECT 245.400 201.940 245.570 202.110 ;
        RECT 246.430 201.950 246.600 202.120 ;
        RECT 247.290 201.940 247.460 202.110 ;
        RECT 345.850 201.760 346.020 201.930 ;
        RECT 346.710 201.750 346.880 201.920 ;
        RECT 347.740 201.760 347.910 201.930 ;
        RECT 348.600 201.750 348.770 201.920 ;
        RECT 23.690 199.590 23.860 199.760 ;
        RECT 24.550 199.580 24.720 199.750 ;
        RECT 25.580 199.590 25.750 199.760 ;
        RECT 26.440 199.580 26.610 199.750 ;
        RECT 125.000 199.400 125.170 199.570 ;
        RECT 125.860 199.390 126.030 199.560 ;
        RECT 126.890 199.400 127.060 199.570 ;
        RECT 127.750 199.390 127.920 199.560 ;
        RECT 260.220 199.530 260.390 199.700 ;
        RECT 261.080 199.520 261.250 199.690 ;
        RECT 262.110 199.530 262.280 199.700 ;
        RECT 262.970 199.520 263.140 199.690 ;
        RECT 361.530 199.340 361.700 199.510 ;
        RECT 362.390 199.330 362.560 199.500 ;
        RECT 363.420 199.340 363.590 199.510 ;
        RECT 364.280 199.330 364.450 199.500 ;
        RECT 73.200 196.220 73.370 196.390 ;
        RECT 74.060 196.210 74.230 196.380 ;
        RECT 75.090 196.220 75.260 196.390 ;
        RECT 75.950 196.210 76.120 196.380 ;
        RECT 8.170 195.610 8.340 195.780 ;
        RECT 9.030 195.600 9.200 195.770 ;
        RECT 10.060 195.610 10.230 195.780 ;
        RECT 10.920 195.600 11.090 195.770 ;
        RECT 174.510 196.030 174.680 196.200 ;
        RECT 175.370 196.020 175.540 196.190 ;
        RECT 176.400 196.030 176.570 196.200 ;
        RECT 177.260 196.020 177.430 196.190 ;
        RECT 309.730 196.160 309.900 196.330 ;
        RECT 310.590 196.150 310.760 196.320 ;
        RECT 311.620 196.160 311.790 196.330 ;
        RECT 312.480 196.150 312.650 196.320 ;
        RECT 109.480 195.420 109.650 195.590 ;
        RECT 110.340 195.410 110.510 195.580 ;
        RECT 111.370 195.420 111.540 195.590 ;
        RECT 112.230 195.410 112.400 195.580 ;
        RECT 244.700 195.550 244.870 195.720 ;
        RECT 245.560 195.540 245.730 195.710 ;
        RECT 246.590 195.550 246.760 195.720 ;
        RECT 247.450 195.540 247.620 195.710 ;
        RECT 411.040 195.970 411.210 196.140 ;
        RECT 411.900 195.960 412.070 196.130 ;
        RECT 412.930 195.970 413.100 196.140 ;
        RECT 413.790 195.960 413.960 196.130 ;
        RECT 346.010 195.360 346.180 195.530 ;
        RECT 346.870 195.350 347.040 195.520 ;
        RECT 347.900 195.360 348.070 195.530 ;
        RECT 348.760 195.350 348.930 195.520 ;
        RECT 7.860 186.580 8.030 186.750 ;
        RECT 8.720 186.570 8.890 186.740 ;
        RECT 9.750 186.580 9.920 186.750 ;
        RECT 10.610 186.570 10.780 186.740 ;
        RECT 109.170 186.390 109.340 186.560 ;
        RECT 110.030 186.380 110.200 186.550 ;
        RECT 111.060 186.390 111.230 186.560 ;
        RECT 111.920 186.380 112.090 186.550 ;
        RECT 244.390 186.520 244.560 186.690 ;
        RECT 245.250 186.510 245.420 186.680 ;
        RECT 246.280 186.520 246.450 186.690 ;
        RECT 247.140 186.510 247.310 186.680 ;
        RECT 345.700 186.330 345.870 186.500 ;
        RECT 346.560 186.320 346.730 186.490 ;
        RECT 347.590 186.330 347.760 186.500 ;
        RECT 348.450 186.320 348.620 186.490 ;
        RECT 23.540 184.160 23.710 184.330 ;
        RECT 24.400 184.150 24.570 184.320 ;
        RECT 25.430 184.160 25.600 184.330 ;
        RECT 26.290 184.150 26.460 184.320 ;
        RECT 124.850 183.970 125.020 184.140 ;
        RECT 125.710 183.960 125.880 184.130 ;
        RECT 126.740 183.970 126.910 184.140 ;
        RECT 127.600 183.960 127.770 184.130 ;
        RECT 260.070 184.100 260.240 184.270 ;
        RECT 260.930 184.090 261.100 184.260 ;
        RECT 261.960 184.100 262.130 184.270 ;
        RECT 262.820 184.090 262.990 184.260 ;
        RECT 361.380 183.910 361.550 184.080 ;
        RECT 362.240 183.900 362.410 184.070 ;
        RECT 363.270 183.910 363.440 184.080 ;
        RECT 364.130 183.900 364.300 184.070 ;
        RECT 8.020 180.180 8.190 180.350 ;
        RECT 8.880 180.170 9.050 180.340 ;
        RECT 9.910 180.180 10.080 180.350 ;
        RECT 10.770 180.170 10.940 180.340 ;
        RECT 109.330 179.990 109.500 180.160 ;
        RECT 110.190 179.980 110.360 180.150 ;
        RECT 111.220 179.990 111.390 180.160 ;
        RECT 112.080 179.980 112.250 180.150 ;
        RECT 244.550 180.120 244.720 180.290 ;
        RECT 245.410 180.110 245.580 180.280 ;
        RECT 246.440 180.120 246.610 180.290 ;
        RECT 247.300 180.110 247.470 180.280 ;
        RECT 345.860 179.930 346.030 180.100 ;
        RECT 346.720 179.920 346.890 180.090 ;
        RECT 347.750 179.930 347.920 180.100 ;
        RECT 348.610 179.920 348.780 180.090 ;
        RECT 41.120 178.610 41.290 178.780 ;
        RECT 41.980 178.600 42.150 178.770 ;
        RECT 43.010 178.610 43.180 178.780 ;
        RECT 43.870 178.600 44.040 178.770 ;
        RECT 142.430 178.420 142.600 178.590 ;
        RECT 143.290 178.410 143.460 178.580 ;
        RECT 144.320 178.420 144.490 178.590 ;
        RECT 145.180 178.410 145.350 178.580 ;
        RECT 277.650 178.550 277.820 178.720 ;
        RECT 278.510 178.540 278.680 178.710 ;
        RECT 279.540 178.550 279.710 178.720 ;
        RECT 280.400 178.540 280.570 178.710 ;
        RECT 378.960 178.360 379.130 178.530 ;
        RECT 379.820 178.350 379.990 178.520 ;
        RECT 380.850 178.360 381.020 178.530 ;
        RECT 381.710 178.350 381.880 178.520 ;
        RECT 7.690 172.160 7.860 172.330 ;
        RECT 8.550 172.150 8.720 172.320 ;
        RECT 9.580 172.160 9.750 172.330 ;
        RECT 10.440 172.150 10.610 172.320 ;
        RECT 109.000 171.970 109.170 172.140 ;
        RECT 109.860 171.960 110.030 172.130 ;
        RECT 110.890 171.970 111.060 172.140 ;
        RECT 111.750 171.960 111.920 172.130 ;
        RECT 244.220 172.100 244.390 172.270 ;
        RECT 245.080 172.090 245.250 172.260 ;
        RECT 246.110 172.100 246.280 172.270 ;
        RECT 246.970 172.090 247.140 172.260 ;
        RECT 345.530 171.910 345.700 172.080 ;
        RECT 346.390 171.900 346.560 172.070 ;
        RECT 347.420 171.910 347.590 172.080 ;
        RECT 348.280 171.900 348.450 172.070 ;
        RECT 23.370 169.740 23.540 169.910 ;
        RECT 24.230 169.730 24.400 169.900 ;
        RECT 25.260 169.740 25.430 169.910 ;
        RECT 26.120 169.730 26.290 169.900 ;
        RECT 124.680 169.550 124.850 169.720 ;
        RECT 125.540 169.540 125.710 169.710 ;
        RECT 126.570 169.550 126.740 169.720 ;
        RECT 127.430 169.540 127.600 169.710 ;
        RECT 259.900 169.680 260.070 169.850 ;
        RECT 260.760 169.670 260.930 169.840 ;
        RECT 261.790 169.680 261.960 169.850 ;
        RECT 262.650 169.670 262.820 169.840 ;
        RECT 361.210 169.490 361.380 169.660 ;
        RECT 362.070 169.480 362.240 169.650 ;
        RECT 363.100 169.490 363.270 169.660 ;
        RECT 363.960 169.480 364.130 169.650 ;
        RECT 7.850 165.760 8.020 165.930 ;
        RECT 8.710 165.750 8.880 165.920 ;
        RECT 9.740 165.760 9.910 165.930 ;
        RECT 10.600 165.750 10.770 165.920 ;
        RECT 109.160 165.570 109.330 165.740 ;
        RECT 110.020 165.560 110.190 165.730 ;
        RECT 111.050 165.570 111.220 165.740 ;
        RECT 111.910 165.560 112.080 165.730 ;
        RECT 244.380 165.700 244.550 165.870 ;
        RECT 245.240 165.690 245.410 165.860 ;
        RECT 246.270 165.700 246.440 165.870 ;
        RECT 247.130 165.690 247.300 165.860 ;
        RECT 345.690 165.510 345.860 165.680 ;
        RECT 346.550 165.500 346.720 165.670 ;
        RECT 347.580 165.510 347.750 165.680 ;
        RECT 348.440 165.500 348.610 165.670 ;
        RECT 58.650 162.590 58.820 162.760 ;
        RECT 59.510 162.580 59.680 162.750 ;
        RECT 60.540 162.590 60.710 162.760 ;
        RECT 61.400 162.580 61.570 162.750 ;
        RECT 159.960 162.400 160.130 162.570 ;
        RECT 160.820 162.390 160.990 162.560 ;
        RECT 161.850 162.400 162.020 162.570 ;
        RECT 162.710 162.390 162.880 162.560 ;
        RECT 295.180 162.530 295.350 162.700 ;
        RECT 296.040 162.520 296.210 162.690 ;
        RECT 297.070 162.530 297.240 162.700 ;
        RECT 297.930 162.520 298.100 162.690 ;
        RECT 396.490 162.340 396.660 162.510 ;
        RECT 397.350 162.330 397.520 162.500 ;
        RECT 398.380 162.340 398.550 162.510 ;
        RECT 399.240 162.330 399.410 162.500 ;
        RECT 7.830 156.510 8.000 156.680 ;
        RECT 8.690 156.500 8.860 156.670 ;
        RECT 9.720 156.510 9.890 156.680 ;
        RECT 10.580 156.500 10.750 156.670 ;
        RECT 109.140 156.320 109.310 156.490 ;
        RECT 110.000 156.310 110.170 156.480 ;
        RECT 111.030 156.320 111.200 156.490 ;
        RECT 111.890 156.310 112.060 156.480 ;
        RECT 244.360 156.450 244.530 156.620 ;
        RECT 245.220 156.440 245.390 156.610 ;
        RECT 246.250 156.450 246.420 156.620 ;
        RECT 247.110 156.440 247.280 156.610 ;
        RECT 345.670 156.260 345.840 156.430 ;
        RECT 346.530 156.250 346.700 156.420 ;
        RECT 347.560 156.260 347.730 156.430 ;
        RECT 348.420 156.250 348.590 156.420 ;
        RECT 23.510 154.090 23.680 154.260 ;
        RECT 24.370 154.080 24.540 154.250 ;
        RECT 25.400 154.090 25.570 154.260 ;
        RECT 26.260 154.080 26.430 154.250 ;
        RECT 124.820 153.900 124.990 154.070 ;
        RECT 125.680 153.890 125.850 154.060 ;
        RECT 126.710 153.900 126.880 154.070 ;
        RECT 127.570 153.890 127.740 154.060 ;
        RECT 260.040 154.030 260.210 154.200 ;
        RECT 260.900 154.020 261.070 154.190 ;
        RECT 261.930 154.030 262.100 154.200 ;
        RECT 262.790 154.020 262.960 154.190 ;
        RECT 361.350 153.840 361.520 154.010 ;
        RECT 362.210 153.830 362.380 154.000 ;
        RECT 363.240 153.840 363.410 154.010 ;
        RECT 364.100 153.830 364.270 154.000 ;
        RECT 7.990 150.110 8.160 150.280 ;
        RECT 8.850 150.100 9.020 150.270 ;
        RECT 9.880 150.110 10.050 150.280 ;
        RECT 10.740 150.100 10.910 150.270 ;
        RECT 109.300 149.920 109.470 150.090 ;
        RECT 110.160 149.910 110.330 150.080 ;
        RECT 111.190 149.920 111.360 150.090 ;
        RECT 112.050 149.910 112.220 150.080 ;
        RECT 244.520 150.050 244.690 150.220 ;
        RECT 245.380 150.040 245.550 150.210 ;
        RECT 246.410 150.050 246.580 150.220 ;
        RECT 247.270 150.040 247.440 150.210 ;
        RECT 345.830 149.860 346.000 150.030 ;
        RECT 346.690 149.850 346.860 150.020 ;
        RECT 347.720 149.860 347.890 150.030 ;
        RECT 348.580 149.850 348.750 150.020 ;
        RECT 41.090 148.540 41.260 148.710 ;
        RECT 41.950 148.530 42.120 148.700 ;
        RECT 42.980 148.540 43.150 148.710 ;
        RECT 43.840 148.530 44.010 148.700 ;
        RECT 142.400 148.350 142.570 148.520 ;
        RECT 143.260 148.340 143.430 148.510 ;
        RECT 144.290 148.350 144.460 148.520 ;
        RECT 145.150 148.340 145.320 148.510 ;
        RECT 277.620 148.480 277.790 148.650 ;
        RECT 278.480 148.470 278.650 148.640 ;
        RECT 279.510 148.480 279.680 148.650 ;
        RECT 280.370 148.470 280.540 148.640 ;
        RECT 378.930 148.290 379.100 148.460 ;
        RECT 379.790 148.280 379.960 148.450 ;
        RECT 380.820 148.290 380.990 148.460 ;
        RECT 381.680 148.280 381.850 148.450 ;
        RECT 7.660 142.090 7.830 142.260 ;
        RECT 8.520 142.080 8.690 142.250 ;
        RECT 9.550 142.090 9.720 142.260 ;
        RECT 10.410 142.080 10.580 142.250 ;
        RECT 108.970 141.900 109.140 142.070 ;
        RECT 109.830 141.890 110.000 142.060 ;
        RECT 110.860 141.900 111.030 142.070 ;
        RECT 111.720 141.890 111.890 142.060 ;
        RECT 244.190 142.030 244.360 142.200 ;
        RECT 245.050 142.020 245.220 142.190 ;
        RECT 246.080 142.030 246.250 142.200 ;
        RECT 246.940 142.020 247.110 142.190 ;
        RECT 345.500 141.840 345.670 142.010 ;
        RECT 346.360 141.830 346.530 142.000 ;
        RECT 347.390 141.840 347.560 142.010 ;
        RECT 348.250 141.830 348.420 142.000 ;
        RECT 23.340 139.670 23.510 139.840 ;
        RECT 24.200 139.660 24.370 139.830 ;
        RECT 25.230 139.670 25.400 139.840 ;
        RECT 26.090 139.660 26.260 139.830 ;
        RECT 124.650 139.480 124.820 139.650 ;
        RECT 125.510 139.470 125.680 139.640 ;
        RECT 126.540 139.480 126.710 139.650 ;
        RECT 127.400 139.470 127.570 139.640 ;
        RECT 259.870 139.610 260.040 139.780 ;
        RECT 260.730 139.600 260.900 139.770 ;
        RECT 261.760 139.610 261.930 139.780 ;
        RECT 262.620 139.600 262.790 139.770 ;
        RECT 361.180 139.420 361.350 139.590 ;
        RECT 362.040 139.410 362.210 139.580 ;
        RECT 363.070 139.420 363.240 139.590 ;
        RECT 363.930 139.410 364.100 139.580 ;
        RECT 7.820 135.690 7.990 135.860 ;
        RECT 8.680 135.680 8.850 135.850 ;
        RECT 9.710 135.690 9.880 135.860 ;
        RECT 10.570 135.680 10.740 135.850 ;
        RECT 109.130 135.500 109.300 135.670 ;
        RECT 109.990 135.490 110.160 135.660 ;
        RECT 111.020 135.500 111.190 135.670 ;
        RECT 111.880 135.490 112.050 135.660 ;
        RECT 244.350 135.630 244.520 135.800 ;
        RECT 245.210 135.620 245.380 135.790 ;
        RECT 246.240 135.630 246.410 135.800 ;
        RECT 247.100 135.620 247.270 135.790 ;
        RECT 217.120 135.220 217.290 135.390 ;
        RECT 217.980 135.210 218.150 135.380 ;
        RECT 219.010 135.220 219.180 135.390 ;
        RECT 219.870 135.210 220.040 135.380 ;
        RECT 345.660 135.440 345.830 135.610 ;
        RECT 346.520 135.430 346.690 135.600 ;
        RECT 347.550 135.440 347.720 135.610 ;
        RECT 348.410 135.430 348.580 135.600 ;
        RECT 453.650 135.160 453.820 135.330 ;
        RECT 454.510 135.150 454.680 135.320 ;
        RECT 455.540 135.160 455.710 135.330 ;
        RECT 456.400 135.150 456.570 135.320 ;
        RECT 89.530 133.080 89.700 133.250 ;
        RECT 90.390 133.070 90.560 133.240 ;
        RECT 91.420 133.080 91.590 133.250 ;
        RECT 92.280 133.070 92.450 133.240 ;
        RECT 190.840 132.890 191.010 133.060 ;
        RECT 191.700 132.880 191.870 133.050 ;
        RECT 192.730 132.890 192.900 133.060 ;
        RECT 193.590 132.880 193.760 133.050 ;
        RECT 326.060 133.020 326.230 133.190 ;
        RECT 326.920 133.010 327.090 133.180 ;
        RECT 327.950 133.020 328.120 133.190 ;
        RECT 328.810 133.010 328.980 133.180 ;
        RECT 427.370 132.830 427.540 133.000 ;
        RECT 428.230 132.820 428.400 132.990 ;
        RECT 429.260 132.830 429.430 133.000 ;
        RECT 430.120 132.820 430.290 132.990 ;
        RECT 470.950 132.810 471.120 132.980 ;
        RECT 471.810 132.800 471.980 132.970 ;
        RECT 472.840 132.810 473.010 132.980 ;
        RECT 473.700 132.800 473.870 132.970 ;
        RECT 7.710 126.260 7.880 126.430 ;
        RECT 8.570 126.250 8.740 126.420 ;
        RECT 9.600 126.260 9.770 126.430 ;
        RECT 10.460 126.250 10.630 126.420 ;
        RECT 109.020 126.070 109.190 126.240 ;
        RECT 109.880 126.060 110.050 126.230 ;
        RECT 110.910 126.070 111.080 126.240 ;
        RECT 111.770 126.060 111.940 126.230 ;
        RECT 244.240 126.200 244.410 126.370 ;
        RECT 245.100 126.190 245.270 126.360 ;
        RECT 246.130 126.200 246.300 126.370 ;
        RECT 246.990 126.190 247.160 126.360 ;
        RECT 345.550 126.010 345.720 126.180 ;
        RECT 346.410 126.000 346.580 126.170 ;
        RECT 347.440 126.010 347.610 126.180 ;
        RECT 348.300 126.000 348.470 126.170 ;
        RECT 23.390 123.840 23.560 124.010 ;
        RECT 24.250 123.830 24.420 124.000 ;
        RECT 25.280 123.840 25.450 124.010 ;
        RECT 26.140 123.830 26.310 124.000 ;
        RECT 124.700 123.650 124.870 123.820 ;
        RECT 125.560 123.640 125.730 123.810 ;
        RECT 126.590 123.650 126.760 123.820 ;
        RECT 127.450 123.640 127.620 123.810 ;
        RECT 259.920 123.780 260.090 123.950 ;
        RECT 260.780 123.770 260.950 123.940 ;
        RECT 261.810 123.780 261.980 123.950 ;
        RECT 262.670 123.770 262.840 123.940 ;
        RECT 361.230 123.590 361.400 123.760 ;
        RECT 362.090 123.580 362.260 123.750 ;
        RECT 363.120 123.590 363.290 123.760 ;
        RECT 363.980 123.580 364.150 123.750 ;
        RECT 7.870 119.860 8.040 120.030 ;
        RECT 8.730 119.850 8.900 120.020 ;
        RECT 9.760 119.860 9.930 120.030 ;
        RECT 10.620 119.850 10.790 120.020 ;
        RECT 109.180 119.670 109.350 119.840 ;
        RECT 110.040 119.660 110.210 119.830 ;
        RECT 111.070 119.670 111.240 119.840 ;
        RECT 111.930 119.660 112.100 119.830 ;
        RECT 244.400 119.800 244.570 119.970 ;
        RECT 245.260 119.790 245.430 119.960 ;
        RECT 246.290 119.800 246.460 119.970 ;
        RECT 247.150 119.790 247.320 119.960 ;
        RECT 345.710 119.610 345.880 119.780 ;
        RECT 346.570 119.600 346.740 119.770 ;
        RECT 347.600 119.610 347.770 119.780 ;
        RECT 348.460 119.600 348.630 119.770 ;
        RECT 40.970 118.290 41.140 118.460 ;
        RECT 41.830 118.280 42.000 118.450 ;
        RECT 42.860 118.290 43.030 118.460 ;
        RECT 43.720 118.280 43.890 118.450 ;
        RECT 142.280 118.100 142.450 118.270 ;
        RECT 143.140 118.090 143.310 118.260 ;
        RECT 144.170 118.100 144.340 118.270 ;
        RECT 145.030 118.090 145.200 118.260 ;
        RECT 277.500 118.230 277.670 118.400 ;
        RECT 278.360 118.220 278.530 118.390 ;
        RECT 279.390 118.230 279.560 118.400 ;
        RECT 280.250 118.220 280.420 118.390 ;
        RECT 378.810 118.040 378.980 118.210 ;
        RECT 379.670 118.030 379.840 118.200 ;
        RECT 380.700 118.040 380.870 118.210 ;
        RECT 381.560 118.030 381.730 118.200 ;
        RECT 7.540 111.840 7.710 112.010 ;
        RECT 8.400 111.830 8.570 112.000 ;
        RECT 9.430 111.840 9.600 112.010 ;
        RECT 10.290 111.830 10.460 112.000 ;
        RECT 108.850 111.650 109.020 111.820 ;
        RECT 109.710 111.640 109.880 111.810 ;
        RECT 110.740 111.650 110.910 111.820 ;
        RECT 111.600 111.640 111.770 111.810 ;
        RECT 244.070 111.780 244.240 111.950 ;
        RECT 244.930 111.770 245.100 111.940 ;
        RECT 245.960 111.780 246.130 111.950 ;
        RECT 246.820 111.770 246.990 111.940 ;
        RECT 345.380 111.590 345.550 111.760 ;
        RECT 346.240 111.580 346.410 111.750 ;
        RECT 347.270 111.590 347.440 111.760 ;
        RECT 348.130 111.580 348.300 111.750 ;
        RECT 23.220 109.420 23.390 109.590 ;
        RECT 24.080 109.410 24.250 109.580 ;
        RECT 25.110 109.420 25.280 109.590 ;
        RECT 25.970 109.410 26.140 109.580 ;
        RECT 124.530 109.230 124.700 109.400 ;
        RECT 125.390 109.220 125.560 109.390 ;
        RECT 126.420 109.230 126.590 109.400 ;
        RECT 127.280 109.220 127.450 109.390 ;
        RECT 259.750 109.360 259.920 109.530 ;
        RECT 260.610 109.350 260.780 109.520 ;
        RECT 261.640 109.360 261.810 109.530 ;
        RECT 262.500 109.350 262.670 109.520 ;
        RECT 361.060 109.170 361.230 109.340 ;
        RECT 361.920 109.160 362.090 109.330 ;
        RECT 362.950 109.170 363.120 109.340 ;
        RECT 363.810 109.160 363.980 109.330 ;
        RECT 7.700 105.440 7.870 105.610 ;
        RECT 8.560 105.430 8.730 105.600 ;
        RECT 9.590 105.440 9.760 105.610 ;
        RECT 10.450 105.430 10.620 105.600 ;
        RECT 109.010 105.250 109.180 105.420 ;
        RECT 109.870 105.240 110.040 105.410 ;
        RECT 110.900 105.250 111.070 105.420 ;
        RECT 111.760 105.240 111.930 105.410 ;
        RECT 244.230 105.380 244.400 105.550 ;
        RECT 245.090 105.370 245.260 105.540 ;
        RECT 246.120 105.380 246.290 105.550 ;
        RECT 246.980 105.370 247.150 105.540 ;
        RECT 345.540 105.190 345.710 105.360 ;
        RECT 346.400 105.180 346.570 105.350 ;
        RECT 347.430 105.190 347.600 105.360 ;
        RECT 348.290 105.180 348.460 105.350 ;
        RECT 58.500 102.270 58.670 102.440 ;
        RECT 59.360 102.260 59.530 102.430 ;
        RECT 60.390 102.270 60.560 102.440 ;
        RECT 61.250 102.260 61.420 102.430 ;
        RECT 159.810 102.080 159.980 102.250 ;
        RECT 160.670 102.070 160.840 102.240 ;
        RECT 161.700 102.080 161.870 102.250 ;
        RECT 162.560 102.070 162.730 102.240 ;
        RECT 295.030 102.210 295.200 102.380 ;
        RECT 295.890 102.200 296.060 102.370 ;
        RECT 296.920 102.210 297.090 102.380 ;
        RECT 297.780 102.200 297.950 102.370 ;
        RECT 396.340 102.020 396.510 102.190 ;
        RECT 397.200 102.010 397.370 102.180 ;
        RECT 398.230 102.020 398.400 102.190 ;
        RECT 399.090 102.010 399.260 102.180 ;
        RECT 7.680 96.190 7.850 96.360 ;
        RECT 8.540 96.180 8.710 96.350 ;
        RECT 9.570 96.190 9.740 96.360 ;
        RECT 10.430 96.180 10.600 96.350 ;
        RECT 108.990 96.000 109.160 96.170 ;
        RECT 109.850 95.990 110.020 96.160 ;
        RECT 110.880 96.000 111.050 96.170 ;
        RECT 111.740 95.990 111.910 96.160 ;
        RECT 244.210 96.130 244.380 96.300 ;
        RECT 245.070 96.120 245.240 96.290 ;
        RECT 246.100 96.130 246.270 96.300 ;
        RECT 246.960 96.120 247.130 96.290 ;
        RECT 345.520 95.940 345.690 96.110 ;
        RECT 346.380 95.930 346.550 96.100 ;
        RECT 347.410 95.940 347.580 96.110 ;
        RECT 348.270 95.930 348.440 96.100 ;
        RECT 23.360 93.770 23.530 93.940 ;
        RECT 24.220 93.760 24.390 93.930 ;
        RECT 25.250 93.770 25.420 93.940 ;
        RECT 26.110 93.760 26.280 93.930 ;
        RECT 124.670 93.580 124.840 93.750 ;
        RECT 125.530 93.570 125.700 93.740 ;
        RECT 126.560 93.580 126.730 93.750 ;
        RECT 127.420 93.570 127.590 93.740 ;
        RECT 259.890 93.710 260.060 93.880 ;
        RECT 260.750 93.700 260.920 93.870 ;
        RECT 261.780 93.710 261.950 93.880 ;
        RECT 262.640 93.700 262.810 93.870 ;
        RECT 361.200 93.520 361.370 93.690 ;
        RECT 362.060 93.510 362.230 93.680 ;
        RECT 363.090 93.520 363.260 93.690 ;
        RECT 363.950 93.510 364.120 93.680 ;
        RECT 7.840 89.790 8.010 89.960 ;
        RECT 8.700 89.780 8.870 89.950 ;
        RECT 9.730 89.790 9.900 89.960 ;
        RECT 10.590 89.780 10.760 89.950 ;
        RECT 109.150 89.600 109.320 89.770 ;
        RECT 110.010 89.590 110.180 89.760 ;
        RECT 111.040 89.600 111.210 89.770 ;
        RECT 111.900 89.590 112.070 89.760 ;
        RECT 244.370 89.730 244.540 89.900 ;
        RECT 245.230 89.720 245.400 89.890 ;
        RECT 246.260 89.730 246.430 89.900 ;
        RECT 247.120 89.720 247.290 89.890 ;
        RECT 345.680 89.540 345.850 89.710 ;
        RECT 346.540 89.530 346.710 89.700 ;
        RECT 347.570 89.540 347.740 89.710 ;
        RECT 348.430 89.530 348.600 89.700 ;
        RECT 40.940 88.220 41.110 88.390 ;
        RECT 41.800 88.210 41.970 88.380 ;
        RECT 42.830 88.220 43.000 88.390 ;
        RECT 43.690 88.210 43.860 88.380 ;
        RECT 142.250 88.030 142.420 88.200 ;
        RECT 143.110 88.020 143.280 88.190 ;
        RECT 144.140 88.030 144.310 88.200 ;
        RECT 145.000 88.020 145.170 88.190 ;
        RECT 277.470 88.160 277.640 88.330 ;
        RECT 278.330 88.150 278.500 88.320 ;
        RECT 279.360 88.160 279.530 88.330 ;
        RECT 280.220 88.150 280.390 88.320 ;
        RECT 378.780 87.970 378.950 88.140 ;
        RECT 379.640 87.960 379.810 88.130 ;
        RECT 380.670 87.970 380.840 88.140 ;
        RECT 381.530 87.960 381.700 88.130 ;
        RECT 7.510 81.770 7.680 81.940 ;
        RECT 8.370 81.760 8.540 81.930 ;
        RECT 9.400 81.770 9.570 81.940 ;
        RECT 10.260 81.760 10.430 81.930 ;
        RECT 108.820 81.580 108.990 81.750 ;
        RECT 109.680 81.570 109.850 81.740 ;
        RECT 110.710 81.580 110.880 81.750 ;
        RECT 111.570 81.570 111.740 81.740 ;
        RECT 244.040 81.710 244.210 81.880 ;
        RECT 244.900 81.700 245.070 81.870 ;
        RECT 245.930 81.710 246.100 81.880 ;
        RECT 246.790 81.700 246.960 81.870 ;
        RECT 345.350 81.520 345.520 81.690 ;
        RECT 346.210 81.510 346.380 81.680 ;
        RECT 347.240 81.520 347.410 81.690 ;
        RECT 348.100 81.510 348.270 81.680 ;
        RECT 23.190 79.350 23.360 79.520 ;
        RECT 24.050 79.340 24.220 79.510 ;
        RECT 25.080 79.350 25.250 79.520 ;
        RECT 25.940 79.340 26.110 79.510 ;
        RECT 124.500 79.160 124.670 79.330 ;
        RECT 125.360 79.150 125.530 79.320 ;
        RECT 126.390 79.160 126.560 79.330 ;
        RECT 127.250 79.150 127.420 79.320 ;
        RECT 259.720 79.290 259.890 79.460 ;
        RECT 260.580 79.280 260.750 79.450 ;
        RECT 261.610 79.290 261.780 79.460 ;
        RECT 262.470 79.280 262.640 79.450 ;
        RECT 361.030 79.100 361.200 79.270 ;
        RECT 361.890 79.090 362.060 79.260 ;
        RECT 362.920 79.100 363.090 79.270 ;
        RECT 363.780 79.090 363.950 79.260 ;
        RECT 72.700 75.980 72.870 76.150 ;
        RECT 73.560 75.970 73.730 76.140 ;
        RECT 74.590 75.980 74.760 76.150 ;
        RECT 75.450 75.970 75.620 76.140 ;
        RECT 7.670 75.370 7.840 75.540 ;
        RECT 8.530 75.360 8.700 75.530 ;
        RECT 9.560 75.370 9.730 75.540 ;
        RECT 10.420 75.360 10.590 75.530 ;
        RECT 174.010 75.790 174.180 75.960 ;
        RECT 174.870 75.780 175.040 75.950 ;
        RECT 175.900 75.790 176.070 75.960 ;
        RECT 176.760 75.780 176.930 75.950 ;
        RECT 309.230 75.920 309.400 76.090 ;
        RECT 310.090 75.910 310.260 76.080 ;
        RECT 311.120 75.920 311.290 76.090 ;
        RECT 311.980 75.910 312.150 76.080 ;
        RECT 108.980 75.180 109.150 75.350 ;
        RECT 109.840 75.170 110.010 75.340 ;
        RECT 110.870 75.180 111.040 75.350 ;
        RECT 111.730 75.170 111.900 75.340 ;
        RECT 244.200 75.310 244.370 75.480 ;
        RECT 245.060 75.300 245.230 75.470 ;
        RECT 246.090 75.310 246.260 75.480 ;
        RECT 246.950 75.300 247.120 75.470 ;
        RECT 410.540 75.730 410.710 75.900 ;
        RECT 411.400 75.720 411.570 75.890 ;
        RECT 412.430 75.730 412.600 75.900 ;
        RECT 413.290 75.720 413.460 75.890 ;
        RECT 345.510 75.120 345.680 75.290 ;
        RECT 346.370 75.110 346.540 75.280 ;
        RECT 347.400 75.120 347.570 75.290 ;
        RECT 348.260 75.110 348.430 75.280 ;
        RECT 7.360 66.340 7.530 66.510 ;
        RECT 8.220 66.330 8.390 66.500 ;
        RECT 9.250 66.340 9.420 66.510 ;
        RECT 10.110 66.330 10.280 66.500 ;
        RECT 108.670 66.150 108.840 66.320 ;
        RECT 109.530 66.140 109.700 66.310 ;
        RECT 110.560 66.150 110.730 66.320 ;
        RECT 111.420 66.140 111.590 66.310 ;
        RECT 243.890 66.280 244.060 66.450 ;
        RECT 244.750 66.270 244.920 66.440 ;
        RECT 245.780 66.280 245.950 66.450 ;
        RECT 246.640 66.270 246.810 66.440 ;
        RECT 345.200 66.090 345.370 66.260 ;
        RECT 346.060 66.080 346.230 66.250 ;
        RECT 347.090 66.090 347.260 66.260 ;
        RECT 347.950 66.080 348.120 66.250 ;
        RECT 23.040 63.920 23.210 64.090 ;
        RECT 23.900 63.910 24.070 64.080 ;
        RECT 24.930 63.920 25.100 64.090 ;
        RECT 25.790 63.910 25.960 64.080 ;
        RECT 124.350 63.730 124.520 63.900 ;
        RECT 125.210 63.720 125.380 63.890 ;
        RECT 126.240 63.730 126.410 63.900 ;
        RECT 127.100 63.720 127.270 63.890 ;
        RECT 259.570 63.860 259.740 64.030 ;
        RECT 260.430 63.850 260.600 64.020 ;
        RECT 261.460 63.860 261.630 64.030 ;
        RECT 262.320 63.850 262.490 64.020 ;
        RECT 360.880 63.670 361.050 63.840 ;
        RECT 361.740 63.660 361.910 63.830 ;
        RECT 362.770 63.670 362.940 63.840 ;
        RECT 363.630 63.660 363.800 63.830 ;
        RECT 7.520 59.940 7.690 60.110 ;
        RECT 8.380 59.930 8.550 60.100 ;
        RECT 9.410 59.940 9.580 60.110 ;
        RECT 10.270 59.930 10.440 60.100 ;
        RECT 108.830 59.750 109.000 59.920 ;
        RECT 109.690 59.740 109.860 59.910 ;
        RECT 110.720 59.750 110.890 59.920 ;
        RECT 111.580 59.740 111.750 59.910 ;
        RECT 244.050 59.880 244.220 60.050 ;
        RECT 244.910 59.870 245.080 60.040 ;
        RECT 245.940 59.880 246.110 60.050 ;
        RECT 246.800 59.870 246.970 60.040 ;
        RECT 345.360 59.690 345.530 59.860 ;
        RECT 346.220 59.680 346.390 59.850 ;
        RECT 347.250 59.690 347.420 59.860 ;
        RECT 348.110 59.680 348.280 59.850 ;
        RECT 40.620 58.370 40.790 58.540 ;
        RECT 41.480 58.360 41.650 58.530 ;
        RECT 42.510 58.370 42.680 58.540 ;
        RECT 43.370 58.360 43.540 58.530 ;
        RECT 141.930 58.180 142.100 58.350 ;
        RECT 142.790 58.170 142.960 58.340 ;
        RECT 143.820 58.180 143.990 58.350 ;
        RECT 144.680 58.170 144.850 58.340 ;
        RECT 277.150 58.310 277.320 58.480 ;
        RECT 278.010 58.300 278.180 58.470 ;
        RECT 279.040 58.310 279.210 58.480 ;
        RECT 279.900 58.300 280.070 58.470 ;
        RECT 378.460 58.120 378.630 58.290 ;
        RECT 379.320 58.110 379.490 58.280 ;
        RECT 380.350 58.120 380.520 58.290 ;
        RECT 381.210 58.110 381.380 58.280 ;
        RECT 7.190 51.920 7.360 52.090 ;
        RECT 8.050 51.910 8.220 52.080 ;
        RECT 9.080 51.920 9.250 52.090 ;
        RECT 9.940 51.910 10.110 52.080 ;
        RECT 108.500 51.730 108.670 51.900 ;
        RECT 109.360 51.720 109.530 51.890 ;
        RECT 110.390 51.730 110.560 51.900 ;
        RECT 111.250 51.720 111.420 51.890 ;
        RECT 243.720 51.860 243.890 52.030 ;
        RECT 244.580 51.850 244.750 52.020 ;
        RECT 245.610 51.860 245.780 52.030 ;
        RECT 246.470 51.850 246.640 52.020 ;
        RECT 345.030 51.670 345.200 51.840 ;
        RECT 345.890 51.660 346.060 51.830 ;
        RECT 346.920 51.670 347.090 51.840 ;
        RECT 347.780 51.660 347.950 51.830 ;
        RECT 22.870 49.500 23.040 49.670 ;
        RECT 23.730 49.490 23.900 49.660 ;
        RECT 24.760 49.500 24.930 49.670 ;
        RECT 25.620 49.490 25.790 49.660 ;
        RECT 124.180 49.310 124.350 49.480 ;
        RECT 125.040 49.300 125.210 49.470 ;
        RECT 126.070 49.310 126.240 49.480 ;
        RECT 126.930 49.300 127.100 49.470 ;
        RECT 259.400 49.440 259.570 49.610 ;
        RECT 260.260 49.430 260.430 49.600 ;
        RECT 261.290 49.440 261.460 49.610 ;
        RECT 262.150 49.430 262.320 49.600 ;
        RECT 360.710 49.250 360.880 49.420 ;
        RECT 361.570 49.240 361.740 49.410 ;
        RECT 362.600 49.250 362.770 49.420 ;
        RECT 363.460 49.240 363.630 49.410 ;
        RECT 7.350 45.520 7.520 45.690 ;
        RECT 8.210 45.510 8.380 45.680 ;
        RECT 9.240 45.520 9.410 45.690 ;
        RECT 10.100 45.510 10.270 45.680 ;
        RECT 108.660 45.330 108.830 45.500 ;
        RECT 109.520 45.320 109.690 45.490 ;
        RECT 110.550 45.330 110.720 45.500 ;
        RECT 111.410 45.320 111.580 45.490 ;
        RECT 243.880 45.460 244.050 45.630 ;
        RECT 244.740 45.450 244.910 45.620 ;
        RECT 245.770 45.460 245.940 45.630 ;
        RECT 246.630 45.450 246.800 45.620 ;
        RECT 345.190 45.270 345.360 45.440 ;
        RECT 346.050 45.260 346.220 45.430 ;
        RECT 347.080 45.270 347.250 45.440 ;
        RECT 347.940 45.260 348.110 45.430 ;
        RECT 58.150 42.350 58.320 42.520 ;
        RECT 59.010 42.340 59.180 42.510 ;
        RECT 60.040 42.350 60.210 42.520 ;
        RECT 60.900 42.340 61.070 42.510 ;
        RECT 159.460 42.160 159.630 42.330 ;
        RECT 160.320 42.150 160.490 42.320 ;
        RECT 161.350 42.160 161.520 42.330 ;
        RECT 162.210 42.150 162.380 42.320 ;
        RECT 294.680 42.290 294.850 42.460 ;
        RECT 295.540 42.280 295.710 42.450 ;
        RECT 296.570 42.290 296.740 42.460 ;
        RECT 297.430 42.280 297.600 42.450 ;
        RECT 395.990 42.100 396.160 42.270 ;
        RECT 396.850 42.090 397.020 42.260 ;
        RECT 397.880 42.100 398.050 42.270 ;
        RECT 398.740 42.090 398.910 42.260 ;
        RECT 7.330 36.270 7.500 36.440 ;
        RECT 8.190 36.260 8.360 36.430 ;
        RECT 9.220 36.270 9.390 36.440 ;
        RECT 10.080 36.260 10.250 36.430 ;
        RECT 108.640 36.080 108.810 36.250 ;
        RECT 109.500 36.070 109.670 36.240 ;
        RECT 110.530 36.080 110.700 36.250 ;
        RECT 111.390 36.070 111.560 36.240 ;
        RECT 243.860 36.210 244.030 36.380 ;
        RECT 244.720 36.200 244.890 36.370 ;
        RECT 245.750 36.210 245.920 36.380 ;
        RECT 246.610 36.200 246.780 36.370 ;
        RECT 345.170 36.020 345.340 36.190 ;
        RECT 346.030 36.010 346.200 36.180 ;
        RECT 347.060 36.020 347.230 36.190 ;
        RECT 347.920 36.010 348.090 36.180 ;
        RECT 23.010 33.850 23.180 34.020 ;
        RECT 23.870 33.840 24.040 34.010 ;
        RECT 24.900 33.850 25.070 34.020 ;
        RECT 25.760 33.840 25.930 34.010 ;
        RECT 124.320 33.660 124.490 33.830 ;
        RECT 125.180 33.650 125.350 33.820 ;
        RECT 126.210 33.660 126.380 33.830 ;
        RECT 127.070 33.650 127.240 33.820 ;
        RECT 259.540 33.790 259.710 33.960 ;
        RECT 260.400 33.780 260.570 33.950 ;
        RECT 261.430 33.790 261.600 33.960 ;
        RECT 262.290 33.780 262.460 33.950 ;
        RECT 360.850 33.600 361.020 33.770 ;
        RECT 361.710 33.590 361.880 33.760 ;
        RECT 362.740 33.600 362.910 33.770 ;
        RECT 363.600 33.590 363.770 33.760 ;
        RECT 7.490 29.870 7.660 30.040 ;
        RECT 8.350 29.860 8.520 30.030 ;
        RECT 9.380 29.870 9.550 30.040 ;
        RECT 10.240 29.860 10.410 30.030 ;
        RECT 108.800 29.680 108.970 29.850 ;
        RECT 109.660 29.670 109.830 29.840 ;
        RECT 110.690 29.680 110.860 29.850 ;
        RECT 111.550 29.670 111.720 29.840 ;
        RECT 244.020 29.810 244.190 29.980 ;
        RECT 244.880 29.800 245.050 29.970 ;
        RECT 245.910 29.810 246.080 29.980 ;
        RECT 246.770 29.800 246.940 29.970 ;
        RECT 345.330 29.620 345.500 29.790 ;
        RECT 346.190 29.610 346.360 29.780 ;
        RECT 347.220 29.620 347.390 29.790 ;
        RECT 348.080 29.610 348.250 29.780 ;
        RECT 40.590 28.300 40.760 28.470 ;
        RECT 41.450 28.290 41.620 28.460 ;
        RECT 42.480 28.300 42.650 28.470 ;
        RECT 43.340 28.290 43.510 28.460 ;
        RECT 141.900 28.110 142.070 28.280 ;
        RECT 142.760 28.100 142.930 28.270 ;
        RECT 143.790 28.110 143.960 28.280 ;
        RECT 144.650 28.100 144.820 28.270 ;
        RECT 277.120 28.240 277.290 28.410 ;
        RECT 277.980 28.230 278.150 28.400 ;
        RECT 279.010 28.240 279.180 28.410 ;
        RECT 279.870 28.230 280.040 28.400 ;
        RECT 378.430 28.050 378.600 28.220 ;
        RECT 379.290 28.040 379.460 28.210 ;
        RECT 380.320 28.050 380.490 28.220 ;
        RECT 381.180 28.040 381.350 28.210 ;
        RECT 7.160 21.850 7.330 22.020 ;
        RECT 8.020 21.840 8.190 22.010 ;
        RECT 9.050 21.850 9.220 22.020 ;
        RECT 9.910 21.840 10.080 22.010 ;
        RECT 108.470 21.660 108.640 21.830 ;
        RECT 109.330 21.650 109.500 21.820 ;
        RECT 110.360 21.660 110.530 21.830 ;
        RECT 111.220 21.650 111.390 21.820 ;
        RECT 243.690 21.790 243.860 21.960 ;
        RECT 244.550 21.780 244.720 21.950 ;
        RECT 245.580 21.790 245.750 21.960 ;
        RECT 246.440 21.780 246.610 21.950 ;
        RECT 345.000 21.600 345.170 21.770 ;
        RECT 345.860 21.590 346.030 21.760 ;
        RECT 346.890 21.600 347.060 21.770 ;
        RECT 347.750 21.590 347.920 21.760 ;
        RECT 22.840 19.430 23.010 19.600 ;
        RECT 23.700 19.420 23.870 19.590 ;
        RECT 24.730 19.430 24.900 19.600 ;
        RECT 25.590 19.420 25.760 19.590 ;
        RECT 124.150 19.240 124.320 19.410 ;
        RECT 125.010 19.230 125.180 19.400 ;
        RECT 126.040 19.240 126.210 19.410 ;
        RECT 126.900 19.230 127.070 19.400 ;
        RECT 259.370 19.370 259.540 19.540 ;
        RECT 260.230 19.360 260.400 19.530 ;
        RECT 261.260 19.370 261.430 19.540 ;
        RECT 262.120 19.360 262.290 19.530 ;
        RECT 360.680 19.180 360.850 19.350 ;
        RECT 361.540 19.170 361.710 19.340 ;
        RECT 362.570 19.180 362.740 19.350 ;
        RECT 363.430 19.170 363.600 19.340 ;
        RECT 7.320 15.450 7.490 15.620 ;
        RECT 8.180 15.440 8.350 15.610 ;
        RECT 9.210 15.450 9.380 15.620 ;
        RECT 10.070 15.440 10.240 15.610 ;
        RECT 108.630 15.260 108.800 15.430 ;
        RECT 109.490 15.250 109.660 15.420 ;
        RECT 110.520 15.260 110.690 15.430 ;
        RECT 111.380 15.250 111.550 15.420 ;
        RECT 243.850 15.390 244.020 15.560 ;
        RECT 244.710 15.380 244.880 15.550 ;
        RECT 245.740 15.390 245.910 15.560 ;
        RECT 246.600 15.380 246.770 15.550 ;
        RECT 345.160 15.200 345.330 15.370 ;
        RECT 346.020 15.190 346.190 15.360 ;
        RECT 347.050 15.200 347.220 15.370 ;
        RECT 347.910 15.190 348.080 15.360 ;
      LAYER met1 ;
        RECT 7.700 246.150 11.290 246.860 ;
        RECT 7.700 246.140 8.000 246.150 ;
        RECT 109.010 245.960 112.600 246.670 ;
        RECT 244.230 246.090 247.820 246.800 ;
        RECT 244.230 246.080 244.530 246.090 ;
        RECT 109.010 245.950 109.310 245.960 ;
        RECT 345.540 245.900 349.130 246.610 ;
        RECT 345.540 245.890 345.840 245.900 ;
        RECT 23.320 244.440 23.730 244.450 ;
        RECT 23.320 243.740 26.970 244.440 ;
        RECT 259.850 244.380 260.260 244.390 ;
        RECT 23.460 243.730 26.970 243.740 ;
        RECT 124.630 244.250 125.040 244.260 ;
        RECT 124.630 243.550 128.280 244.250 ;
        RECT 259.850 243.680 263.500 244.380 ;
        RECT 259.990 243.670 263.500 243.680 ;
        RECT 361.160 244.190 361.570 244.200 ;
        RECT 124.770 243.540 128.280 243.550 ;
        RECT 361.160 243.490 364.810 244.190 ;
        RECT 361.300 243.480 364.810 243.490 ;
        RECT 7.880 240.460 8.180 240.470 ;
        RECT 7.880 239.750 11.450 240.460 ;
        RECT 244.410 240.400 244.710 240.410 ;
        RECT 109.190 240.270 109.490 240.280 ;
        RECT 109.190 239.560 112.760 240.270 ;
        RECT 244.410 239.690 247.980 240.400 ;
        RECT 345.720 240.210 346.020 240.220 ;
        RECT 345.720 239.500 349.290 240.210 ;
        RECT 40.910 238.890 41.290 238.900 ;
        RECT 40.910 238.180 44.550 238.890 ;
        RECT 277.440 238.830 277.820 238.840 ;
        RECT 142.220 238.700 142.600 238.710 ;
        RECT 142.220 237.990 145.860 238.700 ;
        RECT 277.440 238.120 281.080 238.830 ;
        RECT 378.750 238.640 379.130 238.650 ;
        RECT 378.750 237.930 382.390 238.640 ;
        RECT 7.530 231.730 11.120 232.440 ;
        RECT 7.530 231.720 7.830 231.730 ;
        RECT 108.840 231.540 112.430 232.250 ;
        RECT 244.060 231.670 247.650 232.380 ;
        RECT 244.060 231.660 244.360 231.670 ;
        RECT 108.840 231.530 109.140 231.540 ;
        RECT 345.370 231.480 348.960 232.190 ;
        RECT 345.370 231.470 345.670 231.480 ;
        RECT 23.150 230.020 23.560 230.030 ;
        RECT 23.150 229.320 26.800 230.020 ;
        RECT 259.680 229.960 260.090 229.970 ;
        RECT 23.290 229.310 26.800 229.320 ;
        RECT 124.460 229.830 124.870 229.840 ;
        RECT 124.460 229.130 128.110 229.830 ;
        RECT 259.680 229.260 263.330 229.960 ;
        RECT 259.820 229.250 263.330 229.260 ;
        RECT 360.990 229.770 361.400 229.780 ;
        RECT 124.600 229.120 128.110 229.130 ;
        RECT 360.990 229.070 364.640 229.770 ;
        RECT 361.130 229.060 364.640 229.070 ;
        RECT 7.710 226.040 8.010 226.050 ;
        RECT 7.710 225.330 11.280 226.040 ;
        RECT 244.240 225.980 244.540 225.990 ;
        RECT 109.020 225.850 109.320 225.860 ;
        RECT 109.020 225.140 112.590 225.850 ;
        RECT 244.240 225.270 247.810 225.980 ;
        RECT 345.550 225.790 345.850 225.800 ;
        RECT 345.550 225.080 349.120 225.790 ;
        RECT 58.780 222.860 62.080 222.870 ;
        RECT 58.310 222.160 62.080 222.860 ;
        RECT 295.310 222.800 298.610 222.810 ;
        RECT 160.090 222.670 163.390 222.680 ;
        RECT 58.310 222.130 58.890 222.160 ;
        RECT 159.620 221.970 163.390 222.670 ;
        RECT 294.840 222.100 298.610 222.800 ;
        RECT 396.620 222.610 399.920 222.620 ;
        RECT 294.840 222.070 295.420 222.100 ;
        RECT 159.620 221.940 160.200 221.970 ;
        RECT 396.150 221.910 399.920 222.610 ;
        RECT 396.150 221.880 396.730 221.910 ;
        RECT 7.670 216.080 11.260 216.790 ;
        RECT 7.670 216.070 7.970 216.080 ;
        RECT 108.980 215.890 112.570 216.600 ;
        RECT 244.200 216.020 247.790 216.730 ;
        RECT 244.200 216.010 244.500 216.020 ;
        RECT 108.980 215.880 109.280 215.890 ;
        RECT 345.510 215.830 349.100 216.540 ;
        RECT 345.510 215.820 345.810 215.830 ;
        RECT 23.290 214.370 23.700 214.380 ;
        RECT 23.290 213.670 26.940 214.370 ;
        RECT 259.820 214.310 260.230 214.320 ;
        RECT 23.430 213.660 26.940 213.670 ;
        RECT 124.600 214.180 125.010 214.190 ;
        RECT 124.600 213.480 128.250 214.180 ;
        RECT 259.820 213.610 263.470 214.310 ;
        RECT 259.960 213.600 263.470 213.610 ;
        RECT 361.130 214.120 361.540 214.130 ;
        RECT 124.740 213.470 128.250 213.480 ;
        RECT 361.130 213.420 364.780 214.120 ;
        RECT 361.270 213.410 364.780 213.420 ;
        RECT 7.850 210.390 8.150 210.400 ;
        RECT 7.850 209.680 11.420 210.390 ;
        RECT 244.380 210.330 244.680 210.340 ;
        RECT 109.160 210.200 109.460 210.210 ;
        RECT 109.160 209.490 112.730 210.200 ;
        RECT 244.380 209.620 247.950 210.330 ;
        RECT 345.690 210.140 345.990 210.150 ;
        RECT 345.690 209.430 349.260 210.140 ;
        RECT 40.880 208.820 41.260 208.830 ;
        RECT 40.880 208.110 44.520 208.820 ;
        RECT 277.410 208.760 277.790 208.770 ;
        RECT 142.190 208.630 142.570 208.640 ;
        RECT 142.190 207.920 145.830 208.630 ;
        RECT 277.410 208.050 281.050 208.760 ;
        RECT 378.720 208.570 379.100 208.580 ;
        RECT 378.720 207.860 382.360 208.570 ;
        RECT 7.500 201.660 11.090 202.370 ;
        RECT 7.500 201.650 7.800 201.660 ;
        RECT 108.810 201.470 112.400 202.180 ;
        RECT 244.030 201.600 247.620 202.310 ;
        RECT 244.030 201.590 244.330 201.600 ;
        RECT 108.810 201.460 109.110 201.470 ;
        RECT 345.340 201.410 348.930 202.120 ;
        RECT 345.340 201.400 345.640 201.410 ;
        RECT 23.120 199.950 23.530 199.960 ;
        RECT 23.120 199.250 26.770 199.950 ;
        RECT 259.650 199.890 260.060 199.900 ;
        RECT 23.260 199.240 26.770 199.250 ;
        RECT 124.430 199.760 124.840 199.770 ;
        RECT 124.430 199.060 128.080 199.760 ;
        RECT 259.650 199.190 263.300 199.890 ;
        RECT 259.790 199.180 263.300 199.190 ;
        RECT 360.960 199.700 361.370 199.710 ;
        RECT 124.570 199.050 128.080 199.060 ;
        RECT 360.960 199.000 364.610 199.700 ;
        RECT 361.100 198.990 364.610 199.000 ;
        RECT 72.500 196.580 73.060 196.600 ;
        RECT 7.680 195.970 7.980 195.980 ;
        RECT 7.680 195.260 11.250 195.970 ;
        RECT 72.500 195.880 76.280 196.580 ;
        RECT 309.030 196.520 309.590 196.540 ;
        RECT 72.980 195.870 76.280 195.880 ;
        RECT 173.810 196.390 174.370 196.410 ;
        RECT 108.990 195.780 109.290 195.790 ;
        RECT 108.990 195.070 112.560 195.780 ;
        RECT 173.810 195.690 177.590 196.390 ;
        RECT 174.290 195.680 177.590 195.690 ;
        RECT 244.210 195.910 244.510 195.920 ;
        RECT 244.210 195.200 247.780 195.910 ;
        RECT 309.030 195.820 312.810 196.520 ;
        RECT 309.510 195.810 312.810 195.820 ;
        RECT 410.340 196.330 410.900 196.350 ;
        RECT 345.520 195.720 345.820 195.730 ;
        RECT 345.520 195.010 349.090 195.720 ;
        RECT 410.340 195.630 414.120 196.330 ;
        RECT 410.820 195.620 414.120 195.630 ;
        RECT 7.350 186.230 10.940 186.940 ;
        RECT 7.350 186.220 7.650 186.230 ;
        RECT 108.660 186.040 112.250 186.750 ;
        RECT 243.880 186.170 247.470 186.880 ;
        RECT 243.880 186.160 244.180 186.170 ;
        RECT 108.660 186.030 108.960 186.040 ;
        RECT 345.190 185.980 348.780 186.690 ;
        RECT 345.190 185.970 345.490 185.980 ;
        RECT 22.970 184.520 23.380 184.530 ;
        RECT 22.970 183.820 26.620 184.520 ;
        RECT 259.500 184.460 259.910 184.470 ;
        RECT 23.110 183.810 26.620 183.820 ;
        RECT 124.280 184.330 124.690 184.340 ;
        RECT 124.280 183.630 127.930 184.330 ;
        RECT 259.500 183.760 263.150 184.460 ;
        RECT 259.640 183.750 263.150 183.760 ;
        RECT 360.810 184.270 361.220 184.280 ;
        RECT 124.420 183.620 127.930 183.630 ;
        RECT 360.810 183.570 364.460 184.270 ;
        RECT 360.950 183.560 364.460 183.570 ;
        RECT 7.530 180.540 7.830 180.550 ;
        RECT 7.530 179.830 11.100 180.540 ;
        RECT 244.060 180.480 244.360 180.490 ;
        RECT 108.840 180.350 109.140 180.360 ;
        RECT 108.840 179.640 112.410 180.350 ;
        RECT 244.060 179.770 247.630 180.480 ;
        RECT 345.370 180.290 345.670 180.300 ;
        RECT 345.370 179.580 348.940 180.290 ;
        RECT 40.560 178.970 40.940 178.980 ;
        RECT 40.560 178.260 44.200 178.970 ;
        RECT 277.090 178.910 277.470 178.920 ;
        RECT 141.870 178.780 142.250 178.790 ;
        RECT 141.870 178.070 145.510 178.780 ;
        RECT 277.090 178.200 280.730 178.910 ;
        RECT 378.400 178.720 378.780 178.730 ;
        RECT 378.400 178.010 382.040 178.720 ;
        RECT 7.180 171.810 10.770 172.520 ;
        RECT 7.180 171.800 7.480 171.810 ;
        RECT 108.490 171.620 112.080 172.330 ;
        RECT 243.710 171.750 247.300 172.460 ;
        RECT 243.710 171.740 244.010 171.750 ;
        RECT 108.490 171.610 108.790 171.620 ;
        RECT 345.020 171.560 348.610 172.270 ;
        RECT 345.020 171.550 345.320 171.560 ;
        RECT 22.800 170.100 23.210 170.110 ;
        RECT 22.800 169.400 26.450 170.100 ;
        RECT 259.330 170.040 259.740 170.050 ;
        RECT 22.940 169.390 26.450 169.400 ;
        RECT 124.110 169.910 124.520 169.920 ;
        RECT 124.110 169.210 127.760 169.910 ;
        RECT 259.330 169.340 262.980 170.040 ;
        RECT 259.470 169.330 262.980 169.340 ;
        RECT 360.640 169.850 361.050 169.860 ;
        RECT 124.250 169.200 127.760 169.210 ;
        RECT 360.640 169.150 364.290 169.850 ;
        RECT 360.780 169.140 364.290 169.150 ;
        RECT 7.360 166.120 7.660 166.130 ;
        RECT 7.360 165.410 10.930 166.120 ;
        RECT 243.890 166.060 244.190 166.070 ;
        RECT 108.670 165.930 108.970 165.940 ;
        RECT 108.670 165.220 112.240 165.930 ;
        RECT 243.890 165.350 247.460 166.060 ;
        RECT 345.200 165.870 345.500 165.880 ;
        RECT 345.200 165.160 348.770 165.870 ;
        RECT 58.430 162.940 61.730 162.950 ;
        RECT 57.960 162.240 61.730 162.940 ;
        RECT 294.960 162.880 298.260 162.890 ;
        RECT 159.740 162.750 163.040 162.760 ;
        RECT 57.960 162.210 58.540 162.240 ;
        RECT 159.270 162.050 163.040 162.750 ;
        RECT 294.490 162.180 298.260 162.880 ;
        RECT 396.270 162.690 399.570 162.700 ;
        RECT 294.490 162.150 295.070 162.180 ;
        RECT 159.270 162.020 159.850 162.050 ;
        RECT 395.800 161.990 399.570 162.690 ;
        RECT 395.800 161.960 396.380 161.990 ;
        RECT 7.320 156.160 10.910 156.870 ;
        RECT 7.320 156.150 7.620 156.160 ;
        RECT 108.630 155.970 112.220 156.680 ;
        RECT 243.850 156.100 247.440 156.810 ;
        RECT 243.850 156.090 244.150 156.100 ;
        RECT 108.630 155.960 108.930 155.970 ;
        RECT 345.160 155.910 348.750 156.620 ;
        RECT 345.160 155.900 345.460 155.910 ;
        RECT 22.940 154.450 23.350 154.460 ;
        RECT 22.940 153.750 26.590 154.450 ;
        RECT 259.470 154.390 259.880 154.400 ;
        RECT 23.080 153.740 26.590 153.750 ;
        RECT 124.250 154.260 124.660 154.270 ;
        RECT 124.250 153.560 127.900 154.260 ;
        RECT 259.470 153.690 263.120 154.390 ;
        RECT 259.610 153.680 263.120 153.690 ;
        RECT 360.780 154.200 361.190 154.210 ;
        RECT 124.390 153.550 127.900 153.560 ;
        RECT 360.780 153.500 364.430 154.200 ;
        RECT 360.920 153.490 364.430 153.500 ;
        RECT 7.500 150.470 7.800 150.480 ;
        RECT 7.500 149.760 11.070 150.470 ;
        RECT 244.030 150.410 244.330 150.420 ;
        RECT 108.810 150.280 109.110 150.290 ;
        RECT 108.810 149.570 112.380 150.280 ;
        RECT 244.030 149.700 247.600 150.410 ;
        RECT 345.340 150.220 345.640 150.230 ;
        RECT 345.340 149.510 348.910 150.220 ;
        RECT 40.530 148.900 40.910 148.910 ;
        RECT 40.530 148.190 44.170 148.900 ;
        RECT 277.060 148.840 277.440 148.850 ;
        RECT 141.840 148.710 142.220 148.720 ;
        RECT 141.840 148.000 145.480 148.710 ;
        RECT 277.060 148.130 280.700 148.840 ;
        RECT 378.370 148.650 378.750 148.660 ;
        RECT 378.370 147.940 382.010 148.650 ;
        RECT 7.150 141.740 10.740 142.450 ;
        RECT 7.150 141.730 7.450 141.740 ;
        RECT 108.460 141.550 112.050 142.260 ;
        RECT 243.680 141.680 247.270 142.390 ;
        RECT 243.680 141.670 243.980 141.680 ;
        RECT 108.460 141.540 108.760 141.550 ;
        RECT 344.990 141.490 348.580 142.200 ;
        RECT 344.990 141.480 345.290 141.490 ;
        RECT 22.770 140.030 23.180 140.040 ;
        RECT 22.770 139.330 26.420 140.030 ;
        RECT 259.300 139.970 259.710 139.980 ;
        RECT 22.910 139.320 26.420 139.330 ;
        RECT 124.080 139.840 124.490 139.850 ;
        RECT 124.080 139.140 127.730 139.840 ;
        RECT 259.300 139.270 262.950 139.970 ;
        RECT 259.440 139.260 262.950 139.270 ;
        RECT 360.610 139.780 361.020 139.790 ;
        RECT 124.220 139.130 127.730 139.140 ;
        RECT 360.610 139.080 364.260 139.780 ;
        RECT 360.750 139.070 364.260 139.080 ;
        RECT 7.330 136.050 7.630 136.060 ;
        RECT 7.330 135.340 10.900 136.050 ;
        RECT 243.860 135.990 244.160 136.000 ;
        RECT 108.640 135.860 108.940 135.870 ;
        RECT 108.640 135.150 112.210 135.860 ;
        RECT 216.510 135.580 216.930 135.590 ;
        RECT 216.510 134.870 220.200 135.580 ;
        RECT 243.860 135.280 247.430 135.990 ;
        RECT 345.170 135.800 345.470 135.810 ;
        RECT 345.170 135.090 348.740 135.800 ;
        RECT 453.040 135.520 453.460 135.530 ;
        RECT 453.040 134.810 456.730 135.520 ;
        RECT 88.740 132.730 92.610 133.440 ;
        RECT 190.050 132.540 193.920 133.250 ;
        RECT 325.270 132.670 329.140 133.380 ;
        RECT 426.580 132.480 430.450 133.190 ;
        RECT 470.730 133.150 474.030 133.170 ;
        RECT 470.240 132.460 474.030 133.150 ;
        RECT 7.200 125.910 10.790 126.620 ;
        RECT 7.200 125.900 7.500 125.910 ;
        RECT 108.510 125.720 112.100 126.430 ;
        RECT 243.730 125.850 247.320 126.560 ;
        RECT 243.730 125.840 244.030 125.850 ;
        RECT 108.510 125.710 108.810 125.720 ;
        RECT 345.040 125.660 348.630 126.370 ;
        RECT 345.040 125.650 345.340 125.660 ;
        RECT 22.820 124.200 23.230 124.210 ;
        RECT 22.820 123.500 26.470 124.200 ;
        RECT 259.350 124.140 259.760 124.150 ;
        RECT 22.960 123.490 26.470 123.500 ;
        RECT 124.130 124.010 124.540 124.020 ;
        RECT 124.130 123.310 127.780 124.010 ;
        RECT 259.350 123.440 263.000 124.140 ;
        RECT 259.490 123.430 263.000 123.440 ;
        RECT 360.660 123.950 361.070 123.960 ;
        RECT 124.270 123.300 127.780 123.310 ;
        RECT 360.660 123.250 364.310 123.950 ;
        RECT 360.800 123.240 364.310 123.250 ;
        RECT 7.380 120.220 7.680 120.230 ;
        RECT 7.380 119.510 10.950 120.220 ;
        RECT 243.910 120.160 244.210 120.170 ;
        RECT 108.690 120.030 108.990 120.040 ;
        RECT 108.690 119.320 112.260 120.030 ;
        RECT 243.910 119.450 247.480 120.160 ;
        RECT 345.220 119.970 345.520 119.980 ;
        RECT 345.220 119.260 348.790 119.970 ;
        RECT 40.410 118.650 40.790 118.660 ;
        RECT 40.410 117.940 44.050 118.650 ;
        RECT 276.940 118.590 277.320 118.600 ;
        RECT 141.720 118.460 142.100 118.470 ;
        RECT 141.720 117.750 145.360 118.460 ;
        RECT 276.940 117.880 280.580 118.590 ;
        RECT 378.250 118.400 378.630 118.410 ;
        RECT 378.250 117.690 381.890 118.400 ;
        RECT 7.030 111.490 10.620 112.200 ;
        RECT 7.030 111.480 7.330 111.490 ;
        RECT 108.340 111.300 111.930 112.010 ;
        RECT 243.560 111.430 247.150 112.140 ;
        RECT 243.560 111.420 243.860 111.430 ;
        RECT 108.340 111.290 108.640 111.300 ;
        RECT 344.870 111.240 348.460 111.950 ;
        RECT 344.870 111.230 345.170 111.240 ;
        RECT 22.650 109.780 23.060 109.790 ;
        RECT 22.650 109.080 26.300 109.780 ;
        RECT 259.180 109.720 259.590 109.730 ;
        RECT 22.790 109.070 26.300 109.080 ;
        RECT 123.960 109.590 124.370 109.600 ;
        RECT 123.960 108.890 127.610 109.590 ;
        RECT 259.180 109.020 262.830 109.720 ;
        RECT 259.320 109.010 262.830 109.020 ;
        RECT 360.490 109.530 360.900 109.540 ;
        RECT 124.100 108.880 127.610 108.890 ;
        RECT 360.490 108.830 364.140 109.530 ;
        RECT 360.630 108.820 364.140 108.830 ;
        RECT 7.210 105.800 7.510 105.810 ;
        RECT 7.210 105.090 10.780 105.800 ;
        RECT 243.740 105.740 244.040 105.750 ;
        RECT 108.520 105.610 108.820 105.620 ;
        RECT 108.520 104.900 112.090 105.610 ;
        RECT 243.740 105.030 247.310 105.740 ;
        RECT 345.050 105.550 345.350 105.560 ;
        RECT 345.050 104.840 348.620 105.550 ;
        RECT 58.280 102.620 61.580 102.630 ;
        RECT 57.810 101.920 61.580 102.620 ;
        RECT 294.810 102.560 298.110 102.570 ;
        RECT 159.590 102.430 162.890 102.440 ;
        RECT 57.810 101.890 58.390 101.920 ;
        RECT 159.120 101.730 162.890 102.430 ;
        RECT 294.340 101.860 298.110 102.560 ;
        RECT 396.120 102.370 399.420 102.380 ;
        RECT 294.340 101.830 294.920 101.860 ;
        RECT 159.120 101.700 159.700 101.730 ;
        RECT 395.650 101.670 399.420 102.370 ;
        RECT 395.650 101.640 396.230 101.670 ;
        RECT 7.170 95.840 10.760 96.550 ;
        RECT 7.170 95.830 7.470 95.840 ;
        RECT 108.480 95.650 112.070 96.360 ;
        RECT 243.700 95.780 247.290 96.490 ;
        RECT 243.700 95.770 244.000 95.780 ;
        RECT 108.480 95.640 108.780 95.650 ;
        RECT 345.010 95.590 348.600 96.300 ;
        RECT 345.010 95.580 345.310 95.590 ;
        RECT 22.790 94.130 23.200 94.140 ;
        RECT 22.790 93.430 26.440 94.130 ;
        RECT 259.320 94.070 259.730 94.080 ;
        RECT 22.930 93.420 26.440 93.430 ;
        RECT 124.100 93.940 124.510 93.950 ;
        RECT 124.100 93.240 127.750 93.940 ;
        RECT 259.320 93.370 262.970 94.070 ;
        RECT 259.460 93.360 262.970 93.370 ;
        RECT 360.630 93.880 361.040 93.890 ;
        RECT 124.240 93.230 127.750 93.240 ;
        RECT 360.630 93.180 364.280 93.880 ;
        RECT 360.770 93.170 364.280 93.180 ;
        RECT 7.350 90.150 7.650 90.160 ;
        RECT 7.350 89.440 10.920 90.150 ;
        RECT 243.880 90.090 244.180 90.100 ;
        RECT 108.660 89.960 108.960 89.970 ;
        RECT 108.660 89.250 112.230 89.960 ;
        RECT 243.880 89.380 247.450 90.090 ;
        RECT 345.190 89.900 345.490 89.910 ;
        RECT 345.190 89.190 348.760 89.900 ;
        RECT 40.380 88.580 40.760 88.590 ;
        RECT 40.380 87.870 44.020 88.580 ;
        RECT 276.910 88.520 277.290 88.530 ;
        RECT 141.690 88.390 142.070 88.400 ;
        RECT 141.690 87.680 145.330 88.390 ;
        RECT 276.910 87.810 280.550 88.520 ;
        RECT 378.220 88.330 378.600 88.340 ;
        RECT 378.220 87.620 381.860 88.330 ;
        RECT 7.000 81.420 10.590 82.130 ;
        RECT 7.000 81.410 7.300 81.420 ;
        RECT 108.310 81.230 111.900 81.940 ;
        RECT 243.530 81.360 247.120 82.070 ;
        RECT 243.530 81.350 243.830 81.360 ;
        RECT 108.310 81.220 108.610 81.230 ;
        RECT 344.840 81.170 348.430 81.880 ;
        RECT 344.840 81.160 345.140 81.170 ;
        RECT 22.620 79.710 23.030 79.720 ;
        RECT 22.620 79.010 26.270 79.710 ;
        RECT 259.150 79.650 259.560 79.660 ;
        RECT 22.760 79.000 26.270 79.010 ;
        RECT 123.930 79.520 124.340 79.530 ;
        RECT 123.930 78.820 127.580 79.520 ;
        RECT 259.150 78.950 262.800 79.650 ;
        RECT 259.290 78.940 262.800 78.950 ;
        RECT 360.460 79.460 360.870 79.470 ;
        RECT 124.070 78.810 127.580 78.820 ;
        RECT 360.460 78.760 364.110 79.460 ;
        RECT 360.600 78.750 364.110 78.760 ;
        RECT 72.000 76.340 72.560 76.360 ;
        RECT 7.180 75.730 7.480 75.740 ;
        RECT 7.180 75.020 10.750 75.730 ;
        RECT 72.000 75.640 75.780 76.340 ;
        RECT 308.530 76.280 309.090 76.300 ;
        RECT 72.480 75.630 75.780 75.640 ;
        RECT 173.310 76.150 173.870 76.170 ;
        RECT 108.490 75.540 108.790 75.550 ;
        RECT 108.490 74.830 112.060 75.540 ;
        RECT 173.310 75.450 177.090 76.150 ;
        RECT 173.790 75.440 177.090 75.450 ;
        RECT 243.710 75.670 244.010 75.680 ;
        RECT 243.710 74.960 247.280 75.670 ;
        RECT 308.530 75.580 312.310 76.280 ;
        RECT 309.010 75.570 312.310 75.580 ;
        RECT 409.840 76.090 410.400 76.110 ;
        RECT 345.020 75.480 345.320 75.490 ;
        RECT 345.020 74.770 348.590 75.480 ;
        RECT 409.840 75.390 413.620 76.090 ;
        RECT 410.320 75.380 413.620 75.390 ;
        RECT 6.850 65.990 10.440 66.700 ;
        RECT 6.850 65.980 7.150 65.990 ;
        RECT 108.160 65.800 111.750 66.510 ;
        RECT 243.380 65.930 246.970 66.640 ;
        RECT 243.380 65.920 243.680 65.930 ;
        RECT 108.160 65.790 108.460 65.800 ;
        RECT 344.690 65.740 348.280 66.450 ;
        RECT 344.690 65.730 344.990 65.740 ;
        RECT 22.470 64.280 22.880 64.290 ;
        RECT 22.470 63.580 26.120 64.280 ;
        RECT 259.000 64.220 259.410 64.230 ;
        RECT 22.610 63.570 26.120 63.580 ;
        RECT 123.780 64.090 124.190 64.100 ;
        RECT 123.780 63.390 127.430 64.090 ;
        RECT 259.000 63.520 262.650 64.220 ;
        RECT 259.140 63.510 262.650 63.520 ;
        RECT 360.310 64.030 360.720 64.040 ;
        RECT 123.920 63.380 127.430 63.390 ;
        RECT 360.310 63.330 363.960 64.030 ;
        RECT 360.450 63.320 363.960 63.330 ;
        RECT 7.030 60.300 7.330 60.310 ;
        RECT 7.030 59.590 10.600 60.300 ;
        RECT 243.560 60.240 243.860 60.250 ;
        RECT 108.340 60.110 108.640 60.120 ;
        RECT 108.340 59.400 111.910 60.110 ;
        RECT 243.560 59.530 247.130 60.240 ;
        RECT 344.870 60.050 345.170 60.060 ;
        RECT 344.870 59.340 348.440 60.050 ;
        RECT 40.060 58.730 40.440 58.740 ;
        RECT 40.060 58.020 43.700 58.730 ;
        RECT 276.590 58.670 276.970 58.680 ;
        RECT 141.370 58.540 141.750 58.550 ;
        RECT 141.370 57.830 145.010 58.540 ;
        RECT 276.590 57.960 280.230 58.670 ;
        RECT 377.900 58.480 378.280 58.490 ;
        RECT 377.900 57.770 381.540 58.480 ;
        RECT 6.680 51.570 10.270 52.280 ;
        RECT 6.680 51.560 6.980 51.570 ;
        RECT 107.990 51.380 111.580 52.090 ;
        RECT 243.210 51.510 246.800 52.220 ;
        RECT 243.210 51.500 243.510 51.510 ;
        RECT 107.990 51.370 108.290 51.380 ;
        RECT 344.520 51.320 348.110 52.030 ;
        RECT 344.520 51.310 344.820 51.320 ;
        RECT 22.300 49.860 22.710 49.870 ;
        RECT 22.300 49.160 25.950 49.860 ;
        RECT 258.830 49.800 259.240 49.810 ;
        RECT 22.440 49.150 25.950 49.160 ;
        RECT 123.610 49.670 124.020 49.680 ;
        RECT 123.610 48.970 127.260 49.670 ;
        RECT 258.830 49.100 262.480 49.800 ;
        RECT 258.970 49.090 262.480 49.100 ;
        RECT 360.140 49.610 360.550 49.620 ;
        RECT 123.750 48.960 127.260 48.970 ;
        RECT 360.140 48.910 363.790 49.610 ;
        RECT 360.280 48.900 363.790 48.910 ;
        RECT 6.860 45.880 7.160 45.890 ;
        RECT 6.860 45.170 10.430 45.880 ;
        RECT 243.390 45.820 243.690 45.830 ;
        RECT 108.170 45.690 108.470 45.700 ;
        RECT 108.170 44.980 111.740 45.690 ;
        RECT 243.390 45.110 246.960 45.820 ;
        RECT 344.700 45.630 345.000 45.640 ;
        RECT 344.700 44.920 348.270 45.630 ;
        RECT 57.930 42.700 61.230 42.710 ;
        RECT 57.460 42.000 61.230 42.700 ;
        RECT 294.460 42.640 297.760 42.650 ;
        RECT 159.240 42.510 162.540 42.520 ;
        RECT 57.460 41.970 58.040 42.000 ;
        RECT 158.770 41.810 162.540 42.510 ;
        RECT 293.990 41.940 297.760 42.640 ;
        RECT 395.770 42.450 399.070 42.460 ;
        RECT 293.990 41.910 294.570 41.940 ;
        RECT 158.770 41.780 159.350 41.810 ;
        RECT 395.300 41.750 399.070 42.450 ;
        RECT 395.300 41.720 395.880 41.750 ;
        RECT 6.820 35.920 10.410 36.630 ;
        RECT 6.820 35.910 7.120 35.920 ;
        RECT 108.130 35.730 111.720 36.440 ;
        RECT 243.350 35.860 246.940 36.570 ;
        RECT 243.350 35.850 243.650 35.860 ;
        RECT 108.130 35.720 108.430 35.730 ;
        RECT 344.660 35.670 348.250 36.380 ;
        RECT 344.660 35.660 344.960 35.670 ;
        RECT 22.440 34.210 22.850 34.220 ;
        RECT 22.440 33.510 26.090 34.210 ;
        RECT 258.970 34.150 259.380 34.160 ;
        RECT 22.580 33.500 26.090 33.510 ;
        RECT 123.750 34.020 124.160 34.030 ;
        RECT 123.750 33.320 127.400 34.020 ;
        RECT 258.970 33.450 262.620 34.150 ;
        RECT 259.110 33.440 262.620 33.450 ;
        RECT 360.280 33.960 360.690 33.970 ;
        RECT 123.890 33.310 127.400 33.320 ;
        RECT 360.280 33.260 363.930 33.960 ;
        RECT 360.420 33.250 363.930 33.260 ;
        RECT 7.000 30.230 7.300 30.240 ;
        RECT 7.000 29.520 10.570 30.230 ;
        RECT 243.530 30.170 243.830 30.180 ;
        RECT 108.310 30.040 108.610 30.050 ;
        RECT 108.310 29.330 111.880 30.040 ;
        RECT 243.530 29.460 247.100 30.170 ;
        RECT 344.840 29.980 345.140 29.990 ;
        RECT 344.840 29.270 348.410 29.980 ;
        RECT 40.030 28.660 40.410 28.670 ;
        RECT 40.030 27.950 43.670 28.660 ;
        RECT 276.560 28.600 276.940 28.610 ;
        RECT 141.340 28.470 141.720 28.480 ;
        RECT 141.340 27.760 144.980 28.470 ;
        RECT 276.560 27.890 280.200 28.600 ;
        RECT 377.870 28.410 378.250 28.420 ;
        RECT 377.870 27.700 381.510 28.410 ;
        RECT 6.650 21.500 10.240 22.210 ;
        RECT 6.650 21.490 6.950 21.500 ;
        RECT 107.960 21.310 111.550 22.020 ;
        RECT 243.180 21.440 246.770 22.150 ;
        RECT 243.180 21.430 243.480 21.440 ;
        RECT 107.960 21.300 108.260 21.310 ;
        RECT 344.490 21.250 348.080 21.960 ;
        RECT 344.490 21.240 344.790 21.250 ;
        RECT 22.270 19.790 22.680 19.800 ;
        RECT 22.270 19.090 25.920 19.790 ;
        RECT 258.800 19.730 259.210 19.740 ;
        RECT 22.410 19.080 25.920 19.090 ;
        RECT 123.580 19.600 123.990 19.610 ;
        RECT 123.580 18.900 127.230 19.600 ;
        RECT 258.800 19.030 262.450 19.730 ;
        RECT 258.940 19.020 262.450 19.030 ;
        RECT 360.110 19.540 360.520 19.550 ;
        RECT 123.720 18.890 127.230 18.900 ;
        RECT 360.110 18.840 363.760 19.540 ;
        RECT 360.250 18.830 363.760 18.840 ;
        RECT 6.830 15.810 7.130 15.820 ;
        RECT 6.830 15.100 10.400 15.810 ;
        RECT 243.360 15.750 243.660 15.760 ;
        RECT 108.140 15.620 108.440 15.630 ;
        RECT 108.140 14.910 111.710 15.620 ;
        RECT 243.360 15.040 246.930 15.750 ;
        RECT 344.670 15.560 344.970 15.570 ;
        RECT 344.670 14.850 348.240 15.560 ;
      LAYER via ;
        RECT 7.715 246.365 7.975 246.625 ;
        RECT 109.025 246.175 109.285 246.435 ;
        RECT 244.245 246.305 244.505 246.565 ;
        RECT 345.555 246.115 345.815 246.375 ;
        RECT 23.365 243.865 23.625 244.125 ;
        RECT 124.675 243.675 124.935 243.935 ;
        RECT 259.895 243.805 260.155 244.065 ;
        RECT 361.205 243.615 361.465 243.875 ;
        RECT 7.885 239.955 8.145 240.215 ;
        RECT 109.195 239.765 109.455 240.025 ;
        RECT 244.415 239.895 244.675 240.155 ;
        RECT 345.725 239.705 345.985 239.965 ;
        RECT 40.980 238.360 41.240 238.620 ;
        RECT 142.290 238.170 142.550 238.430 ;
        RECT 277.510 238.300 277.770 238.560 ;
        RECT 378.820 238.110 379.080 238.370 ;
        RECT 7.545 231.945 7.805 232.205 ;
        RECT 108.855 231.755 109.115 232.015 ;
        RECT 244.075 231.885 244.335 232.145 ;
        RECT 345.385 231.695 345.645 231.955 ;
        RECT 23.195 229.445 23.455 229.705 ;
        RECT 124.505 229.255 124.765 229.515 ;
        RECT 259.725 229.385 259.985 229.645 ;
        RECT 361.035 229.195 361.295 229.455 ;
        RECT 7.715 225.535 7.975 225.795 ;
        RECT 109.025 225.345 109.285 225.605 ;
        RECT 244.245 225.475 244.505 225.735 ;
        RECT 345.555 225.285 345.815 225.545 ;
        RECT 58.330 222.220 58.590 222.480 ;
        RECT 159.640 222.030 159.900 222.290 ;
        RECT 294.860 222.160 295.120 222.420 ;
        RECT 396.170 221.970 396.430 222.230 ;
        RECT 7.685 216.295 7.945 216.555 ;
        RECT 108.995 216.105 109.255 216.365 ;
        RECT 244.215 216.235 244.475 216.495 ;
        RECT 345.525 216.045 345.785 216.305 ;
        RECT 23.335 213.795 23.595 214.055 ;
        RECT 124.645 213.605 124.905 213.865 ;
        RECT 259.865 213.735 260.125 213.995 ;
        RECT 361.175 213.545 361.435 213.805 ;
        RECT 7.855 209.885 8.115 210.145 ;
        RECT 109.165 209.695 109.425 209.955 ;
        RECT 244.385 209.825 244.645 210.085 ;
        RECT 345.695 209.635 345.955 209.895 ;
        RECT 40.950 208.290 41.210 208.550 ;
        RECT 142.260 208.100 142.520 208.360 ;
        RECT 277.480 208.230 277.740 208.490 ;
        RECT 378.790 208.040 379.050 208.300 ;
        RECT 7.515 201.875 7.775 202.135 ;
        RECT 108.825 201.685 109.085 201.945 ;
        RECT 244.045 201.815 244.305 202.075 ;
        RECT 345.355 201.625 345.615 201.885 ;
        RECT 23.165 199.375 23.425 199.635 ;
        RECT 124.475 199.185 124.735 199.445 ;
        RECT 259.695 199.315 259.955 199.575 ;
        RECT 361.005 199.125 361.265 199.385 ;
        RECT 72.580 196.010 72.840 196.270 ;
        RECT 173.890 195.820 174.150 196.080 ;
        RECT 309.110 195.950 309.370 196.210 ;
        RECT 7.685 195.465 7.945 195.725 ;
        RECT 108.995 195.275 109.255 195.535 ;
        RECT 410.420 195.760 410.680 196.020 ;
        RECT 244.215 195.405 244.475 195.665 ;
        RECT 345.525 195.215 345.785 195.475 ;
        RECT 7.365 186.445 7.625 186.705 ;
        RECT 108.675 186.255 108.935 186.515 ;
        RECT 243.895 186.385 244.155 186.645 ;
        RECT 345.205 186.195 345.465 186.455 ;
        RECT 23.015 183.945 23.275 184.205 ;
        RECT 124.325 183.755 124.585 184.015 ;
        RECT 259.545 183.885 259.805 184.145 ;
        RECT 360.855 183.695 361.115 183.955 ;
        RECT 7.535 180.035 7.795 180.295 ;
        RECT 108.845 179.845 109.105 180.105 ;
        RECT 244.065 179.975 244.325 180.235 ;
        RECT 345.375 179.785 345.635 180.045 ;
        RECT 40.630 178.440 40.890 178.700 ;
        RECT 141.940 178.250 142.200 178.510 ;
        RECT 277.160 178.380 277.420 178.640 ;
        RECT 378.470 178.190 378.730 178.450 ;
        RECT 7.195 172.025 7.455 172.285 ;
        RECT 108.505 171.835 108.765 172.095 ;
        RECT 243.725 171.965 243.985 172.225 ;
        RECT 345.035 171.775 345.295 172.035 ;
        RECT 22.845 169.525 23.105 169.785 ;
        RECT 124.155 169.335 124.415 169.595 ;
        RECT 259.375 169.465 259.635 169.725 ;
        RECT 360.685 169.275 360.945 169.535 ;
        RECT 7.365 165.615 7.625 165.875 ;
        RECT 108.675 165.425 108.935 165.685 ;
        RECT 243.895 165.555 244.155 165.815 ;
        RECT 345.205 165.365 345.465 165.625 ;
        RECT 57.980 162.300 58.240 162.560 ;
        RECT 159.290 162.110 159.550 162.370 ;
        RECT 294.510 162.240 294.770 162.500 ;
        RECT 395.820 162.050 396.080 162.310 ;
        RECT 7.335 156.375 7.595 156.635 ;
        RECT 108.645 156.185 108.905 156.445 ;
        RECT 243.865 156.315 244.125 156.575 ;
        RECT 345.175 156.125 345.435 156.385 ;
        RECT 22.985 153.875 23.245 154.135 ;
        RECT 124.295 153.685 124.555 153.945 ;
        RECT 259.515 153.815 259.775 154.075 ;
        RECT 360.825 153.625 361.085 153.885 ;
        RECT 7.505 149.965 7.765 150.225 ;
        RECT 108.815 149.775 109.075 150.035 ;
        RECT 244.035 149.905 244.295 150.165 ;
        RECT 345.345 149.715 345.605 149.975 ;
        RECT 40.600 148.370 40.860 148.630 ;
        RECT 141.910 148.180 142.170 148.440 ;
        RECT 277.130 148.310 277.390 148.570 ;
        RECT 378.440 148.120 378.700 148.380 ;
        RECT 7.165 141.955 7.425 142.215 ;
        RECT 108.475 141.765 108.735 142.025 ;
        RECT 243.695 141.895 243.955 142.155 ;
        RECT 345.005 141.705 345.265 141.965 ;
        RECT 22.815 139.455 23.075 139.715 ;
        RECT 124.125 139.265 124.385 139.525 ;
        RECT 259.345 139.395 259.605 139.655 ;
        RECT 360.655 139.205 360.915 139.465 ;
        RECT 7.335 135.545 7.595 135.805 ;
        RECT 108.645 135.355 108.905 135.615 ;
        RECT 216.575 135.060 216.835 135.320 ;
        RECT 243.865 135.485 244.125 135.745 ;
        RECT 345.175 135.295 345.435 135.555 ;
        RECT 453.105 135.000 453.365 135.260 ;
        RECT 88.885 132.875 89.145 133.135 ;
        RECT 190.195 132.685 190.455 132.945 ;
        RECT 325.415 132.815 325.675 133.075 ;
        RECT 426.725 132.625 426.985 132.885 ;
        RECT 470.365 132.630 470.625 132.890 ;
        RECT 7.215 126.125 7.475 126.385 ;
        RECT 108.525 125.935 108.785 126.195 ;
        RECT 243.745 126.065 244.005 126.325 ;
        RECT 345.055 125.875 345.315 126.135 ;
        RECT 22.865 123.625 23.125 123.885 ;
        RECT 124.175 123.435 124.435 123.695 ;
        RECT 259.395 123.565 259.655 123.825 ;
        RECT 360.705 123.375 360.965 123.635 ;
        RECT 7.385 119.715 7.645 119.975 ;
        RECT 108.695 119.525 108.955 119.785 ;
        RECT 243.915 119.655 244.175 119.915 ;
        RECT 345.225 119.465 345.485 119.725 ;
        RECT 40.480 118.120 40.740 118.380 ;
        RECT 141.790 117.930 142.050 118.190 ;
        RECT 277.010 118.060 277.270 118.320 ;
        RECT 378.320 117.870 378.580 118.130 ;
        RECT 7.045 111.705 7.305 111.965 ;
        RECT 108.355 111.515 108.615 111.775 ;
        RECT 243.575 111.645 243.835 111.905 ;
        RECT 344.885 111.455 345.145 111.715 ;
        RECT 22.695 109.205 22.955 109.465 ;
        RECT 124.005 109.015 124.265 109.275 ;
        RECT 259.225 109.145 259.485 109.405 ;
        RECT 360.535 108.955 360.795 109.215 ;
        RECT 7.215 105.295 7.475 105.555 ;
        RECT 108.525 105.105 108.785 105.365 ;
        RECT 243.745 105.235 244.005 105.495 ;
        RECT 345.055 105.045 345.315 105.305 ;
        RECT 57.830 101.980 58.090 102.240 ;
        RECT 159.140 101.790 159.400 102.050 ;
        RECT 294.360 101.920 294.620 102.180 ;
        RECT 395.670 101.730 395.930 101.990 ;
        RECT 7.185 96.055 7.445 96.315 ;
        RECT 108.495 95.865 108.755 96.125 ;
        RECT 243.715 95.995 243.975 96.255 ;
        RECT 345.025 95.805 345.285 96.065 ;
        RECT 22.835 93.555 23.095 93.815 ;
        RECT 124.145 93.365 124.405 93.625 ;
        RECT 259.365 93.495 259.625 93.755 ;
        RECT 360.675 93.305 360.935 93.565 ;
        RECT 7.355 89.645 7.615 89.905 ;
        RECT 108.665 89.455 108.925 89.715 ;
        RECT 243.885 89.585 244.145 89.845 ;
        RECT 345.195 89.395 345.455 89.655 ;
        RECT 40.450 88.050 40.710 88.310 ;
        RECT 141.760 87.860 142.020 88.120 ;
        RECT 276.980 87.990 277.240 88.250 ;
        RECT 378.290 87.800 378.550 88.060 ;
        RECT 7.015 81.635 7.275 81.895 ;
        RECT 108.325 81.445 108.585 81.705 ;
        RECT 243.545 81.575 243.805 81.835 ;
        RECT 344.855 81.385 345.115 81.645 ;
        RECT 22.665 79.135 22.925 79.395 ;
        RECT 123.975 78.945 124.235 79.205 ;
        RECT 259.195 79.075 259.455 79.335 ;
        RECT 360.505 78.885 360.765 79.145 ;
        RECT 72.080 75.770 72.340 76.030 ;
        RECT 173.390 75.580 173.650 75.840 ;
        RECT 308.610 75.710 308.870 75.970 ;
        RECT 7.185 75.225 7.445 75.485 ;
        RECT 108.495 75.035 108.755 75.295 ;
        RECT 409.920 75.520 410.180 75.780 ;
        RECT 243.715 75.165 243.975 75.425 ;
        RECT 345.025 74.975 345.285 75.235 ;
        RECT 6.865 66.205 7.125 66.465 ;
        RECT 108.175 66.015 108.435 66.275 ;
        RECT 243.395 66.145 243.655 66.405 ;
        RECT 344.705 65.955 344.965 66.215 ;
        RECT 22.515 63.705 22.775 63.965 ;
        RECT 123.825 63.515 124.085 63.775 ;
        RECT 259.045 63.645 259.305 63.905 ;
        RECT 360.355 63.455 360.615 63.715 ;
        RECT 7.035 59.795 7.295 60.055 ;
        RECT 108.345 59.605 108.605 59.865 ;
        RECT 243.565 59.735 243.825 59.995 ;
        RECT 344.875 59.545 345.135 59.805 ;
        RECT 40.130 58.200 40.390 58.460 ;
        RECT 141.440 58.010 141.700 58.270 ;
        RECT 276.660 58.140 276.920 58.400 ;
        RECT 377.970 57.950 378.230 58.210 ;
        RECT 6.695 51.785 6.955 52.045 ;
        RECT 108.005 51.595 108.265 51.855 ;
        RECT 243.225 51.725 243.485 51.985 ;
        RECT 344.535 51.535 344.795 51.795 ;
        RECT 22.345 49.285 22.605 49.545 ;
        RECT 123.655 49.095 123.915 49.355 ;
        RECT 258.875 49.225 259.135 49.485 ;
        RECT 360.185 49.035 360.445 49.295 ;
        RECT 6.865 45.375 7.125 45.635 ;
        RECT 108.175 45.185 108.435 45.445 ;
        RECT 243.395 45.315 243.655 45.575 ;
        RECT 344.705 45.125 344.965 45.385 ;
        RECT 57.480 42.060 57.740 42.320 ;
        RECT 158.790 41.870 159.050 42.130 ;
        RECT 294.010 42.000 294.270 42.260 ;
        RECT 395.320 41.810 395.580 42.070 ;
        RECT 6.835 36.135 7.095 36.395 ;
        RECT 108.145 35.945 108.405 36.205 ;
        RECT 243.365 36.075 243.625 36.335 ;
        RECT 344.675 35.885 344.935 36.145 ;
        RECT 22.485 33.635 22.745 33.895 ;
        RECT 123.795 33.445 124.055 33.705 ;
        RECT 259.015 33.575 259.275 33.835 ;
        RECT 360.325 33.385 360.585 33.645 ;
        RECT 7.005 29.725 7.265 29.985 ;
        RECT 108.315 29.535 108.575 29.795 ;
        RECT 243.535 29.665 243.795 29.925 ;
        RECT 344.845 29.475 345.105 29.735 ;
        RECT 40.100 28.130 40.360 28.390 ;
        RECT 141.410 27.940 141.670 28.200 ;
        RECT 276.630 28.070 276.890 28.330 ;
        RECT 377.940 27.880 378.200 28.140 ;
        RECT 6.665 21.715 6.925 21.975 ;
        RECT 107.975 21.525 108.235 21.785 ;
        RECT 243.195 21.655 243.455 21.915 ;
        RECT 344.505 21.465 344.765 21.725 ;
        RECT 22.315 19.215 22.575 19.475 ;
        RECT 123.625 19.025 123.885 19.285 ;
        RECT 258.845 19.155 259.105 19.415 ;
        RECT 360.155 18.965 360.415 19.225 ;
        RECT 6.835 15.305 7.095 15.565 ;
        RECT 108.145 15.115 108.405 15.375 ;
        RECT 243.365 15.245 243.625 15.505 ;
        RECT 344.675 15.055 344.935 15.315 ;
      LAYER met2 ;
        RECT 96.950 254.600 121.780 254.630 ;
        RECT 83.010 254.580 125.760 254.600 ;
        RECT 55.100 254.550 125.760 254.580 ;
        RECT 55.100 254.530 291.410 254.550 ;
        RECT 333.480 254.540 358.310 254.570 ;
        RECT 55.100 254.520 292.000 254.530 ;
        RECT 319.540 254.520 358.310 254.540 ;
        RECT 55.100 254.270 358.310 254.520 ;
        RECT 55.100 254.250 291.410 254.270 ;
        RECT 55.100 254.200 121.780 254.250 ;
        RECT 125.600 254.240 291.410 254.250 ;
        RECT 55.100 254.170 97.190 254.200 ;
        RECT 55.100 254.150 83.240 254.170 ;
        RECT 7.530 246.280 8.010 246.680 ;
        RECT 7.530 240.310 7.720 246.280 ;
        RECT 23.170 244.180 23.380 244.190 ;
        RECT 22.720 244.140 23.640 244.180 ;
        RECT 22.670 244.100 23.640 244.140 ;
        RECT 22.670 243.830 23.650 244.100 ;
        RECT 22.670 243.800 23.640 243.830 ;
        RECT 22.670 241.570 22.910 243.800 ;
        RECT 23.170 243.790 23.380 243.800 ;
        RECT 22.670 240.420 22.920 241.570 ;
        RECT 7.530 240.280 7.780 240.310 ;
        RECT 7.530 239.880 8.180 240.280 ;
        RECT 7.540 238.740 7.780 239.880 ;
        RECT 20.400 238.740 20.650 238.790 ;
        RECT 22.680 238.740 22.920 240.420 ;
        RECT 7.540 238.570 22.920 238.740 ;
        RECT 40.260 238.710 41.310 238.730 ;
        RECT 7.540 238.500 22.650 238.570 ;
        RECT 20.400 232.410 20.650 238.500 ;
        RECT 40.250 238.210 41.310 238.710 ;
        RECT 40.250 237.460 40.570 238.210 ;
        RECT 40.250 235.890 40.560 237.460 ;
        RECT 7.360 231.860 7.840 232.260 ;
        RECT 7.360 225.890 7.550 231.860 ;
        RECT 7.360 225.860 7.610 225.890 ;
        RECT 7.360 225.460 8.010 225.860 ;
        RECT 7.370 224.320 7.610 225.460 ;
        RECT 20.370 224.320 20.670 232.410 ;
        RECT 23.000 229.760 23.210 229.770 ;
        RECT 22.550 229.720 23.470 229.760 ;
        RECT 22.500 229.680 23.470 229.720 ;
        RECT 22.500 229.410 23.480 229.680 ;
        RECT 22.500 229.380 23.470 229.410 ;
        RECT 22.500 227.150 22.740 229.380 ;
        RECT 23.000 229.370 23.210 229.380 ;
        RECT 22.500 226.000 22.750 227.150 ;
        RECT 22.510 224.550 22.750 226.000 ;
        RECT 40.220 224.990 40.580 235.890 ;
        RECT 55.100 230.270 55.420 254.150 ;
        RECT 121.560 254.090 121.780 254.200 ;
        RECT 291.630 254.140 358.310 254.270 ;
        RECT 291.630 254.110 333.720 254.140 ;
        RECT 291.630 254.090 319.770 254.110 ;
        RECT 121.560 251.090 121.840 254.090 ;
        RECT 108.840 246.090 109.320 246.490 ;
        RECT 108.840 240.120 109.030 246.090 ;
        RECT 121.560 244.820 121.890 251.090 ;
        RECT 244.060 246.220 244.540 246.620 ;
        RECT 121.560 244.630 121.920 244.820 ;
        RECT 108.840 240.090 109.090 240.120 ;
        RECT 108.840 239.690 109.490 240.090 ;
        RECT 108.850 238.550 109.090 239.690 ;
        RECT 121.590 238.600 121.920 244.630 ;
        RECT 124.480 243.990 124.690 244.000 ;
        RECT 124.030 243.950 124.950 243.990 ;
        RECT 123.980 243.910 124.950 243.950 ;
        RECT 123.980 243.640 124.960 243.910 ;
        RECT 123.980 243.610 124.950 243.640 ;
        RECT 123.980 241.380 124.220 243.610 ;
        RECT 124.480 243.600 124.690 243.610 ;
        RECT 123.980 240.230 124.230 241.380 ;
        RECT 121.590 238.550 121.960 238.600 ;
        RECT 123.990 238.550 124.230 240.230 ;
        RECT 244.060 240.250 244.250 246.220 ;
        RECT 259.700 244.120 259.910 244.130 ;
        RECT 259.250 244.080 260.170 244.120 ;
        RECT 259.200 244.040 260.170 244.080 ;
        RECT 259.200 243.770 260.180 244.040 ;
        RECT 259.200 243.740 260.170 243.770 ;
        RECT 259.200 241.510 259.440 243.740 ;
        RECT 259.700 243.730 259.910 243.740 ;
        RECT 259.200 240.360 259.450 241.510 ;
        RECT 244.060 240.220 244.310 240.250 ;
        RECT 244.060 239.820 244.710 240.220 ;
        RECT 108.850 238.380 124.230 238.550 ;
        RECT 244.070 238.680 244.310 239.820 ;
        RECT 256.930 238.680 257.180 238.730 ;
        RECT 259.210 238.680 259.450 240.360 ;
        RECT 141.570 238.520 142.620 238.540 ;
        RECT 108.850 238.310 123.960 238.380 ;
        RECT 121.710 232.220 121.960 238.310 ;
        RECT 141.560 238.020 142.620 238.520 ;
        RECT 244.070 238.510 259.450 238.680 ;
        RECT 276.790 238.650 277.840 238.670 ;
        RECT 244.070 238.440 259.180 238.510 ;
        RECT 141.560 237.270 141.880 238.020 ;
        RECT 141.560 235.700 141.870 237.270 ;
        RECT 108.670 231.670 109.150 232.070 ;
        RECT 55.100 229.870 55.530 230.270 ;
        RECT 28.460 224.620 37.230 224.630 ;
        RECT 40.220 224.620 40.550 224.990 ;
        RECT 28.460 224.570 40.550 224.620 ;
        RECT 27.600 224.560 40.550 224.570 ;
        RECT 24.580 224.550 40.550 224.560 ;
        RECT 22.510 224.340 40.550 224.550 ;
        RECT 22.510 224.330 28.670 224.340 ;
        RECT 22.510 224.320 27.680 224.330 ;
        RECT 7.370 224.310 24.610 224.320 ;
        RECT 7.370 224.150 22.750 224.310 ;
        RECT 7.370 224.080 22.480 224.150 ;
        RECT 20.370 224.030 20.670 224.080 ;
        RECT 35.510 222.440 35.700 224.340 ;
        RECT 36.930 224.330 40.550 224.340 ;
        RECT 55.150 222.520 55.530 229.870 ;
        RECT 108.670 225.700 108.860 231.670 ;
        RECT 108.670 225.670 108.920 225.700 ;
        RECT 108.670 225.270 109.320 225.670 ;
        RECT 108.680 224.130 108.920 225.270 ;
        RECT 121.680 224.130 121.980 232.220 ;
        RECT 124.310 229.570 124.520 229.580 ;
        RECT 123.860 229.530 124.780 229.570 ;
        RECT 123.810 229.490 124.780 229.530 ;
        RECT 123.810 229.220 124.790 229.490 ;
        RECT 123.810 229.190 124.780 229.220 ;
        RECT 123.810 226.960 124.050 229.190 ;
        RECT 124.310 229.180 124.520 229.190 ;
        RECT 123.810 225.810 124.060 226.960 ;
        RECT 123.820 224.360 124.060 225.810 ;
        RECT 141.530 224.800 141.890 235.700 ;
        RECT 256.930 232.350 257.180 238.440 ;
        RECT 276.780 238.150 277.840 238.650 ;
        RECT 276.780 237.400 277.100 238.150 ;
        RECT 276.780 235.830 277.090 237.400 ;
        RECT 243.890 231.800 244.370 232.200 ;
        RECT 243.890 225.830 244.080 231.800 ;
        RECT 243.890 225.800 244.140 225.830 ;
        RECT 243.890 225.400 244.540 225.800 ;
        RECT 129.770 224.430 138.540 224.440 ;
        RECT 141.530 224.430 141.860 224.800 ;
        RECT 129.770 224.380 141.860 224.430 ;
        RECT 128.910 224.370 141.860 224.380 ;
        RECT 125.890 224.360 141.860 224.370 ;
        RECT 123.820 224.150 141.860 224.360 ;
        RECT 123.820 224.140 129.980 224.150 ;
        RECT 123.820 224.130 128.990 224.140 ;
        RECT 108.680 224.120 125.920 224.130 ;
        RECT 108.680 223.960 124.060 224.120 ;
        RECT 108.680 223.890 123.790 223.960 ;
        RECT 121.680 223.840 121.980 223.890 ;
        RECT 55.120 222.440 55.570 222.520 ;
        RECT 58.300 222.440 58.670 222.560 ;
        RECT 35.510 222.200 58.670 222.440 ;
        RECT 136.820 222.250 137.010 224.150 ;
        RECT 138.240 224.140 141.860 224.150 ;
        RECT 243.900 224.260 244.140 225.400 ;
        RECT 256.900 224.260 257.200 232.350 ;
        RECT 259.530 229.700 259.740 229.710 ;
        RECT 259.080 229.660 260.000 229.700 ;
        RECT 259.030 229.620 260.000 229.660 ;
        RECT 259.030 229.350 260.010 229.620 ;
        RECT 259.030 229.320 260.000 229.350 ;
        RECT 259.030 227.090 259.270 229.320 ;
        RECT 259.530 229.310 259.740 229.320 ;
        RECT 259.030 225.940 259.280 227.090 ;
        RECT 259.040 224.490 259.280 225.940 ;
        RECT 276.750 224.930 277.110 235.830 ;
        RECT 291.630 230.210 291.950 254.090 ;
        RECT 358.090 254.030 358.310 254.140 ;
        RECT 358.090 251.030 358.370 254.030 ;
        RECT 345.370 246.030 345.850 246.430 ;
        RECT 345.370 240.060 345.560 246.030 ;
        RECT 358.090 244.760 358.420 251.030 ;
        RECT 358.090 244.570 358.450 244.760 ;
        RECT 345.370 240.030 345.620 240.060 ;
        RECT 345.370 239.630 346.020 240.030 ;
        RECT 345.380 238.490 345.620 239.630 ;
        RECT 358.120 238.540 358.450 244.570 ;
        RECT 361.010 243.930 361.220 243.940 ;
        RECT 360.560 243.890 361.480 243.930 ;
        RECT 360.510 243.850 361.480 243.890 ;
        RECT 360.510 243.580 361.490 243.850 ;
        RECT 360.510 243.550 361.480 243.580 ;
        RECT 360.510 241.320 360.750 243.550 ;
        RECT 361.010 243.540 361.220 243.550 ;
        RECT 360.510 240.170 360.760 241.320 ;
        RECT 358.120 238.490 358.490 238.540 ;
        RECT 360.520 238.490 360.760 240.170 ;
        RECT 345.380 238.320 360.760 238.490 ;
        RECT 378.100 238.460 379.150 238.480 ;
        RECT 345.380 238.250 360.490 238.320 ;
        RECT 358.240 232.160 358.490 238.250 ;
        RECT 378.090 237.960 379.150 238.460 ;
        RECT 378.090 237.210 378.410 237.960 ;
        RECT 378.090 235.640 378.400 237.210 ;
        RECT 345.200 231.610 345.680 232.010 ;
        RECT 291.630 229.810 292.060 230.210 ;
        RECT 264.990 224.560 273.760 224.570 ;
        RECT 276.750 224.560 277.080 224.930 ;
        RECT 264.990 224.510 277.080 224.560 ;
        RECT 264.130 224.500 277.080 224.510 ;
        RECT 261.110 224.490 277.080 224.500 ;
        RECT 259.040 224.280 277.080 224.490 ;
        RECT 259.040 224.270 265.200 224.280 ;
        RECT 259.040 224.260 264.210 224.270 ;
        RECT 243.900 224.250 261.140 224.260 ;
        RECT 243.900 224.090 259.280 224.250 ;
        RECT 243.900 224.020 259.010 224.090 ;
        RECT 256.900 223.970 257.200 224.020 ;
        RECT 272.040 222.380 272.230 224.280 ;
        RECT 273.460 224.270 277.080 224.280 ;
        RECT 291.680 222.460 292.060 229.810 ;
        RECT 345.200 225.640 345.390 231.610 ;
        RECT 345.200 225.610 345.450 225.640 ;
        RECT 345.200 225.210 345.850 225.610 ;
        RECT 345.210 224.070 345.450 225.210 ;
        RECT 358.210 224.070 358.510 232.160 ;
        RECT 360.840 229.510 361.050 229.520 ;
        RECT 360.390 229.470 361.310 229.510 ;
        RECT 360.340 229.430 361.310 229.470 ;
        RECT 360.340 229.160 361.320 229.430 ;
        RECT 360.340 229.130 361.310 229.160 ;
        RECT 360.340 226.900 360.580 229.130 ;
        RECT 360.840 229.120 361.050 229.130 ;
        RECT 360.340 225.750 360.590 226.900 ;
        RECT 360.350 224.300 360.590 225.750 ;
        RECT 378.060 224.740 378.420 235.640 ;
        RECT 366.300 224.370 375.070 224.380 ;
        RECT 378.060 224.370 378.390 224.740 ;
        RECT 366.300 224.320 378.390 224.370 ;
        RECT 365.440 224.310 378.390 224.320 ;
        RECT 362.420 224.300 378.390 224.310 ;
        RECT 360.350 224.090 378.390 224.300 ;
        RECT 360.350 224.080 366.510 224.090 ;
        RECT 360.350 224.070 365.520 224.080 ;
        RECT 345.210 224.060 362.450 224.070 ;
        RECT 345.210 223.900 360.590 224.060 ;
        RECT 345.210 223.830 360.320 223.900 ;
        RECT 358.210 223.780 358.510 223.830 ;
        RECT 291.650 222.380 292.100 222.460 ;
        RECT 294.830 222.380 295.200 222.500 ;
        RECT 156.430 222.250 156.880 222.330 ;
        RECT 159.610 222.250 159.980 222.370 ;
        RECT 7.500 216.210 7.980 216.610 ;
        RECT 7.500 210.240 7.690 216.210 ;
        RECT 23.140 214.110 23.350 214.120 ;
        RECT 22.690 214.070 23.610 214.110 ;
        RECT 22.640 214.030 23.610 214.070 ;
        RECT 22.640 213.760 23.620 214.030 ;
        RECT 22.640 213.730 23.610 213.760 ;
        RECT 22.640 211.500 22.880 213.730 ;
        RECT 23.140 213.720 23.350 213.730 ;
        RECT 22.640 210.350 22.890 211.500 ;
        RECT 7.500 210.210 7.750 210.240 ;
        RECT 7.500 209.810 8.150 210.210 ;
        RECT 7.510 208.670 7.750 209.810 ;
        RECT 20.370 208.670 20.620 208.720 ;
        RECT 22.650 208.670 22.890 210.350 ;
        RECT 7.510 208.500 22.890 208.670 ;
        RECT 7.510 208.430 22.620 208.500 ;
        RECT 20.370 202.340 20.620 208.430 ;
        RECT 7.330 201.790 7.810 202.190 ;
        RECT 7.330 195.820 7.520 201.790 ;
        RECT 7.330 195.790 7.580 195.820 ;
        RECT 7.330 195.390 7.980 195.790 ;
        RECT 7.340 194.250 7.580 195.390 ;
        RECT 20.340 194.250 20.640 202.340 ;
        RECT 22.970 199.690 23.180 199.700 ;
        RECT 22.520 199.650 23.440 199.690 ;
        RECT 22.470 199.610 23.440 199.650 ;
        RECT 22.470 199.340 23.450 199.610 ;
        RECT 22.470 199.310 23.440 199.340 ;
        RECT 22.470 197.080 22.710 199.310 ;
        RECT 22.970 199.300 23.180 199.310 ;
        RECT 22.470 195.930 22.720 197.080 ;
        RECT 22.480 194.480 22.720 195.930 ;
        RECT 35.510 194.560 35.700 222.200 ;
        RECT 55.120 217.670 55.570 222.200 ;
        RECT 136.820 222.010 159.980 222.250 ;
        RECT 272.040 222.140 295.200 222.380 ;
        RECT 373.350 222.190 373.540 224.090 ;
        RECT 374.770 224.080 378.390 224.090 ;
        RECT 392.960 222.190 393.410 222.270 ;
        RECT 396.140 222.190 396.510 222.310 ;
        RECT 55.120 217.610 69.940 217.670 ;
        RECT 55.120 217.150 70.240 217.610 ;
        RECT 40.230 208.640 41.280 208.660 ;
        RECT 40.220 208.140 41.280 208.640 ;
        RECT 40.220 207.390 40.540 208.140 ;
        RECT 40.220 205.820 40.530 207.390 ;
        RECT 40.190 194.920 40.550 205.820 ;
        RECT 69.790 196.130 70.240 217.150 ;
        RECT 108.810 216.020 109.290 216.420 ;
        RECT 108.810 210.050 109.000 216.020 ;
        RECT 124.450 213.920 124.660 213.930 ;
        RECT 124.000 213.880 124.920 213.920 ;
        RECT 123.950 213.840 124.920 213.880 ;
        RECT 123.950 213.570 124.930 213.840 ;
        RECT 123.950 213.540 124.920 213.570 ;
        RECT 123.950 211.310 124.190 213.540 ;
        RECT 124.450 213.530 124.660 213.540 ;
        RECT 123.950 210.160 124.200 211.310 ;
        RECT 108.810 210.020 109.060 210.050 ;
        RECT 108.810 209.620 109.460 210.020 ;
        RECT 108.820 208.480 109.060 209.620 ;
        RECT 121.680 208.480 121.930 208.530 ;
        RECT 123.960 208.480 124.200 210.160 ;
        RECT 108.820 208.310 124.200 208.480 ;
        RECT 108.820 208.240 123.930 208.310 ;
        RECT 121.680 202.150 121.930 208.240 ;
        RECT 108.640 201.600 109.120 202.000 ;
        RECT 72.510 196.130 72.870 196.440 ;
        RECT 69.770 195.870 72.870 196.130 ;
        RECT 28.430 194.550 37.200 194.560 ;
        RECT 40.190 194.550 40.520 194.920 ;
        RECT 28.430 194.500 40.520 194.550 ;
        RECT 27.570 194.490 40.520 194.500 ;
        RECT 24.550 194.480 40.520 194.490 ;
        RECT 22.480 194.270 40.520 194.480 ;
        RECT 22.480 194.260 28.640 194.270 ;
        RECT 22.480 194.250 27.650 194.260 ;
        RECT 7.340 194.240 24.580 194.250 ;
        RECT 7.340 194.080 22.720 194.240 ;
        RECT 35.510 194.180 35.700 194.270 ;
        RECT 36.900 194.260 40.520 194.270 ;
        RECT 7.340 194.010 22.450 194.080 ;
        RECT 20.340 193.960 20.640 194.010 ;
        RECT 69.790 192.420 70.240 195.870 ;
        RECT 108.640 195.630 108.830 201.600 ;
        RECT 108.640 195.600 108.890 195.630 ;
        RECT 108.640 195.200 109.290 195.600 ;
        RECT 108.650 194.060 108.890 195.200 ;
        RECT 121.650 194.060 121.950 202.150 ;
        RECT 124.280 199.500 124.490 199.510 ;
        RECT 123.830 199.460 124.750 199.500 ;
        RECT 123.780 199.420 124.750 199.460 ;
        RECT 123.780 199.150 124.760 199.420 ;
        RECT 123.780 199.120 124.750 199.150 ;
        RECT 123.780 196.890 124.020 199.120 ;
        RECT 124.280 199.110 124.490 199.120 ;
        RECT 123.780 195.740 124.030 196.890 ;
        RECT 123.790 194.290 124.030 195.740 ;
        RECT 136.820 194.370 137.010 222.010 ;
        RECT 156.430 217.480 156.880 222.010 ;
        RECT 156.430 217.420 171.250 217.480 ;
        RECT 156.430 216.960 171.550 217.420 ;
        RECT 141.540 208.450 142.590 208.470 ;
        RECT 141.530 207.950 142.590 208.450 ;
        RECT 141.530 207.200 141.850 207.950 ;
        RECT 141.530 205.630 141.840 207.200 ;
        RECT 141.500 194.730 141.860 205.630 ;
        RECT 171.100 195.940 171.550 216.960 ;
        RECT 244.030 216.150 244.510 216.550 ;
        RECT 244.030 210.180 244.220 216.150 ;
        RECT 259.670 214.050 259.880 214.060 ;
        RECT 259.220 214.010 260.140 214.050 ;
        RECT 259.170 213.970 260.140 214.010 ;
        RECT 259.170 213.700 260.150 213.970 ;
        RECT 259.170 213.670 260.140 213.700 ;
        RECT 259.170 211.440 259.410 213.670 ;
        RECT 259.670 213.660 259.880 213.670 ;
        RECT 259.170 210.290 259.420 211.440 ;
        RECT 244.030 210.150 244.280 210.180 ;
        RECT 244.030 209.750 244.680 210.150 ;
        RECT 244.040 208.610 244.280 209.750 ;
        RECT 256.900 208.610 257.150 208.660 ;
        RECT 259.180 208.610 259.420 210.290 ;
        RECT 244.040 208.440 259.420 208.610 ;
        RECT 244.040 208.370 259.150 208.440 ;
        RECT 256.900 202.280 257.150 208.370 ;
        RECT 243.860 201.730 244.340 202.130 ;
        RECT 173.820 195.940 174.180 196.250 ;
        RECT 171.080 195.680 174.180 195.940 ;
        RECT 243.860 195.760 244.050 201.730 ;
        RECT 243.860 195.730 244.110 195.760 ;
        RECT 129.740 194.360 138.510 194.370 ;
        RECT 141.500 194.360 141.830 194.730 ;
        RECT 129.740 194.310 141.830 194.360 ;
        RECT 128.880 194.300 141.830 194.310 ;
        RECT 125.860 194.290 141.830 194.300 ;
        RECT 123.790 194.080 141.830 194.290 ;
        RECT 123.790 194.070 129.950 194.080 ;
        RECT 123.790 194.060 128.960 194.070 ;
        RECT 108.650 194.050 125.890 194.060 ;
        RECT 108.650 193.890 124.030 194.050 ;
        RECT 136.820 193.990 137.010 194.080 ;
        RECT 138.210 194.070 141.830 194.080 ;
        RECT 108.650 193.820 123.760 193.890 ;
        RECT 121.650 193.770 121.950 193.820 ;
        RECT 69.760 192.010 70.240 192.420 ;
        RECT 171.100 192.230 171.550 195.680 ;
        RECT 243.860 195.330 244.510 195.730 ;
        RECT 243.870 194.190 244.110 195.330 ;
        RECT 256.870 194.190 257.170 202.280 ;
        RECT 259.500 199.630 259.710 199.640 ;
        RECT 259.050 199.590 259.970 199.630 ;
        RECT 259.000 199.550 259.970 199.590 ;
        RECT 259.000 199.280 259.980 199.550 ;
        RECT 259.000 199.250 259.970 199.280 ;
        RECT 259.000 197.020 259.240 199.250 ;
        RECT 259.500 199.240 259.710 199.250 ;
        RECT 259.000 195.870 259.250 197.020 ;
        RECT 259.010 194.420 259.250 195.870 ;
        RECT 272.040 194.500 272.230 222.140 ;
        RECT 291.650 217.610 292.100 222.140 ;
        RECT 373.350 221.950 396.510 222.190 ;
        RECT 291.650 217.550 306.470 217.610 ;
        RECT 291.650 217.090 306.770 217.550 ;
        RECT 276.760 208.580 277.810 208.600 ;
        RECT 276.750 208.080 277.810 208.580 ;
        RECT 276.750 207.330 277.070 208.080 ;
        RECT 276.750 205.760 277.060 207.330 ;
        RECT 276.720 194.860 277.080 205.760 ;
        RECT 306.320 196.070 306.770 217.090 ;
        RECT 345.340 215.960 345.820 216.360 ;
        RECT 345.340 209.990 345.530 215.960 ;
        RECT 360.980 213.860 361.190 213.870 ;
        RECT 360.530 213.820 361.450 213.860 ;
        RECT 360.480 213.780 361.450 213.820 ;
        RECT 360.480 213.510 361.460 213.780 ;
        RECT 360.480 213.480 361.450 213.510 ;
        RECT 360.480 211.250 360.720 213.480 ;
        RECT 360.980 213.470 361.190 213.480 ;
        RECT 360.480 210.100 360.730 211.250 ;
        RECT 345.340 209.960 345.590 209.990 ;
        RECT 345.340 209.560 345.990 209.960 ;
        RECT 345.350 208.420 345.590 209.560 ;
        RECT 358.210 208.420 358.460 208.470 ;
        RECT 360.490 208.420 360.730 210.100 ;
        RECT 345.350 208.250 360.730 208.420 ;
        RECT 345.350 208.180 360.460 208.250 ;
        RECT 358.210 202.090 358.460 208.180 ;
        RECT 345.170 201.540 345.650 201.940 ;
        RECT 309.040 196.070 309.400 196.380 ;
        RECT 306.300 195.810 309.400 196.070 ;
        RECT 264.960 194.490 273.730 194.500 ;
        RECT 276.720 194.490 277.050 194.860 ;
        RECT 264.960 194.440 277.050 194.490 ;
        RECT 264.100 194.430 277.050 194.440 ;
        RECT 261.080 194.420 277.050 194.430 ;
        RECT 259.010 194.210 277.050 194.420 ;
        RECT 259.010 194.200 265.170 194.210 ;
        RECT 259.010 194.190 264.180 194.200 ;
        RECT 243.870 194.180 261.110 194.190 ;
        RECT 243.870 194.020 259.250 194.180 ;
        RECT 272.040 194.120 272.230 194.210 ;
        RECT 273.430 194.200 277.050 194.210 ;
        RECT 243.870 193.950 258.980 194.020 ;
        RECT 256.870 193.900 257.170 193.950 ;
        RECT 306.320 192.360 306.770 195.810 ;
        RECT 345.170 195.570 345.360 201.540 ;
        RECT 345.170 195.540 345.420 195.570 ;
        RECT 345.170 195.140 345.820 195.540 ;
        RECT 345.180 194.000 345.420 195.140 ;
        RECT 358.180 194.000 358.480 202.090 ;
        RECT 360.810 199.440 361.020 199.450 ;
        RECT 360.360 199.400 361.280 199.440 ;
        RECT 360.310 199.360 361.280 199.400 ;
        RECT 360.310 199.090 361.290 199.360 ;
        RECT 360.310 199.060 361.280 199.090 ;
        RECT 360.310 196.830 360.550 199.060 ;
        RECT 360.810 199.050 361.020 199.060 ;
        RECT 360.310 195.680 360.560 196.830 ;
        RECT 360.320 194.230 360.560 195.680 ;
        RECT 373.350 194.310 373.540 221.950 ;
        RECT 392.960 217.420 393.410 221.950 ;
        RECT 392.960 217.360 407.780 217.420 ;
        RECT 392.960 216.900 408.080 217.360 ;
        RECT 378.070 208.390 379.120 208.410 ;
        RECT 378.060 207.890 379.120 208.390 ;
        RECT 378.060 207.140 378.380 207.890 ;
        RECT 378.060 205.570 378.370 207.140 ;
        RECT 378.030 194.670 378.390 205.570 ;
        RECT 407.630 195.880 408.080 216.900 ;
        RECT 410.350 195.880 410.710 196.190 ;
        RECT 407.610 195.620 410.710 195.880 ;
        RECT 366.270 194.300 375.040 194.310 ;
        RECT 378.030 194.300 378.360 194.670 ;
        RECT 366.270 194.250 378.360 194.300 ;
        RECT 365.410 194.240 378.360 194.250 ;
        RECT 362.390 194.230 378.360 194.240 ;
        RECT 360.320 194.020 378.360 194.230 ;
        RECT 360.320 194.010 366.480 194.020 ;
        RECT 360.320 194.000 365.490 194.010 ;
        RECT 345.180 193.990 362.420 194.000 ;
        RECT 345.180 193.830 360.560 193.990 ;
        RECT 373.350 193.930 373.540 194.020 ;
        RECT 374.740 194.010 378.360 194.020 ;
        RECT 345.180 193.760 360.290 193.830 ;
        RECT 358.180 193.710 358.480 193.760 ;
        RECT 7.180 186.360 7.660 186.760 ;
        RECT 7.180 180.390 7.370 186.360 ;
        RECT 22.820 184.260 23.030 184.270 ;
        RECT 22.370 184.220 23.290 184.260 ;
        RECT 22.320 184.180 23.290 184.220 ;
        RECT 22.320 183.910 23.300 184.180 ;
        RECT 22.320 183.880 23.290 183.910 ;
        RECT 22.320 181.650 22.560 183.880 ;
        RECT 22.820 183.870 23.030 183.880 ;
        RECT 22.320 180.500 22.570 181.650 ;
        RECT 7.180 180.360 7.430 180.390 ;
        RECT 7.180 179.960 7.830 180.360 ;
        RECT 7.190 178.820 7.430 179.960 ;
        RECT 20.050 178.820 20.300 178.870 ;
        RECT 22.330 178.820 22.570 180.500 ;
        RECT 7.190 178.650 22.570 178.820 ;
        RECT 39.910 178.790 40.960 178.810 ;
        RECT 7.190 178.580 22.300 178.650 ;
        RECT 20.050 172.490 20.300 178.580 ;
        RECT 39.900 178.290 40.960 178.790 ;
        RECT 39.900 177.540 40.220 178.290 ;
        RECT 39.900 175.970 40.210 177.540 ;
        RECT 7.010 171.940 7.490 172.340 ;
        RECT 7.010 165.970 7.200 171.940 ;
        RECT 7.010 165.940 7.260 165.970 ;
        RECT 7.010 165.540 7.660 165.940 ;
        RECT 7.020 164.400 7.260 165.540 ;
        RECT 20.020 164.400 20.320 172.490 ;
        RECT 22.650 169.840 22.860 169.850 ;
        RECT 22.200 169.800 23.120 169.840 ;
        RECT 22.150 169.760 23.120 169.800 ;
        RECT 22.150 169.490 23.130 169.760 ;
        RECT 22.150 169.460 23.120 169.490 ;
        RECT 22.150 167.230 22.390 169.460 ;
        RECT 22.650 169.450 22.860 169.460 ;
        RECT 22.150 166.080 22.400 167.230 ;
        RECT 22.160 164.630 22.400 166.080 ;
        RECT 39.870 165.070 40.230 175.970 ;
        RECT 69.760 169.770 70.210 192.010 ;
        RECT 171.070 191.820 171.550 192.230 ;
        RECT 306.290 191.950 306.770 192.360 ;
        RECT 407.630 192.170 408.080 195.620 ;
        RECT 108.490 186.170 108.970 186.570 ;
        RECT 108.490 180.200 108.680 186.170 ;
        RECT 124.130 184.070 124.340 184.080 ;
        RECT 123.680 184.030 124.600 184.070 ;
        RECT 123.630 183.990 124.600 184.030 ;
        RECT 123.630 183.720 124.610 183.990 ;
        RECT 123.630 183.690 124.600 183.720 ;
        RECT 123.630 181.460 123.870 183.690 ;
        RECT 124.130 183.680 124.340 183.690 ;
        RECT 123.630 180.310 123.880 181.460 ;
        RECT 108.490 180.170 108.740 180.200 ;
        RECT 108.490 179.770 109.140 180.170 ;
        RECT 108.500 178.630 108.740 179.770 ;
        RECT 121.360 178.630 121.610 178.680 ;
        RECT 123.640 178.630 123.880 180.310 ;
        RECT 108.500 178.460 123.880 178.630 ;
        RECT 141.220 178.600 142.270 178.620 ;
        RECT 108.500 178.390 123.610 178.460 ;
        RECT 121.360 172.300 121.610 178.390 ;
        RECT 141.210 178.100 142.270 178.600 ;
        RECT 141.210 177.350 141.530 178.100 ;
        RECT 141.210 175.780 141.520 177.350 ;
        RECT 108.320 171.750 108.800 172.150 ;
        RECT 69.760 169.550 70.240 169.770 ;
        RECT 28.110 164.700 36.880 164.710 ;
        RECT 39.870 164.700 40.200 165.070 ;
        RECT 28.110 164.650 40.200 164.700 ;
        RECT 27.250 164.640 40.200 164.650 ;
        RECT 24.230 164.630 40.200 164.640 ;
        RECT 22.160 164.420 40.200 164.630 ;
        RECT 22.160 164.410 28.320 164.420 ;
        RECT 22.160 164.400 27.330 164.410 ;
        RECT 7.020 164.390 24.260 164.400 ;
        RECT 7.020 164.230 22.400 164.390 ;
        RECT 7.020 164.160 22.130 164.230 ;
        RECT 20.020 164.110 20.320 164.160 ;
        RECT 35.160 162.520 35.350 164.420 ;
        RECT 36.580 164.410 40.200 164.420 ;
        RECT 56.610 162.520 57.020 162.530 ;
        RECT 57.950 162.520 58.320 162.640 ;
        RECT 35.160 162.280 58.320 162.520 ;
        RECT 7.150 156.290 7.630 156.690 ;
        RECT 7.150 150.320 7.340 156.290 ;
        RECT 22.790 154.190 23.000 154.200 ;
        RECT 22.340 154.150 23.260 154.190 ;
        RECT 22.290 154.110 23.260 154.150 ;
        RECT 22.290 153.840 23.270 154.110 ;
        RECT 22.290 153.810 23.260 153.840 ;
        RECT 22.290 151.580 22.530 153.810 ;
        RECT 22.790 153.800 23.000 153.810 ;
        RECT 22.290 150.430 22.540 151.580 ;
        RECT 7.150 150.290 7.400 150.320 ;
        RECT 7.150 149.890 7.800 150.290 ;
        RECT 7.160 148.750 7.400 149.890 ;
        RECT 20.020 148.750 20.270 148.800 ;
        RECT 22.300 148.750 22.540 150.430 ;
        RECT 7.160 148.580 22.540 148.750 ;
        RECT 7.160 148.510 22.270 148.580 ;
        RECT 20.020 142.420 20.270 148.510 ;
        RECT 6.980 141.870 7.460 142.270 ;
        RECT 6.980 135.900 7.170 141.870 ;
        RECT 6.980 135.870 7.230 135.900 ;
        RECT 6.980 135.470 7.630 135.870 ;
        RECT 6.990 134.330 7.230 135.470 ;
        RECT 19.990 134.330 20.290 142.420 ;
        RECT 22.620 139.770 22.830 139.780 ;
        RECT 22.170 139.730 23.090 139.770 ;
        RECT 22.120 139.690 23.090 139.730 ;
        RECT 22.120 139.420 23.100 139.690 ;
        RECT 22.120 139.390 23.090 139.420 ;
        RECT 22.120 137.160 22.360 139.390 ;
        RECT 22.620 139.380 22.830 139.390 ;
        RECT 22.120 136.010 22.370 137.160 ;
        RECT 22.130 134.560 22.370 136.010 ;
        RECT 35.160 134.640 35.350 162.280 ;
        RECT 56.610 158.620 57.020 162.280 ;
        RECT 69.790 158.750 70.240 169.550 ;
        RECT 108.320 165.780 108.510 171.750 ;
        RECT 108.320 165.750 108.570 165.780 ;
        RECT 108.320 165.350 108.970 165.750 ;
        RECT 108.330 164.210 108.570 165.350 ;
        RECT 121.330 164.210 121.630 172.300 ;
        RECT 123.960 169.650 124.170 169.660 ;
        RECT 123.510 169.610 124.430 169.650 ;
        RECT 123.460 169.570 124.430 169.610 ;
        RECT 123.460 169.300 124.440 169.570 ;
        RECT 123.460 169.270 124.430 169.300 ;
        RECT 123.460 167.040 123.700 169.270 ;
        RECT 123.960 169.260 124.170 169.270 ;
        RECT 123.460 165.890 123.710 167.040 ;
        RECT 123.470 164.440 123.710 165.890 ;
        RECT 141.180 164.880 141.540 175.780 ;
        RECT 171.070 169.580 171.520 191.820 ;
        RECT 243.710 186.300 244.190 186.700 ;
        RECT 243.710 180.330 243.900 186.300 ;
        RECT 259.350 184.200 259.560 184.210 ;
        RECT 258.900 184.160 259.820 184.200 ;
        RECT 258.850 184.120 259.820 184.160 ;
        RECT 258.850 183.850 259.830 184.120 ;
        RECT 258.850 183.820 259.820 183.850 ;
        RECT 258.850 181.590 259.090 183.820 ;
        RECT 259.350 183.810 259.560 183.820 ;
        RECT 258.850 180.440 259.100 181.590 ;
        RECT 243.710 180.300 243.960 180.330 ;
        RECT 243.710 179.900 244.360 180.300 ;
        RECT 243.720 178.760 243.960 179.900 ;
        RECT 256.580 178.760 256.830 178.810 ;
        RECT 258.860 178.760 259.100 180.440 ;
        RECT 243.720 178.590 259.100 178.760 ;
        RECT 276.440 178.730 277.490 178.750 ;
        RECT 243.720 178.520 258.830 178.590 ;
        RECT 256.580 172.430 256.830 178.520 ;
        RECT 276.430 178.230 277.490 178.730 ;
        RECT 276.430 177.480 276.750 178.230 ;
        RECT 276.430 175.910 276.740 177.480 ;
        RECT 243.540 171.880 244.020 172.280 ;
        RECT 171.070 169.360 171.550 169.580 ;
        RECT 129.420 164.510 138.190 164.520 ;
        RECT 141.180 164.510 141.510 164.880 ;
        RECT 129.420 164.460 141.510 164.510 ;
        RECT 128.560 164.450 141.510 164.460 ;
        RECT 125.540 164.440 141.510 164.450 ;
        RECT 123.470 164.230 141.510 164.440 ;
        RECT 123.470 164.220 129.630 164.230 ;
        RECT 123.470 164.210 128.640 164.220 ;
        RECT 108.330 164.200 125.570 164.210 ;
        RECT 108.330 164.040 123.710 164.200 ;
        RECT 108.330 163.970 123.440 164.040 ;
        RECT 121.330 163.920 121.630 163.970 ;
        RECT 136.470 162.330 136.660 164.230 ;
        RECT 137.890 164.220 141.510 164.230 ;
        RECT 157.920 162.330 158.330 162.340 ;
        RECT 159.260 162.330 159.630 162.450 ;
        RECT 136.470 162.090 159.630 162.330 ;
        RECT 56.540 158.600 64.620 158.620 ;
        RECT 69.720 158.600 86.450 158.750 ;
        RECT 56.540 158.250 86.450 158.600 ;
        RECT 56.610 158.230 57.020 158.250 ;
        RECT 63.360 158.230 86.450 158.250 ;
        RECT 69.720 158.220 86.450 158.230 ;
        RECT 69.790 158.170 70.240 158.220 ;
        RECT 39.880 148.720 40.930 148.740 ;
        RECT 39.870 148.220 40.930 148.720 ;
        RECT 39.870 147.470 40.190 148.220 ;
        RECT 39.870 145.900 40.180 147.470 ;
        RECT 39.840 135.000 40.200 145.900 ;
        RECT 28.080 134.630 36.850 134.640 ;
        RECT 39.840 134.630 40.170 135.000 ;
        RECT 28.080 134.580 40.170 134.630 ;
        RECT 27.220 134.570 40.170 134.580 ;
        RECT 24.200 134.560 40.170 134.570 ;
        RECT 22.130 134.350 40.170 134.560 ;
        RECT 22.130 134.340 28.290 134.350 ;
        RECT 22.130 134.330 27.300 134.340 ;
        RECT 6.990 134.320 24.230 134.330 ;
        RECT 6.990 134.160 22.370 134.320 ;
        RECT 35.160 134.260 35.350 134.350 ;
        RECT 36.550 134.340 40.170 134.350 ;
        RECT 6.990 134.090 22.100 134.160 ;
        RECT 19.990 134.040 20.290 134.090 ;
        RECT 85.910 133.180 86.410 158.220 ;
        RECT 108.460 156.100 108.940 156.500 ;
        RECT 108.460 150.130 108.650 156.100 ;
        RECT 124.100 154.000 124.310 154.010 ;
        RECT 123.650 153.960 124.570 154.000 ;
        RECT 123.600 153.920 124.570 153.960 ;
        RECT 123.600 153.650 124.580 153.920 ;
        RECT 123.600 153.620 124.570 153.650 ;
        RECT 123.600 151.390 123.840 153.620 ;
        RECT 124.100 153.610 124.310 153.620 ;
        RECT 123.600 150.240 123.850 151.390 ;
        RECT 108.460 150.100 108.710 150.130 ;
        RECT 108.460 149.700 109.110 150.100 ;
        RECT 108.470 148.560 108.710 149.700 ;
        RECT 121.330 148.560 121.580 148.610 ;
        RECT 123.610 148.560 123.850 150.240 ;
        RECT 108.470 148.390 123.850 148.560 ;
        RECT 108.470 148.320 123.580 148.390 ;
        RECT 121.330 142.230 121.580 148.320 ;
        RECT 108.290 141.680 108.770 142.080 ;
        RECT 108.290 135.710 108.480 141.680 ;
        RECT 108.290 135.680 108.540 135.710 ;
        RECT 108.290 135.280 108.940 135.680 ;
        RECT 108.300 134.140 108.540 135.280 ;
        RECT 121.300 134.140 121.600 142.230 ;
        RECT 123.930 139.580 124.140 139.590 ;
        RECT 123.480 139.540 124.400 139.580 ;
        RECT 123.430 139.500 124.400 139.540 ;
        RECT 123.430 139.230 124.410 139.500 ;
        RECT 123.430 139.200 124.400 139.230 ;
        RECT 123.430 136.970 123.670 139.200 ;
        RECT 123.930 139.190 124.140 139.200 ;
        RECT 123.430 135.820 123.680 136.970 ;
        RECT 123.440 134.370 123.680 135.820 ;
        RECT 136.470 134.450 136.660 162.090 ;
        RECT 157.920 158.430 158.330 162.090 ;
        RECT 171.100 158.560 171.550 169.360 ;
        RECT 243.540 165.910 243.730 171.880 ;
        RECT 243.540 165.880 243.790 165.910 ;
        RECT 243.540 165.480 244.190 165.880 ;
        RECT 243.550 164.340 243.790 165.480 ;
        RECT 256.550 164.340 256.850 172.430 ;
        RECT 259.180 169.780 259.390 169.790 ;
        RECT 258.730 169.740 259.650 169.780 ;
        RECT 258.680 169.700 259.650 169.740 ;
        RECT 258.680 169.430 259.660 169.700 ;
        RECT 258.680 169.400 259.650 169.430 ;
        RECT 258.680 167.170 258.920 169.400 ;
        RECT 259.180 169.390 259.390 169.400 ;
        RECT 258.680 166.020 258.930 167.170 ;
        RECT 258.690 164.570 258.930 166.020 ;
        RECT 276.400 165.010 276.760 175.910 ;
        RECT 306.290 169.710 306.740 191.950 ;
        RECT 407.600 191.760 408.080 192.170 ;
        RECT 345.020 186.110 345.500 186.510 ;
        RECT 345.020 180.140 345.210 186.110 ;
        RECT 360.660 184.010 360.870 184.020 ;
        RECT 360.210 183.970 361.130 184.010 ;
        RECT 360.160 183.930 361.130 183.970 ;
        RECT 360.160 183.660 361.140 183.930 ;
        RECT 360.160 183.630 361.130 183.660 ;
        RECT 360.160 181.400 360.400 183.630 ;
        RECT 360.660 183.620 360.870 183.630 ;
        RECT 360.160 180.250 360.410 181.400 ;
        RECT 345.020 180.110 345.270 180.140 ;
        RECT 345.020 179.710 345.670 180.110 ;
        RECT 345.030 178.570 345.270 179.710 ;
        RECT 357.890 178.570 358.140 178.620 ;
        RECT 360.170 178.570 360.410 180.250 ;
        RECT 345.030 178.400 360.410 178.570 ;
        RECT 377.750 178.540 378.800 178.560 ;
        RECT 345.030 178.330 360.140 178.400 ;
        RECT 357.890 172.240 358.140 178.330 ;
        RECT 377.740 178.040 378.800 178.540 ;
        RECT 377.740 177.290 378.060 178.040 ;
        RECT 377.740 175.720 378.050 177.290 ;
        RECT 344.850 171.690 345.330 172.090 ;
        RECT 306.290 169.490 306.770 169.710 ;
        RECT 264.640 164.640 273.410 164.650 ;
        RECT 276.400 164.640 276.730 165.010 ;
        RECT 264.640 164.590 276.730 164.640 ;
        RECT 263.780 164.580 276.730 164.590 ;
        RECT 260.760 164.570 276.730 164.580 ;
        RECT 258.690 164.360 276.730 164.570 ;
        RECT 258.690 164.350 264.850 164.360 ;
        RECT 258.690 164.340 263.860 164.350 ;
        RECT 243.550 164.330 260.790 164.340 ;
        RECT 243.550 164.170 258.930 164.330 ;
        RECT 243.550 164.100 258.660 164.170 ;
        RECT 256.550 164.050 256.850 164.100 ;
        RECT 271.690 162.460 271.880 164.360 ;
        RECT 273.110 164.350 276.730 164.360 ;
        RECT 293.140 162.460 293.550 162.470 ;
        RECT 294.480 162.460 294.850 162.580 ;
        RECT 271.690 162.220 294.850 162.460 ;
        RECT 157.850 158.410 165.930 158.430 ;
        RECT 171.030 158.410 187.760 158.560 ;
        RECT 157.850 158.060 187.760 158.410 ;
        RECT 157.920 158.040 158.330 158.060 ;
        RECT 164.670 158.040 187.760 158.060 ;
        RECT 171.030 158.030 187.760 158.040 ;
        RECT 171.100 157.980 171.550 158.030 ;
        RECT 141.190 148.530 142.240 148.550 ;
        RECT 141.180 148.030 142.240 148.530 ;
        RECT 141.180 147.280 141.500 148.030 ;
        RECT 141.180 145.710 141.490 147.280 ;
        RECT 141.150 134.810 141.510 145.710 ;
        RECT 129.390 134.440 138.160 134.450 ;
        RECT 141.150 134.440 141.480 134.810 ;
        RECT 129.390 134.390 141.480 134.440 ;
        RECT 128.530 134.380 141.480 134.390 ;
        RECT 125.510 134.370 141.480 134.380 ;
        RECT 123.440 134.160 141.480 134.370 ;
        RECT 123.440 134.150 129.600 134.160 ;
        RECT 123.440 134.140 128.610 134.150 ;
        RECT 108.300 134.130 125.540 134.140 ;
        RECT 108.300 133.970 123.680 134.130 ;
        RECT 136.470 134.070 136.660 134.160 ;
        RECT 137.860 134.150 141.480 134.160 ;
        RECT 108.300 133.900 123.410 133.970 ;
        RECT 121.300 133.850 121.600 133.900 ;
        RECT 88.840 133.180 89.250 133.190 ;
        RECT 85.910 132.930 89.250 133.180 ;
        RECT 7.030 126.040 7.510 126.440 ;
        RECT 7.030 120.070 7.220 126.040 ;
        RECT 22.670 123.940 22.880 123.950 ;
        RECT 22.220 123.900 23.140 123.940 ;
        RECT 22.170 123.860 23.140 123.900 ;
        RECT 22.170 123.590 23.150 123.860 ;
        RECT 22.170 123.560 23.140 123.590 ;
        RECT 22.170 121.330 22.410 123.560 ;
        RECT 22.670 123.550 22.880 123.560 ;
        RECT 22.170 120.180 22.420 121.330 ;
        RECT 7.030 120.040 7.280 120.070 ;
        RECT 7.030 119.640 7.680 120.040 ;
        RECT 7.040 118.500 7.280 119.640 ;
        RECT 19.900 118.500 20.150 118.550 ;
        RECT 22.180 118.500 22.420 120.180 ;
        RECT 7.040 118.330 22.420 118.500 ;
        RECT 39.760 118.470 40.810 118.490 ;
        RECT 7.040 118.260 22.150 118.330 ;
        RECT 19.900 112.170 20.150 118.260 ;
        RECT 39.750 117.970 40.810 118.470 ;
        RECT 39.750 117.220 40.070 117.970 ;
        RECT 39.750 115.650 40.060 117.220 ;
        RECT 6.860 111.620 7.340 112.020 ;
        RECT 6.860 105.650 7.050 111.620 ;
        RECT 6.860 105.620 7.110 105.650 ;
        RECT 6.860 105.220 7.510 105.620 ;
        RECT 6.870 104.080 7.110 105.220 ;
        RECT 19.870 104.080 20.170 112.170 ;
        RECT 22.500 109.520 22.710 109.530 ;
        RECT 22.050 109.480 22.970 109.520 ;
        RECT 22.000 109.440 22.970 109.480 ;
        RECT 22.000 109.170 22.980 109.440 ;
        RECT 22.000 109.140 22.970 109.170 ;
        RECT 22.000 106.910 22.240 109.140 ;
        RECT 22.500 109.130 22.710 109.140 ;
        RECT 22.000 105.760 22.250 106.910 ;
        RECT 22.010 104.310 22.250 105.760 ;
        RECT 39.720 104.750 40.080 115.650 ;
        RECT 85.910 111.210 86.410 132.930 ;
        RECT 88.840 132.790 89.250 132.930 ;
        RECT 187.220 132.990 187.720 158.030 ;
        RECT 243.680 156.230 244.160 156.630 ;
        RECT 243.680 150.260 243.870 156.230 ;
        RECT 259.320 154.130 259.530 154.140 ;
        RECT 258.870 154.090 259.790 154.130 ;
        RECT 258.820 154.050 259.790 154.090 ;
        RECT 258.820 153.780 259.800 154.050 ;
        RECT 258.820 153.750 259.790 153.780 ;
        RECT 258.820 151.520 259.060 153.750 ;
        RECT 259.320 153.740 259.530 153.750 ;
        RECT 258.820 150.370 259.070 151.520 ;
        RECT 243.680 150.230 243.930 150.260 ;
        RECT 243.680 149.830 244.330 150.230 ;
        RECT 243.690 148.690 243.930 149.830 ;
        RECT 256.550 148.690 256.800 148.740 ;
        RECT 258.830 148.690 259.070 150.370 ;
        RECT 243.690 148.520 259.070 148.690 ;
        RECT 243.690 148.450 258.800 148.520 ;
        RECT 256.550 142.360 256.800 148.450 ;
        RECT 243.510 141.810 243.990 142.210 ;
        RECT 243.510 135.840 243.700 141.810 ;
        RECT 243.510 135.810 243.760 135.840 ;
        RECT 243.510 135.410 244.160 135.810 ;
        RECT 216.010 135.380 216.900 135.400 ;
        RECT 215.980 134.910 216.900 135.380 ;
        RECT 190.150 132.990 190.560 133.000 ;
        RECT 187.220 132.740 190.560 132.990 ;
        RECT 187.220 131.290 187.720 132.740 ;
        RECT 190.150 132.600 190.560 132.740 ;
        RECT 215.980 131.450 216.160 134.910 ;
        RECT 243.520 134.270 243.760 135.410 ;
        RECT 256.520 134.270 256.820 142.360 ;
        RECT 259.150 139.710 259.360 139.720 ;
        RECT 258.700 139.670 259.620 139.710 ;
        RECT 258.650 139.630 259.620 139.670 ;
        RECT 258.650 139.360 259.630 139.630 ;
        RECT 258.650 139.330 259.620 139.360 ;
        RECT 258.650 137.100 258.890 139.330 ;
        RECT 259.150 139.320 259.360 139.330 ;
        RECT 258.650 135.950 258.900 137.100 ;
        RECT 258.660 134.500 258.900 135.950 ;
        RECT 271.690 134.580 271.880 162.220 ;
        RECT 293.140 158.560 293.550 162.220 ;
        RECT 306.320 158.690 306.770 169.490 ;
        RECT 344.850 165.720 345.040 171.690 ;
        RECT 344.850 165.690 345.100 165.720 ;
        RECT 344.850 165.290 345.500 165.690 ;
        RECT 344.860 164.150 345.100 165.290 ;
        RECT 357.860 164.150 358.160 172.240 ;
        RECT 360.490 169.590 360.700 169.600 ;
        RECT 360.040 169.550 360.960 169.590 ;
        RECT 359.990 169.510 360.960 169.550 ;
        RECT 359.990 169.240 360.970 169.510 ;
        RECT 359.990 169.210 360.960 169.240 ;
        RECT 359.990 166.980 360.230 169.210 ;
        RECT 360.490 169.200 360.700 169.210 ;
        RECT 359.990 165.830 360.240 166.980 ;
        RECT 360.000 164.380 360.240 165.830 ;
        RECT 377.710 164.820 378.070 175.720 ;
        RECT 407.600 169.520 408.050 191.760 ;
        RECT 407.600 169.300 408.080 169.520 ;
        RECT 365.950 164.450 374.720 164.460 ;
        RECT 377.710 164.450 378.040 164.820 ;
        RECT 365.950 164.400 378.040 164.450 ;
        RECT 365.090 164.390 378.040 164.400 ;
        RECT 362.070 164.380 378.040 164.390 ;
        RECT 360.000 164.170 378.040 164.380 ;
        RECT 360.000 164.160 366.160 164.170 ;
        RECT 360.000 164.150 365.170 164.160 ;
        RECT 344.860 164.140 362.100 164.150 ;
        RECT 344.860 163.980 360.240 164.140 ;
        RECT 344.860 163.910 359.970 163.980 ;
        RECT 357.860 163.860 358.160 163.910 ;
        RECT 373.000 162.270 373.190 164.170 ;
        RECT 374.420 164.160 378.040 164.170 ;
        RECT 394.450 162.270 394.860 162.280 ;
        RECT 395.790 162.270 396.160 162.390 ;
        RECT 373.000 162.030 396.160 162.270 ;
        RECT 293.070 158.540 301.150 158.560 ;
        RECT 306.250 158.540 322.980 158.690 ;
        RECT 293.070 158.190 322.980 158.540 ;
        RECT 293.140 158.170 293.550 158.190 ;
        RECT 299.890 158.170 322.980 158.190 ;
        RECT 306.250 158.160 322.980 158.170 ;
        RECT 306.320 158.110 306.770 158.160 ;
        RECT 276.410 148.660 277.460 148.680 ;
        RECT 276.400 148.160 277.460 148.660 ;
        RECT 276.400 147.410 276.720 148.160 ;
        RECT 276.400 145.840 276.710 147.410 ;
        RECT 276.370 134.940 276.730 145.840 ;
        RECT 264.610 134.570 273.380 134.580 ;
        RECT 276.370 134.570 276.700 134.940 ;
        RECT 264.610 134.520 276.700 134.570 ;
        RECT 263.750 134.510 276.700 134.520 ;
        RECT 260.730 134.500 276.700 134.510 ;
        RECT 258.660 134.290 276.700 134.500 ;
        RECT 258.660 134.280 264.820 134.290 ;
        RECT 258.660 134.270 263.830 134.280 ;
        RECT 243.520 134.260 260.760 134.270 ;
        RECT 243.520 134.100 258.900 134.260 ;
        RECT 271.690 134.200 271.880 134.290 ;
        RECT 273.080 134.280 276.700 134.290 ;
        RECT 243.520 134.030 258.630 134.100 ;
        RECT 256.520 133.980 256.820 134.030 ;
        RECT 322.440 133.120 322.940 158.160 ;
        RECT 344.990 156.040 345.470 156.440 ;
        RECT 344.990 150.070 345.180 156.040 ;
        RECT 360.630 153.940 360.840 153.950 ;
        RECT 360.180 153.900 361.100 153.940 ;
        RECT 360.130 153.860 361.100 153.900 ;
        RECT 360.130 153.590 361.110 153.860 ;
        RECT 360.130 153.560 361.100 153.590 ;
        RECT 360.130 151.330 360.370 153.560 ;
        RECT 360.630 153.550 360.840 153.560 ;
        RECT 360.130 150.180 360.380 151.330 ;
        RECT 344.990 150.040 345.240 150.070 ;
        RECT 344.990 149.640 345.640 150.040 ;
        RECT 345.000 148.500 345.240 149.640 ;
        RECT 357.860 148.500 358.110 148.550 ;
        RECT 360.140 148.500 360.380 150.180 ;
        RECT 345.000 148.330 360.380 148.500 ;
        RECT 345.000 148.260 360.110 148.330 ;
        RECT 357.860 142.170 358.110 148.260 ;
        RECT 344.820 141.620 345.300 142.020 ;
        RECT 344.820 135.650 345.010 141.620 ;
        RECT 344.820 135.620 345.070 135.650 ;
        RECT 344.820 135.220 345.470 135.620 ;
        RECT 344.830 134.080 345.070 135.220 ;
        RECT 357.830 134.080 358.130 142.170 ;
        RECT 360.460 139.520 360.670 139.530 ;
        RECT 360.010 139.480 360.930 139.520 ;
        RECT 359.960 139.440 360.930 139.480 ;
        RECT 359.960 139.170 360.940 139.440 ;
        RECT 359.960 139.140 360.930 139.170 ;
        RECT 359.960 136.910 360.200 139.140 ;
        RECT 360.460 139.130 360.670 139.140 ;
        RECT 359.960 135.760 360.210 136.910 ;
        RECT 359.970 134.310 360.210 135.760 ;
        RECT 373.000 134.390 373.190 162.030 ;
        RECT 394.450 158.370 394.860 162.030 ;
        RECT 407.630 158.500 408.080 169.300 ;
        RECT 394.380 158.350 402.460 158.370 ;
        RECT 407.560 158.350 424.290 158.500 ;
        RECT 394.380 158.000 424.290 158.350 ;
        RECT 394.450 157.980 394.860 158.000 ;
        RECT 401.200 157.980 424.290 158.000 ;
        RECT 407.560 157.970 424.290 157.980 ;
        RECT 407.630 157.920 408.080 157.970 ;
        RECT 377.720 148.470 378.770 148.490 ;
        RECT 377.710 147.970 378.770 148.470 ;
        RECT 377.710 147.220 378.030 147.970 ;
        RECT 377.710 145.650 378.020 147.220 ;
        RECT 377.680 134.750 378.040 145.650 ;
        RECT 365.920 134.380 374.690 134.390 ;
        RECT 377.680 134.380 378.010 134.750 ;
        RECT 365.920 134.330 378.010 134.380 ;
        RECT 365.060 134.320 378.010 134.330 ;
        RECT 362.040 134.310 378.010 134.320 ;
        RECT 359.970 134.100 378.010 134.310 ;
        RECT 359.970 134.090 366.130 134.100 ;
        RECT 359.970 134.080 365.140 134.090 ;
        RECT 344.830 134.070 362.070 134.080 ;
        RECT 344.830 133.910 360.210 134.070 ;
        RECT 373.000 134.010 373.190 134.100 ;
        RECT 374.390 134.090 378.010 134.100 ;
        RECT 344.830 133.840 359.940 133.910 ;
        RECT 357.830 133.790 358.130 133.840 ;
        RECT 325.370 133.120 325.780 133.130 ;
        RECT 322.440 132.870 325.780 133.120 ;
        RECT 187.220 131.230 211.110 131.290 ;
        RECT 215.980 131.230 216.140 131.450 ;
        RECT 187.220 131.060 216.140 131.230 ;
        RECT 108.340 125.850 108.820 126.250 ;
        RECT 108.340 119.880 108.530 125.850 ;
        RECT 123.980 123.750 124.190 123.760 ;
        RECT 123.530 123.710 124.450 123.750 ;
        RECT 123.480 123.670 124.450 123.710 ;
        RECT 123.480 123.400 124.460 123.670 ;
        RECT 123.480 123.370 124.450 123.400 ;
        RECT 123.480 121.140 123.720 123.370 ;
        RECT 123.980 123.360 124.190 123.370 ;
        RECT 123.480 119.990 123.730 121.140 ;
        RECT 108.340 119.850 108.590 119.880 ;
        RECT 108.340 119.450 108.990 119.850 ;
        RECT 108.350 118.310 108.590 119.450 ;
        RECT 121.210 118.310 121.460 118.360 ;
        RECT 123.490 118.310 123.730 119.990 ;
        RECT 108.350 118.140 123.730 118.310 ;
        RECT 141.070 118.280 142.120 118.300 ;
        RECT 108.350 118.070 123.460 118.140 ;
        RECT 121.210 111.980 121.460 118.070 ;
        RECT 141.060 117.780 142.120 118.280 ;
        RECT 141.060 117.030 141.380 117.780 ;
        RECT 141.060 115.460 141.370 117.030 ;
        RECT 108.170 111.430 108.650 111.830 ;
        RECT 27.960 104.380 36.730 104.390 ;
        RECT 39.720 104.380 40.050 104.750 ;
        RECT 27.960 104.330 40.050 104.380 ;
        RECT 27.100 104.320 40.050 104.330 ;
        RECT 24.080 104.310 40.050 104.320 ;
        RECT 22.010 104.100 40.050 104.310 ;
        RECT 22.010 104.090 28.170 104.100 ;
        RECT 22.010 104.080 27.180 104.090 ;
        RECT 6.870 104.070 24.110 104.080 ;
        RECT 6.870 103.910 22.250 104.070 ;
        RECT 6.870 103.840 21.980 103.910 ;
        RECT 19.870 103.790 20.170 103.840 ;
        RECT 35.010 102.200 35.200 104.100 ;
        RECT 36.430 104.090 40.050 104.100 ;
        RECT 54.620 102.200 55.070 102.280 ;
        RECT 57.800 102.200 58.170 102.320 ;
        RECT 35.010 101.960 58.170 102.200 ;
        RECT 7.000 95.970 7.480 96.370 ;
        RECT 7.000 90.000 7.190 95.970 ;
        RECT 22.640 93.870 22.850 93.880 ;
        RECT 22.190 93.830 23.110 93.870 ;
        RECT 22.140 93.790 23.110 93.830 ;
        RECT 22.140 93.520 23.120 93.790 ;
        RECT 22.140 93.490 23.110 93.520 ;
        RECT 22.140 91.260 22.380 93.490 ;
        RECT 22.640 93.480 22.850 93.490 ;
        RECT 22.140 90.110 22.390 91.260 ;
        RECT 7.000 89.970 7.250 90.000 ;
        RECT 7.000 89.570 7.650 89.970 ;
        RECT 7.010 88.430 7.250 89.570 ;
        RECT 19.870 88.430 20.120 88.480 ;
        RECT 22.150 88.430 22.390 90.110 ;
        RECT 7.010 88.260 22.390 88.430 ;
        RECT 7.010 88.190 22.120 88.260 ;
        RECT 19.870 82.100 20.120 88.190 ;
        RECT 6.830 81.550 7.310 81.950 ;
        RECT 6.830 75.580 7.020 81.550 ;
        RECT 6.830 75.550 7.080 75.580 ;
        RECT 6.830 75.150 7.480 75.550 ;
        RECT 6.840 74.010 7.080 75.150 ;
        RECT 19.840 74.010 20.140 82.100 ;
        RECT 22.470 79.450 22.680 79.460 ;
        RECT 22.020 79.410 22.940 79.450 ;
        RECT 21.970 79.370 22.940 79.410 ;
        RECT 21.970 79.100 22.950 79.370 ;
        RECT 21.970 79.070 22.940 79.100 ;
        RECT 21.970 76.840 22.210 79.070 ;
        RECT 22.470 79.060 22.680 79.070 ;
        RECT 21.970 75.690 22.220 76.840 ;
        RECT 21.980 74.240 22.220 75.690 ;
        RECT 35.010 74.320 35.200 101.960 ;
        RECT 54.620 97.430 55.070 101.960 ;
        RECT 85.880 98.640 86.450 111.210 ;
        RECT 108.170 105.460 108.360 111.430 ;
        RECT 108.170 105.430 108.420 105.460 ;
        RECT 108.170 105.030 108.820 105.430 ;
        RECT 108.180 103.890 108.420 105.030 ;
        RECT 121.180 103.890 121.480 111.980 ;
        RECT 123.810 109.330 124.020 109.340 ;
        RECT 123.360 109.290 124.280 109.330 ;
        RECT 123.310 109.250 124.280 109.290 ;
        RECT 123.310 108.980 124.290 109.250 ;
        RECT 123.310 108.950 124.280 108.980 ;
        RECT 123.310 106.720 123.550 108.950 ;
        RECT 123.810 108.940 124.020 108.950 ;
        RECT 123.310 105.570 123.560 106.720 ;
        RECT 123.320 104.120 123.560 105.570 ;
        RECT 141.030 104.560 141.390 115.460 ;
        RECT 187.220 111.020 187.720 131.060 ;
        RECT 215.980 131.050 216.140 131.060 ;
        RECT 243.560 125.980 244.040 126.380 ;
        RECT 243.560 120.010 243.750 125.980 ;
        RECT 259.200 123.880 259.410 123.890 ;
        RECT 258.750 123.840 259.670 123.880 ;
        RECT 258.700 123.800 259.670 123.840 ;
        RECT 258.700 123.530 259.680 123.800 ;
        RECT 258.700 123.500 259.670 123.530 ;
        RECT 258.700 121.270 258.940 123.500 ;
        RECT 259.200 123.490 259.410 123.500 ;
        RECT 258.700 120.120 258.950 121.270 ;
        RECT 243.560 119.980 243.810 120.010 ;
        RECT 243.560 119.580 244.210 119.980 ;
        RECT 243.570 118.440 243.810 119.580 ;
        RECT 256.430 118.440 256.680 118.490 ;
        RECT 258.710 118.440 258.950 120.120 ;
        RECT 243.570 118.270 258.950 118.440 ;
        RECT 276.290 118.410 277.340 118.430 ;
        RECT 243.570 118.200 258.680 118.270 ;
        RECT 256.430 112.110 256.680 118.200 ;
        RECT 276.280 117.910 277.340 118.410 ;
        RECT 276.280 117.160 276.600 117.910 ;
        RECT 276.280 115.590 276.590 117.160 ;
        RECT 243.390 111.560 243.870 111.960 ;
        RECT 129.270 104.190 138.040 104.200 ;
        RECT 141.030 104.190 141.360 104.560 ;
        RECT 129.270 104.140 141.360 104.190 ;
        RECT 128.410 104.130 141.360 104.140 ;
        RECT 125.390 104.120 141.360 104.130 ;
        RECT 123.320 103.910 141.360 104.120 ;
        RECT 123.320 103.900 129.480 103.910 ;
        RECT 123.320 103.890 128.490 103.900 ;
        RECT 108.180 103.880 125.420 103.890 ;
        RECT 108.180 103.720 123.560 103.880 ;
        RECT 108.180 103.650 123.290 103.720 ;
        RECT 121.180 103.600 121.480 103.650 ;
        RECT 136.320 102.010 136.510 103.910 ;
        RECT 137.740 103.900 141.360 103.910 ;
        RECT 155.930 102.010 156.380 102.090 ;
        RECT 159.110 102.010 159.480 102.130 ;
        RECT 136.320 101.770 159.480 102.010 ;
        RECT 85.880 98.070 86.520 98.640 ;
        RECT 54.620 97.370 69.440 97.430 ;
        RECT 54.620 96.910 69.740 97.370 ;
        RECT 69.290 96.260 69.740 96.910 ;
        RECT 85.910 96.260 86.520 98.070 ;
        RECT 69.290 95.730 86.520 96.260 ;
        RECT 39.730 88.400 40.780 88.420 ;
        RECT 39.720 87.900 40.780 88.400 ;
        RECT 39.720 87.150 40.040 87.900 ;
        RECT 39.720 85.580 40.030 87.150 ;
        RECT 39.690 74.680 40.050 85.580 ;
        RECT 69.290 75.890 69.740 95.730 ;
        RECT 85.910 95.590 86.520 95.730 ;
        RECT 108.310 95.780 108.790 96.180 ;
        RECT 108.310 89.810 108.500 95.780 ;
        RECT 123.950 93.680 124.160 93.690 ;
        RECT 123.500 93.640 124.420 93.680 ;
        RECT 123.450 93.600 124.420 93.640 ;
        RECT 123.450 93.330 124.430 93.600 ;
        RECT 123.450 93.300 124.420 93.330 ;
        RECT 123.450 91.070 123.690 93.300 ;
        RECT 123.950 93.290 124.160 93.300 ;
        RECT 123.450 89.920 123.700 91.070 ;
        RECT 108.310 89.780 108.560 89.810 ;
        RECT 108.310 89.380 108.960 89.780 ;
        RECT 108.320 88.240 108.560 89.380 ;
        RECT 121.180 88.240 121.430 88.290 ;
        RECT 123.460 88.240 123.700 89.920 ;
        RECT 108.320 88.070 123.700 88.240 ;
        RECT 108.320 88.000 123.430 88.070 ;
        RECT 121.180 81.910 121.430 88.000 ;
        RECT 108.140 81.360 108.620 81.760 ;
        RECT 72.010 75.890 72.370 76.200 ;
        RECT 69.270 75.630 72.370 75.890 ;
        RECT 27.930 74.310 36.700 74.320 ;
        RECT 39.690 74.310 40.020 74.680 ;
        RECT 27.930 74.260 40.020 74.310 ;
        RECT 27.070 74.250 40.020 74.260 ;
        RECT 24.050 74.240 40.020 74.250 ;
        RECT 21.980 74.030 40.020 74.240 ;
        RECT 21.980 74.020 28.140 74.030 ;
        RECT 21.980 74.010 27.150 74.020 ;
        RECT 6.840 74.000 24.080 74.010 ;
        RECT 6.840 73.840 22.220 74.000 ;
        RECT 35.010 73.940 35.200 74.030 ;
        RECT 36.400 74.020 40.020 74.030 ;
        RECT 6.840 73.770 21.950 73.840 ;
        RECT 19.840 73.720 20.140 73.770 ;
        RECT 69.290 72.180 69.740 75.630 ;
        RECT 108.140 75.390 108.330 81.360 ;
        RECT 108.140 75.360 108.390 75.390 ;
        RECT 108.140 74.960 108.790 75.360 ;
        RECT 108.150 73.820 108.390 74.960 ;
        RECT 121.150 73.820 121.450 81.910 ;
        RECT 123.780 79.260 123.990 79.270 ;
        RECT 123.330 79.220 124.250 79.260 ;
        RECT 123.280 79.180 124.250 79.220 ;
        RECT 123.280 78.910 124.260 79.180 ;
        RECT 123.280 78.880 124.250 78.910 ;
        RECT 123.280 76.650 123.520 78.880 ;
        RECT 123.780 78.870 123.990 78.880 ;
        RECT 123.280 75.500 123.530 76.650 ;
        RECT 123.290 74.050 123.530 75.500 ;
        RECT 136.320 74.130 136.510 101.770 ;
        RECT 155.930 97.240 156.380 101.770 ;
        RECT 187.190 98.450 187.760 111.020 ;
        RECT 243.390 105.590 243.580 111.560 ;
        RECT 243.390 105.560 243.640 105.590 ;
        RECT 243.390 105.160 244.040 105.560 ;
        RECT 243.400 104.020 243.640 105.160 ;
        RECT 256.400 104.020 256.700 112.110 ;
        RECT 259.030 109.460 259.240 109.470 ;
        RECT 258.580 109.420 259.500 109.460 ;
        RECT 258.530 109.380 259.500 109.420 ;
        RECT 258.530 109.110 259.510 109.380 ;
        RECT 258.530 109.080 259.500 109.110 ;
        RECT 258.530 106.850 258.770 109.080 ;
        RECT 259.030 109.070 259.240 109.080 ;
        RECT 258.530 105.700 258.780 106.850 ;
        RECT 258.540 104.250 258.780 105.700 ;
        RECT 276.250 104.690 276.610 115.590 ;
        RECT 322.440 111.150 322.940 132.870 ;
        RECT 325.370 132.730 325.780 132.870 ;
        RECT 423.750 132.930 424.250 157.970 ;
        RECT 452.540 135.320 453.430 135.340 ;
        RECT 452.510 134.850 453.430 135.320 ;
        RECT 426.680 132.930 427.090 132.940 ;
        RECT 423.750 132.680 427.090 132.930 ;
        RECT 423.750 131.230 424.250 132.680 ;
        RECT 426.680 132.540 427.090 132.680 ;
        RECT 452.510 131.390 452.690 134.850 ;
        RECT 469.670 132.930 470.730 132.960 ;
        RECT 469.570 132.500 470.730 132.930 ;
        RECT 423.750 131.170 447.640 131.230 ;
        RECT 452.510 131.190 452.670 131.390 ;
        RECT 469.570 131.200 469.770 132.500 ;
        RECT 455.060 131.190 469.790 131.200 ;
        RECT 452.500 131.170 469.790 131.190 ;
        RECT 423.750 131.010 469.790 131.170 ;
        RECT 423.750 131.000 460.150 131.010 ;
        RECT 344.870 125.790 345.350 126.190 ;
        RECT 344.870 119.820 345.060 125.790 ;
        RECT 360.510 123.690 360.720 123.700 ;
        RECT 360.060 123.650 360.980 123.690 ;
        RECT 360.010 123.610 360.980 123.650 ;
        RECT 360.010 123.340 360.990 123.610 ;
        RECT 360.010 123.310 360.980 123.340 ;
        RECT 360.010 121.080 360.250 123.310 ;
        RECT 360.510 123.300 360.720 123.310 ;
        RECT 360.010 119.930 360.260 121.080 ;
        RECT 344.870 119.790 345.120 119.820 ;
        RECT 344.870 119.390 345.520 119.790 ;
        RECT 344.880 118.250 345.120 119.390 ;
        RECT 357.740 118.250 357.990 118.300 ;
        RECT 360.020 118.250 360.260 119.930 ;
        RECT 344.880 118.080 360.260 118.250 ;
        RECT 377.600 118.220 378.650 118.240 ;
        RECT 344.880 118.010 359.990 118.080 ;
        RECT 357.740 111.920 357.990 118.010 ;
        RECT 377.590 117.720 378.650 118.220 ;
        RECT 377.590 116.970 377.910 117.720 ;
        RECT 377.590 115.400 377.900 116.970 ;
        RECT 344.700 111.370 345.180 111.770 ;
        RECT 264.490 104.320 273.260 104.330 ;
        RECT 276.250 104.320 276.580 104.690 ;
        RECT 264.490 104.270 276.580 104.320 ;
        RECT 263.630 104.260 276.580 104.270 ;
        RECT 260.610 104.250 276.580 104.260 ;
        RECT 258.540 104.040 276.580 104.250 ;
        RECT 258.540 104.030 264.700 104.040 ;
        RECT 258.540 104.020 263.710 104.030 ;
        RECT 243.400 104.010 260.640 104.020 ;
        RECT 243.400 103.850 258.780 104.010 ;
        RECT 243.400 103.780 258.510 103.850 ;
        RECT 256.400 103.730 256.700 103.780 ;
        RECT 271.540 102.140 271.730 104.040 ;
        RECT 272.960 104.030 276.580 104.040 ;
        RECT 291.150 102.140 291.600 102.220 ;
        RECT 294.330 102.140 294.700 102.260 ;
        RECT 271.540 101.900 294.700 102.140 ;
        RECT 187.190 97.880 187.830 98.450 ;
        RECT 155.930 97.180 170.750 97.240 ;
        RECT 155.930 96.720 171.050 97.180 ;
        RECT 170.600 96.070 171.050 96.720 ;
        RECT 187.220 96.070 187.830 97.880 ;
        RECT 170.600 95.540 187.830 96.070 ;
        RECT 141.040 88.210 142.090 88.230 ;
        RECT 141.030 87.710 142.090 88.210 ;
        RECT 141.030 86.960 141.350 87.710 ;
        RECT 141.030 85.390 141.340 86.960 ;
        RECT 141.000 74.490 141.360 85.390 ;
        RECT 170.600 75.700 171.050 95.540 ;
        RECT 187.220 95.400 187.830 95.540 ;
        RECT 243.530 95.910 244.010 96.310 ;
        RECT 243.530 89.940 243.720 95.910 ;
        RECT 259.170 93.810 259.380 93.820 ;
        RECT 258.720 93.770 259.640 93.810 ;
        RECT 258.670 93.730 259.640 93.770 ;
        RECT 258.670 93.460 259.650 93.730 ;
        RECT 258.670 93.430 259.640 93.460 ;
        RECT 258.670 91.200 258.910 93.430 ;
        RECT 259.170 93.420 259.380 93.430 ;
        RECT 258.670 90.050 258.920 91.200 ;
        RECT 243.530 89.910 243.780 89.940 ;
        RECT 243.530 89.510 244.180 89.910 ;
        RECT 243.540 88.370 243.780 89.510 ;
        RECT 256.400 88.370 256.650 88.420 ;
        RECT 258.680 88.370 258.920 90.050 ;
        RECT 243.540 88.200 258.920 88.370 ;
        RECT 243.540 88.130 258.650 88.200 ;
        RECT 256.400 82.040 256.650 88.130 ;
        RECT 243.360 81.490 243.840 81.890 ;
        RECT 173.320 75.700 173.680 76.010 ;
        RECT 170.580 75.440 173.680 75.700 ;
        RECT 243.360 75.520 243.550 81.490 ;
        RECT 243.360 75.490 243.610 75.520 ;
        RECT 129.240 74.120 138.010 74.130 ;
        RECT 141.000 74.120 141.330 74.490 ;
        RECT 129.240 74.070 141.330 74.120 ;
        RECT 128.380 74.060 141.330 74.070 ;
        RECT 125.360 74.050 141.330 74.060 ;
        RECT 123.290 73.840 141.330 74.050 ;
        RECT 123.290 73.830 129.450 73.840 ;
        RECT 123.290 73.820 128.460 73.830 ;
        RECT 108.150 73.810 125.390 73.820 ;
        RECT 108.150 73.650 123.530 73.810 ;
        RECT 136.320 73.750 136.510 73.840 ;
        RECT 137.710 73.830 141.330 73.840 ;
        RECT 108.150 73.580 123.260 73.650 ;
        RECT 121.150 73.530 121.450 73.580 ;
        RECT 69.260 71.770 69.740 72.180 ;
        RECT 170.600 71.990 171.050 75.440 ;
        RECT 243.360 75.090 244.010 75.490 ;
        RECT 243.370 73.950 243.610 75.090 ;
        RECT 256.370 73.950 256.670 82.040 ;
        RECT 259.000 79.390 259.210 79.400 ;
        RECT 258.550 79.350 259.470 79.390 ;
        RECT 258.500 79.310 259.470 79.350 ;
        RECT 258.500 79.040 259.480 79.310 ;
        RECT 258.500 79.010 259.470 79.040 ;
        RECT 258.500 76.780 258.740 79.010 ;
        RECT 259.000 79.000 259.210 79.010 ;
        RECT 258.500 75.630 258.750 76.780 ;
        RECT 258.510 74.180 258.750 75.630 ;
        RECT 271.540 74.260 271.730 101.900 ;
        RECT 291.150 97.370 291.600 101.900 ;
        RECT 322.410 98.580 322.980 111.150 ;
        RECT 344.700 105.400 344.890 111.370 ;
        RECT 344.700 105.370 344.950 105.400 ;
        RECT 344.700 104.970 345.350 105.370 ;
        RECT 344.710 103.830 344.950 104.970 ;
        RECT 357.710 103.830 358.010 111.920 ;
        RECT 360.340 109.270 360.550 109.280 ;
        RECT 359.890 109.230 360.810 109.270 ;
        RECT 359.840 109.190 360.810 109.230 ;
        RECT 359.840 108.920 360.820 109.190 ;
        RECT 359.840 108.890 360.810 108.920 ;
        RECT 359.840 106.660 360.080 108.890 ;
        RECT 360.340 108.880 360.550 108.890 ;
        RECT 359.840 105.510 360.090 106.660 ;
        RECT 359.850 104.060 360.090 105.510 ;
        RECT 377.560 104.500 377.920 115.400 ;
        RECT 423.750 110.960 424.250 131.000 ;
        RECT 452.500 130.990 455.070 131.000 ;
        RECT 365.800 104.130 374.570 104.140 ;
        RECT 377.560 104.130 377.890 104.500 ;
        RECT 365.800 104.080 377.890 104.130 ;
        RECT 364.940 104.070 377.890 104.080 ;
        RECT 361.920 104.060 377.890 104.070 ;
        RECT 359.850 103.850 377.890 104.060 ;
        RECT 359.850 103.840 366.010 103.850 ;
        RECT 359.850 103.830 365.020 103.840 ;
        RECT 344.710 103.820 361.950 103.830 ;
        RECT 344.710 103.660 360.090 103.820 ;
        RECT 344.710 103.590 359.820 103.660 ;
        RECT 357.710 103.540 358.010 103.590 ;
        RECT 372.850 101.950 373.040 103.850 ;
        RECT 374.270 103.840 377.890 103.850 ;
        RECT 392.460 101.950 392.910 102.030 ;
        RECT 395.640 101.950 396.010 102.070 ;
        RECT 372.850 101.710 396.010 101.950 ;
        RECT 322.410 98.010 323.050 98.580 ;
        RECT 291.150 97.310 305.970 97.370 ;
        RECT 291.150 96.850 306.270 97.310 ;
        RECT 305.820 96.200 306.270 96.850 ;
        RECT 322.440 96.200 323.050 98.010 ;
        RECT 305.820 95.670 323.050 96.200 ;
        RECT 276.260 88.340 277.310 88.360 ;
        RECT 276.250 87.840 277.310 88.340 ;
        RECT 276.250 87.090 276.570 87.840 ;
        RECT 276.250 85.520 276.560 87.090 ;
        RECT 276.220 74.620 276.580 85.520 ;
        RECT 305.820 75.830 306.270 95.670 ;
        RECT 322.440 95.530 323.050 95.670 ;
        RECT 344.840 95.720 345.320 96.120 ;
        RECT 344.840 89.750 345.030 95.720 ;
        RECT 360.480 93.620 360.690 93.630 ;
        RECT 360.030 93.580 360.950 93.620 ;
        RECT 359.980 93.540 360.950 93.580 ;
        RECT 359.980 93.270 360.960 93.540 ;
        RECT 359.980 93.240 360.950 93.270 ;
        RECT 359.980 91.010 360.220 93.240 ;
        RECT 360.480 93.230 360.690 93.240 ;
        RECT 359.980 89.860 360.230 91.010 ;
        RECT 344.840 89.720 345.090 89.750 ;
        RECT 344.840 89.320 345.490 89.720 ;
        RECT 344.850 88.180 345.090 89.320 ;
        RECT 357.710 88.180 357.960 88.230 ;
        RECT 359.990 88.180 360.230 89.860 ;
        RECT 344.850 88.010 360.230 88.180 ;
        RECT 344.850 87.940 359.960 88.010 ;
        RECT 357.710 81.850 357.960 87.940 ;
        RECT 344.670 81.300 345.150 81.700 ;
        RECT 308.540 75.830 308.900 76.140 ;
        RECT 305.800 75.570 308.900 75.830 ;
        RECT 264.460 74.250 273.230 74.260 ;
        RECT 276.220 74.250 276.550 74.620 ;
        RECT 264.460 74.200 276.550 74.250 ;
        RECT 263.600 74.190 276.550 74.200 ;
        RECT 260.580 74.180 276.550 74.190 ;
        RECT 258.510 73.970 276.550 74.180 ;
        RECT 258.510 73.960 264.670 73.970 ;
        RECT 258.510 73.950 263.680 73.960 ;
        RECT 243.370 73.940 260.610 73.950 ;
        RECT 243.370 73.780 258.750 73.940 ;
        RECT 271.540 73.880 271.730 73.970 ;
        RECT 272.930 73.960 276.550 73.970 ;
        RECT 243.370 73.710 258.480 73.780 ;
        RECT 256.370 73.660 256.670 73.710 ;
        RECT 305.820 72.120 306.270 75.570 ;
        RECT 344.670 75.330 344.860 81.300 ;
        RECT 344.670 75.300 344.920 75.330 ;
        RECT 344.670 74.900 345.320 75.300 ;
        RECT 344.680 73.760 344.920 74.900 ;
        RECT 357.680 73.760 357.980 81.850 ;
        RECT 360.310 79.200 360.520 79.210 ;
        RECT 359.860 79.160 360.780 79.200 ;
        RECT 359.810 79.120 360.780 79.160 ;
        RECT 359.810 78.850 360.790 79.120 ;
        RECT 359.810 78.820 360.780 78.850 ;
        RECT 359.810 76.590 360.050 78.820 ;
        RECT 360.310 78.810 360.520 78.820 ;
        RECT 359.810 75.440 360.060 76.590 ;
        RECT 359.820 73.990 360.060 75.440 ;
        RECT 372.850 74.070 373.040 101.710 ;
        RECT 392.460 97.180 392.910 101.710 ;
        RECT 423.720 98.390 424.290 110.960 ;
        RECT 423.720 97.820 424.360 98.390 ;
        RECT 392.460 97.120 407.280 97.180 ;
        RECT 392.460 96.660 407.580 97.120 ;
        RECT 407.130 96.010 407.580 96.660 ;
        RECT 423.750 96.010 424.360 97.820 ;
        RECT 407.130 95.480 424.360 96.010 ;
        RECT 377.570 88.150 378.620 88.170 ;
        RECT 377.560 87.650 378.620 88.150 ;
        RECT 377.560 86.900 377.880 87.650 ;
        RECT 377.560 85.330 377.870 86.900 ;
        RECT 377.530 74.430 377.890 85.330 ;
        RECT 407.130 75.640 407.580 95.480 ;
        RECT 423.750 95.340 424.360 95.480 ;
        RECT 409.850 75.640 410.210 75.950 ;
        RECT 407.110 75.380 410.210 75.640 ;
        RECT 365.770 74.060 374.540 74.070 ;
        RECT 377.530 74.060 377.860 74.430 ;
        RECT 365.770 74.010 377.860 74.060 ;
        RECT 364.910 74.000 377.860 74.010 ;
        RECT 361.890 73.990 377.860 74.000 ;
        RECT 359.820 73.780 377.860 73.990 ;
        RECT 359.820 73.770 365.980 73.780 ;
        RECT 359.820 73.760 364.990 73.770 ;
        RECT 344.680 73.750 361.920 73.760 ;
        RECT 344.680 73.590 360.060 73.750 ;
        RECT 372.850 73.690 373.040 73.780 ;
        RECT 374.240 73.770 377.860 73.780 ;
        RECT 344.680 73.520 359.790 73.590 ;
        RECT 357.680 73.470 357.980 73.520 ;
        RECT 6.680 66.120 7.160 66.520 ;
        RECT 6.680 60.150 6.870 66.120 ;
        RECT 22.320 64.020 22.530 64.030 ;
        RECT 21.870 63.980 22.790 64.020 ;
        RECT 21.820 63.940 22.790 63.980 ;
        RECT 21.820 63.670 22.800 63.940 ;
        RECT 21.820 63.640 22.790 63.670 ;
        RECT 21.820 61.410 22.060 63.640 ;
        RECT 22.320 63.630 22.530 63.640 ;
        RECT 21.820 60.260 22.070 61.410 ;
        RECT 6.680 60.120 6.930 60.150 ;
        RECT 6.680 59.720 7.330 60.120 ;
        RECT 6.690 58.580 6.930 59.720 ;
        RECT 19.550 58.580 19.800 58.630 ;
        RECT 21.830 58.580 22.070 60.260 ;
        RECT 6.690 58.410 22.070 58.580 ;
        RECT 39.410 58.550 40.460 58.570 ;
        RECT 6.690 58.340 21.800 58.410 ;
        RECT 19.550 52.250 19.800 58.340 ;
        RECT 39.400 58.050 40.460 58.550 ;
        RECT 39.400 57.300 39.720 58.050 ;
        RECT 39.400 55.730 39.710 57.300 ;
        RECT 6.510 51.700 6.990 52.100 ;
        RECT 6.510 45.730 6.700 51.700 ;
        RECT 6.510 45.700 6.760 45.730 ;
        RECT 6.510 45.300 7.160 45.700 ;
        RECT 6.520 44.160 6.760 45.300 ;
        RECT 19.520 44.160 19.820 52.250 ;
        RECT 22.150 49.600 22.360 49.610 ;
        RECT 21.700 49.560 22.620 49.600 ;
        RECT 21.650 49.520 22.620 49.560 ;
        RECT 21.650 49.250 22.630 49.520 ;
        RECT 21.650 49.220 22.620 49.250 ;
        RECT 21.650 46.990 21.890 49.220 ;
        RECT 22.150 49.210 22.360 49.220 ;
        RECT 21.650 45.840 21.900 46.990 ;
        RECT 21.660 44.390 21.900 45.840 ;
        RECT 39.370 44.830 39.730 55.730 ;
        RECT 69.260 49.530 69.710 71.770 ;
        RECT 170.570 71.580 171.050 71.990 ;
        RECT 305.790 71.710 306.270 72.120 ;
        RECT 407.130 71.930 407.580 75.380 ;
        RECT 107.990 65.930 108.470 66.330 ;
        RECT 107.990 59.960 108.180 65.930 ;
        RECT 123.630 63.830 123.840 63.840 ;
        RECT 123.180 63.790 124.100 63.830 ;
        RECT 123.130 63.750 124.100 63.790 ;
        RECT 123.130 63.480 124.110 63.750 ;
        RECT 123.130 63.450 124.100 63.480 ;
        RECT 123.130 61.220 123.370 63.450 ;
        RECT 123.630 63.440 123.840 63.450 ;
        RECT 123.130 60.070 123.380 61.220 ;
        RECT 107.990 59.930 108.240 59.960 ;
        RECT 107.990 59.530 108.640 59.930 ;
        RECT 108.000 58.390 108.240 59.530 ;
        RECT 120.860 58.390 121.110 58.440 ;
        RECT 123.140 58.390 123.380 60.070 ;
        RECT 108.000 58.220 123.380 58.390 ;
        RECT 140.720 58.360 141.770 58.380 ;
        RECT 108.000 58.150 123.110 58.220 ;
        RECT 120.860 52.060 121.110 58.150 ;
        RECT 140.710 57.860 141.770 58.360 ;
        RECT 140.710 57.110 141.030 57.860 ;
        RECT 140.710 55.540 141.020 57.110 ;
        RECT 107.820 51.510 108.300 51.910 ;
        RECT 69.260 49.310 69.740 49.530 ;
        RECT 27.610 44.460 36.380 44.470 ;
        RECT 39.370 44.460 39.700 44.830 ;
        RECT 27.610 44.410 39.700 44.460 ;
        RECT 26.750 44.400 39.700 44.410 ;
        RECT 23.730 44.390 39.700 44.400 ;
        RECT 21.660 44.180 39.700 44.390 ;
        RECT 21.660 44.170 27.820 44.180 ;
        RECT 21.660 44.160 26.830 44.170 ;
        RECT 6.520 44.150 23.760 44.160 ;
        RECT 6.520 43.990 21.900 44.150 ;
        RECT 6.520 43.920 21.630 43.990 ;
        RECT 19.520 43.870 19.820 43.920 ;
        RECT 34.660 42.280 34.850 44.180 ;
        RECT 36.080 44.170 39.700 44.180 ;
        RECT 56.110 42.280 56.520 42.290 ;
        RECT 57.450 42.280 57.820 42.400 ;
        RECT 34.660 42.040 57.820 42.280 ;
        RECT 6.650 36.050 7.130 36.450 ;
        RECT 6.650 30.080 6.840 36.050 ;
        RECT 22.290 33.950 22.500 33.960 ;
        RECT 21.840 33.910 22.760 33.950 ;
        RECT 21.790 33.870 22.760 33.910 ;
        RECT 21.790 33.600 22.770 33.870 ;
        RECT 21.790 33.570 22.760 33.600 ;
        RECT 21.790 31.340 22.030 33.570 ;
        RECT 22.290 33.560 22.500 33.570 ;
        RECT 21.790 30.190 22.040 31.340 ;
        RECT 6.650 30.050 6.900 30.080 ;
        RECT 6.650 29.650 7.300 30.050 ;
        RECT 6.660 28.510 6.900 29.650 ;
        RECT 19.520 28.510 19.770 28.560 ;
        RECT 21.800 28.510 22.040 30.190 ;
        RECT 6.660 28.340 22.040 28.510 ;
        RECT 6.660 28.270 21.770 28.340 ;
        RECT 19.520 22.180 19.770 28.270 ;
        RECT 6.480 21.630 6.960 22.030 ;
        RECT 6.480 15.660 6.670 21.630 ;
        RECT 6.480 15.630 6.730 15.660 ;
        RECT 6.480 15.230 7.130 15.630 ;
        RECT 6.490 14.090 6.730 15.230 ;
        RECT 19.490 14.090 19.790 22.180 ;
        RECT 22.120 19.530 22.330 19.540 ;
        RECT 21.670 19.490 22.590 19.530 ;
        RECT 21.620 19.450 22.590 19.490 ;
        RECT 21.620 19.180 22.600 19.450 ;
        RECT 21.620 19.150 22.590 19.180 ;
        RECT 21.620 16.920 21.860 19.150 ;
        RECT 22.120 19.140 22.330 19.150 ;
        RECT 21.620 15.770 21.870 16.920 ;
        RECT 21.630 14.320 21.870 15.770 ;
        RECT 34.660 14.400 34.850 42.040 ;
        RECT 56.110 38.380 56.520 42.040 ;
        RECT 56.040 38.360 64.120 38.380 ;
        RECT 69.290 38.360 69.740 49.310 ;
        RECT 107.820 45.540 108.010 51.510 ;
        RECT 107.820 45.510 108.070 45.540 ;
        RECT 107.820 45.110 108.470 45.510 ;
        RECT 107.830 43.970 108.070 45.110 ;
        RECT 120.830 43.970 121.130 52.060 ;
        RECT 123.460 49.410 123.670 49.420 ;
        RECT 123.010 49.370 123.930 49.410 ;
        RECT 122.960 49.330 123.930 49.370 ;
        RECT 122.960 49.060 123.940 49.330 ;
        RECT 122.960 49.030 123.930 49.060 ;
        RECT 122.960 46.800 123.200 49.030 ;
        RECT 123.460 49.020 123.670 49.030 ;
        RECT 122.960 45.650 123.210 46.800 ;
        RECT 122.970 44.200 123.210 45.650 ;
        RECT 140.680 44.640 141.040 55.540 ;
        RECT 170.570 49.340 171.020 71.580 ;
        RECT 243.210 66.060 243.690 66.460 ;
        RECT 243.210 60.090 243.400 66.060 ;
        RECT 258.850 63.960 259.060 63.970 ;
        RECT 258.400 63.920 259.320 63.960 ;
        RECT 258.350 63.880 259.320 63.920 ;
        RECT 258.350 63.610 259.330 63.880 ;
        RECT 258.350 63.580 259.320 63.610 ;
        RECT 258.350 61.350 258.590 63.580 ;
        RECT 258.850 63.570 259.060 63.580 ;
        RECT 258.350 60.200 258.600 61.350 ;
        RECT 243.210 60.060 243.460 60.090 ;
        RECT 243.210 59.660 243.860 60.060 ;
        RECT 243.220 58.520 243.460 59.660 ;
        RECT 256.080 58.520 256.330 58.570 ;
        RECT 258.360 58.520 258.600 60.200 ;
        RECT 243.220 58.350 258.600 58.520 ;
        RECT 275.940 58.490 276.990 58.510 ;
        RECT 243.220 58.280 258.330 58.350 ;
        RECT 256.080 52.190 256.330 58.280 ;
        RECT 275.930 57.990 276.990 58.490 ;
        RECT 275.930 57.240 276.250 57.990 ;
        RECT 275.930 55.670 276.240 57.240 ;
        RECT 243.040 51.640 243.520 52.040 ;
        RECT 170.570 49.120 171.050 49.340 ;
        RECT 128.920 44.270 137.690 44.280 ;
        RECT 140.680 44.270 141.010 44.640 ;
        RECT 128.920 44.220 141.010 44.270 ;
        RECT 128.060 44.210 141.010 44.220 ;
        RECT 125.040 44.200 141.010 44.210 ;
        RECT 122.970 43.990 141.010 44.200 ;
        RECT 122.970 43.980 129.130 43.990 ;
        RECT 122.970 43.970 128.140 43.980 ;
        RECT 107.830 43.960 125.070 43.970 ;
        RECT 107.830 43.800 123.210 43.960 ;
        RECT 107.830 43.730 122.940 43.800 ;
        RECT 120.830 43.680 121.130 43.730 ;
        RECT 135.970 42.090 136.160 43.990 ;
        RECT 137.390 43.980 141.010 43.990 ;
        RECT 157.420 42.090 157.830 42.100 ;
        RECT 158.760 42.090 159.130 42.210 ;
        RECT 135.970 41.850 159.130 42.090 ;
        RECT 56.040 38.010 69.750 38.360 ;
        RECT 56.110 37.990 56.520 38.010 ;
        RECT 62.860 37.990 69.750 38.010 ;
        RECT 69.290 37.930 69.740 37.990 ;
        RECT 107.960 35.860 108.440 36.260 ;
        RECT 107.960 29.890 108.150 35.860 ;
        RECT 123.600 33.760 123.810 33.770 ;
        RECT 123.150 33.720 124.070 33.760 ;
        RECT 123.100 33.680 124.070 33.720 ;
        RECT 123.100 33.410 124.080 33.680 ;
        RECT 123.100 33.380 124.070 33.410 ;
        RECT 123.100 31.150 123.340 33.380 ;
        RECT 123.600 33.370 123.810 33.380 ;
        RECT 123.100 30.000 123.350 31.150 ;
        RECT 107.960 29.860 108.210 29.890 ;
        RECT 107.960 29.460 108.610 29.860 ;
        RECT 39.380 28.480 40.430 28.500 ;
        RECT 39.370 27.980 40.430 28.480 ;
        RECT 107.970 28.320 108.210 29.460 ;
        RECT 120.830 28.320 121.080 28.370 ;
        RECT 123.110 28.320 123.350 30.000 ;
        RECT 107.970 28.150 123.350 28.320 ;
        RECT 107.970 28.080 123.080 28.150 ;
        RECT 39.370 27.230 39.690 27.980 ;
        RECT 39.370 25.660 39.680 27.230 ;
        RECT 39.340 14.760 39.700 25.660 ;
        RECT 120.830 21.990 121.080 28.080 ;
        RECT 107.790 21.440 108.270 21.840 ;
        RECT 107.790 15.470 107.980 21.440 ;
        RECT 107.790 15.440 108.040 15.470 ;
        RECT 107.790 15.040 108.440 15.440 ;
        RECT 27.580 14.390 36.350 14.400 ;
        RECT 39.340 14.390 39.670 14.760 ;
        RECT 27.580 14.340 39.670 14.390 ;
        RECT 26.720 14.330 39.670 14.340 ;
        RECT 23.700 14.320 39.670 14.330 ;
        RECT 21.630 14.110 39.670 14.320 ;
        RECT 21.630 14.100 27.790 14.110 ;
        RECT 21.630 14.090 26.800 14.100 ;
        RECT 6.490 14.080 23.730 14.090 ;
        RECT 6.490 13.920 21.870 14.080 ;
        RECT 34.660 14.020 34.850 14.110 ;
        RECT 36.050 14.100 39.670 14.110 ;
        RECT 6.490 13.850 21.600 13.920 ;
        RECT 107.800 13.900 108.040 15.040 ;
        RECT 120.800 13.900 121.100 21.990 ;
        RECT 123.430 19.340 123.640 19.350 ;
        RECT 122.980 19.300 123.900 19.340 ;
        RECT 122.930 19.260 123.900 19.300 ;
        RECT 122.930 18.990 123.910 19.260 ;
        RECT 122.930 18.960 123.900 18.990 ;
        RECT 122.930 16.730 123.170 18.960 ;
        RECT 123.430 18.950 123.640 18.960 ;
        RECT 122.930 15.580 123.180 16.730 ;
        RECT 122.940 14.130 123.180 15.580 ;
        RECT 135.970 14.210 136.160 41.850 ;
        RECT 157.420 38.190 157.830 41.850 ;
        RECT 157.350 38.170 165.430 38.190 ;
        RECT 170.600 38.170 171.050 49.120 ;
        RECT 243.040 45.670 243.230 51.640 ;
        RECT 243.040 45.640 243.290 45.670 ;
        RECT 243.040 45.240 243.690 45.640 ;
        RECT 243.050 44.100 243.290 45.240 ;
        RECT 256.050 44.100 256.350 52.190 ;
        RECT 258.680 49.540 258.890 49.550 ;
        RECT 258.230 49.500 259.150 49.540 ;
        RECT 258.180 49.460 259.150 49.500 ;
        RECT 258.180 49.190 259.160 49.460 ;
        RECT 258.180 49.160 259.150 49.190 ;
        RECT 258.180 46.930 258.420 49.160 ;
        RECT 258.680 49.150 258.890 49.160 ;
        RECT 258.180 45.780 258.430 46.930 ;
        RECT 258.190 44.330 258.430 45.780 ;
        RECT 275.900 44.770 276.260 55.670 ;
        RECT 305.790 49.470 306.240 71.710 ;
        RECT 407.100 71.520 407.580 71.930 ;
        RECT 344.520 65.870 345.000 66.270 ;
        RECT 344.520 59.900 344.710 65.870 ;
        RECT 360.160 63.770 360.370 63.780 ;
        RECT 359.710 63.730 360.630 63.770 ;
        RECT 359.660 63.690 360.630 63.730 ;
        RECT 359.660 63.420 360.640 63.690 ;
        RECT 359.660 63.390 360.630 63.420 ;
        RECT 359.660 61.160 359.900 63.390 ;
        RECT 360.160 63.380 360.370 63.390 ;
        RECT 359.660 60.010 359.910 61.160 ;
        RECT 344.520 59.870 344.770 59.900 ;
        RECT 344.520 59.470 345.170 59.870 ;
        RECT 344.530 58.330 344.770 59.470 ;
        RECT 357.390 58.330 357.640 58.380 ;
        RECT 359.670 58.330 359.910 60.010 ;
        RECT 344.530 58.160 359.910 58.330 ;
        RECT 377.250 58.300 378.300 58.320 ;
        RECT 344.530 58.090 359.640 58.160 ;
        RECT 357.390 52.000 357.640 58.090 ;
        RECT 377.240 57.800 378.300 58.300 ;
        RECT 377.240 57.050 377.560 57.800 ;
        RECT 377.240 55.480 377.550 57.050 ;
        RECT 344.350 51.450 344.830 51.850 ;
        RECT 305.790 49.250 306.270 49.470 ;
        RECT 264.140 44.400 272.910 44.410 ;
        RECT 275.900 44.400 276.230 44.770 ;
        RECT 264.140 44.350 276.230 44.400 ;
        RECT 263.280 44.340 276.230 44.350 ;
        RECT 260.260 44.330 276.230 44.340 ;
        RECT 258.190 44.120 276.230 44.330 ;
        RECT 258.190 44.110 264.350 44.120 ;
        RECT 258.190 44.100 263.360 44.110 ;
        RECT 243.050 44.090 260.290 44.100 ;
        RECT 243.050 43.930 258.430 44.090 ;
        RECT 243.050 43.860 258.160 43.930 ;
        RECT 256.050 43.810 256.350 43.860 ;
        RECT 271.190 42.220 271.380 44.120 ;
        RECT 272.610 44.110 276.230 44.120 ;
        RECT 292.640 42.220 293.050 42.230 ;
        RECT 293.980 42.220 294.350 42.340 ;
        RECT 271.190 41.980 294.350 42.220 ;
        RECT 157.350 37.820 171.060 38.170 ;
        RECT 157.420 37.800 157.830 37.820 ;
        RECT 164.170 37.800 171.060 37.820 ;
        RECT 170.600 37.740 171.050 37.800 ;
        RECT 243.180 35.990 243.660 36.390 ;
        RECT 243.180 30.020 243.370 35.990 ;
        RECT 258.820 33.890 259.030 33.900 ;
        RECT 258.370 33.850 259.290 33.890 ;
        RECT 258.320 33.810 259.290 33.850 ;
        RECT 258.320 33.540 259.300 33.810 ;
        RECT 258.320 33.510 259.290 33.540 ;
        RECT 258.320 31.280 258.560 33.510 ;
        RECT 258.820 33.500 259.030 33.510 ;
        RECT 258.320 30.130 258.570 31.280 ;
        RECT 243.180 29.990 243.430 30.020 ;
        RECT 243.180 29.590 243.830 29.990 ;
        RECT 243.190 28.450 243.430 29.590 ;
        RECT 256.050 28.450 256.300 28.500 ;
        RECT 258.330 28.450 258.570 30.130 ;
        RECT 140.690 28.290 141.740 28.310 ;
        RECT 140.680 27.790 141.740 28.290 ;
        RECT 243.190 28.280 258.570 28.450 ;
        RECT 243.190 28.210 258.300 28.280 ;
        RECT 140.680 27.040 141.000 27.790 ;
        RECT 140.680 25.470 140.990 27.040 ;
        RECT 140.650 14.570 141.010 25.470 ;
        RECT 256.050 22.120 256.300 28.210 ;
        RECT 243.010 21.570 243.490 21.970 ;
        RECT 243.010 15.600 243.200 21.570 ;
        RECT 243.010 15.570 243.260 15.600 ;
        RECT 243.010 15.170 243.660 15.570 ;
        RECT 128.890 14.200 137.660 14.210 ;
        RECT 140.650 14.200 140.980 14.570 ;
        RECT 128.890 14.150 140.980 14.200 ;
        RECT 128.030 14.140 140.980 14.150 ;
        RECT 125.010 14.130 140.980 14.140 ;
        RECT 122.940 13.920 140.980 14.130 ;
        RECT 122.940 13.910 129.100 13.920 ;
        RECT 122.940 13.900 128.110 13.910 ;
        RECT 107.800 13.890 125.040 13.900 ;
        RECT 19.490 13.800 19.790 13.850 ;
        RECT 107.800 13.730 123.180 13.890 ;
        RECT 135.970 13.830 136.160 13.920 ;
        RECT 137.360 13.910 140.980 13.920 ;
        RECT 243.020 14.030 243.260 15.170 ;
        RECT 256.020 14.030 256.320 22.120 ;
        RECT 258.650 19.470 258.860 19.480 ;
        RECT 258.200 19.430 259.120 19.470 ;
        RECT 258.150 19.390 259.120 19.430 ;
        RECT 258.150 19.120 259.130 19.390 ;
        RECT 258.150 19.090 259.120 19.120 ;
        RECT 258.150 16.860 258.390 19.090 ;
        RECT 258.650 19.080 258.860 19.090 ;
        RECT 258.150 15.710 258.400 16.860 ;
        RECT 258.160 14.260 258.400 15.710 ;
        RECT 271.190 14.340 271.380 41.980 ;
        RECT 292.640 38.320 293.050 41.980 ;
        RECT 292.570 38.300 300.650 38.320 ;
        RECT 305.820 38.300 306.270 49.250 ;
        RECT 344.350 45.480 344.540 51.450 ;
        RECT 344.350 45.450 344.600 45.480 ;
        RECT 344.350 45.050 345.000 45.450 ;
        RECT 344.360 43.910 344.600 45.050 ;
        RECT 357.360 43.910 357.660 52.000 ;
        RECT 359.990 49.350 360.200 49.360 ;
        RECT 359.540 49.310 360.460 49.350 ;
        RECT 359.490 49.270 360.460 49.310 ;
        RECT 359.490 49.000 360.470 49.270 ;
        RECT 359.490 48.970 360.460 49.000 ;
        RECT 359.490 46.740 359.730 48.970 ;
        RECT 359.990 48.960 360.200 48.970 ;
        RECT 359.490 45.590 359.740 46.740 ;
        RECT 359.500 44.140 359.740 45.590 ;
        RECT 377.210 44.580 377.570 55.480 ;
        RECT 407.100 49.280 407.550 71.520 ;
        RECT 407.100 49.060 407.580 49.280 ;
        RECT 365.450 44.210 374.220 44.220 ;
        RECT 377.210 44.210 377.540 44.580 ;
        RECT 365.450 44.160 377.540 44.210 ;
        RECT 364.590 44.150 377.540 44.160 ;
        RECT 361.570 44.140 377.540 44.150 ;
        RECT 359.500 43.930 377.540 44.140 ;
        RECT 359.500 43.920 365.660 43.930 ;
        RECT 359.500 43.910 364.670 43.920 ;
        RECT 344.360 43.900 361.600 43.910 ;
        RECT 344.360 43.740 359.740 43.900 ;
        RECT 344.360 43.670 359.470 43.740 ;
        RECT 357.360 43.620 357.660 43.670 ;
        RECT 372.500 42.030 372.690 43.930 ;
        RECT 373.920 43.920 377.540 43.930 ;
        RECT 393.950 42.030 394.360 42.040 ;
        RECT 395.290 42.030 395.660 42.150 ;
        RECT 372.500 41.790 395.660 42.030 ;
        RECT 292.570 37.950 306.280 38.300 ;
        RECT 292.640 37.930 293.050 37.950 ;
        RECT 299.390 37.930 306.280 37.950 ;
        RECT 305.820 37.870 306.270 37.930 ;
        RECT 344.490 35.800 344.970 36.200 ;
        RECT 344.490 29.830 344.680 35.800 ;
        RECT 360.130 33.700 360.340 33.710 ;
        RECT 359.680 33.660 360.600 33.700 ;
        RECT 359.630 33.620 360.600 33.660 ;
        RECT 359.630 33.350 360.610 33.620 ;
        RECT 359.630 33.320 360.600 33.350 ;
        RECT 359.630 31.090 359.870 33.320 ;
        RECT 360.130 33.310 360.340 33.320 ;
        RECT 359.630 29.940 359.880 31.090 ;
        RECT 344.490 29.800 344.740 29.830 ;
        RECT 344.490 29.400 345.140 29.800 ;
        RECT 275.910 28.420 276.960 28.440 ;
        RECT 275.900 27.920 276.960 28.420 ;
        RECT 344.500 28.260 344.740 29.400 ;
        RECT 357.360 28.260 357.610 28.310 ;
        RECT 359.640 28.260 359.880 29.940 ;
        RECT 344.500 28.090 359.880 28.260 ;
        RECT 344.500 28.020 359.610 28.090 ;
        RECT 275.900 27.170 276.220 27.920 ;
        RECT 275.900 25.600 276.210 27.170 ;
        RECT 275.870 14.700 276.230 25.600 ;
        RECT 357.360 21.930 357.610 28.020 ;
        RECT 344.320 21.380 344.800 21.780 ;
        RECT 344.320 15.410 344.510 21.380 ;
        RECT 344.320 15.380 344.570 15.410 ;
        RECT 344.320 14.980 344.970 15.380 ;
        RECT 264.110 14.330 272.880 14.340 ;
        RECT 275.870 14.330 276.200 14.700 ;
        RECT 264.110 14.280 276.200 14.330 ;
        RECT 263.250 14.270 276.200 14.280 ;
        RECT 260.230 14.260 276.200 14.270 ;
        RECT 258.160 14.050 276.200 14.260 ;
        RECT 258.160 14.040 264.320 14.050 ;
        RECT 258.160 14.030 263.330 14.040 ;
        RECT 243.020 14.020 260.260 14.030 ;
        RECT 243.020 13.860 258.400 14.020 ;
        RECT 271.190 13.960 271.380 14.050 ;
        RECT 272.580 14.040 276.200 14.050 ;
        RECT 243.020 13.790 258.130 13.860 ;
        RECT 344.330 13.840 344.570 14.980 ;
        RECT 357.330 13.840 357.630 21.930 ;
        RECT 359.960 19.280 360.170 19.290 ;
        RECT 359.510 19.240 360.430 19.280 ;
        RECT 359.460 19.200 360.430 19.240 ;
        RECT 359.460 18.930 360.440 19.200 ;
        RECT 359.460 18.900 360.430 18.930 ;
        RECT 359.460 16.670 359.700 18.900 ;
        RECT 359.960 18.890 360.170 18.900 ;
        RECT 359.460 15.520 359.710 16.670 ;
        RECT 359.470 14.070 359.710 15.520 ;
        RECT 372.500 14.150 372.690 41.790 ;
        RECT 393.950 38.130 394.360 41.790 ;
        RECT 393.880 38.110 401.960 38.130 ;
        RECT 407.130 38.110 407.580 49.060 ;
        RECT 393.880 37.760 407.590 38.110 ;
        RECT 393.950 37.740 394.360 37.760 ;
        RECT 400.700 37.740 407.590 37.760 ;
        RECT 407.130 37.680 407.580 37.740 ;
        RECT 377.220 28.230 378.270 28.250 ;
        RECT 377.210 27.730 378.270 28.230 ;
        RECT 377.210 26.980 377.530 27.730 ;
        RECT 377.210 25.410 377.520 26.980 ;
        RECT 377.180 14.510 377.540 25.410 ;
        RECT 365.420 14.140 374.190 14.150 ;
        RECT 377.180 14.140 377.510 14.510 ;
        RECT 365.420 14.090 377.510 14.140 ;
        RECT 364.560 14.080 377.510 14.090 ;
        RECT 361.540 14.070 377.510 14.080 ;
        RECT 359.470 13.860 377.510 14.070 ;
        RECT 359.470 13.850 365.630 13.860 ;
        RECT 359.470 13.840 364.640 13.850 ;
        RECT 344.330 13.830 361.570 13.840 ;
        RECT 256.020 13.740 256.320 13.790 ;
        RECT 107.800 13.660 122.910 13.730 ;
        RECT 344.330 13.670 359.710 13.830 ;
        RECT 372.500 13.770 372.690 13.860 ;
        RECT 373.890 13.850 377.510 13.860 ;
        RECT 120.800 13.610 121.100 13.660 ;
        RECT 344.330 13.600 359.440 13.670 ;
        RECT 357.330 13.550 357.630 13.600 ;
      LAYER via2 ;
        RECT 55.250 254.250 55.530 254.530 ;
        RECT 55.560 254.250 55.840 254.530 ;
        RECT 55.860 254.250 56.140 254.530 ;
        RECT 56.170 254.250 56.450 254.530 ;
        RECT 56.495 254.250 56.775 254.530 ;
        RECT 56.805 254.250 57.085 254.530 ;
        RECT 57.105 254.250 57.385 254.530 ;
        RECT 57.415 254.250 57.695 254.530 ;
        RECT 57.760 254.250 58.040 254.530 ;
        RECT 58.070 254.250 58.350 254.530 ;
        RECT 58.370 254.250 58.650 254.530 ;
        RECT 58.680 254.250 58.960 254.530 ;
        RECT 59.005 254.250 59.285 254.530 ;
        RECT 59.315 254.250 59.595 254.530 ;
        RECT 59.615 254.250 59.895 254.530 ;
        RECT 59.925 254.250 60.205 254.530 ;
      LAYER met3 ;
        RECT 55.100 254.200 60.350 257.005 ;
      LAYER via3 ;
        RECT 59.415 256.915 60.090 256.920 ;
        RECT 59.090 256.910 60.090 256.915 ;
        RECT 58.700 256.905 60.090 256.910 ;
        RECT 58.045 256.900 60.090 256.905 ;
        RECT 57.365 256.895 60.090 256.900 ;
        RECT 57.040 256.890 60.090 256.895 ;
        RECT 56.650 256.885 60.090 256.890 ;
        RECT 55.970 256.880 60.090 256.885 ;
        RECT 55.250 256.600 60.090 256.880 ;
        RECT 55.250 256.535 60.085 256.600 ;
        RECT 55.245 256.255 60.085 256.535 ;
        RECT 55.245 256.200 60.080 256.255 ;
        RECT 55.240 255.920 60.080 256.200 ;
        RECT 55.240 255.915 59.400 255.920 ;
        RECT 55.240 255.910 59.010 255.915 ;
        RECT 55.240 255.905 58.685 255.910 ;
        RECT 55.240 255.900 58.030 255.905 ;
        RECT 55.240 255.895 57.350 255.900 ;
        RECT 55.240 255.890 56.960 255.895 ;
        RECT 55.240 255.885 56.635 255.890 ;
        RECT 55.240 255.880 55.955 255.885 ;
      LAYER met4 ;
        RECT 55.030 255.695 60.350 276.250 ;
    END
  END gnd
  OBS
      LAYER nwell ;
        RECT 12.880 250.740 13.730 250.850 ;
      LAYER pwell ;
        RECT 3.100 248.270 4.000 249.210 ;
      LAYER nwell ;
        RECT 12.660 248.510 14.570 250.740 ;
        RECT 249.410 250.680 250.260 250.790 ;
        RECT 114.190 250.550 115.040 250.660 ;
      LAYER pwell ;
        RECT 16.300 249.210 17.610 250.070 ;
        RECT 3.090 248.010 4.000 248.270 ;
        RECT 3.090 247.110 3.990 248.010 ;
        RECT 3.060 246.030 3.960 246.970 ;
        RECT 13.000 246.810 14.310 247.670 ;
      LAYER nwell ;
        RECT 15.910 246.100 17.830 248.360 ;
        RECT 28.560 248.320 29.410 248.430 ;
      LAYER pwell ;
        RECT 3.050 245.770 3.960 246.030 ;
      LAYER nwell ;
        RECT 16.880 246.010 17.730 246.100 ;
        RECT 28.340 246.090 30.250 248.320 ;
      LAYER pwell ;
        RECT 104.410 248.080 105.310 249.020 ;
      LAYER nwell ;
        RECT 113.970 248.320 115.880 250.550 ;
      LAYER pwell ;
        RECT 117.610 249.020 118.920 249.880 ;
        RECT 104.400 247.820 105.310 248.080 ;
        RECT 31.980 246.790 33.290 247.650 ;
        RECT 104.400 246.920 105.300 247.820 ;
        RECT 3.050 244.870 3.950 245.770 ;
      LAYER nwell ;
        RECT 13.040 244.340 13.890 244.450 ;
      LAYER pwell ;
        RECT 28.680 244.390 29.990 245.250 ;
        RECT 3.060 242.870 3.960 243.810 ;
        RECT 3.050 242.610 3.960 242.870 ;
        RECT 3.050 241.710 3.950 242.610 ;
      LAYER nwell ;
        RECT 12.820 242.110 14.730 244.340 ;
        RECT 31.590 243.680 33.510 245.940 ;
      LAYER pwell ;
        RECT 104.370 245.840 105.270 246.780 ;
        RECT 114.310 246.620 115.620 247.480 ;
      LAYER nwell ;
        RECT 117.220 245.910 119.140 248.170 ;
        RECT 129.870 248.130 130.720 248.240 ;
      LAYER pwell ;
        RECT 239.630 248.210 240.530 249.150 ;
      LAYER nwell ;
        RECT 249.190 248.450 251.100 250.680 ;
        RECT 350.720 250.490 351.570 250.600 ;
      LAYER pwell ;
        RECT 252.830 249.150 254.140 250.010 ;
        RECT 104.360 245.580 105.270 245.840 ;
      LAYER nwell ;
        RECT 118.190 245.820 119.040 245.910 ;
        RECT 129.650 245.900 131.560 248.130 ;
      LAYER pwell ;
        RECT 239.620 247.950 240.530 248.210 ;
        RECT 133.290 246.600 134.600 247.460 ;
        RECT 239.620 247.050 240.520 247.950 ;
        RECT 239.590 245.970 240.490 246.910 ;
        RECT 249.530 246.750 250.840 247.610 ;
      LAYER nwell ;
        RECT 252.440 246.040 254.360 248.300 ;
        RECT 265.090 248.260 265.940 248.370 ;
      LAYER pwell ;
        RECT 104.360 244.680 105.260 245.580 ;
      LAYER nwell ;
        RECT 114.350 244.150 115.200 244.260 ;
      LAYER pwell ;
        RECT 129.990 244.200 131.300 245.060 ;
        RECT 16.460 242.810 17.770 243.670 ;
      LAYER nwell ;
        RECT 32.560 243.590 33.410 243.680 ;
        RECT 46.140 242.770 46.990 242.880 ;
      LAYER pwell ;
        RECT 3.320 239.460 4.220 240.990 ;
        RECT 13.160 240.410 14.470 241.270 ;
      LAYER nwell ;
        RECT 16.070 239.700 17.990 241.960 ;
        RECT 45.920 240.540 47.830 242.770 ;
      LAYER pwell ;
        RECT 104.370 242.680 105.270 243.620 ;
        RECT 104.360 242.420 105.270 242.680 ;
        RECT 49.560 241.240 50.870 242.100 ;
        RECT 104.360 241.520 105.260 242.420 ;
      LAYER nwell ;
        RECT 114.130 241.920 116.040 244.150 ;
        RECT 132.900 243.490 134.820 245.750 ;
      LAYER pwell ;
        RECT 239.580 245.710 240.490 245.970 ;
      LAYER nwell ;
        RECT 253.410 245.950 254.260 246.040 ;
        RECT 264.870 246.030 266.780 248.260 ;
      LAYER pwell ;
        RECT 340.940 248.020 341.840 248.960 ;
      LAYER nwell ;
        RECT 350.500 248.260 352.410 250.490 ;
      LAYER pwell ;
        RECT 354.140 248.960 355.450 249.820 ;
        RECT 340.930 247.760 341.840 248.020 ;
        RECT 268.510 246.730 269.820 247.590 ;
        RECT 340.930 246.860 341.830 247.760 ;
        RECT 239.580 244.810 240.480 245.710 ;
      LAYER nwell ;
        RECT 249.570 244.280 250.420 244.390 ;
      LAYER pwell ;
        RECT 265.210 244.330 266.520 245.190 ;
        RECT 117.770 242.620 119.080 243.480 ;
      LAYER nwell ;
        RECT 133.870 243.400 134.720 243.490 ;
      LAYER pwell ;
        RECT 239.590 242.810 240.490 243.750 ;
      LAYER nwell ;
        RECT 147.450 242.580 148.300 242.690 ;
        RECT 17.040 239.610 17.890 239.700 ;
      LAYER pwell ;
        RECT 3.320 239.450 3.740 239.460 ;
        RECT 46.260 238.840 47.570 239.700 ;
      LAYER nwell ;
        RECT 49.170 238.130 51.090 240.390 ;
      LAYER pwell ;
        RECT 104.630 239.270 105.530 240.800 ;
        RECT 114.470 240.220 115.780 241.080 ;
      LAYER nwell ;
        RECT 117.380 239.510 119.300 241.770 ;
        RECT 147.230 240.350 149.140 242.580 ;
      LAYER pwell ;
        RECT 239.580 242.550 240.490 242.810 ;
        RECT 150.870 241.050 152.180 241.910 ;
        RECT 239.580 241.650 240.480 242.550 ;
      LAYER nwell ;
        RECT 249.350 242.050 251.260 244.280 ;
        RECT 268.120 243.620 270.040 245.880 ;
      LAYER pwell ;
        RECT 340.900 245.780 341.800 246.720 ;
        RECT 350.840 246.560 352.150 247.420 ;
      LAYER nwell ;
        RECT 353.750 245.850 355.670 248.110 ;
        RECT 366.400 248.070 367.250 248.180 ;
      LAYER pwell ;
        RECT 340.890 245.520 341.800 245.780 ;
      LAYER nwell ;
        RECT 354.720 245.760 355.570 245.850 ;
        RECT 366.180 245.840 368.090 248.070 ;
      LAYER pwell ;
        RECT 369.820 246.540 371.130 247.400 ;
        RECT 340.890 244.620 341.790 245.520 ;
      LAYER nwell ;
        RECT 350.880 244.090 351.730 244.200 ;
      LAYER pwell ;
        RECT 366.520 244.140 367.830 245.000 ;
        RECT 252.990 242.750 254.300 243.610 ;
      LAYER nwell ;
        RECT 269.090 243.530 269.940 243.620 ;
        RECT 282.670 242.710 283.520 242.820 ;
        RECT 118.350 239.420 119.200 239.510 ;
      LAYER pwell ;
        RECT 104.630 239.260 105.050 239.270 ;
        RECT 147.570 238.650 148.880 239.510 ;
      LAYER nwell ;
        RECT 50.140 238.040 50.990 238.130 ;
      LAYER pwell ;
        RECT 3.050 236.420 3.950 237.950 ;
      LAYER nwell ;
        RECT 150.480 237.940 152.400 240.200 ;
      LAYER pwell ;
        RECT 239.850 239.400 240.750 240.930 ;
        RECT 249.690 240.350 251.000 241.210 ;
      LAYER nwell ;
        RECT 252.600 239.640 254.520 241.900 ;
        RECT 282.450 240.480 284.360 242.710 ;
      LAYER pwell ;
        RECT 340.900 242.620 341.800 243.560 ;
        RECT 340.890 242.360 341.800 242.620 ;
        RECT 286.090 241.180 287.400 242.040 ;
        RECT 340.890 241.460 341.790 242.360 ;
      LAYER nwell ;
        RECT 350.660 241.860 352.570 244.090 ;
        RECT 369.430 243.430 371.350 245.690 ;
      LAYER pwell ;
        RECT 354.300 242.560 355.610 243.420 ;
      LAYER nwell ;
        RECT 370.400 243.340 371.250 243.430 ;
        RECT 383.980 242.520 384.830 242.630 ;
        RECT 253.570 239.550 254.420 239.640 ;
      LAYER pwell ;
        RECT 239.850 239.390 240.270 239.400 ;
        RECT 282.790 238.780 284.100 239.640 ;
      LAYER nwell ;
        RECT 285.700 238.070 287.620 240.330 ;
      LAYER pwell ;
        RECT 341.160 239.210 342.060 240.740 ;
        RECT 351.000 240.160 352.310 241.020 ;
      LAYER nwell ;
        RECT 353.910 239.450 355.830 241.710 ;
        RECT 383.760 240.290 385.670 242.520 ;
      LAYER pwell ;
        RECT 387.400 240.990 388.710 241.850 ;
      LAYER nwell ;
        RECT 354.880 239.360 355.730 239.450 ;
      LAYER pwell ;
        RECT 341.160 239.200 341.580 239.210 ;
        RECT 384.100 238.590 385.410 239.450 ;
      LAYER nwell ;
        RECT 286.670 237.980 287.520 238.070 ;
        RECT 151.450 237.850 152.300 237.940 ;
      LAYER pwell ;
        RECT 3.050 236.410 3.470 236.420 ;
      LAYER nwell ;
        RECT 12.710 236.320 13.560 236.430 ;
      LAYER pwell ;
        RECT 2.930 233.850 3.830 234.790 ;
      LAYER nwell ;
        RECT 12.490 234.090 14.400 236.320 ;
      LAYER pwell ;
        RECT 104.360 236.230 105.260 237.760 ;
        RECT 239.580 236.360 240.480 237.890 ;
      LAYER nwell ;
        RECT 387.010 237.880 388.930 240.140 ;
        RECT 387.980 237.790 388.830 237.880 ;
      LAYER pwell ;
        RECT 239.580 236.350 240.000 236.360 ;
      LAYER nwell ;
        RECT 249.240 236.260 250.090 236.370 ;
      LAYER pwell ;
        RECT 104.360 236.220 104.780 236.230 ;
      LAYER nwell ;
        RECT 114.020 236.130 114.870 236.240 ;
      LAYER pwell ;
        RECT 16.130 234.790 17.440 235.650 ;
        RECT 2.920 233.590 3.830 233.850 ;
        RECT 2.920 232.690 3.820 233.590 ;
        RECT 2.890 231.610 3.790 232.550 ;
        RECT 12.830 232.390 14.140 233.250 ;
      LAYER nwell ;
        RECT 15.740 231.680 17.660 233.940 ;
        RECT 28.390 233.900 29.240 234.010 ;
      LAYER pwell ;
        RECT 2.880 231.350 3.790 231.610 ;
      LAYER nwell ;
        RECT 16.710 231.590 17.560 231.680 ;
        RECT 28.170 231.670 30.080 233.900 ;
      LAYER pwell ;
        RECT 104.240 233.660 105.140 234.600 ;
      LAYER nwell ;
        RECT 113.800 233.900 115.710 236.130 ;
      LAYER pwell ;
        RECT 117.440 234.600 118.750 235.460 ;
        RECT 104.230 233.400 105.140 233.660 ;
        RECT 31.810 232.370 33.120 233.230 ;
        RECT 104.230 232.500 105.130 233.400 ;
        RECT 2.880 230.450 3.780 231.350 ;
      LAYER nwell ;
        RECT 12.870 229.920 13.720 230.030 ;
      LAYER pwell ;
        RECT 28.510 229.970 29.820 230.830 ;
        RECT 2.890 228.450 3.790 229.390 ;
        RECT 2.880 228.190 3.790 228.450 ;
        RECT 2.880 227.290 3.780 228.190 ;
      LAYER nwell ;
        RECT 12.650 227.690 14.560 229.920 ;
        RECT 31.420 229.260 33.340 231.520 ;
      LAYER pwell ;
        RECT 104.200 231.420 105.100 232.360 ;
        RECT 114.140 232.200 115.450 233.060 ;
      LAYER nwell ;
        RECT 117.050 231.490 118.970 233.750 ;
        RECT 129.700 233.710 130.550 233.820 ;
      LAYER pwell ;
        RECT 239.460 233.790 240.360 234.730 ;
      LAYER nwell ;
        RECT 249.020 234.030 250.930 236.260 ;
      LAYER pwell ;
        RECT 340.890 236.170 341.790 237.700 ;
        RECT 340.890 236.160 341.310 236.170 ;
      LAYER nwell ;
        RECT 350.550 236.070 351.400 236.180 ;
      LAYER pwell ;
        RECT 252.660 234.730 253.970 235.590 ;
        RECT 104.190 231.160 105.100 231.420 ;
      LAYER nwell ;
        RECT 118.020 231.400 118.870 231.490 ;
        RECT 129.480 231.480 131.390 233.710 ;
      LAYER pwell ;
        RECT 239.450 233.530 240.360 233.790 ;
        RECT 133.120 232.180 134.430 233.040 ;
        RECT 239.450 232.630 240.350 233.530 ;
        RECT 239.420 231.550 240.320 232.490 ;
        RECT 249.360 232.330 250.670 233.190 ;
      LAYER nwell ;
        RECT 252.270 231.620 254.190 233.880 ;
        RECT 264.920 233.840 265.770 233.950 ;
      LAYER pwell ;
        RECT 104.190 230.260 105.090 231.160 ;
      LAYER nwell ;
        RECT 114.180 229.730 115.030 229.840 ;
      LAYER pwell ;
        RECT 129.820 229.780 131.130 230.640 ;
        RECT 16.290 228.390 17.600 229.250 ;
      LAYER nwell ;
        RECT 32.390 229.170 33.240 229.260 ;
      LAYER pwell ;
        RECT 104.200 228.260 105.100 229.200 ;
        RECT 104.190 228.000 105.100 228.260 ;
        RECT 3.150 225.040 4.050 226.570 ;
        RECT 12.990 225.990 14.300 226.850 ;
      LAYER nwell ;
        RECT 15.900 225.280 17.820 227.540 ;
      LAYER pwell ;
        RECT 104.190 227.100 105.090 228.000 ;
      LAYER nwell ;
        RECT 113.960 227.500 115.870 229.730 ;
        RECT 132.730 229.070 134.650 231.330 ;
      LAYER pwell ;
        RECT 239.410 231.290 240.320 231.550 ;
      LAYER nwell ;
        RECT 253.240 231.530 254.090 231.620 ;
        RECT 264.700 231.610 266.610 233.840 ;
      LAYER pwell ;
        RECT 340.770 233.600 341.670 234.540 ;
      LAYER nwell ;
        RECT 350.330 233.840 352.240 236.070 ;
      LAYER pwell ;
        RECT 353.970 234.540 355.280 235.400 ;
        RECT 340.760 233.340 341.670 233.600 ;
        RECT 268.340 232.310 269.650 233.170 ;
        RECT 340.760 232.440 341.660 233.340 ;
        RECT 239.410 230.390 240.310 231.290 ;
      LAYER nwell ;
        RECT 249.400 229.860 250.250 229.970 ;
      LAYER pwell ;
        RECT 265.040 229.910 266.350 230.770 ;
        RECT 117.600 228.200 118.910 229.060 ;
      LAYER nwell ;
        RECT 133.700 228.980 134.550 229.070 ;
      LAYER pwell ;
        RECT 239.420 228.390 240.320 229.330 ;
        RECT 239.410 228.130 240.320 228.390 ;
      LAYER nwell ;
        RECT 63.670 226.750 64.520 226.860 ;
        RECT 16.870 225.190 17.720 225.280 ;
      LAYER pwell ;
        RECT 3.150 225.030 3.570 225.040 ;
      LAYER nwell ;
        RECT 63.450 224.520 65.360 226.750 ;
      LAYER pwell ;
        RECT 67.090 225.220 68.400 226.080 ;
        RECT 104.460 224.850 105.360 226.380 ;
        RECT 114.300 225.800 115.610 226.660 ;
      LAYER nwell ;
        RECT 117.210 225.090 119.130 227.350 ;
      LAYER pwell ;
        RECT 239.410 227.230 240.310 228.130 ;
      LAYER nwell ;
        RECT 249.180 227.630 251.090 229.860 ;
        RECT 267.950 229.200 269.870 231.460 ;
      LAYER pwell ;
        RECT 340.730 231.360 341.630 232.300 ;
        RECT 350.670 232.140 351.980 233.000 ;
      LAYER nwell ;
        RECT 353.580 231.430 355.500 233.690 ;
        RECT 366.230 233.650 367.080 233.760 ;
      LAYER pwell ;
        RECT 340.720 231.100 341.630 231.360 ;
      LAYER nwell ;
        RECT 354.550 231.340 355.400 231.430 ;
        RECT 366.010 231.420 367.920 233.650 ;
      LAYER pwell ;
        RECT 369.650 232.120 370.960 232.980 ;
        RECT 340.720 230.200 341.620 231.100 ;
      LAYER nwell ;
        RECT 350.710 229.670 351.560 229.780 ;
      LAYER pwell ;
        RECT 366.350 229.720 367.660 230.580 ;
        RECT 252.820 228.330 254.130 229.190 ;
      LAYER nwell ;
        RECT 268.920 229.110 269.770 229.200 ;
      LAYER pwell ;
        RECT 340.730 228.200 341.630 229.140 ;
        RECT 340.720 227.940 341.630 228.200 ;
      LAYER nwell ;
        RECT 164.980 226.560 165.830 226.670 ;
        RECT 118.180 225.000 119.030 225.090 ;
      LAYER pwell ;
        RECT 104.460 224.840 104.880 224.850 ;
        RECT 63.790 222.820 65.100 223.680 ;
        RECT 3.740 222.720 4.160 222.730 ;
        RECT 3.260 221.190 4.160 222.720 ;
      LAYER nwell ;
        RECT 66.700 222.110 68.620 224.370 ;
        RECT 164.760 224.330 166.670 226.560 ;
      LAYER pwell ;
        RECT 168.400 225.030 169.710 225.890 ;
        RECT 239.680 224.980 240.580 226.510 ;
        RECT 249.520 225.930 250.830 226.790 ;
      LAYER nwell ;
        RECT 252.430 225.220 254.350 227.480 ;
      LAYER pwell ;
        RECT 340.720 227.040 341.620 227.940 ;
      LAYER nwell ;
        RECT 350.490 227.440 352.400 229.670 ;
        RECT 369.260 229.010 371.180 231.270 ;
      LAYER pwell ;
        RECT 354.130 228.140 355.440 229.000 ;
      LAYER nwell ;
        RECT 370.230 228.920 371.080 229.010 ;
        RECT 300.200 226.690 301.050 226.800 ;
        RECT 253.400 225.130 254.250 225.220 ;
      LAYER pwell ;
        RECT 239.680 224.970 240.100 224.980 ;
      LAYER nwell ;
        RECT 299.980 224.460 301.890 226.690 ;
      LAYER pwell ;
        RECT 303.620 225.160 304.930 226.020 ;
        RECT 340.990 224.790 341.890 226.320 ;
        RECT 350.830 225.740 352.140 226.600 ;
      LAYER nwell ;
        RECT 353.740 225.030 355.660 227.290 ;
        RECT 401.510 226.500 402.360 226.610 ;
        RECT 354.710 224.940 355.560 225.030 ;
      LAYER pwell ;
        RECT 340.990 224.780 341.410 224.790 ;
        RECT 165.100 222.630 166.410 223.490 ;
        RECT 105.050 222.530 105.470 222.540 ;
      LAYER nwell ;
        RECT 67.670 222.020 68.520 222.110 ;
      LAYER pwell ;
        RECT 104.570 221.000 105.470 222.530 ;
      LAYER nwell ;
        RECT 168.010 221.920 169.930 224.180 ;
      LAYER pwell ;
        RECT 300.320 222.760 301.630 223.620 ;
        RECT 240.270 222.660 240.690 222.670 ;
      LAYER nwell ;
        RECT 168.980 221.830 169.830 221.920 ;
      LAYER pwell ;
        RECT 239.790 221.130 240.690 222.660 ;
      LAYER nwell ;
        RECT 303.230 222.050 305.150 224.310 ;
        RECT 401.290 224.270 403.200 226.500 ;
      LAYER pwell ;
        RECT 404.930 224.970 406.240 225.830 ;
        RECT 401.630 222.570 402.940 223.430 ;
        RECT 341.580 222.470 342.000 222.480 ;
      LAYER nwell ;
        RECT 304.200 221.960 305.050 222.050 ;
      LAYER pwell ;
        RECT 341.100 220.940 342.000 222.470 ;
      LAYER nwell ;
        RECT 404.540 221.860 406.460 224.120 ;
        RECT 405.510 221.770 406.360 221.860 ;
        RECT 12.850 220.670 13.700 220.780 ;
      LAYER pwell ;
        RECT 3.070 218.200 3.970 219.140 ;
      LAYER nwell ;
        RECT 12.630 218.440 14.540 220.670 ;
        RECT 249.380 220.610 250.230 220.720 ;
        RECT 114.160 220.480 115.010 220.590 ;
      LAYER pwell ;
        RECT 16.270 219.140 17.580 220.000 ;
        RECT 3.060 217.940 3.970 218.200 ;
        RECT 3.060 217.040 3.960 217.940 ;
        RECT 3.030 215.960 3.930 216.900 ;
        RECT 12.970 216.740 14.280 217.600 ;
      LAYER nwell ;
        RECT 15.880 216.030 17.800 218.290 ;
        RECT 28.530 218.250 29.380 218.360 ;
      LAYER pwell ;
        RECT 3.020 215.700 3.930 215.960 ;
      LAYER nwell ;
        RECT 16.850 215.940 17.700 216.030 ;
        RECT 28.310 216.020 30.220 218.250 ;
      LAYER pwell ;
        RECT 104.380 218.010 105.280 218.950 ;
      LAYER nwell ;
        RECT 113.940 218.250 115.850 220.480 ;
      LAYER pwell ;
        RECT 117.580 218.950 118.890 219.810 ;
        RECT 104.370 217.750 105.280 218.010 ;
        RECT 31.950 216.720 33.260 217.580 ;
        RECT 104.370 216.850 105.270 217.750 ;
        RECT 3.020 214.800 3.920 215.700 ;
      LAYER nwell ;
        RECT 13.010 214.270 13.860 214.380 ;
      LAYER pwell ;
        RECT 28.650 214.320 29.960 215.180 ;
        RECT 3.030 212.800 3.930 213.740 ;
        RECT 3.020 212.540 3.930 212.800 ;
        RECT 3.020 211.640 3.920 212.540 ;
      LAYER nwell ;
        RECT 12.790 212.040 14.700 214.270 ;
        RECT 31.560 213.610 33.480 215.870 ;
      LAYER pwell ;
        RECT 104.340 215.770 105.240 216.710 ;
        RECT 114.280 216.550 115.590 217.410 ;
      LAYER nwell ;
        RECT 117.190 215.840 119.110 218.100 ;
        RECT 129.840 218.060 130.690 218.170 ;
      LAYER pwell ;
        RECT 239.600 218.140 240.500 219.080 ;
      LAYER nwell ;
        RECT 249.160 218.380 251.070 220.610 ;
        RECT 350.690 220.420 351.540 220.530 ;
      LAYER pwell ;
        RECT 252.800 219.080 254.110 219.940 ;
        RECT 104.330 215.510 105.240 215.770 ;
      LAYER nwell ;
        RECT 118.160 215.750 119.010 215.840 ;
        RECT 129.620 215.830 131.530 218.060 ;
      LAYER pwell ;
        RECT 239.590 217.880 240.500 218.140 ;
        RECT 133.260 216.530 134.570 217.390 ;
        RECT 239.590 216.980 240.490 217.880 ;
        RECT 239.560 215.900 240.460 216.840 ;
        RECT 249.500 216.680 250.810 217.540 ;
      LAYER nwell ;
        RECT 252.410 215.970 254.330 218.230 ;
        RECT 265.060 218.190 265.910 218.300 ;
      LAYER pwell ;
        RECT 104.330 214.610 105.230 215.510 ;
      LAYER nwell ;
        RECT 114.320 214.080 115.170 214.190 ;
      LAYER pwell ;
        RECT 129.960 214.130 131.270 214.990 ;
        RECT 16.430 212.740 17.740 213.600 ;
      LAYER nwell ;
        RECT 32.530 213.520 33.380 213.610 ;
        RECT 46.110 212.700 46.960 212.810 ;
      LAYER pwell ;
        RECT 3.290 209.390 4.190 210.920 ;
        RECT 13.130 210.340 14.440 211.200 ;
      LAYER nwell ;
        RECT 16.040 209.630 17.960 211.890 ;
        RECT 45.890 210.470 47.800 212.700 ;
      LAYER pwell ;
        RECT 104.340 212.610 105.240 213.550 ;
        RECT 104.330 212.350 105.240 212.610 ;
        RECT 49.530 211.170 50.840 212.030 ;
        RECT 104.330 211.450 105.230 212.350 ;
      LAYER nwell ;
        RECT 114.100 211.850 116.010 214.080 ;
        RECT 132.870 213.420 134.790 215.680 ;
      LAYER pwell ;
        RECT 239.550 215.640 240.460 215.900 ;
      LAYER nwell ;
        RECT 253.380 215.880 254.230 215.970 ;
        RECT 264.840 215.960 266.750 218.190 ;
      LAYER pwell ;
        RECT 340.910 217.950 341.810 218.890 ;
      LAYER nwell ;
        RECT 350.470 218.190 352.380 220.420 ;
      LAYER pwell ;
        RECT 354.110 218.890 355.420 219.750 ;
        RECT 340.900 217.690 341.810 217.950 ;
        RECT 268.480 216.660 269.790 217.520 ;
        RECT 340.900 216.790 341.800 217.690 ;
        RECT 239.550 214.740 240.450 215.640 ;
      LAYER nwell ;
        RECT 249.540 214.210 250.390 214.320 ;
      LAYER pwell ;
        RECT 265.180 214.260 266.490 215.120 ;
        RECT 117.740 212.550 119.050 213.410 ;
      LAYER nwell ;
        RECT 133.840 213.330 134.690 213.420 ;
      LAYER pwell ;
        RECT 239.560 212.740 240.460 213.680 ;
      LAYER nwell ;
        RECT 147.420 212.510 148.270 212.620 ;
        RECT 17.010 209.540 17.860 209.630 ;
      LAYER pwell ;
        RECT 3.290 209.380 3.710 209.390 ;
        RECT 46.230 208.770 47.540 209.630 ;
      LAYER nwell ;
        RECT 49.140 208.060 51.060 210.320 ;
      LAYER pwell ;
        RECT 104.600 209.200 105.500 210.730 ;
        RECT 114.440 210.150 115.750 211.010 ;
      LAYER nwell ;
        RECT 117.350 209.440 119.270 211.700 ;
        RECT 147.200 210.280 149.110 212.510 ;
      LAYER pwell ;
        RECT 239.550 212.480 240.460 212.740 ;
        RECT 150.840 210.980 152.150 211.840 ;
        RECT 239.550 211.580 240.450 212.480 ;
      LAYER nwell ;
        RECT 249.320 211.980 251.230 214.210 ;
        RECT 268.090 213.550 270.010 215.810 ;
      LAYER pwell ;
        RECT 340.870 215.710 341.770 216.650 ;
        RECT 350.810 216.490 352.120 217.350 ;
      LAYER nwell ;
        RECT 353.720 215.780 355.640 218.040 ;
        RECT 366.370 218.000 367.220 218.110 ;
      LAYER pwell ;
        RECT 340.860 215.450 341.770 215.710 ;
      LAYER nwell ;
        RECT 354.690 215.690 355.540 215.780 ;
        RECT 366.150 215.770 368.060 218.000 ;
      LAYER pwell ;
        RECT 369.790 216.470 371.100 217.330 ;
        RECT 340.860 214.550 341.760 215.450 ;
      LAYER nwell ;
        RECT 350.850 214.020 351.700 214.130 ;
      LAYER pwell ;
        RECT 366.490 214.070 367.800 214.930 ;
        RECT 252.960 212.680 254.270 213.540 ;
      LAYER nwell ;
        RECT 269.060 213.460 269.910 213.550 ;
        RECT 282.640 212.640 283.490 212.750 ;
        RECT 118.320 209.350 119.170 209.440 ;
      LAYER pwell ;
        RECT 104.600 209.190 105.020 209.200 ;
        RECT 147.540 208.580 148.850 209.440 ;
      LAYER nwell ;
        RECT 50.110 207.970 50.960 208.060 ;
      LAYER pwell ;
        RECT 3.020 206.350 3.920 207.880 ;
      LAYER nwell ;
        RECT 150.450 207.870 152.370 210.130 ;
      LAYER pwell ;
        RECT 239.820 209.330 240.720 210.860 ;
        RECT 249.660 210.280 250.970 211.140 ;
      LAYER nwell ;
        RECT 252.570 209.570 254.490 211.830 ;
        RECT 282.420 210.410 284.330 212.640 ;
      LAYER pwell ;
        RECT 340.870 212.550 341.770 213.490 ;
        RECT 340.860 212.290 341.770 212.550 ;
        RECT 286.060 211.110 287.370 211.970 ;
        RECT 340.860 211.390 341.760 212.290 ;
      LAYER nwell ;
        RECT 350.630 211.790 352.540 214.020 ;
        RECT 369.400 213.360 371.320 215.620 ;
      LAYER pwell ;
        RECT 354.270 212.490 355.580 213.350 ;
      LAYER nwell ;
        RECT 370.370 213.270 371.220 213.360 ;
        RECT 383.950 212.450 384.800 212.560 ;
        RECT 253.540 209.480 254.390 209.570 ;
      LAYER pwell ;
        RECT 239.820 209.320 240.240 209.330 ;
        RECT 282.760 208.710 284.070 209.570 ;
      LAYER nwell ;
        RECT 285.670 208.000 287.590 210.260 ;
      LAYER pwell ;
        RECT 341.130 209.140 342.030 210.670 ;
        RECT 350.970 210.090 352.280 210.950 ;
      LAYER nwell ;
        RECT 353.880 209.380 355.800 211.640 ;
        RECT 383.730 210.220 385.640 212.450 ;
      LAYER pwell ;
        RECT 387.370 210.920 388.680 211.780 ;
      LAYER nwell ;
        RECT 354.850 209.290 355.700 209.380 ;
      LAYER pwell ;
        RECT 341.130 209.130 341.550 209.140 ;
        RECT 384.070 208.520 385.380 209.380 ;
      LAYER nwell ;
        RECT 286.640 207.910 287.490 208.000 ;
        RECT 151.420 207.780 152.270 207.870 ;
      LAYER pwell ;
        RECT 3.020 206.340 3.440 206.350 ;
      LAYER nwell ;
        RECT 12.680 206.250 13.530 206.360 ;
      LAYER pwell ;
        RECT 2.900 203.780 3.800 204.720 ;
      LAYER nwell ;
        RECT 12.460 204.020 14.370 206.250 ;
      LAYER pwell ;
        RECT 104.330 206.160 105.230 207.690 ;
        RECT 239.550 206.290 240.450 207.820 ;
      LAYER nwell ;
        RECT 386.980 207.810 388.900 210.070 ;
        RECT 387.950 207.720 388.800 207.810 ;
      LAYER pwell ;
        RECT 239.550 206.280 239.970 206.290 ;
      LAYER nwell ;
        RECT 249.210 206.190 250.060 206.300 ;
      LAYER pwell ;
        RECT 104.330 206.150 104.750 206.160 ;
      LAYER nwell ;
        RECT 113.990 206.060 114.840 206.170 ;
      LAYER pwell ;
        RECT 16.100 204.720 17.410 205.580 ;
        RECT 2.890 203.520 3.800 203.780 ;
        RECT 2.890 202.620 3.790 203.520 ;
        RECT 2.860 201.540 3.760 202.480 ;
        RECT 12.800 202.320 14.110 203.180 ;
      LAYER nwell ;
        RECT 15.710 201.610 17.630 203.870 ;
        RECT 28.360 203.830 29.210 203.940 ;
      LAYER pwell ;
        RECT 2.850 201.280 3.760 201.540 ;
      LAYER nwell ;
        RECT 16.680 201.520 17.530 201.610 ;
        RECT 28.140 201.600 30.050 203.830 ;
      LAYER pwell ;
        RECT 104.210 203.590 105.110 204.530 ;
      LAYER nwell ;
        RECT 113.770 203.830 115.680 206.060 ;
      LAYER pwell ;
        RECT 117.410 204.530 118.720 205.390 ;
        RECT 104.200 203.330 105.110 203.590 ;
        RECT 31.780 202.300 33.090 203.160 ;
        RECT 104.200 202.430 105.100 203.330 ;
        RECT 2.850 200.380 3.750 201.280 ;
      LAYER nwell ;
        RECT 12.840 199.850 13.690 199.960 ;
      LAYER pwell ;
        RECT 28.480 199.900 29.790 200.760 ;
        RECT 2.860 198.380 3.760 199.320 ;
        RECT 2.850 198.120 3.760 198.380 ;
        RECT 2.850 197.220 3.750 198.120 ;
      LAYER nwell ;
        RECT 12.620 197.620 14.530 199.850 ;
        RECT 31.390 199.190 33.310 201.450 ;
      LAYER pwell ;
        RECT 104.170 201.350 105.070 202.290 ;
        RECT 114.110 202.130 115.420 202.990 ;
      LAYER nwell ;
        RECT 117.020 201.420 118.940 203.680 ;
        RECT 129.670 203.640 130.520 203.750 ;
      LAYER pwell ;
        RECT 239.430 203.720 240.330 204.660 ;
      LAYER nwell ;
        RECT 248.990 203.960 250.900 206.190 ;
      LAYER pwell ;
        RECT 340.860 206.100 341.760 207.630 ;
        RECT 340.860 206.090 341.280 206.100 ;
      LAYER nwell ;
        RECT 350.520 206.000 351.370 206.110 ;
      LAYER pwell ;
        RECT 252.630 204.660 253.940 205.520 ;
        RECT 104.160 201.090 105.070 201.350 ;
      LAYER nwell ;
        RECT 117.990 201.330 118.840 201.420 ;
        RECT 129.450 201.410 131.360 203.640 ;
      LAYER pwell ;
        RECT 239.420 203.460 240.330 203.720 ;
        RECT 133.090 202.110 134.400 202.970 ;
        RECT 239.420 202.560 240.320 203.460 ;
        RECT 239.390 201.480 240.290 202.420 ;
        RECT 249.330 202.260 250.640 203.120 ;
      LAYER nwell ;
        RECT 252.240 201.550 254.160 203.810 ;
        RECT 264.890 203.770 265.740 203.880 ;
        RECT 77.870 200.460 78.720 200.570 ;
      LAYER pwell ;
        RECT 16.260 198.320 17.570 199.180 ;
      LAYER nwell ;
        RECT 32.360 199.100 33.210 199.190 ;
        RECT 77.650 198.230 79.560 200.460 ;
      LAYER pwell ;
        RECT 104.160 200.190 105.060 201.090 ;
        RECT 81.290 198.930 82.600 199.790 ;
      LAYER nwell ;
        RECT 114.150 199.660 115.000 199.770 ;
      LAYER pwell ;
        RECT 129.790 199.710 131.100 200.570 ;
        RECT 104.170 198.190 105.070 199.130 ;
        RECT 3.120 194.970 4.020 196.500 ;
        RECT 12.960 195.920 14.270 196.780 ;
      LAYER nwell ;
        RECT 15.870 195.210 17.790 197.470 ;
      LAYER pwell ;
        RECT 77.990 196.530 79.300 197.390 ;
      LAYER nwell ;
        RECT 80.900 195.820 82.820 198.080 ;
      LAYER pwell ;
        RECT 104.160 197.930 105.070 198.190 ;
        RECT 104.160 197.030 105.060 197.930 ;
      LAYER nwell ;
        RECT 113.930 197.430 115.840 199.660 ;
        RECT 132.700 199.000 134.620 201.260 ;
      LAYER pwell ;
        RECT 239.380 201.220 240.290 201.480 ;
      LAYER nwell ;
        RECT 253.210 201.460 254.060 201.550 ;
        RECT 264.670 201.540 266.580 203.770 ;
      LAYER pwell ;
        RECT 340.740 203.530 341.640 204.470 ;
      LAYER nwell ;
        RECT 350.300 203.770 352.210 206.000 ;
      LAYER pwell ;
        RECT 353.940 204.470 355.250 205.330 ;
        RECT 340.730 203.270 341.640 203.530 ;
        RECT 268.310 202.240 269.620 203.100 ;
        RECT 340.730 202.370 341.630 203.270 ;
      LAYER nwell ;
        RECT 179.180 200.270 180.030 200.380 ;
      LAYER pwell ;
        RECT 239.380 200.320 240.280 201.220 ;
        RECT 117.570 198.130 118.880 198.990 ;
      LAYER nwell ;
        RECT 133.670 198.910 134.520 199.000 ;
        RECT 178.960 198.040 180.870 200.270 ;
        RECT 249.370 199.790 250.220 199.900 ;
      LAYER pwell ;
        RECT 265.010 199.840 266.320 200.700 ;
        RECT 182.600 198.740 183.910 199.600 ;
        RECT 239.390 198.320 240.290 199.260 ;
        RECT 239.380 198.060 240.290 198.320 ;
      LAYER nwell ;
        RECT 81.870 195.730 82.720 195.820 ;
        RECT 16.840 195.120 17.690 195.210 ;
      LAYER pwell ;
        RECT 3.120 194.960 3.540 194.970 ;
        RECT 104.430 194.780 105.330 196.310 ;
        RECT 114.270 195.730 115.580 196.590 ;
      LAYER nwell ;
        RECT 117.180 195.020 119.100 197.280 ;
      LAYER pwell ;
        RECT 179.300 196.340 180.610 197.200 ;
      LAYER nwell ;
        RECT 182.210 195.630 184.130 197.890 ;
      LAYER pwell ;
        RECT 239.380 197.160 240.280 198.060 ;
      LAYER nwell ;
        RECT 249.150 197.560 251.060 199.790 ;
        RECT 267.920 199.130 269.840 201.390 ;
      LAYER pwell ;
        RECT 340.700 201.290 341.600 202.230 ;
        RECT 350.640 202.070 351.950 202.930 ;
      LAYER nwell ;
        RECT 353.550 201.360 355.470 203.620 ;
        RECT 366.200 203.580 367.050 203.690 ;
      LAYER pwell ;
        RECT 340.690 201.030 341.600 201.290 ;
      LAYER nwell ;
        RECT 354.520 201.270 355.370 201.360 ;
        RECT 365.980 201.350 367.890 203.580 ;
      LAYER pwell ;
        RECT 369.620 202.050 370.930 202.910 ;
      LAYER nwell ;
        RECT 314.400 200.400 315.250 200.510 ;
      LAYER pwell ;
        RECT 252.790 198.260 254.100 199.120 ;
      LAYER nwell ;
        RECT 268.890 199.040 269.740 199.130 ;
        RECT 314.180 198.170 316.090 200.400 ;
      LAYER pwell ;
        RECT 340.690 200.130 341.590 201.030 ;
        RECT 317.820 198.870 319.130 199.730 ;
      LAYER nwell ;
        RECT 350.680 199.600 351.530 199.710 ;
      LAYER pwell ;
        RECT 366.320 199.650 367.630 200.510 ;
        RECT 340.700 198.130 341.600 199.070 ;
      LAYER nwell ;
        RECT 183.180 195.540 184.030 195.630 ;
        RECT 118.150 194.930 119.000 195.020 ;
      LAYER pwell ;
        RECT 239.650 194.910 240.550 196.440 ;
        RECT 249.490 195.860 250.800 196.720 ;
      LAYER nwell ;
        RECT 252.400 195.150 254.320 197.410 ;
      LAYER pwell ;
        RECT 314.520 196.470 315.830 197.330 ;
      LAYER nwell ;
        RECT 317.430 195.760 319.350 198.020 ;
      LAYER pwell ;
        RECT 340.690 197.870 341.600 198.130 ;
        RECT 340.690 196.970 341.590 197.870 ;
      LAYER nwell ;
        RECT 350.460 197.370 352.370 199.600 ;
        RECT 369.230 198.940 371.150 201.200 ;
        RECT 415.710 200.210 416.560 200.320 ;
      LAYER pwell ;
        RECT 354.100 198.070 355.410 198.930 ;
      LAYER nwell ;
        RECT 370.200 198.850 371.050 198.940 ;
        RECT 415.490 197.980 417.400 200.210 ;
      LAYER pwell ;
        RECT 419.130 198.680 420.440 199.540 ;
      LAYER nwell ;
        RECT 318.400 195.670 319.250 195.760 ;
        RECT 253.370 195.060 254.220 195.150 ;
      LAYER pwell ;
        RECT 239.650 194.900 240.070 194.910 ;
        RECT 104.430 194.770 104.850 194.780 ;
        RECT 340.960 194.720 341.860 196.250 ;
        RECT 350.800 195.670 352.110 196.530 ;
      LAYER nwell ;
        RECT 353.710 194.960 355.630 197.220 ;
      LAYER pwell ;
        RECT 415.830 196.280 417.140 197.140 ;
      LAYER nwell ;
        RECT 418.740 195.570 420.660 197.830 ;
        RECT 419.710 195.480 420.560 195.570 ;
        RECT 354.680 194.870 355.530 194.960 ;
      LAYER pwell ;
        RECT 340.960 194.710 341.380 194.720 ;
        RECT 2.680 191.840 4.210 192.320 ;
        RECT 2.680 191.420 4.220 191.840 ;
        RECT 103.990 191.650 105.520 192.130 ;
        RECT 239.210 191.780 240.740 192.260 ;
        RECT 103.990 191.230 105.530 191.650 ;
        RECT 239.210 191.360 240.750 191.780 ;
        RECT 340.520 191.590 342.050 192.070 ;
        RECT 340.520 191.170 342.060 191.590 ;
      LAYER nwell ;
        RECT 12.530 190.820 13.380 190.930 ;
      LAYER pwell ;
        RECT 2.750 188.350 3.650 189.290 ;
      LAYER nwell ;
        RECT 12.310 188.590 14.220 190.820 ;
        RECT 249.060 190.760 249.910 190.870 ;
        RECT 113.840 190.630 114.690 190.740 ;
      LAYER pwell ;
        RECT 15.950 189.290 17.260 190.150 ;
        RECT 2.740 188.090 3.650 188.350 ;
        RECT 2.740 187.190 3.640 188.090 ;
        RECT 2.710 186.110 3.610 187.050 ;
        RECT 12.650 186.890 13.960 187.750 ;
      LAYER nwell ;
        RECT 15.560 186.180 17.480 188.440 ;
        RECT 28.210 188.400 29.060 188.510 ;
      LAYER pwell ;
        RECT 2.700 185.850 3.610 186.110 ;
      LAYER nwell ;
        RECT 16.530 186.090 17.380 186.180 ;
        RECT 27.990 186.170 29.900 188.400 ;
      LAYER pwell ;
        RECT 104.060 188.160 104.960 189.100 ;
      LAYER nwell ;
        RECT 113.620 188.400 115.530 190.630 ;
      LAYER pwell ;
        RECT 117.260 189.100 118.570 189.960 ;
        RECT 104.050 187.900 104.960 188.160 ;
        RECT 31.630 186.870 32.940 187.730 ;
        RECT 104.050 187.000 104.950 187.900 ;
        RECT 2.700 184.950 3.600 185.850 ;
      LAYER nwell ;
        RECT 12.690 184.420 13.540 184.530 ;
      LAYER pwell ;
        RECT 28.330 184.470 29.640 185.330 ;
        RECT 2.710 182.950 3.610 183.890 ;
        RECT 2.700 182.690 3.610 182.950 ;
        RECT 2.700 181.790 3.600 182.690 ;
      LAYER nwell ;
        RECT 12.470 182.190 14.380 184.420 ;
        RECT 31.240 183.760 33.160 186.020 ;
      LAYER pwell ;
        RECT 104.020 185.920 104.920 186.860 ;
        RECT 113.960 186.700 115.270 187.560 ;
      LAYER nwell ;
        RECT 116.870 185.990 118.790 188.250 ;
        RECT 129.520 188.210 130.370 188.320 ;
      LAYER pwell ;
        RECT 239.280 188.290 240.180 189.230 ;
      LAYER nwell ;
        RECT 248.840 188.530 250.750 190.760 ;
        RECT 350.370 190.570 351.220 190.680 ;
      LAYER pwell ;
        RECT 252.480 189.230 253.790 190.090 ;
        RECT 104.010 185.660 104.920 185.920 ;
      LAYER nwell ;
        RECT 117.840 185.900 118.690 185.990 ;
        RECT 129.300 185.980 131.210 188.210 ;
      LAYER pwell ;
        RECT 239.270 188.030 240.180 188.290 ;
        RECT 132.940 186.680 134.250 187.540 ;
        RECT 239.270 187.130 240.170 188.030 ;
        RECT 239.240 186.050 240.140 186.990 ;
        RECT 249.180 186.830 250.490 187.690 ;
      LAYER nwell ;
        RECT 252.090 186.120 254.010 188.380 ;
        RECT 264.740 188.340 265.590 188.450 ;
      LAYER pwell ;
        RECT 104.010 184.760 104.910 185.660 ;
      LAYER nwell ;
        RECT 114.000 184.230 114.850 184.340 ;
      LAYER pwell ;
        RECT 129.640 184.280 130.950 185.140 ;
        RECT 16.110 182.890 17.420 183.750 ;
      LAYER nwell ;
        RECT 32.210 183.670 33.060 183.760 ;
        RECT 45.790 182.850 46.640 182.960 ;
      LAYER pwell ;
        RECT 2.970 179.540 3.870 181.070 ;
        RECT 12.810 180.490 14.120 181.350 ;
      LAYER nwell ;
        RECT 15.720 179.780 17.640 182.040 ;
        RECT 45.570 180.620 47.480 182.850 ;
      LAYER pwell ;
        RECT 104.020 182.760 104.920 183.700 ;
        RECT 104.010 182.500 104.920 182.760 ;
        RECT 49.210 181.320 50.520 182.180 ;
        RECT 104.010 181.600 104.910 182.500 ;
      LAYER nwell ;
        RECT 113.780 182.000 115.690 184.230 ;
        RECT 132.550 183.570 134.470 185.830 ;
      LAYER pwell ;
        RECT 239.230 185.790 240.140 186.050 ;
      LAYER nwell ;
        RECT 253.060 186.030 253.910 186.120 ;
        RECT 264.520 186.110 266.430 188.340 ;
      LAYER pwell ;
        RECT 340.590 188.100 341.490 189.040 ;
      LAYER nwell ;
        RECT 350.150 188.340 352.060 190.570 ;
      LAYER pwell ;
        RECT 353.790 189.040 355.100 189.900 ;
        RECT 340.580 187.840 341.490 188.100 ;
        RECT 268.160 186.810 269.470 187.670 ;
        RECT 340.580 186.940 341.480 187.840 ;
        RECT 239.230 184.890 240.130 185.790 ;
      LAYER nwell ;
        RECT 249.220 184.360 250.070 184.470 ;
      LAYER pwell ;
        RECT 264.860 184.410 266.170 185.270 ;
        RECT 117.420 182.700 118.730 183.560 ;
      LAYER nwell ;
        RECT 133.520 183.480 134.370 183.570 ;
      LAYER pwell ;
        RECT 239.240 182.890 240.140 183.830 ;
      LAYER nwell ;
        RECT 147.100 182.660 147.950 182.770 ;
        RECT 16.690 179.690 17.540 179.780 ;
      LAYER pwell ;
        RECT 2.970 179.530 3.390 179.540 ;
        RECT 45.910 178.920 47.220 179.780 ;
      LAYER nwell ;
        RECT 48.820 178.210 50.740 180.470 ;
      LAYER pwell ;
        RECT 104.280 179.350 105.180 180.880 ;
        RECT 114.120 180.300 115.430 181.160 ;
      LAYER nwell ;
        RECT 117.030 179.590 118.950 181.850 ;
        RECT 146.880 180.430 148.790 182.660 ;
      LAYER pwell ;
        RECT 239.230 182.630 240.140 182.890 ;
        RECT 150.520 181.130 151.830 181.990 ;
        RECT 239.230 181.730 240.130 182.630 ;
      LAYER nwell ;
        RECT 249.000 182.130 250.910 184.360 ;
        RECT 267.770 183.700 269.690 185.960 ;
      LAYER pwell ;
        RECT 340.550 185.860 341.450 186.800 ;
        RECT 350.490 186.640 351.800 187.500 ;
      LAYER nwell ;
        RECT 353.400 185.930 355.320 188.190 ;
        RECT 366.050 188.150 366.900 188.260 ;
      LAYER pwell ;
        RECT 340.540 185.600 341.450 185.860 ;
      LAYER nwell ;
        RECT 354.370 185.840 355.220 185.930 ;
        RECT 365.830 185.920 367.740 188.150 ;
      LAYER pwell ;
        RECT 369.470 186.620 370.780 187.480 ;
        RECT 340.540 184.700 341.440 185.600 ;
      LAYER nwell ;
        RECT 350.530 184.170 351.380 184.280 ;
      LAYER pwell ;
        RECT 366.170 184.220 367.480 185.080 ;
        RECT 252.640 182.830 253.950 183.690 ;
      LAYER nwell ;
        RECT 268.740 183.610 269.590 183.700 ;
        RECT 282.320 182.790 283.170 182.900 ;
        RECT 118.000 179.500 118.850 179.590 ;
      LAYER pwell ;
        RECT 104.280 179.340 104.700 179.350 ;
        RECT 147.220 178.730 148.530 179.590 ;
      LAYER nwell ;
        RECT 49.790 178.120 50.640 178.210 ;
      LAYER pwell ;
        RECT 2.700 176.500 3.600 178.030 ;
      LAYER nwell ;
        RECT 150.130 178.020 152.050 180.280 ;
      LAYER pwell ;
        RECT 239.500 179.480 240.400 181.010 ;
        RECT 249.340 180.430 250.650 181.290 ;
      LAYER nwell ;
        RECT 252.250 179.720 254.170 181.980 ;
        RECT 282.100 180.560 284.010 182.790 ;
      LAYER pwell ;
        RECT 340.550 182.700 341.450 183.640 ;
        RECT 340.540 182.440 341.450 182.700 ;
        RECT 285.740 181.260 287.050 182.120 ;
        RECT 340.540 181.540 341.440 182.440 ;
      LAYER nwell ;
        RECT 350.310 181.940 352.220 184.170 ;
        RECT 369.080 183.510 371.000 185.770 ;
      LAYER pwell ;
        RECT 353.950 182.640 355.260 183.500 ;
      LAYER nwell ;
        RECT 370.050 183.420 370.900 183.510 ;
        RECT 383.630 182.600 384.480 182.710 ;
        RECT 253.220 179.630 254.070 179.720 ;
      LAYER pwell ;
        RECT 239.500 179.470 239.920 179.480 ;
        RECT 282.440 178.860 283.750 179.720 ;
      LAYER nwell ;
        RECT 285.350 178.150 287.270 180.410 ;
      LAYER pwell ;
        RECT 340.810 179.290 341.710 180.820 ;
        RECT 350.650 180.240 351.960 181.100 ;
      LAYER nwell ;
        RECT 353.560 179.530 355.480 181.790 ;
        RECT 383.410 180.370 385.320 182.600 ;
      LAYER pwell ;
        RECT 387.050 181.070 388.360 181.930 ;
      LAYER nwell ;
        RECT 354.530 179.440 355.380 179.530 ;
      LAYER pwell ;
        RECT 340.810 179.280 341.230 179.290 ;
        RECT 383.750 178.670 385.060 179.530 ;
      LAYER nwell ;
        RECT 286.320 178.060 287.170 178.150 ;
        RECT 151.100 177.930 151.950 178.020 ;
      LAYER pwell ;
        RECT 2.700 176.490 3.120 176.500 ;
      LAYER nwell ;
        RECT 12.360 176.400 13.210 176.510 ;
      LAYER pwell ;
        RECT 2.580 173.930 3.480 174.870 ;
      LAYER nwell ;
        RECT 12.140 174.170 14.050 176.400 ;
      LAYER pwell ;
        RECT 104.010 176.310 104.910 177.840 ;
        RECT 239.230 176.440 240.130 177.970 ;
      LAYER nwell ;
        RECT 386.660 177.960 388.580 180.220 ;
        RECT 387.630 177.870 388.480 177.960 ;
      LAYER pwell ;
        RECT 239.230 176.430 239.650 176.440 ;
      LAYER nwell ;
        RECT 248.890 176.340 249.740 176.450 ;
      LAYER pwell ;
        RECT 104.010 176.300 104.430 176.310 ;
      LAYER nwell ;
        RECT 113.670 176.210 114.520 176.320 ;
      LAYER pwell ;
        RECT 15.780 174.870 17.090 175.730 ;
        RECT 2.570 173.670 3.480 173.930 ;
        RECT 2.570 172.770 3.470 173.670 ;
        RECT 2.540 171.690 3.440 172.630 ;
        RECT 12.480 172.470 13.790 173.330 ;
      LAYER nwell ;
        RECT 15.390 171.760 17.310 174.020 ;
        RECT 28.040 173.980 28.890 174.090 ;
      LAYER pwell ;
        RECT 2.530 171.430 3.440 171.690 ;
      LAYER nwell ;
        RECT 16.360 171.670 17.210 171.760 ;
        RECT 27.820 171.750 29.730 173.980 ;
      LAYER pwell ;
        RECT 103.890 173.740 104.790 174.680 ;
      LAYER nwell ;
        RECT 113.450 173.980 115.360 176.210 ;
      LAYER pwell ;
        RECT 117.090 174.680 118.400 175.540 ;
        RECT 103.880 173.480 104.790 173.740 ;
        RECT 31.460 172.450 32.770 173.310 ;
        RECT 103.880 172.580 104.780 173.480 ;
        RECT 2.530 170.530 3.430 171.430 ;
      LAYER nwell ;
        RECT 12.520 170.000 13.370 170.110 ;
      LAYER pwell ;
        RECT 28.160 170.050 29.470 170.910 ;
        RECT 2.540 168.530 3.440 169.470 ;
        RECT 2.530 168.270 3.440 168.530 ;
        RECT 2.530 167.370 3.430 168.270 ;
      LAYER nwell ;
        RECT 12.300 167.770 14.210 170.000 ;
        RECT 31.070 169.340 32.990 171.600 ;
      LAYER pwell ;
        RECT 103.850 171.500 104.750 172.440 ;
        RECT 113.790 172.280 115.100 173.140 ;
      LAYER nwell ;
        RECT 116.700 171.570 118.620 173.830 ;
        RECT 129.350 173.790 130.200 173.900 ;
      LAYER pwell ;
        RECT 239.110 173.870 240.010 174.810 ;
      LAYER nwell ;
        RECT 248.670 174.110 250.580 176.340 ;
      LAYER pwell ;
        RECT 340.540 176.250 341.440 177.780 ;
        RECT 340.540 176.240 340.960 176.250 ;
      LAYER nwell ;
        RECT 350.200 176.150 351.050 176.260 ;
      LAYER pwell ;
        RECT 252.310 174.810 253.620 175.670 ;
        RECT 103.840 171.240 104.750 171.500 ;
      LAYER nwell ;
        RECT 117.670 171.480 118.520 171.570 ;
        RECT 129.130 171.560 131.040 173.790 ;
      LAYER pwell ;
        RECT 239.100 173.610 240.010 173.870 ;
        RECT 132.770 172.260 134.080 173.120 ;
        RECT 239.100 172.710 240.000 173.610 ;
        RECT 239.070 171.630 239.970 172.570 ;
        RECT 249.010 172.410 250.320 173.270 ;
      LAYER nwell ;
        RECT 251.920 171.700 253.840 173.960 ;
        RECT 264.570 173.920 265.420 174.030 ;
      LAYER pwell ;
        RECT 103.840 170.340 104.740 171.240 ;
      LAYER nwell ;
        RECT 113.830 169.810 114.680 169.920 ;
      LAYER pwell ;
        RECT 129.470 169.860 130.780 170.720 ;
        RECT 15.940 168.470 17.250 169.330 ;
      LAYER nwell ;
        RECT 32.040 169.250 32.890 169.340 ;
      LAYER pwell ;
        RECT 103.850 168.340 104.750 169.280 ;
        RECT 103.840 168.080 104.750 168.340 ;
        RECT 2.800 165.120 3.700 166.650 ;
        RECT 12.640 166.070 13.950 166.930 ;
      LAYER nwell ;
        RECT 15.550 165.360 17.470 167.620 ;
      LAYER pwell ;
        RECT 103.840 167.180 104.740 168.080 ;
      LAYER nwell ;
        RECT 113.610 167.580 115.520 169.810 ;
        RECT 132.380 169.150 134.300 171.410 ;
      LAYER pwell ;
        RECT 239.060 171.370 239.970 171.630 ;
      LAYER nwell ;
        RECT 252.890 171.610 253.740 171.700 ;
        RECT 264.350 171.690 266.260 173.920 ;
      LAYER pwell ;
        RECT 340.420 173.680 341.320 174.620 ;
      LAYER nwell ;
        RECT 349.980 173.920 351.890 176.150 ;
      LAYER pwell ;
        RECT 353.620 174.620 354.930 175.480 ;
        RECT 340.410 173.420 341.320 173.680 ;
        RECT 267.990 172.390 269.300 173.250 ;
        RECT 340.410 172.520 341.310 173.420 ;
        RECT 239.060 170.470 239.960 171.370 ;
      LAYER nwell ;
        RECT 249.050 169.940 249.900 170.050 ;
      LAYER pwell ;
        RECT 264.690 169.990 266.000 170.850 ;
        RECT 117.250 168.280 118.560 169.140 ;
      LAYER nwell ;
        RECT 133.350 169.060 134.200 169.150 ;
      LAYER pwell ;
        RECT 239.070 168.470 239.970 169.410 ;
        RECT 239.060 168.210 239.970 168.470 ;
      LAYER nwell ;
        RECT 63.320 166.830 64.170 166.940 ;
        RECT 16.520 165.270 17.370 165.360 ;
      LAYER pwell ;
        RECT 2.800 165.110 3.220 165.120 ;
      LAYER nwell ;
        RECT 63.100 164.600 65.010 166.830 ;
      LAYER pwell ;
        RECT 66.740 165.300 68.050 166.160 ;
        RECT 104.110 164.930 105.010 166.460 ;
        RECT 113.950 165.880 115.260 166.740 ;
      LAYER nwell ;
        RECT 116.860 165.170 118.780 167.430 ;
      LAYER pwell ;
        RECT 239.060 167.310 239.960 168.210 ;
      LAYER nwell ;
        RECT 248.830 167.710 250.740 169.940 ;
        RECT 267.600 169.280 269.520 171.540 ;
      LAYER pwell ;
        RECT 340.380 171.440 341.280 172.380 ;
        RECT 350.320 172.220 351.630 173.080 ;
      LAYER nwell ;
        RECT 353.230 171.510 355.150 173.770 ;
        RECT 365.880 173.730 366.730 173.840 ;
      LAYER pwell ;
        RECT 340.370 171.180 341.280 171.440 ;
      LAYER nwell ;
        RECT 354.200 171.420 355.050 171.510 ;
        RECT 365.660 171.500 367.570 173.730 ;
      LAYER pwell ;
        RECT 369.300 172.200 370.610 173.060 ;
        RECT 340.370 170.280 341.270 171.180 ;
      LAYER nwell ;
        RECT 350.360 169.750 351.210 169.860 ;
      LAYER pwell ;
        RECT 366.000 169.800 367.310 170.660 ;
        RECT 252.470 168.410 253.780 169.270 ;
      LAYER nwell ;
        RECT 268.570 169.190 269.420 169.280 ;
      LAYER pwell ;
        RECT 340.380 168.280 341.280 169.220 ;
        RECT 340.370 168.020 341.280 168.280 ;
      LAYER nwell ;
        RECT 164.630 166.640 165.480 166.750 ;
        RECT 117.830 165.080 118.680 165.170 ;
      LAYER pwell ;
        RECT 104.110 164.920 104.530 164.930 ;
        RECT 63.440 162.900 64.750 163.760 ;
        RECT 3.390 162.800 3.810 162.810 ;
        RECT 2.910 161.270 3.810 162.800 ;
      LAYER nwell ;
        RECT 66.350 162.190 68.270 164.450 ;
        RECT 164.410 164.410 166.320 166.640 ;
      LAYER pwell ;
        RECT 168.050 165.110 169.360 165.970 ;
        RECT 239.330 165.060 240.230 166.590 ;
        RECT 249.170 166.010 250.480 166.870 ;
      LAYER nwell ;
        RECT 252.080 165.300 254.000 167.560 ;
      LAYER pwell ;
        RECT 340.370 167.120 341.270 168.020 ;
      LAYER nwell ;
        RECT 350.140 167.520 352.050 169.750 ;
        RECT 368.910 169.090 370.830 171.350 ;
      LAYER pwell ;
        RECT 353.780 168.220 355.090 169.080 ;
      LAYER nwell ;
        RECT 369.880 169.000 370.730 169.090 ;
        RECT 299.850 166.770 300.700 166.880 ;
        RECT 253.050 165.210 253.900 165.300 ;
      LAYER pwell ;
        RECT 239.330 165.050 239.750 165.060 ;
      LAYER nwell ;
        RECT 299.630 164.540 301.540 166.770 ;
      LAYER pwell ;
        RECT 303.270 165.240 304.580 166.100 ;
        RECT 340.640 164.870 341.540 166.400 ;
        RECT 350.480 165.820 351.790 166.680 ;
      LAYER nwell ;
        RECT 353.390 165.110 355.310 167.370 ;
        RECT 401.160 166.580 402.010 166.690 ;
        RECT 354.360 165.020 355.210 165.110 ;
      LAYER pwell ;
        RECT 340.640 164.860 341.060 164.870 ;
        RECT 164.750 162.710 166.060 163.570 ;
        RECT 104.700 162.610 105.120 162.620 ;
      LAYER nwell ;
        RECT 67.320 162.100 68.170 162.190 ;
      LAYER pwell ;
        RECT 104.220 161.080 105.120 162.610 ;
      LAYER nwell ;
        RECT 167.660 162.000 169.580 164.260 ;
      LAYER pwell ;
        RECT 299.970 162.840 301.280 163.700 ;
        RECT 239.920 162.740 240.340 162.750 ;
      LAYER nwell ;
        RECT 168.630 161.910 169.480 162.000 ;
      LAYER pwell ;
        RECT 239.440 161.210 240.340 162.740 ;
      LAYER nwell ;
        RECT 302.880 162.130 304.800 164.390 ;
        RECT 400.940 164.350 402.850 166.580 ;
      LAYER pwell ;
        RECT 404.580 165.050 405.890 165.910 ;
        RECT 401.280 162.650 402.590 163.510 ;
        RECT 341.230 162.550 341.650 162.560 ;
      LAYER nwell ;
        RECT 303.850 162.040 304.700 162.130 ;
      LAYER pwell ;
        RECT 340.750 161.020 341.650 162.550 ;
      LAYER nwell ;
        RECT 404.190 161.940 406.110 164.200 ;
        RECT 405.160 161.850 406.010 161.940 ;
        RECT 12.500 160.750 13.350 160.860 ;
      LAYER pwell ;
        RECT 2.720 158.280 3.620 159.220 ;
      LAYER nwell ;
        RECT 12.280 158.520 14.190 160.750 ;
        RECT 249.030 160.690 249.880 160.800 ;
        RECT 113.810 160.560 114.660 160.670 ;
      LAYER pwell ;
        RECT 15.920 159.220 17.230 160.080 ;
        RECT 2.710 158.020 3.620 158.280 ;
        RECT 2.710 157.120 3.610 158.020 ;
        RECT 2.680 156.040 3.580 156.980 ;
        RECT 12.620 156.820 13.930 157.680 ;
      LAYER nwell ;
        RECT 15.530 156.110 17.450 158.370 ;
        RECT 28.180 158.330 29.030 158.440 ;
      LAYER pwell ;
        RECT 2.670 155.780 3.580 156.040 ;
      LAYER nwell ;
        RECT 16.500 156.020 17.350 156.110 ;
        RECT 27.960 156.100 29.870 158.330 ;
      LAYER pwell ;
        RECT 104.030 158.090 104.930 159.030 ;
      LAYER nwell ;
        RECT 113.590 158.330 115.500 160.560 ;
      LAYER pwell ;
        RECT 117.230 159.030 118.540 159.890 ;
        RECT 104.020 157.830 104.930 158.090 ;
        RECT 31.600 156.800 32.910 157.660 ;
        RECT 104.020 156.930 104.920 157.830 ;
        RECT 2.670 154.880 3.570 155.780 ;
      LAYER nwell ;
        RECT 12.660 154.350 13.510 154.460 ;
      LAYER pwell ;
        RECT 28.300 154.400 29.610 155.260 ;
        RECT 2.680 152.880 3.580 153.820 ;
        RECT 2.670 152.620 3.580 152.880 ;
        RECT 2.670 151.720 3.570 152.620 ;
      LAYER nwell ;
        RECT 12.440 152.120 14.350 154.350 ;
        RECT 31.210 153.690 33.130 155.950 ;
      LAYER pwell ;
        RECT 103.990 155.850 104.890 156.790 ;
        RECT 113.930 156.630 115.240 157.490 ;
      LAYER nwell ;
        RECT 116.840 155.920 118.760 158.180 ;
        RECT 129.490 158.140 130.340 158.250 ;
      LAYER pwell ;
        RECT 239.250 158.220 240.150 159.160 ;
      LAYER nwell ;
        RECT 248.810 158.460 250.720 160.690 ;
        RECT 350.340 160.500 351.190 160.610 ;
      LAYER pwell ;
        RECT 252.450 159.160 253.760 160.020 ;
        RECT 103.980 155.590 104.890 155.850 ;
      LAYER nwell ;
        RECT 117.810 155.830 118.660 155.920 ;
        RECT 129.270 155.910 131.180 158.140 ;
      LAYER pwell ;
        RECT 239.240 157.960 240.150 158.220 ;
        RECT 132.910 156.610 134.220 157.470 ;
        RECT 239.240 157.060 240.140 157.960 ;
        RECT 239.210 155.980 240.110 156.920 ;
        RECT 249.150 156.760 250.460 157.620 ;
      LAYER nwell ;
        RECT 252.060 156.050 253.980 158.310 ;
        RECT 264.710 158.270 265.560 158.380 ;
      LAYER pwell ;
        RECT 103.980 154.690 104.880 155.590 ;
      LAYER nwell ;
        RECT 113.970 154.160 114.820 154.270 ;
      LAYER pwell ;
        RECT 129.610 154.210 130.920 155.070 ;
        RECT 16.080 152.820 17.390 153.680 ;
      LAYER nwell ;
        RECT 32.180 153.600 33.030 153.690 ;
        RECT 45.760 152.780 46.610 152.890 ;
      LAYER pwell ;
        RECT 2.940 149.470 3.840 151.000 ;
        RECT 12.780 150.420 14.090 151.280 ;
      LAYER nwell ;
        RECT 15.690 149.710 17.610 151.970 ;
        RECT 45.540 150.550 47.450 152.780 ;
      LAYER pwell ;
        RECT 103.990 152.690 104.890 153.630 ;
        RECT 103.980 152.430 104.890 152.690 ;
        RECT 49.180 151.250 50.490 152.110 ;
        RECT 103.980 151.530 104.880 152.430 ;
      LAYER nwell ;
        RECT 113.750 151.930 115.660 154.160 ;
        RECT 132.520 153.500 134.440 155.760 ;
      LAYER pwell ;
        RECT 239.200 155.720 240.110 155.980 ;
      LAYER nwell ;
        RECT 253.030 155.960 253.880 156.050 ;
        RECT 264.490 156.040 266.400 158.270 ;
      LAYER pwell ;
        RECT 340.560 158.030 341.460 158.970 ;
      LAYER nwell ;
        RECT 350.120 158.270 352.030 160.500 ;
      LAYER pwell ;
        RECT 353.760 158.970 355.070 159.830 ;
        RECT 340.550 157.770 341.460 158.030 ;
        RECT 268.130 156.740 269.440 157.600 ;
        RECT 340.550 156.870 341.450 157.770 ;
        RECT 239.200 154.820 240.100 155.720 ;
      LAYER nwell ;
        RECT 249.190 154.290 250.040 154.400 ;
      LAYER pwell ;
        RECT 264.830 154.340 266.140 155.200 ;
        RECT 117.390 152.630 118.700 153.490 ;
      LAYER nwell ;
        RECT 133.490 153.410 134.340 153.500 ;
      LAYER pwell ;
        RECT 239.210 152.820 240.110 153.760 ;
      LAYER nwell ;
        RECT 147.070 152.590 147.920 152.700 ;
        RECT 16.660 149.620 17.510 149.710 ;
      LAYER pwell ;
        RECT 2.940 149.460 3.360 149.470 ;
        RECT 45.880 148.850 47.190 149.710 ;
      LAYER nwell ;
        RECT 48.790 148.140 50.710 150.400 ;
      LAYER pwell ;
        RECT 104.250 149.280 105.150 150.810 ;
        RECT 114.090 150.230 115.400 151.090 ;
      LAYER nwell ;
        RECT 117.000 149.520 118.920 151.780 ;
        RECT 146.850 150.360 148.760 152.590 ;
      LAYER pwell ;
        RECT 239.200 152.560 240.110 152.820 ;
        RECT 150.490 151.060 151.800 151.920 ;
        RECT 239.200 151.660 240.100 152.560 ;
      LAYER nwell ;
        RECT 248.970 152.060 250.880 154.290 ;
        RECT 267.740 153.630 269.660 155.890 ;
      LAYER pwell ;
        RECT 340.520 155.790 341.420 156.730 ;
        RECT 350.460 156.570 351.770 157.430 ;
      LAYER nwell ;
        RECT 353.370 155.860 355.290 158.120 ;
        RECT 366.020 158.080 366.870 158.190 ;
      LAYER pwell ;
        RECT 340.510 155.530 341.420 155.790 ;
      LAYER nwell ;
        RECT 354.340 155.770 355.190 155.860 ;
        RECT 365.800 155.850 367.710 158.080 ;
      LAYER pwell ;
        RECT 369.440 156.550 370.750 157.410 ;
        RECT 340.510 154.630 341.410 155.530 ;
      LAYER nwell ;
        RECT 350.500 154.100 351.350 154.210 ;
      LAYER pwell ;
        RECT 366.140 154.150 367.450 155.010 ;
        RECT 252.610 152.760 253.920 153.620 ;
      LAYER nwell ;
        RECT 268.710 153.540 269.560 153.630 ;
        RECT 282.290 152.720 283.140 152.830 ;
        RECT 117.970 149.430 118.820 149.520 ;
      LAYER pwell ;
        RECT 104.250 149.270 104.670 149.280 ;
        RECT 147.190 148.660 148.500 149.520 ;
      LAYER nwell ;
        RECT 49.760 148.050 50.610 148.140 ;
      LAYER pwell ;
        RECT 2.670 146.430 3.570 147.960 ;
      LAYER nwell ;
        RECT 150.100 147.950 152.020 150.210 ;
      LAYER pwell ;
        RECT 239.470 149.410 240.370 150.940 ;
        RECT 249.310 150.360 250.620 151.220 ;
      LAYER nwell ;
        RECT 252.220 149.650 254.140 151.910 ;
        RECT 282.070 150.490 283.980 152.720 ;
      LAYER pwell ;
        RECT 340.520 152.630 341.420 153.570 ;
        RECT 340.510 152.370 341.420 152.630 ;
        RECT 285.710 151.190 287.020 152.050 ;
        RECT 340.510 151.470 341.410 152.370 ;
      LAYER nwell ;
        RECT 350.280 151.870 352.190 154.100 ;
        RECT 369.050 153.440 370.970 155.700 ;
      LAYER pwell ;
        RECT 353.920 152.570 355.230 153.430 ;
      LAYER nwell ;
        RECT 370.020 153.350 370.870 153.440 ;
        RECT 383.600 152.530 384.450 152.640 ;
        RECT 253.190 149.560 254.040 149.650 ;
      LAYER pwell ;
        RECT 239.470 149.400 239.890 149.410 ;
        RECT 282.410 148.790 283.720 149.650 ;
      LAYER nwell ;
        RECT 285.320 148.080 287.240 150.340 ;
      LAYER pwell ;
        RECT 340.780 149.220 341.680 150.750 ;
        RECT 350.620 150.170 351.930 151.030 ;
      LAYER nwell ;
        RECT 353.530 149.460 355.450 151.720 ;
        RECT 383.380 150.300 385.290 152.530 ;
      LAYER pwell ;
        RECT 387.020 151.000 388.330 151.860 ;
      LAYER nwell ;
        RECT 354.500 149.370 355.350 149.460 ;
      LAYER pwell ;
        RECT 340.780 149.210 341.200 149.220 ;
        RECT 383.720 148.600 385.030 149.460 ;
      LAYER nwell ;
        RECT 286.290 147.990 287.140 148.080 ;
        RECT 151.070 147.860 151.920 147.950 ;
      LAYER pwell ;
        RECT 2.670 146.420 3.090 146.430 ;
      LAYER nwell ;
        RECT 12.330 146.330 13.180 146.440 ;
      LAYER pwell ;
        RECT 2.550 143.860 3.450 144.800 ;
      LAYER nwell ;
        RECT 12.110 144.100 14.020 146.330 ;
      LAYER pwell ;
        RECT 103.980 146.240 104.880 147.770 ;
        RECT 239.200 146.370 240.100 147.900 ;
      LAYER nwell ;
        RECT 386.630 147.890 388.550 150.150 ;
        RECT 387.600 147.800 388.450 147.890 ;
      LAYER pwell ;
        RECT 239.200 146.360 239.620 146.370 ;
      LAYER nwell ;
        RECT 248.860 146.270 249.710 146.380 ;
      LAYER pwell ;
        RECT 103.980 146.230 104.400 146.240 ;
      LAYER nwell ;
        RECT 113.640 146.140 114.490 146.250 ;
      LAYER pwell ;
        RECT 15.750 144.800 17.060 145.660 ;
        RECT 2.540 143.600 3.450 143.860 ;
        RECT 2.540 142.700 3.440 143.600 ;
        RECT 2.510 141.620 3.410 142.560 ;
        RECT 12.450 142.400 13.760 143.260 ;
      LAYER nwell ;
        RECT 15.360 141.690 17.280 143.950 ;
        RECT 28.010 143.910 28.860 144.020 ;
      LAYER pwell ;
        RECT 2.500 141.360 3.410 141.620 ;
      LAYER nwell ;
        RECT 16.330 141.600 17.180 141.690 ;
        RECT 27.790 141.680 29.700 143.910 ;
      LAYER pwell ;
        RECT 103.860 143.670 104.760 144.610 ;
      LAYER nwell ;
        RECT 113.420 143.910 115.330 146.140 ;
      LAYER pwell ;
        RECT 117.060 144.610 118.370 145.470 ;
        RECT 103.850 143.410 104.760 143.670 ;
        RECT 31.430 142.380 32.740 143.240 ;
        RECT 103.850 142.510 104.750 143.410 ;
        RECT 2.500 140.460 3.400 141.360 ;
      LAYER nwell ;
        RECT 12.490 139.930 13.340 140.040 ;
      LAYER pwell ;
        RECT 28.130 139.980 29.440 140.840 ;
        RECT 2.510 138.460 3.410 139.400 ;
        RECT 2.500 138.200 3.410 138.460 ;
        RECT 2.500 137.300 3.400 138.200 ;
      LAYER nwell ;
        RECT 12.270 137.700 14.180 139.930 ;
        RECT 31.040 139.270 32.960 141.530 ;
      LAYER pwell ;
        RECT 103.820 141.430 104.720 142.370 ;
        RECT 113.760 142.210 115.070 143.070 ;
      LAYER nwell ;
        RECT 116.670 141.500 118.590 143.760 ;
        RECT 129.320 143.720 130.170 143.830 ;
      LAYER pwell ;
        RECT 239.080 143.800 239.980 144.740 ;
      LAYER nwell ;
        RECT 248.640 144.040 250.550 146.270 ;
      LAYER pwell ;
        RECT 340.510 146.180 341.410 147.710 ;
        RECT 340.510 146.170 340.930 146.180 ;
      LAYER nwell ;
        RECT 350.170 146.080 351.020 146.190 ;
      LAYER pwell ;
        RECT 252.280 144.740 253.590 145.600 ;
        RECT 103.810 141.170 104.720 141.430 ;
      LAYER nwell ;
        RECT 117.640 141.410 118.490 141.500 ;
        RECT 129.100 141.490 131.010 143.720 ;
      LAYER pwell ;
        RECT 239.070 143.540 239.980 143.800 ;
        RECT 132.740 142.190 134.050 143.050 ;
        RECT 239.070 142.640 239.970 143.540 ;
        RECT 239.040 141.560 239.940 142.500 ;
        RECT 248.980 142.340 250.290 143.200 ;
      LAYER nwell ;
        RECT 251.890 141.630 253.810 143.890 ;
        RECT 264.540 143.850 265.390 143.960 ;
      LAYER pwell ;
        RECT 103.810 140.270 104.710 141.170 ;
      LAYER nwell ;
        RECT 113.800 139.740 114.650 139.850 ;
      LAYER pwell ;
        RECT 129.440 139.790 130.750 140.650 ;
        RECT 15.910 138.400 17.220 139.260 ;
      LAYER nwell ;
        RECT 32.010 139.180 32.860 139.270 ;
      LAYER pwell ;
        RECT 103.820 138.270 104.720 139.210 ;
        RECT 103.810 138.010 104.720 138.270 ;
        RECT 2.770 135.050 3.670 136.580 ;
        RECT 12.610 136.000 13.920 136.860 ;
      LAYER nwell ;
        RECT 15.520 135.290 17.440 137.550 ;
        RECT 94.200 137.320 95.050 137.430 ;
        RECT 16.490 135.200 17.340 135.290 ;
        RECT 93.980 135.090 95.890 137.320 ;
      LAYER pwell ;
        RECT 103.810 137.110 104.710 138.010 ;
      LAYER nwell ;
        RECT 113.580 137.510 115.490 139.740 ;
        RECT 132.350 139.080 134.270 141.340 ;
      LAYER pwell ;
        RECT 239.030 141.300 239.940 141.560 ;
      LAYER nwell ;
        RECT 252.860 141.540 253.710 141.630 ;
        RECT 264.320 141.620 266.230 143.850 ;
      LAYER pwell ;
        RECT 340.390 143.610 341.290 144.550 ;
      LAYER nwell ;
        RECT 349.950 143.850 351.860 146.080 ;
      LAYER pwell ;
        RECT 353.590 144.550 354.900 145.410 ;
        RECT 340.380 143.350 341.290 143.610 ;
        RECT 267.960 142.320 269.270 143.180 ;
        RECT 340.380 142.450 341.280 143.350 ;
        RECT 239.030 140.400 239.930 141.300 ;
      LAYER nwell ;
        RECT 249.020 139.870 249.870 139.980 ;
      LAYER pwell ;
        RECT 264.660 139.920 265.970 140.780 ;
      LAYER nwell ;
        RECT 221.790 139.460 222.640 139.570 ;
      LAYER pwell ;
        RECT 117.220 138.210 118.530 139.070 ;
      LAYER nwell ;
        RECT 133.320 138.990 134.170 139.080 ;
      LAYER pwell ;
        RECT 97.620 135.790 98.930 136.650 ;
        RECT 2.770 135.040 3.190 135.050 ;
        RECT 94.320 133.390 95.630 134.250 ;
      LAYER nwell ;
        RECT 97.230 132.680 99.150 134.940 ;
      LAYER pwell ;
        RECT 104.080 134.860 104.980 136.390 ;
        RECT 113.920 135.810 115.230 136.670 ;
      LAYER nwell ;
        RECT 116.830 135.100 118.750 137.360 ;
        RECT 195.510 137.130 196.360 137.240 ;
        RECT 221.570 137.230 223.480 139.460 ;
      LAYER pwell ;
        RECT 225.210 137.930 226.520 138.790 ;
        RECT 239.040 138.400 239.940 139.340 ;
        RECT 239.030 138.140 239.940 138.400 ;
        RECT 239.030 137.240 239.930 138.140 ;
      LAYER nwell ;
        RECT 248.800 137.640 250.710 139.870 ;
        RECT 267.570 139.210 269.490 141.470 ;
      LAYER pwell ;
        RECT 340.350 141.370 341.250 142.310 ;
        RECT 350.290 142.150 351.600 143.010 ;
      LAYER nwell ;
        RECT 353.200 141.440 355.120 143.700 ;
        RECT 365.850 143.660 366.700 143.770 ;
      LAYER pwell ;
        RECT 340.340 141.110 341.250 141.370 ;
      LAYER nwell ;
        RECT 354.170 141.350 355.020 141.440 ;
        RECT 365.630 141.430 367.540 143.660 ;
      LAYER pwell ;
        RECT 369.270 142.130 370.580 142.990 ;
        RECT 340.340 140.210 341.240 141.110 ;
      LAYER nwell ;
        RECT 350.330 139.680 351.180 139.790 ;
      LAYER pwell ;
        RECT 365.970 139.730 367.280 140.590 ;
        RECT 252.440 138.340 253.750 139.200 ;
      LAYER nwell ;
        RECT 268.540 139.120 269.390 139.210 ;
      LAYER pwell ;
        RECT 340.350 138.210 341.250 139.150 ;
        RECT 340.340 137.950 341.250 138.210 ;
      LAYER nwell ;
        RECT 117.800 135.010 118.650 135.100 ;
        RECT 195.290 134.900 197.200 137.130 ;
      LAYER pwell ;
        RECT 198.930 135.600 200.240 136.460 ;
        RECT 221.910 135.530 223.220 136.390 ;
        RECT 104.080 134.850 104.500 134.860 ;
      LAYER nwell ;
        RECT 224.820 134.820 226.740 137.080 ;
      LAYER pwell ;
        RECT 239.300 134.990 240.200 136.520 ;
        RECT 249.140 135.940 250.450 136.800 ;
      LAYER nwell ;
        RECT 252.050 135.230 253.970 137.490 ;
        RECT 330.730 137.260 331.580 137.370 ;
        RECT 253.020 135.140 253.870 135.230 ;
        RECT 330.510 135.030 332.420 137.260 ;
      LAYER pwell ;
        RECT 340.340 137.050 341.240 137.950 ;
      LAYER nwell ;
        RECT 350.110 137.450 352.020 139.680 ;
        RECT 368.880 139.020 370.800 141.280 ;
        RECT 458.320 139.400 459.170 139.510 ;
      LAYER pwell ;
        RECT 353.750 138.150 355.060 139.010 ;
      LAYER nwell ;
        RECT 369.850 138.930 370.700 139.020 ;
      LAYER pwell ;
        RECT 334.150 135.730 335.460 136.590 ;
        RECT 239.300 134.980 239.720 134.990 ;
        RECT 195.630 133.200 196.940 134.060 ;
      LAYER nwell ;
        RECT 98.200 132.590 99.050 132.680 ;
        RECT 198.540 132.490 200.460 134.750 ;
        RECT 225.790 134.730 226.640 134.820 ;
      LAYER pwell ;
        RECT 330.850 133.330 332.160 134.190 ;
      LAYER nwell ;
        RECT 333.760 132.620 335.680 134.880 ;
      LAYER pwell ;
        RECT 340.610 134.800 341.510 136.330 ;
        RECT 350.450 135.750 351.760 136.610 ;
      LAYER nwell ;
        RECT 353.360 135.040 355.280 137.300 ;
        RECT 432.040 137.070 432.890 137.180 ;
        RECT 458.100 137.170 460.010 139.400 ;
      LAYER pwell ;
        RECT 461.740 137.870 463.050 138.730 ;
      LAYER nwell ;
        RECT 354.330 134.950 355.180 135.040 ;
        RECT 431.820 134.840 433.730 137.070 ;
      LAYER pwell ;
        RECT 435.460 135.540 436.770 136.400 ;
        RECT 458.440 135.470 459.750 136.330 ;
        RECT 340.610 134.790 341.030 134.800 ;
      LAYER nwell ;
        RECT 461.350 134.760 463.270 137.020 ;
      LAYER pwell ;
        RECT 479.040 135.520 480.350 136.380 ;
        RECT 432.160 133.140 433.470 134.000 ;
      LAYER nwell ;
        RECT 334.730 132.530 335.580 132.620 ;
        RECT 199.510 132.400 200.360 132.490 ;
        RECT 435.070 132.430 436.990 134.690 ;
        RECT 462.320 134.670 463.170 134.760 ;
      LAYER pwell ;
        RECT 475.740 133.120 477.050 133.980 ;
      LAYER nwell ;
        RECT 436.040 132.340 436.890 132.430 ;
      LAYER pwell ;
        RECT 1.180 131.470 2.710 131.950 ;
        RECT 1.180 131.050 2.720 131.470 ;
        RECT 102.490 131.280 104.020 131.760 ;
        RECT 237.710 131.410 239.240 131.890 ;
        RECT 102.490 130.860 104.030 131.280 ;
        RECT 237.710 130.990 239.250 131.410 ;
        RECT 339.020 131.220 340.550 131.700 ;
        RECT 339.020 130.800 340.560 131.220 ;
      LAYER nwell ;
        RECT 12.380 130.500 13.230 130.610 ;
      LAYER pwell ;
        RECT 2.600 128.030 3.500 128.970 ;
      LAYER nwell ;
        RECT 12.160 128.270 14.070 130.500 ;
        RECT 248.910 130.440 249.760 130.550 ;
        RECT 113.690 130.310 114.540 130.420 ;
      LAYER pwell ;
        RECT 15.800 128.970 17.110 129.830 ;
        RECT 2.590 127.770 3.500 128.030 ;
        RECT 2.590 126.870 3.490 127.770 ;
        RECT 2.560 125.790 3.460 126.730 ;
        RECT 12.500 126.570 13.810 127.430 ;
      LAYER nwell ;
        RECT 15.410 125.860 17.330 128.120 ;
        RECT 28.060 128.080 28.910 128.190 ;
      LAYER pwell ;
        RECT 2.550 125.530 3.460 125.790 ;
      LAYER nwell ;
        RECT 16.380 125.770 17.230 125.860 ;
        RECT 27.840 125.850 29.750 128.080 ;
      LAYER pwell ;
        RECT 103.910 127.840 104.810 128.780 ;
      LAYER nwell ;
        RECT 113.470 128.080 115.380 130.310 ;
      LAYER pwell ;
        RECT 117.110 128.780 118.420 129.640 ;
        RECT 103.900 127.580 104.810 127.840 ;
        RECT 31.480 126.550 32.790 127.410 ;
        RECT 103.900 126.680 104.800 127.580 ;
        RECT 2.550 124.630 3.450 125.530 ;
      LAYER nwell ;
        RECT 12.540 124.100 13.390 124.210 ;
      LAYER pwell ;
        RECT 28.180 124.150 29.490 125.010 ;
        RECT 2.560 122.630 3.460 123.570 ;
        RECT 2.550 122.370 3.460 122.630 ;
        RECT 2.550 121.470 3.450 122.370 ;
      LAYER nwell ;
        RECT 12.320 121.870 14.230 124.100 ;
        RECT 31.090 123.440 33.010 125.700 ;
      LAYER pwell ;
        RECT 103.870 125.600 104.770 126.540 ;
        RECT 113.810 126.380 115.120 127.240 ;
      LAYER nwell ;
        RECT 116.720 125.670 118.640 127.930 ;
        RECT 129.370 127.890 130.220 128.000 ;
      LAYER pwell ;
        RECT 239.130 127.970 240.030 128.910 ;
      LAYER nwell ;
        RECT 248.690 128.210 250.600 130.440 ;
        RECT 350.220 130.250 351.070 130.360 ;
      LAYER pwell ;
        RECT 252.330 128.910 253.640 129.770 ;
        RECT 103.860 125.340 104.770 125.600 ;
      LAYER nwell ;
        RECT 117.690 125.580 118.540 125.670 ;
        RECT 129.150 125.660 131.060 127.890 ;
      LAYER pwell ;
        RECT 239.120 127.710 240.030 127.970 ;
        RECT 132.790 126.360 134.100 127.220 ;
        RECT 239.120 126.810 240.020 127.710 ;
        RECT 239.090 125.730 239.990 126.670 ;
        RECT 249.030 126.510 250.340 127.370 ;
      LAYER nwell ;
        RECT 251.940 125.800 253.860 128.060 ;
        RECT 264.590 128.020 265.440 128.130 ;
      LAYER pwell ;
        RECT 103.860 124.440 104.760 125.340 ;
      LAYER nwell ;
        RECT 113.850 123.910 114.700 124.020 ;
      LAYER pwell ;
        RECT 129.490 123.960 130.800 124.820 ;
        RECT 15.960 122.570 17.270 123.430 ;
      LAYER nwell ;
        RECT 32.060 123.350 32.910 123.440 ;
        RECT 45.640 122.530 46.490 122.640 ;
      LAYER pwell ;
        RECT 2.820 119.220 3.720 120.750 ;
        RECT 12.660 120.170 13.970 121.030 ;
      LAYER nwell ;
        RECT 15.570 119.460 17.490 121.720 ;
        RECT 45.420 120.300 47.330 122.530 ;
      LAYER pwell ;
        RECT 103.870 122.440 104.770 123.380 ;
        RECT 103.860 122.180 104.770 122.440 ;
        RECT 49.060 121.000 50.370 121.860 ;
        RECT 103.860 121.280 104.760 122.180 ;
      LAYER nwell ;
        RECT 113.630 121.680 115.540 123.910 ;
        RECT 132.400 123.250 134.320 125.510 ;
      LAYER pwell ;
        RECT 239.080 125.470 239.990 125.730 ;
      LAYER nwell ;
        RECT 252.910 125.710 253.760 125.800 ;
        RECT 264.370 125.790 266.280 128.020 ;
      LAYER pwell ;
        RECT 340.440 127.780 341.340 128.720 ;
      LAYER nwell ;
        RECT 350.000 128.020 351.910 130.250 ;
      LAYER pwell ;
        RECT 353.640 128.720 354.950 129.580 ;
        RECT 340.430 127.520 341.340 127.780 ;
        RECT 268.010 126.490 269.320 127.350 ;
        RECT 340.430 126.620 341.330 127.520 ;
        RECT 239.080 124.570 239.980 125.470 ;
      LAYER nwell ;
        RECT 249.070 124.040 249.920 124.150 ;
      LAYER pwell ;
        RECT 264.710 124.090 266.020 124.950 ;
        RECT 117.270 122.380 118.580 123.240 ;
      LAYER nwell ;
        RECT 133.370 123.160 134.220 123.250 ;
      LAYER pwell ;
        RECT 239.090 122.570 239.990 123.510 ;
      LAYER nwell ;
        RECT 146.950 122.340 147.800 122.450 ;
        RECT 16.540 119.370 17.390 119.460 ;
      LAYER pwell ;
        RECT 2.820 119.210 3.240 119.220 ;
        RECT 45.760 118.600 47.070 119.460 ;
      LAYER nwell ;
        RECT 48.670 117.890 50.590 120.150 ;
      LAYER pwell ;
        RECT 104.130 119.030 105.030 120.560 ;
        RECT 113.970 119.980 115.280 120.840 ;
      LAYER nwell ;
        RECT 116.880 119.270 118.800 121.530 ;
        RECT 146.730 120.110 148.640 122.340 ;
      LAYER pwell ;
        RECT 239.080 122.310 239.990 122.570 ;
        RECT 150.370 120.810 151.680 121.670 ;
        RECT 239.080 121.410 239.980 122.310 ;
      LAYER nwell ;
        RECT 248.850 121.810 250.760 124.040 ;
        RECT 267.620 123.380 269.540 125.640 ;
      LAYER pwell ;
        RECT 340.400 125.540 341.300 126.480 ;
        RECT 350.340 126.320 351.650 127.180 ;
      LAYER nwell ;
        RECT 353.250 125.610 355.170 127.870 ;
        RECT 365.900 127.830 366.750 127.940 ;
      LAYER pwell ;
        RECT 340.390 125.280 341.300 125.540 ;
      LAYER nwell ;
        RECT 354.220 125.520 355.070 125.610 ;
        RECT 365.680 125.600 367.590 127.830 ;
      LAYER pwell ;
        RECT 369.320 126.300 370.630 127.160 ;
        RECT 340.390 124.380 341.290 125.280 ;
      LAYER nwell ;
        RECT 350.380 123.850 351.230 123.960 ;
      LAYER pwell ;
        RECT 366.020 123.900 367.330 124.760 ;
        RECT 252.490 122.510 253.800 123.370 ;
      LAYER nwell ;
        RECT 268.590 123.290 269.440 123.380 ;
        RECT 282.170 122.470 283.020 122.580 ;
        RECT 117.850 119.180 118.700 119.270 ;
      LAYER pwell ;
        RECT 104.130 119.020 104.550 119.030 ;
        RECT 147.070 118.410 148.380 119.270 ;
      LAYER nwell ;
        RECT 49.640 117.800 50.490 117.890 ;
      LAYER pwell ;
        RECT 2.550 116.180 3.450 117.710 ;
      LAYER nwell ;
        RECT 149.980 117.700 151.900 119.960 ;
      LAYER pwell ;
        RECT 239.350 119.160 240.250 120.690 ;
        RECT 249.190 120.110 250.500 120.970 ;
      LAYER nwell ;
        RECT 252.100 119.400 254.020 121.660 ;
        RECT 281.950 120.240 283.860 122.470 ;
      LAYER pwell ;
        RECT 340.400 122.380 341.300 123.320 ;
        RECT 340.390 122.120 341.300 122.380 ;
        RECT 285.590 120.940 286.900 121.800 ;
        RECT 340.390 121.220 341.290 122.120 ;
      LAYER nwell ;
        RECT 350.160 121.620 352.070 123.850 ;
        RECT 368.930 123.190 370.850 125.450 ;
      LAYER pwell ;
        RECT 353.800 122.320 355.110 123.180 ;
      LAYER nwell ;
        RECT 369.900 123.100 370.750 123.190 ;
        RECT 383.480 122.280 384.330 122.390 ;
        RECT 253.070 119.310 253.920 119.400 ;
      LAYER pwell ;
        RECT 239.350 119.150 239.770 119.160 ;
        RECT 282.290 118.540 283.600 119.400 ;
      LAYER nwell ;
        RECT 285.200 117.830 287.120 120.090 ;
      LAYER pwell ;
        RECT 340.660 118.970 341.560 120.500 ;
        RECT 350.500 119.920 351.810 120.780 ;
      LAYER nwell ;
        RECT 353.410 119.210 355.330 121.470 ;
        RECT 383.260 120.050 385.170 122.280 ;
      LAYER pwell ;
        RECT 386.900 120.750 388.210 121.610 ;
      LAYER nwell ;
        RECT 354.380 119.120 355.230 119.210 ;
      LAYER pwell ;
        RECT 340.660 118.960 341.080 118.970 ;
        RECT 383.600 118.350 384.910 119.210 ;
      LAYER nwell ;
        RECT 286.170 117.740 287.020 117.830 ;
        RECT 150.950 117.610 151.800 117.700 ;
      LAYER pwell ;
        RECT 2.550 116.170 2.970 116.180 ;
      LAYER nwell ;
        RECT 12.210 116.080 13.060 116.190 ;
      LAYER pwell ;
        RECT 2.430 113.610 3.330 114.550 ;
      LAYER nwell ;
        RECT 11.990 113.850 13.900 116.080 ;
      LAYER pwell ;
        RECT 103.860 115.990 104.760 117.520 ;
        RECT 239.080 116.120 239.980 117.650 ;
      LAYER nwell ;
        RECT 386.510 117.640 388.430 119.900 ;
        RECT 387.480 117.550 388.330 117.640 ;
      LAYER pwell ;
        RECT 239.080 116.110 239.500 116.120 ;
      LAYER nwell ;
        RECT 248.740 116.020 249.590 116.130 ;
      LAYER pwell ;
        RECT 103.860 115.980 104.280 115.990 ;
      LAYER nwell ;
        RECT 113.520 115.890 114.370 116.000 ;
      LAYER pwell ;
        RECT 15.630 114.550 16.940 115.410 ;
        RECT 2.420 113.350 3.330 113.610 ;
        RECT 2.420 112.450 3.320 113.350 ;
        RECT 2.390 111.370 3.290 112.310 ;
        RECT 12.330 112.150 13.640 113.010 ;
      LAYER nwell ;
        RECT 15.240 111.440 17.160 113.700 ;
        RECT 27.890 113.660 28.740 113.770 ;
      LAYER pwell ;
        RECT 2.380 111.110 3.290 111.370 ;
      LAYER nwell ;
        RECT 16.210 111.350 17.060 111.440 ;
        RECT 27.670 111.430 29.580 113.660 ;
      LAYER pwell ;
        RECT 103.740 113.420 104.640 114.360 ;
      LAYER nwell ;
        RECT 113.300 113.660 115.210 115.890 ;
      LAYER pwell ;
        RECT 116.940 114.360 118.250 115.220 ;
        RECT 103.730 113.160 104.640 113.420 ;
        RECT 31.310 112.130 32.620 112.990 ;
        RECT 103.730 112.260 104.630 113.160 ;
        RECT 2.380 110.210 3.280 111.110 ;
      LAYER nwell ;
        RECT 12.370 109.680 13.220 109.790 ;
      LAYER pwell ;
        RECT 28.010 109.730 29.320 110.590 ;
        RECT 2.390 108.210 3.290 109.150 ;
        RECT 2.380 107.950 3.290 108.210 ;
        RECT 2.380 107.050 3.280 107.950 ;
      LAYER nwell ;
        RECT 12.150 107.450 14.060 109.680 ;
        RECT 30.920 109.020 32.840 111.280 ;
      LAYER pwell ;
        RECT 103.700 111.180 104.600 112.120 ;
        RECT 113.640 111.960 114.950 112.820 ;
      LAYER nwell ;
        RECT 116.550 111.250 118.470 113.510 ;
        RECT 129.200 113.470 130.050 113.580 ;
      LAYER pwell ;
        RECT 238.960 113.550 239.860 114.490 ;
      LAYER nwell ;
        RECT 248.520 113.790 250.430 116.020 ;
      LAYER pwell ;
        RECT 340.390 115.930 341.290 117.460 ;
        RECT 340.390 115.920 340.810 115.930 ;
      LAYER nwell ;
        RECT 350.050 115.830 350.900 115.940 ;
      LAYER pwell ;
        RECT 252.160 114.490 253.470 115.350 ;
        RECT 103.690 110.920 104.600 111.180 ;
      LAYER nwell ;
        RECT 117.520 111.160 118.370 111.250 ;
        RECT 128.980 111.240 130.890 113.470 ;
      LAYER pwell ;
        RECT 238.950 113.290 239.860 113.550 ;
        RECT 132.620 111.940 133.930 112.800 ;
        RECT 238.950 112.390 239.850 113.290 ;
        RECT 238.920 111.310 239.820 112.250 ;
        RECT 248.860 112.090 250.170 112.950 ;
      LAYER nwell ;
        RECT 251.770 111.380 253.690 113.640 ;
        RECT 264.420 113.600 265.270 113.710 ;
      LAYER pwell ;
        RECT 103.690 110.020 104.590 110.920 ;
      LAYER nwell ;
        RECT 113.680 109.490 114.530 109.600 ;
      LAYER pwell ;
        RECT 129.320 109.540 130.630 110.400 ;
        RECT 15.790 108.150 17.100 109.010 ;
      LAYER nwell ;
        RECT 31.890 108.930 32.740 109.020 ;
      LAYER pwell ;
        RECT 103.700 108.020 104.600 108.960 ;
        RECT 103.690 107.760 104.600 108.020 ;
        RECT 2.650 104.800 3.550 106.330 ;
        RECT 12.490 105.750 13.800 106.610 ;
      LAYER nwell ;
        RECT 15.400 105.040 17.320 107.300 ;
      LAYER pwell ;
        RECT 103.690 106.860 104.590 107.760 ;
      LAYER nwell ;
        RECT 113.460 107.260 115.370 109.490 ;
        RECT 132.230 108.830 134.150 111.090 ;
      LAYER pwell ;
        RECT 238.910 111.050 239.820 111.310 ;
      LAYER nwell ;
        RECT 252.740 111.290 253.590 111.380 ;
        RECT 264.200 111.370 266.110 113.600 ;
      LAYER pwell ;
        RECT 340.270 113.360 341.170 114.300 ;
      LAYER nwell ;
        RECT 349.830 113.600 351.740 115.830 ;
      LAYER pwell ;
        RECT 353.470 114.300 354.780 115.160 ;
        RECT 340.260 113.100 341.170 113.360 ;
        RECT 267.840 112.070 269.150 112.930 ;
        RECT 340.260 112.200 341.160 113.100 ;
        RECT 238.910 110.150 239.810 111.050 ;
      LAYER nwell ;
        RECT 248.900 109.620 249.750 109.730 ;
      LAYER pwell ;
        RECT 264.540 109.670 265.850 110.530 ;
        RECT 117.100 107.960 118.410 108.820 ;
      LAYER nwell ;
        RECT 133.200 108.740 134.050 108.830 ;
      LAYER pwell ;
        RECT 238.920 108.150 239.820 109.090 ;
        RECT 238.910 107.890 239.820 108.150 ;
      LAYER nwell ;
        RECT 63.170 106.510 64.020 106.620 ;
        RECT 16.370 104.950 17.220 105.040 ;
      LAYER pwell ;
        RECT 2.650 104.790 3.070 104.800 ;
      LAYER nwell ;
        RECT 62.950 104.280 64.860 106.510 ;
      LAYER pwell ;
        RECT 66.590 104.980 67.900 105.840 ;
        RECT 103.960 104.610 104.860 106.140 ;
        RECT 113.800 105.560 115.110 106.420 ;
      LAYER nwell ;
        RECT 116.710 104.850 118.630 107.110 ;
      LAYER pwell ;
        RECT 238.910 106.990 239.810 107.890 ;
      LAYER nwell ;
        RECT 248.680 107.390 250.590 109.620 ;
        RECT 267.450 108.960 269.370 111.220 ;
      LAYER pwell ;
        RECT 340.230 111.120 341.130 112.060 ;
        RECT 350.170 111.900 351.480 112.760 ;
      LAYER nwell ;
        RECT 353.080 111.190 355.000 113.450 ;
        RECT 365.730 113.410 366.580 113.520 ;
      LAYER pwell ;
        RECT 340.220 110.860 341.130 111.120 ;
      LAYER nwell ;
        RECT 354.050 111.100 354.900 111.190 ;
        RECT 365.510 111.180 367.420 113.410 ;
      LAYER pwell ;
        RECT 369.150 111.880 370.460 112.740 ;
        RECT 340.220 109.960 341.120 110.860 ;
      LAYER nwell ;
        RECT 350.210 109.430 351.060 109.540 ;
      LAYER pwell ;
        RECT 365.850 109.480 367.160 110.340 ;
        RECT 252.320 108.090 253.630 108.950 ;
      LAYER nwell ;
        RECT 268.420 108.870 269.270 108.960 ;
      LAYER pwell ;
        RECT 340.230 107.960 341.130 108.900 ;
        RECT 340.220 107.700 341.130 107.960 ;
      LAYER nwell ;
        RECT 164.480 106.320 165.330 106.430 ;
        RECT 117.680 104.760 118.530 104.850 ;
      LAYER pwell ;
        RECT 103.960 104.600 104.380 104.610 ;
        RECT 63.290 102.580 64.600 103.440 ;
        RECT 3.240 102.480 3.660 102.490 ;
        RECT 2.760 100.950 3.660 102.480 ;
      LAYER nwell ;
        RECT 66.200 101.870 68.120 104.130 ;
        RECT 164.260 104.090 166.170 106.320 ;
      LAYER pwell ;
        RECT 167.900 104.790 169.210 105.650 ;
        RECT 239.180 104.740 240.080 106.270 ;
        RECT 249.020 105.690 250.330 106.550 ;
      LAYER nwell ;
        RECT 251.930 104.980 253.850 107.240 ;
      LAYER pwell ;
        RECT 340.220 106.800 341.120 107.700 ;
      LAYER nwell ;
        RECT 349.990 107.200 351.900 109.430 ;
        RECT 368.760 108.770 370.680 111.030 ;
      LAYER pwell ;
        RECT 353.630 107.900 354.940 108.760 ;
      LAYER nwell ;
        RECT 369.730 108.680 370.580 108.770 ;
        RECT 299.700 106.450 300.550 106.560 ;
        RECT 252.900 104.890 253.750 104.980 ;
      LAYER pwell ;
        RECT 239.180 104.730 239.600 104.740 ;
      LAYER nwell ;
        RECT 299.480 104.220 301.390 106.450 ;
      LAYER pwell ;
        RECT 303.120 104.920 304.430 105.780 ;
        RECT 340.490 104.550 341.390 106.080 ;
        RECT 350.330 105.500 351.640 106.360 ;
      LAYER nwell ;
        RECT 353.240 104.790 355.160 107.050 ;
        RECT 401.010 106.260 401.860 106.370 ;
        RECT 354.210 104.700 355.060 104.790 ;
      LAYER pwell ;
        RECT 340.490 104.540 340.910 104.550 ;
        RECT 164.600 102.390 165.910 103.250 ;
        RECT 104.550 102.290 104.970 102.300 ;
      LAYER nwell ;
        RECT 67.170 101.780 68.020 101.870 ;
      LAYER pwell ;
        RECT 104.070 100.760 104.970 102.290 ;
      LAYER nwell ;
        RECT 167.510 101.680 169.430 103.940 ;
      LAYER pwell ;
        RECT 299.820 102.520 301.130 103.380 ;
        RECT 239.770 102.420 240.190 102.430 ;
      LAYER nwell ;
        RECT 168.480 101.590 169.330 101.680 ;
      LAYER pwell ;
        RECT 239.290 100.890 240.190 102.420 ;
      LAYER nwell ;
        RECT 302.730 101.810 304.650 104.070 ;
        RECT 400.790 104.030 402.700 106.260 ;
      LAYER pwell ;
        RECT 404.430 104.730 405.740 105.590 ;
        RECT 401.130 102.330 402.440 103.190 ;
        RECT 341.080 102.230 341.500 102.240 ;
      LAYER nwell ;
        RECT 303.700 101.720 304.550 101.810 ;
      LAYER pwell ;
        RECT 340.600 100.700 341.500 102.230 ;
      LAYER nwell ;
        RECT 404.040 101.620 405.960 103.880 ;
        RECT 405.010 101.530 405.860 101.620 ;
        RECT 12.350 100.430 13.200 100.540 ;
      LAYER pwell ;
        RECT 2.570 97.960 3.470 98.900 ;
      LAYER nwell ;
        RECT 12.130 98.200 14.040 100.430 ;
        RECT 248.880 100.370 249.730 100.480 ;
        RECT 113.660 100.240 114.510 100.350 ;
      LAYER pwell ;
        RECT 15.770 98.900 17.080 99.760 ;
        RECT 2.560 97.700 3.470 97.960 ;
        RECT 2.560 96.800 3.460 97.700 ;
        RECT 2.530 95.720 3.430 96.660 ;
        RECT 12.470 96.500 13.780 97.360 ;
      LAYER nwell ;
        RECT 15.380 95.790 17.300 98.050 ;
        RECT 28.030 98.010 28.880 98.120 ;
      LAYER pwell ;
        RECT 2.520 95.460 3.430 95.720 ;
      LAYER nwell ;
        RECT 16.350 95.700 17.200 95.790 ;
        RECT 27.810 95.780 29.720 98.010 ;
      LAYER pwell ;
        RECT 103.880 97.770 104.780 98.710 ;
      LAYER nwell ;
        RECT 113.440 98.010 115.350 100.240 ;
      LAYER pwell ;
        RECT 117.080 98.710 118.390 99.570 ;
        RECT 103.870 97.510 104.780 97.770 ;
        RECT 31.450 96.480 32.760 97.340 ;
        RECT 103.870 96.610 104.770 97.510 ;
        RECT 2.520 94.560 3.420 95.460 ;
      LAYER nwell ;
        RECT 12.510 94.030 13.360 94.140 ;
      LAYER pwell ;
        RECT 28.150 94.080 29.460 94.940 ;
        RECT 2.530 92.560 3.430 93.500 ;
        RECT 2.520 92.300 3.430 92.560 ;
        RECT 2.520 91.400 3.420 92.300 ;
      LAYER nwell ;
        RECT 12.290 91.800 14.200 94.030 ;
        RECT 31.060 93.370 32.980 95.630 ;
      LAYER pwell ;
        RECT 103.840 95.530 104.740 96.470 ;
        RECT 113.780 96.310 115.090 97.170 ;
      LAYER nwell ;
        RECT 116.690 95.600 118.610 97.860 ;
        RECT 129.340 97.820 130.190 97.930 ;
      LAYER pwell ;
        RECT 239.100 97.900 240.000 98.840 ;
      LAYER nwell ;
        RECT 248.660 98.140 250.570 100.370 ;
        RECT 350.190 100.180 351.040 100.290 ;
      LAYER pwell ;
        RECT 252.300 98.840 253.610 99.700 ;
        RECT 103.830 95.270 104.740 95.530 ;
      LAYER nwell ;
        RECT 117.660 95.510 118.510 95.600 ;
        RECT 129.120 95.590 131.030 97.820 ;
      LAYER pwell ;
        RECT 239.090 97.640 240.000 97.900 ;
        RECT 132.760 96.290 134.070 97.150 ;
        RECT 239.090 96.740 239.990 97.640 ;
        RECT 239.060 95.660 239.960 96.600 ;
        RECT 249.000 96.440 250.310 97.300 ;
      LAYER nwell ;
        RECT 251.910 95.730 253.830 97.990 ;
        RECT 264.560 97.950 265.410 98.060 ;
      LAYER pwell ;
        RECT 103.830 94.370 104.730 95.270 ;
      LAYER nwell ;
        RECT 113.820 93.840 114.670 93.950 ;
      LAYER pwell ;
        RECT 129.460 93.890 130.770 94.750 ;
        RECT 15.930 92.500 17.240 93.360 ;
      LAYER nwell ;
        RECT 32.030 93.280 32.880 93.370 ;
        RECT 45.610 92.460 46.460 92.570 ;
      LAYER pwell ;
        RECT 2.790 89.150 3.690 90.680 ;
        RECT 12.630 90.100 13.940 90.960 ;
      LAYER nwell ;
        RECT 15.540 89.390 17.460 91.650 ;
        RECT 45.390 90.230 47.300 92.460 ;
      LAYER pwell ;
        RECT 103.840 92.370 104.740 93.310 ;
        RECT 103.830 92.110 104.740 92.370 ;
        RECT 49.030 90.930 50.340 91.790 ;
        RECT 103.830 91.210 104.730 92.110 ;
      LAYER nwell ;
        RECT 113.600 91.610 115.510 93.840 ;
        RECT 132.370 93.180 134.290 95.440 ;
      LAYER pwell ;
        RECT 239.050 95.400 239.960 95.660 ;
      LAYER nwell ;
        RECT 252.880 95.640 253.730 95.730 ;
        RECT 264.340 95.720 266.250 97.950 ;
      LAYER pwell ;
        RECT 340.410 97.710 341.310 98.650 ;
      LAYER nwell ;
        RECT 349.970 97.950 351.880 100.180 ;
      LAYER pwell ;
        RECT 353.610 98.650 354.920 99.510 ;
        RECT 340.400 97.450 341.310 97.710 ;
        RECT 267.980 96.420 269.290 97.280 ;
        RECT 340.400 96.550 341.300 97.450 ;
        RECT 239.050 94.500 239.950 95.400 ;
      LAYER nwell ;
        RECT 249.040 93.970 249.890 94.080 ;
      LAYER pwell ;
        RECT 264.680 94.020 265.990 94.880 ;
        RECT 117.240 92.310 118.550 93.170 ;
      LAYER nwell ;
        RECT 133.340 93.090 134.190 93.180 ;
      LAYER pwell ;
        RECT 239.060 92.500 239.960 93.440 ;
      LAYER nwell ;
        RECT 146.920 92.270 147.770 92.380 ;
        RECT 16.510 89.300 17.360 89.390 ;
      LAYER pwell ;
        RECT 2.790 89.140 3.210 89.150 ;
        RECT 45.730 88.530 47.040 89.390 ;
      LAYER nwell ;
        RECT 48.640 87.820 50.560 90.080 ;
      LAYER pwell ;
        RECT 104.100 88.960 105.000 90.490 ;
        RECT 113.940 89.910 115.250 90.770 ;
      LAYER nwell ;
        RECT 116.850 89.200 118.770 91.460 ;
        RECT 146.700 90.040 148.610 92.270 ;
      LAYER pwell ;
        RECT 239.050 92.240 239.960 92.500 ;
        RECT 150.340 90.740 151.650 91.600 ;
        RECT 239.050 91.340 239.950 92.240 ;
      LAYER nwell ;
        RECT 248.820 91.740 250.730 93.970 ;
        RECT 267.590 93.310 269.510 95.570 ;
      LAYER pwell ;
        RECT 340.370 95.470 341.270 96.410 ;
        RECT 350.310 96.250 351.620 97.110 ;
      LAYER nwell ;
        RECT 353.220 95.540 355.140 97.800 ;
        RECT 365.870 97.760 366.720 97.870 ;
      LAYER pwell ;
        RECT 340.360 95.210 341.270 95.470 ;
      LAYER nwell ;
        RECT 354.190 95.450 355.040 95.540 ;
        RECT 365.650 95.530 367.560 97.760 ;
      LAYER pwell ;
        RECT 369.290 96.230 370.600 97.090 ;
        RECT 340.360 94.310 341.260 95.210 ;
      LAYER nwell ;
        RECT 350.350 93.780 351.200 93.890 ;
      LAYER pwell ;
        RECT 365.990 93.830 367.300 94.690 ;
        RECT 252.460 92.440 253.770 93.300 ;
      LAYER nwell ;
        RECT 268.560 93.220 269.410 93.310 ;
        RECT 282.140 92.400 282.990 92.510 ;
        RECT 117.820 89.110 118.670 89.200 ;
      LAYER pwell ;
        RECT 104.100 88.950 104.520 88.960 ;
        RECT 147.040 88.340 148.350 89.200 ;
      LAYER nwell ;
        RECT 49.610 87.730 50.460 87.820 ;
      LAYER pwell ;
        RECT 2.520 86.110 3.420 87.640 ;
      LAYER nwell ;
        RECT 149.950 87.630 151.870 89.890 ;
      LAYER pwell ;
        RECT 239.320 89.090 240.220 90.620 ;
        RECT 249.160 90.040 250.470 90.900 ;
      LAYER nwell ;
        RECT 252.070 89.330 253.990 91.590 ;
        RECT 281.920 90.170 283.830 92.400 ;
      LAYER pwell ;
        RECT 340.370 92.310 341.270 93.250 ;
        RECT 340.360 92.050 341.270 92.310 ;
        RECT 285.560 90.870 286.870 91.730 ;
        RECT 340.360 91.150 341.260 92.050 ;
      LAYER nwell ;
        RECT 350.130 91.550 352.040 93.780 ;
        RECT 368.900 93.120 370.820 95.380 ;
      LAYER pwell ;
        RECT 353.770 92.250 355.080 93.110 ;
      LAYER nwell ;
        RECT 369.870 93.030 370.720 93.120 ;
        RECT 383.450 92.210 384.300 92.320 ;
        RECT 253.040 89.240 253.890 89.330 ;
      LAYER pwell ;
        RECT 239.320 89.080 239.740 89.090 ;
        RECT 282.260 88.470 283.570 89.330 ;
      LAYER nwell ;
        RECT 285.170 87.760 287.090 90.020 ;
      LAYER pwell ;
        RECT 340.630 88.900 341.530 90.430 ;
        RECT 350.470 89.850 351.780 90.710 ;
      LAYER nwell ;
        RECT 353.380 89.140 355.300 91.400 ;
        RECT 383.230 89.980 385.140 92.210 ;
      LAYER pwell ;
        RECT 386.870 90.680 388.180 91.540 ;
      LAYER nwell ;
        RECT 354.350 89.050 355.200 89.140 ;
      LAYER pwell ;
        RECT 340.630 88.890 341.050 88.900 ;
        RECT 383.570 88.280 384.880 89.140 ;
      LAYER nwell ;
        RECT 286.140 87.670 286.990 87.760 ;
        RECT 150.920 87.540 151.770 87.630 ;
      LAYER pwell ;
        RECT 2.520 86.100 2.940 86.110 ;
      LAYER nwell ;
        RECT 12.180 86.010 13.030 86.120 ;
      LAYER pwell ;
        RECT 2.400 83.540 3.300 84.480 ;
      LAYER nwell ;
        RECT 11.960 83.780 13.870 86.010 ;
      LAYER pwell ;
        RECT 103.830 85.920 104.730 87.450 ;
        RECT 239.050 86.050 239.950 87.580 ;
      LAYER nwell ;
        RECT 386.480 87.570 388.400 89.830 ;
        RECT 387.450 87.480 388.300 87.570 ;
      LAYER pwell ;
        RECT 239.050 86.040 239.470 86.050 ;
      LAYER nwell ;
        RECT 248.710 85.950 249.560 86.060 ;
      LAYER pwell ;
        RECT 103.830 85.910 104.250 85.920 ;
      LAYER nwell ;
        RECT 113.490 85.820 114.340 85.930 ;
      LAYER pwell ;
        RECT 15.600 84.480 16.910 85.340 ;
        RECT 2.390 83.280 3.300 83.540 ;
        RECT 2.390 82.380 3.290 83.280 ;
        RECT 2.360 81.300 3.260 82.240 ;
        RECT 12.300 82.080 13.610 82.940 ;
      LAYER nwell ;
        RECT 15.210 81.370 17.130 83.630 ;
        RECT 27.860 83.590 28.710 83.700 ;
      LAYER pwell ;
        RECT 2.350 81.040 3.260 81.300 ;
      LAYER nwell ;
        RECT 16.180 81.280 17.030 81.370 ;
        RECT 27.640 81.360 29.550 83.590 ;
      LAYER pwell ;
        RECT 103.710 83.350 104.610 84.290 ;
      LAYER nwell ;
        RECT 113.270 83.590 115.180 85.820 ;
      LAYER pwell ;
        RECT 116.910 84.290 118.220 85.150 ;
        RECT 103.700 83.090 104.610 83.350 ;
        RECT 31.280 82.060 32.590 82.920 ;
        RECT 103.700 82.190 104.600 83.090 ;
        RECT 2.350 80.140 3.250 81.040 ;
      LAYER nwell ;
        RECT 12.340 79.610 13.190 79.720 ;
      LAYER pwell ;
        RECT 27.980 79.660 29.290 80.520 ;
        RECT 2.360 78.140 3.260 79.080 ;
        RECT 2.350 77.880 3.260 78.140 ;
        RECT 2.350 76.980 3.250 77.880 ;
      LAYER nwell ;
        RECT 12.120 77.380 14.030 79.610 ;
        RECT 30.890 78.950 32.810 81.210 ;
      LAYER pwell ;
        RECT 103.670 81.110 104.570 82.050 ;
        RECT 113.610 81.890 114.920 82.750 ;
      LAYER nwell ;
        RECT 116.520 81.180 118.440 83.440 ;
        RECT 129.170 83.400 130.020 83.510 ;
      LAYER pwell ;
        RECT 238.930 83.480 239.830 84.420 ;
      LAYER nwell ;
        RECT 248.490 83.720 250.400 85.950 ;
      LAYER pwell ;
        RECT 340.360 85.860 341.260 87.390 ;
        RECT 340.360 85.850 340.780 85.860 ;
      LAYER nwell ;
        RECT 350.020 85.760 350.870 85.870 ;
      LAYER pwell ;
        RECT 252.130 84.420 253.440 85.280 ;
        RECT 103.660 80.850 104.570 81.110 ;
      LAYER nwell ;
        RECT 117.490 81.090 118.340 81.180 ;
        RECT 128.950 81.170 130.860 83.400 ;
      LAYER pwell ;
        RECT 238.920 83.220 239.830 83.480 ;
        RECT 132.590 81.870 133.900 82.730 ;
        RECT 238.920 82.320 239.820 83.220 ;
        RECT 238.890 81.240 239.790 82.180 ;
        RECT 248.830 82.020 250.140 82.880 ;
      LAYER nwell ;
        RECT 251.740 81.310 253.660 83.570 ;
        RECT 264.390 83.530 265.240 83.640 ;
        RECT 77.370 80.220 78.220 80.330 ;
      LAYER pwell ;
        RECT 15.760 78.080 17.070 78.940 ;
      LAYER nwell ;
        RECT 31.860 78.860 32.710 78.950 ;
        RECT 77.150 77.990 79.060 80.220 ;
      LAYER pwell ;
        RECT 103.660 79.950 104.560 80.850 ;
        RECT 80.790 78.690 82.100 79.550 ;
      LAYER nwell ;
        RECT 113.650 79.420 114.500 79.530 ;
      LAYER pwell ;
        RECT 129.290 79.470 130.600 80.330 ;
        RECT 103.670 77.950 104.570 78.890 ;
        RECT 2.620 74.730 3.520 76.260 ;
        RECT 12.460 75.680 13.770 76.540 ;
      LAYER nwell ;
        RECT 15.370 74.970 17.290 77.230 ;
      LAYER pwell ;
        RECT 77.490 76.290 78.800 77.150 ;
      LAYER nwell ;
        RECT 80.400 75.580 82.320 77.840 ;
      LAYER pwell ;
        RECT 103.660 77.690 104.570 77.950 ;
        RECT 103.660 76.790 104.560 77.690 ;
      LAYER nwell ;
        RECT 113.430 77.190 115.340 79.420 ;
        RECT 132.200 78.760 134.120 81.020 ;
      LAYER pwell ;
        RECT 238.880 80.980 239.790 81.240 ;
      LAYER nwell ;
        RECT 252.710 81.220 253.560 81.310 ;
        RECT 264.170 81.300 266.080 83.530 ;
      LAYER pwell ;
        RECT 340.240 83.290 341.140 84.230 ;
      LAYER nwell ;
        RECT 349.800 83.530 351.710 85.760 ;
      LAYER pwell ;
        RECT 353.440 84.230 354.750 85.090 ;
        RECT 340.230 83.030 341.140 83.290 ;
        RECT 267.810 82.000 269.120 82.860 ;
        RECT 340.230 82.130 341.130 83.030 ;
      LAYER nwell ;
        RECT 178.680 80.030 179.530 80.140 ;
      LAYER pwell ;
        RECT 238.880 80.080 239.780 80.980 ;
        RECT 117.070 77.890 118.380 78.750 ;
      LAYER nwell ;
        RECT 133.170 78.670 134.020 78.760 ;
        RECT 178.460 77.800 180.370 80.030 ;
        RECT 248.870 79.550 249.720 79.660 ;
      LAYER pwell ;
        RECT 264.510 79.600 265.820 80.460 ;
        RECT 182.100 78.500 183.410 79.360 ;
        RECT 238.890 78.080 239.790 79.020 ;
        RECT 238.880 77.820 239.790 78.080 ;
      LAYER nwell ;
        RECT 81.370 75.490 82.220 75.580 ;
        RECT 16.340 74.880 17.190 74.970 ;
      LAYER pwell ;
        RECT 2.620 74.720 3.040 74.730 ;
        RECT 103.930 74.540 104.830 76.070 ;
        RECT 113.770 75.490 115.080 76.350 ;
      LAYER nwell ;
        RECT 116.680 74.780 118.600 77.040 ;
      LAYER pwell ;
        RECT 178.800 76.100 180.110 76.960 ;
      LAYER nwell ;
        RECT 181.710 75.390 183.630 77.650 ;
      LAYER pwell ;
        RECT 238.880 76.920 239.780 77.820 ;
      LAYER nwell ;
        RECT 248.650 77.320 250.560 79.550 ;
        RECT 267.420 78.890 269.340 81.150 ;
      LAYER pwell ;
        RECT 340.200 81.050 341.100 81.990 ;
        RECT 350.140 81.830 351.450 82.690 ;
      LAYER nwell ;
        RECT 353.050 81.120 354.970 83.380 ;
        RECT 365.700 83.340 366.550 83.450 ;
      LAYER pwell ;
        RECT 340.190 80.790 341.100 81.050 ;
      LAYER nwell ;
        RECT 354.020 81.030 354.870 81.120 ;
        RECT 365.480 81.110 367.390 83.340 ;
      LAYER pwell ;
        RECT 369.120 81.810 370.430 82.670 ;
      LAYER nwell ;
        RECT 313.900 80.160 314.750 80.270 ;
      LAYER pwell ;
        RECT 252.290 78.020 253.600 78.880 ;
      LAYER nwell ;
        RECT 268.390 78.800 269.240 78.890 ;
        RECT 313.680 77.930 315.590 80.160 ;
      LAYER pwell ;
        RECT 340.190 79.890 341.090 80.790 ;
        RECT 317.320 78.630 318.630 79.490 ;
      LAYER nwell ;
        RECT 350.180 79.360 351.030 79.470 ;
      LAYER pwell ;
        RECT 365.820 79.410 367.130 80.270 ;
        RECT 340.200 77.890 341.100 78.830 ;
      LAYER nwell ;
        RECT 182.680 75.300 183.530 75.390 ;
        RECT 117.650 74.690 118.500 74.780 ;
      LAYER pwell ;
        RECT 239.150 74.670 240.050 76.200 ;
        RECT 248.990 75.620 250.300 76.480 ;
      LAYER nwell ;
        RECT 251.900 74.910 253.820 77.170 ;
      LAYER pwell ;
        RECT 314.020 76.230 315.330 77.090 ;
      LAYER nwell ;
        RECT 316.930 75.520 318.850 77.780 ;
      LAYER pwell ;
        RECT 340.190 77.630 341.100 77.890 ;
        RECT 340.190 76.730 341.090 77.630 ;
      LAYER nwell ;
        RECT 349.960 77.130 351.870 79.360 ;
        RECT 368.730 78.700 370.650 80.960 ;
        RECT 415.210 79.970 416.060 80.080 ;
      LAYER pwell ;
        RECT 353.600 77.830 354.910 78.690 ;
      LAYER nwell ;
        RECT 369.700 78.610 370.550 78.700 ;
        RECT 414.990 77.740 416.900 79.970 ;
      LAYER pwell ;
        RECT 418.630 78.440 419.940 79.300 ;
      LAYER nwell ;
        RECT 317.900 75.430 318.750 75.520 ;
        RECT 252.870 74.820 253.720 74.910 ;
      LAYER pwell ;
        RECT 239.150 74.660 239.570 74.670 ;
        RECT 103.930 74.530 104.350 74.540 ;
        RECT 340.460 74.480 341.360 76.010 ;
        RECT 350.300 75.430 351.610 76.290 ;
      LAYER nwell ;
        RECT 353.210 74.720 355.130 76.980 ;
      LAYER pwell ;
        RECT 415.330 76.040 416.640 76.900 ;
      LAYER nwell ;
        RECT 418.240 75.330 420.160 77.590 ;
        RECT 419.210 75.240 420.060 75.330 ;
        RECT 354.180 74.630 355.030 74.720 ;
      LAYER pwell ;
        RECT 340.460 74.470 340.880 74.480 ;
        RECT 2.180 71.600 3.710 72.080 ;
        RECT 2.180 71.180 3.720 71.600 ;
        RECT 103.490 71.410 105.020 71.890 ;
        RECT 238.710 71.540 240.240 72.020 ;
        RECT 103.490 70.990 105.030 71.410 ;
        RECT 238.710 71.120 240.250 71.540 ;
        RECT 340.020 71.350 341.550 71.830 ;
        RECT 340.020 70.930 341.560 71.350 ;
      LAYER nwell ;
        RECT 12.030 70.580 12.880 70.690 ;
      LAYER pwell ;
        RECT 2.250 68.110 3.150 69.050 ;
      LAYER nwell ;
        RECT 11.810 68.350 13.720 70.580 ;
        RECT 248.560 70.520 249.410 70.630 ;
        RECT 113.340 70.390 114.190 70.500 ;
      LAYER pwell ;
        RECT 15.450 69.050 16.760 69.910 ;
        RECT 2.240 67.850 3.150 68.110 ;
        RECT 2.240 66.950 3.140 67.850 ;
        RECT 2.210 65.870 3.110 66.810 ;
        RECT 12.150 66.650 13.460 67.510 ;
      LAYER nwell ;
        RECT 15.060 65.940 16.980 68.200 ;
        RECT 27.710 68.160 28.560 68.270 ;
      LAYER pwell ;
        RECT 2.200 65.610 3.110 65.870 ;
      LAYER nwell ;
        RECT 16.030 65.850 16.880 65.940 ;
        RECT 27.490 65.930 29.400 68.160 ;
      LAYER pwell ;
        RECT 103.560 67.920 104.460 68.860 ;
      LAYER nwell ;
        RECT 113.120 68.160 115.030 70.390 ;
      LAYER pwell ;
        RECT 116.760 68.860 118.070 69.720 ;
        RECT 103.550 67.660 104.460 67.920 ;
        RECT 31.130 66.630 32.440 67.490 ;
        RECT 103.550 66.760 104.450 67.660 ;
        RECT 2.200 64.710 3.100 65.610 ;
      LAYER nwell ;
        RECT 12.190 64.180 13.040 64.290 ;
      LAYER pwell ;
        RECT 27.830 64.230 29.140 65.090 ;
        RECT 2.210 62.710 3.110 63.650 ;
        RECT 2.200 62.450 3.110 62.710 ;
        RECT 2.200 61.550 3.100 62.450 ;
      LAYER nwell ;
        RECT 11.970 61.950 13.880 64.180 ;
        RECT 30.740 63.520 32.660 65.780 ;
      LAYER pwell ;
        RECT 103.520 65.680 104.420 66.620 ;
        RECT 113.460 66.460 114.770 67.320 ;
      LAYER nwell ;
        RECT 116.370 65.750 118.290 68.010 ;
        RECT 129.020 67.970 129.870 68.080 ;
      LAYER pwell ;
        RECT 238.780 68.050 239.680 68.990 ;
      LAYER nwell ;
        RECT 248.340 68.290 250.250 70.520 ;
        RECT 349.870 70.330 350.720 70.440 ;
      LAYER pwell ;
        RECT 251.980 68.990 253.290 69.850 ;
        RECT 103.510 65.420 104.420 65.680 ;
      LAYER nwell ;
        RECT 117.340 65.660 118.190 65.750 ;
        RECT 128.800 65.740 130.710 67.970 ;
      LAYER pwell ;
        RECT 238.770 67.790 239.680 68.050 ;
        RECT 132.440 66.440 133.750 67.300 ;
        RECT 238.770 66.890 239.670 67.790 ;
        RECT 238.740 65.810 239.640 66.750 ;
        RECT 248.680 66.590 249.990 67.450 ;
      LAYER nwell ;
        RECT 251.590 65.880 253.510 68.140 ;
        RECT 264.240 68.100 265.090 68.210 ;
      LAYER pwell ;
        RECT 103.510 64.520 104.410 65.420 ;
      LAYER nwell ;
        RECT 113.500 63.990 114.350 64.100 ;
      LAYER pwell ;
        RECT 129.140 64.040 130.450 64.900 ;
        RECT 15.610 62.650 16.920 63.510 ;
      LAYER nwell ;
        RECT 31.710 63.430 32.560 63.520 ;
        RECT 45.290 62.610 46.140 62.720 ;
      LAYER pwell ;
        RECT 2.470 59.300 3.370 60.830 ;
        RECT 12.310 60.250 13.620 61.110 ;
      LAYER nwell ;
        RECT 15.220 59.540 17.140 61.800 ;
        RECT 45.070 60.380 46.980 62.610 ;
      LAYER pwell ;
        RECT 103.520 62.520 104.420 63.460 ;
        RECT 103.510 62.260 104.420 62.520 ;
        RECT 48.710 61.080 50.020 61.940 ;
        RECT 103.510 61.360 104.410 62.260 ;
      LAYER nwell ;
        RECT 113.280 61.760 115.190 63.990 ;
        RECT 132.050 63.330 133.970 65.590 ;
      LAYER pwell ;
        RECT 238.730 65.550 239.640 65.810 ;
      LAYER nwell ;
        RECT 252.560 65.790 253.410 65.880 ;
        RECT 264.020 65.870 265.930 68.100 ;
      LAYER pwell ;
        RECT 340.090 67.860 340.990 68.800 ;
      LAYER nwell ;
        RECT 349.650 68.100 351.560 70.330 ;
      LAYER pwell ;
        RECT 353.290 68.800 354.600 69.660 ;
        RECT 340.080 67.600 340.990 67.860 ;
        RECT 267.660 66.570 268.970 67.430 ;
        RECT 340.080 66.700 340.980 67.600 ;
        RECT 238.730 64.650 239.630 65.550 ;
      LAYER nwell ;
        RECT 248.720 64.120 249.570 64.230 ;
      LAYER pwell ;
        RECT 264.360 64.170 265.670 65.030 ;
        RECT 116.920 62.460 118.230 63.320 ;
      LAYER nwell ;
        RECT 133.020 63.240 133.870 63.330 ;
      LAYER pwell ;
        RECT 238.740 62.650 239.640 63.590 ;
      LAYER nwell ;
        RECT 146.600 62.420 147.450 62.530 ;
        RECT 16.190 59.450 17.040 59.540 ;
      LAYER pwell ;
        RECT 2.470 59.290 2.890 59.300 ;
        RECT 45.410 58.680 46.720 59.540 ;
      LAYER nwell ;
        RECT 48.320 57.970 50.240 60.230 ;
      LAYER pwell ;
        RECT 103.780 59.110 104.680 60.640 ;
        RECT 113.620 60.060 114.930 60.920 ;
      LAYER nwell ;
        RECT 116.530 59.350 118.450 61.610 ;
        RECT 146.380 60.190 148.290 62.420 ;
      LAYER pwell ;
        RECT 238.730 62.390 239.640 62.650 ;
        RECT 150.020 60.890 151.330 61.750 ;
        RECT 238.730 61.490 239.630 62.390 ;
      LAYER nwell ;
        RECT 248.500 61.890 250.410 64.120 ;
        RECT 267.270 63.460 269.190 65.720 ;
      LAYER pwell ;
        RECT 340.050 65.620 340.950 66.560 ;
        RECT 349.990 66.400 351.300 67.260 ;
      LAYER nwell ;
        RECT 352.900 65.690 354.820 67.950 ;
        RECT 365.550 67.910 366.400 68.020 ;
      LAYER pwell ;
        RECT 340.040 65.360 340.950 65.620 ;
      LAYER nwell ;
        RECT 353.870 65.600 354.720 65.690 ;
        RECT 365.330 65.680 367.240 67.910 ;
      LAYER pwell ;
        RECT 368.970 66.380 370.280 67.240 ;
        RECT 340.040 64.460 340.940 65.360 ;
      LAYER nwell ;
        RECT 350.030 63.930 350.880 64.040 ;
      LAYER pwell ;
        RECT 365.670 63.980 366.980 64.840 ;
        RECT 252.140 62.590 253.450 63.450 ;
      LAYER nwell ;
        RECT 268.240 63.370 269.090 63.460 ;
        RECT 281.820 62.550 282.670 62.660 ;
        RECT 117.500 59.260 118.350 59.350 ;
      LAYER pwell ;
        RECT 103.780 59.100 104.200 59.110 ;
        RECT 146.720 58.490 148.030 59.350 ;
      LAYER nwell ;
        RECT 49.290 57.880 50.140 57.970 ;
      LAYER pwell ;
        RECT 2.200 56.260 3.100 57.790 ;
      LAYER nwell ;
        RECT 149.630 57.780 151.550 60.040 ;
      LAYER pwell ;
        RECT 239.000 59.240 239.900 60.770 ;
        RECT 248.840 60.190 250.150 61.050 ;
      LAYER nwell ;
        RECT 251.750 59.480 253.670 61.740 ;
        RECT 281.600 60.320 283.510 62.550 ;
      LAYER pwell ;
        RECT 340.050 62.460 340.950 63.400 ;
        RECT 340.040 62.200 340.950 62.460 ;
        RECT 285.240 61.020 286.550 61.880 ;
        RECT 340.040 61.300 340.940 62.200 ;
      LAYER nwell ;
        RECT 349.810 61.700 351.720 63.930 ;
        RECT 368.580 63.270 370.500 65.530 ;
      LAYER pwell ;
        RECT 353.450 62.400 354.760 63.260 ;
      LAYER nwell ;
        RECT 369.550 63.180 370.400 63.270 ;
        RECT 383.130 62.360 383.980 62.470 ;
        RECT 252.720 59.390 253.570 59.480 ;
      LAYER pwell ;
        RECT 239.000 59.230 239.420 59.240 ;
        RECT 281.940 58.620 283.250 59.480 ;
      LAYER nwell ;
        RECT 284.850 57.910 286.770 60.170 ;
      LAYER pwell ;
        RECT 340.310 59.050 341.210 60.580 ;
        RECT 350.150 60.000 351.460 60.860 ;
      LAYER nwell ;
        RECT 353.060 59.290 354.980 61.550 ;
        RECT 382.910 60.130 384.820 62.360 ;
      LAYER pwell ;
        RECT 386.550 60.830 387.860 61.690 ;
      LAYER nwell ;
        RECT 354.030 59.200 354.880 59.290 ;
      LAYER pwell ;
        RECT 340.310 59.040 340.730 59.050 ;
        RECT 383.250 58.430 384.560 59.290 ;
      LAYER nwell ;
        RECT 285.820 57.820 286.670 57.910 ;
        RECT 150.600 57.690 151.450 57.780 ;
      LAYER pwell ;
        RECT 2.200 56.250 2.620 56.260 ;
      LAYER nwell ;
        RECT 11.860 56.160 12.710 56.270 ;
      LAYER pwell ;
        RECT 2.080 53.690 2.980 54.630 ;
      LAYER nwell ;
        RECT 11.640 53.930 13.550 56.160 ;
      LAYER pwell ;
        RECT 103.510 56.070 104.410 57.600 ;
        RECT 238.730 56.200 239.630 57.730 ;
      LAYER nwell ;
        RECT 386.160 57.720 388.080 59.980 ;
        RECT 387.130 57.630 387.980 57.720 ;
      LAYER pwell ;
        RECT 238.730 56.190 239.150 56.200 ;
      LAYER nwell ;
        RECT 248.390 56.100 249.240 56.210 ;
      LAYER pwell ;
        RECT 103.510 56.060 103.930 56.070 ;
      LAYER nwell ;
        RECT 113.170 55.970 114.020 56.080 ;
      LAYER pwell ;
        RECT 15.280 54.630 16.590 55.490 ;
        RECT 2.070 53.430 2.980 53.690 ;
        RECT 2.070 52.530 2.970 53.430 ;
        RECT 2.040 51.450 2.940 52.390 ;
        RECT 11.980 52.230 13.290 53.090 ;
      LAYER nwell ;
        RECT 14.890 51.520 16.810 53.780 ;
        RECT 27.540 53.740 28.390 53.850 ;
      LAYER pwell ;
        RECT 2.030 51.190 2.940 51.450 ;
      LAYER nwell ;
        RECT 15.860 51.430 16.710 51.520 ;
        RECT 27.320 51.510 29.230 53.740 ;
      LAYER pwell ;
        RECT 103.390 53.500 104.290 54.440 ;
      LAYER nwell ;
        RECT 112.950 53.740 114.860 55.970 ;
      LAYER pwell ;
        RECT 116.590 54.440 117.900 55.300 ;
        RECT 103.380 53.240 104.290 53.500 ;
        RECT 30.960 52.210 32.270 53.070 ;
        RECT 103.380 52.340 104.280 53.240 ;
        RECT 2.030 50.290 2.930 51.190 ;
      LAYER nwell ;
        RECT 12.020 49.760 12.870 49.870 ;
      LAYER pwell ;
        RECT 27.660 49.810 28.970 50.670 ;
        RECT 2.040 48.290 2.940 49.230 ;
        RECT 2.030 48.030 2.940 48.290 ;
        RECT 2.030 47.130 2.930 48.030 ;
      LAYER nwell ;
        RECT 11.800 47.530 13.710 49.760 ;
        RECT 30.570 49.100 32.490 51.360 ;
      LAYER pwell ;
        RECT 103.350 51.260 104.250 52.200 ;
        RECT 113.290 52.040 114.600 52.900 ;
      LAYER nwell ;
        RECT 116.200 51.330 118.120 53.590 ;
        RECT 128.850 53.550 129.700 53.660 ;
      LAYER pwell ;
        RECT 238.610 53.630 239.510 54.570 ;
      LAYER nwell ;
        RECT 248.170 53.870 250.080 56.100 ;
      LAYER pwell ;
        RECT 340.040 56.010 340.940 57.540 ;
        RECT 340.040 56.000 340.460 56.010 ;
      LAYER nwell ;
        RECT 349.700 55.910 350.550 56.020 ;
      LAYER pwell ;
        RECT 251.810 54.570 253.120 55.430 ;
        RECT 103.340 51.000 104.250 51.260 ;
      LAYER nwell ;
        RECT 117.170 51.240 118.020 51.330 ;
        RECT 128.630 51.320 130.540 53.550 ;
      LAYER pwell ;
        RECT 238.600 53.370 239.510 53.630 ;
        RECT 132.270 52.020 133.580 52.880 ;
        RECT 238.600 52.470 239.500 53.370 ;
        RECT 238.570 51.390 239.470 52.330 ;
        RECT 248.510 52.170 249.820 53.030 ;
      LAYER nwell ;
        RECT 251.420 51.460 253.340 53.720 ;
        RECT 264.070 53.680 264.920 53.790 ;
      LAYER pwell ;
        RECT 103.340 50.100 104.240 51.000 ;
      LAYER nwell ;
        RECT 113.330 49.570 114.180 49.680 ;
      LAYER pwell ;
        RECT 128.970 49.620 130.280 50.480 ;
        RECT 15.440 48.230 16.750 49.090 ;
      LAYER nwell ;
        RECT 31.540 49.010 32.390 49.100 ;
      LAYER pwell ;
        RECT 103.350 48.100 104.250 49.040 ;
        RECT 103.340 47.840 104.250 48.100 ;
        RECT 2.300 44.880 3.200 46.410 ;
        RECT 12.140 45.830 13.450 46.690 ;
      LAYER nwell ;
        RECT 15.050 45.120 16.970 47.380 ;
      LAYER pwell ;
        RECT 103.340 46.940 104.240 47.840 ;
      LAYER nwell ;
        RECT 113.110 47.340 115.020 49.570 ;
        RECT 131.880 48.910 133.800 51.170 ;
      LAYER pwell ;
        RECT 238.560 51.130 239.470 51.390 ;
      LAYER nwell ;
        RECT 252.390 51.370 253.240 51.460 ;
        RECT 263.850 51.450 265.760 53.680 ;
      LAYER pwell ;
        RECT 339.920 53.440 340.820 54.380 ;
      LAYER nwell ;
        RECT 349.480 53.680 351.390 55.910 ;
      LAYER pwell ;
        RECT 353.120 54.380 354.430 55.240 ;
        RECT 339.910 53.180 340.820 53.440 ;
        RECT 267.490 52.150 268.800 53.010 ;
        RECT 339.910 52.280 340.810 53.180 ;
        RECT 238.560 50.230 239.460 51.130 ;
      LAYER nwell ;
        RECT 248.550 49.700 249.400 49.810 ;
      LAYER pwell ;
        RECT 264.190 49.750 265.500 50.610 ;
        RECT 116.750 48.040 118.060 48.900 ;
      LAYER nwell ;
        RECT 132.850 48.820 133.700 48.910 ;
      LAYER pwell ;
        RECT 238.570 48.230 239.470 49.170 ;
        RECT 238.560 47.970 239.470 48.230 ;
      LAYER nwell ;
        RECT 62.820 46.590 63.670 46.700 ;
        RECT 16.020 45.030 16.870 45.120 ;
      LAYER pwell ;
        RECT 2.300 44.870 2.720 44.880 ;
      LAYER nwell ;
        RECT 62.600 44.360 64.510 46.590 ;
      LAYER pwell ;
        RECT 66.240 45.060 67.550 45.920 ;
        RECT 103.610 44.690 104.510 46.220 ;
        RECT 113.450 45.640 114.760 46.500 ;
      LAYER nwell ;
        RECT 116.360 44.930 118.280 47.190 ;
      LAYER pwell ;
        RECT 238.560 47.070 239.460 47.970 ;
      LAYER nwell ;
        RECT 248.330 47.470 250.240 49.700 ;
        RECT 267.100 49.040 269.020 51.300 ;
      LAYER pwell ;
        RECT 339.880 51.200 340.780 52.140 ;
        RECT 349.820 51.980 351.130 52.840 ;
      LAYER nwell ;
        RECT 352.730 51.270 354.650 53.530 ;
        RECT 365.380 53.490 366.230 53.600 ;
      LAYER pwell ;
        RECT 339.870 50.940 340.780 51.200 ;
      LAYER nwell ;
        RECT 353.700 51.180 354.550 51.270 ;
        RECT 365.160 51.260 367.070 53.490 ;
      LAYER pwell ;
        RECT 368.800 51.960 370.110 52.820 ;
        RECT 339.870 50.040 340.770 50.940 ;
      LAYER nwell ;
        RECT 349.860 49.510 350.710 49.620 ;
      LAYER pwell ;
        RECT 365.500 49.560 366.810 50.420 ;
        RECT 251.970 48.170 253.280 49.030 ;
      LAYER nwell ;
        RECT 268.070 48.950 268.920 49.040 ;
      LAYER pwell ;
        RECT 339.880 48.040 340.780 48.980 ;
        RECT 339.870 47.780 340.780 48.040 ;
      LAYER nwell ;
        RECT 164.130 46.400 164.980 46.510 ;
        RECT 117.330 44.840 118.180 44.930 ;
      LAYER pwell ;
        RECT 103.610 44.680 104.030 44.690 ;
        RECT 62.940 42.660 64.250 43.520 ;
        RECT 2.890 42.560 3.310 42.570 ;
        RECT 2.410 41.030 3.310 42.560 ;
      LAYER nwell ;
        RECT 65.850 41.950 67.770 44.210 ;
        RECT 163.910 44.170 165.820 46.400 ;
      LAYER pwell ;
        RECT 167.550 44.870 168.860 45.730 ;
        RECT 238.830 44.820 239.730 46.350 ;
        RECT 248.670 45.770 249.980 46.630 ;
      LAYER nwell ;
        RECT 251.580 45.060 253.500 47.320 ;
      LAYER pwell ;
        RECT 339.870 46.880 340.770 47.780 ;
      LAYER nwell ;
        RECT 349.640 47.280 351.550 49.510 ;
        RECT 368.410 48.850 370.330 51.110 ;
      LAYER pwell ;
        RECT 353.280 47.980 354.590 48.840 ;
      LAYER nwell ;
        RECT 369.380 48.760 370.230 48.850 ;
        RECT 299.350 46.530 300.200 46.640 ;
        RECT 252.550 44.970 253.400 45.060 ;
      LAYER pwell ;
        RECT 238.830 44.810 239.250 44.820 ;
      LAYER nwell ;
        RECT 299.130 44.300 301.040 46.530 ;
      LAYER pwell ;
        RECT 302.770 45.000 304.080 45.860 ;
        RECT 340.140 44.630 341.040 46.160 ;
        RECT 349.980 45.580 351.290 46.440 ;
      LAYER nwell ;
        RECT 352.890 44.870 354.810 47.130 ;
        RECT 400.660 46.340 401.510 46.450 ;
        RECT 353.860 44.780 354.710 44.870 ;
      LAYER pwell ;
        RECT 340.140 44.620 340.560 44.630 ;
        RECT 164.250 42.470 165.560 43.330 ;
        RECT 104.200 42.370 104.620 42.380 ;
      LAYER nwell ;
        RECT 66.820 41.860 67.670 41.950 ;
      LAYER pwell ;
        RECT 103.720 40.840 104.620 42.370 ;
      LAYER nwell ;
        RECT 167.160 41.760 169.080 44.020 ;
      LAYER pwell ;
        RECT 299.470 42.600 300.780 43.460 ;
        RECT 239.420 42.500 239.840 42.510 ;
      LAYER nwell ;
        RECT 168.130 41.670 168.980 41.760 ;
      LAYER pwell ;
        RECT 238.940 40.970 239.840 42.500 ;
      LAYER nwell ;
        RECT 302.380 41.890 304.300 44.150 ;
        RECT 400.440 44.110 402.350 46.340 ;
      LAYER pwell ;
        RECT 404.080 44.810 405.390 45.670 ;
        RECT 400.780 42.410 402.090 43.270 ;
        RECT 340.730 42.310 341.150 42.320 ;
      LAYER nwell ;
        RECT 303.350 41.800 304.200 41.890 ;
      LAYER pwell ;
        RECT 340.250 40.780 341.150 42.310 ;
      LAYER nwell ;
        RECT 403.690 41.700 405.610 43.960 ;
        RECT 404.660 41.610 405.510 41.700 ;
        RECT 12.000 40.510 12.850 40.620 ;
      LAYER pwell ;
        RECT 2.220 38.040 3.120 38.980 ;
      LAYER nwell ;
        RECT 11.780 38.280 13.690 40.510 ;
        RECT 248.530 40.450 249.380 40.560 ;
        RECT 113.310 40.320 114.160 40.430 ;
      LAYER pwell ;
        RECT 15.420 38.980 16.730 39.840 ;
        RECT 2.210 37.780 3.120 38.040 ;
        RECT 2.210 36.880 3.110 37.780 ;
        RECT 2.180 35.800 3.080 36.740 ;
        RECT 12.120 36.580 13.430 37.440 ;
      LAYER nwell ;
        RECT 15.030 35.870 16.950 38.130 ;
        RECT 27.680 38.090 28.530 38.200 ;
      LAYER pwell ;
        RECT 2.170 35.540 3.080 35.800 ;
      LAYER nwell ;
        RECT 16.000 35.780 16.850 35.870 ;
        RECT 27.460 35.860 29.370 38.090 ;
      LAYER pwell ;
        RECT 103.530 37.850 104.430 38.790 ;
      LAYER nwell ;
        RECT 113.090 38.090 115.000 40.320 ;
      LAYER pwell ;
        RECT 116.730 38.790 118.040 39.650 ;
        RECT 103.520 37.590 104.430 37.850 ;
        RECT 31.100 36.560 32.410 37.420 ;
        RECT 103.520 36.690 104.420 37.590 ;
        RECT 2.170 34.640 3.070 35.540 ;
      LAYER nwell ;
        RECT 12.160 34.110 13.010 34.220 ;
      LAYER pwell ;
        RECT 27.800 34.160 29.110 35.020 ;
        RECT 2.180 32.640 3.080 33.580 ;
        RECT 2.170 32.380 3.080 32.640 ;
        RECT 2.170 31.480 3.070 32.380 ;
      LAYER nwell ;
        RECT 11.940 31.880 13.850 34.110 ;
        RECT 30.710 33.450 32.630 35.710 ;
      LAYER pwell ;
        RECT 103.490 35.610 104.390 36.550 ;
        RECT 113.430 36.390 114.740 37.250 ;
      LAYER nwell ;
        RECT 116.340 35.680 118.260 37.940 ;
        RECT 128.990 37.900 129.840 38.010 ;
      LAYER pwell ;
        RECT 238.750 37.980 239.650 38.920 ;
      LAYER nwell ;
        RECT 248.310 38.220 250.220 40.450 ;
        RECT 349.840 40.260 350.690 40.370 ;
      LAYER pwell ;
        RECT 251.950 38.920 253.260 39.780 ;
        RECT 103.480 35.350 104.390 35.610 ;
      LAYER nwell ;
        RECT 117.310 35.590 118.160 35.680 ;
        RECT 128.770 35.670 130.680 37.900 ;
      LAYER pwell ;
        RECT 238.740 37.720 239.650 37.980 ;
        RECT 132.410 36.370 133.720 37.230 ;
        RECT 238.740 36.820 239.640 37.720 ;
        RECT 238.710 35.740 239.610 36.680 ;
        RECT 248.650 36.520 249.960 37.380 ;
      LAYER nwell ;
        RECT 251.560 35.810 253.480 38.070 ;
        RECT 264.210 38.030 265.060 38.140 ;
      LAYER pwell ;
        RECT 103.480 34.450 104.380 35.350 ;
      LAYER nwell ;
        RECT 113.470 33.920 114.320 34.030 ;
      LAYER pwell ;
        RECT 129.110 33.970 130.420 34.830 ;
        RECT 15.580 32.580 16.890 33.440 ;
      LAYER nwell ;
        RECT 31.680 33.360 32.530 33.450 ;
        RECT 45.260 32.540 46.110 32.650 ;
      LAYER pwell ;
        RECT 2.440 29.230 3.340 30.760 ;
        RECT 12.280 30.180 13.590 31.040 ;
      LAYER nwell ;
        RECT 15.190 29.470 17.110 31.730 ;
        RECT 45.040 30.310 46.950 32.540 ;
      LAYER pwell ;
        RECT 103.490 32.450 104.390 33.390 ;
        RECT 103.480 32.190 104.390 32.450 ;
        RECT 48.680 31.010 49.990 31.870 ;
        RECT 103.480 31.290 104.380 32.190 ;
      LAYER nwell ;
        RECT 113.250 31.690 115.160 33.920 ;
        RECT 132.020 33.260 133.940 35.520 ;
      LAYER pwell ;
        RECT 238.700 35.480 239.610 35.740 ;
      LAYER nwell ;
        RECT 252.530 35.720 253.380 35.810 ;
        RECT 263.990 35.800 265.900 38.030 ;
      LAYER pwell ;
        RECT 340.060 37.790 340.960 38.730 ;
      LAYER nwell ;
        RECT 349.620 38.030 351.530 40.260 ;
      LAYER pwell ;
        RECT 353.260 38.730 354.570 39.590 ;
        RECT 340.050 37.530 340.960 37.790 ;
        RECT 267.630 36.500 268.940 37.360 ;
        RECT 340.050 36.630 340.950 37.530 ;
        RECT 238.700 34.580 239.600 35.480 ;
      LAYER nwell ;
        RECT 248.690 34.050 249.540 34.160 ;
      LAYER pwell ;
        RECT 264.330 34.100 265.640 34.960 ;
        RECT 116.890 32.390 118.200 33.250 ;
      LAYER nwell ;
        RECT 132.990 33.170 133.840 33.260 ;
      LAYER pwell ;
        RECT 238.710 32.580 239.610 33.520 ;
      LAYER nwell ;
        RECT 146.570 32.350 147.420 32.460 ;
        RECT 16.160 29.380 17.010 29.470 ;
      LAYER pwell ;
        RECT 2.440 29.220 2.860 29.230 ;
        RECT 45.380 28.610 46.690 29.470 ;
      LAYER nwell ;
        RECT 48.290 27.900 50.210 30.160 ;
      LAYER pwell ;
        RECT 103.750 29.040 104.650 30.570 ;
        RECT 113.590 29.990 114.900 30.850 ;
      LAYER nwell ;
        RECT 116.500 29.280 118.420 31.540 ;
        RECT 146.350 30.120 148.260 32.350 ;
      LAYER pwell ;
        RECT 238.700 32.320 239.610 32.580 ;
        RECT 149.990 30.820 151.300 31.680 ;
        RECT 238.700 31.420 239.600 32.320 ;
      LAYER nwell ;
        RECT 248.470 31.820 250.380 34.050 ;
        RECT 267.240 33.390 269.160 35.650 ;
      LAYER pwell ;
        RECT 340.020 35.550 340.920 36.490 ;
        RECT 349.960 36.330 351.270 37.190 ;
      LAYER nwell ;
        RECT 352.870 35.620 354.790 37.880 ;
        RECT 365.520 37.840 366.370 37.950 ;
      LAYER pwell ;
        RECT 340.010 35.290 340.920 35.550 ;
      LAYER nwell ;
        RECT 353.840 35.530 354.690 35.620 ;
        RECT 365.300 35.610 367.210 37.840 ;
      LAYER pwell ;
        RECT 368.940 36.310 370.250 37.170 ;
        RECT 340.010 34.390 340.910 35.290 ;
      LAYER nwell ;
        RECT 350.000 33.860 350.850 33.970 ;
      LAYER pwell ;
        RECT 365.640 33.910 366.950 34.770 ;
        RECT 252.110 32.520 253.420 33.380 ;
      LAYER nwell ;
        RECT 268.210 33.300 269.060 33.390 ;
        RECT 281.790 32.480 282.640 32.590 ;
        RECT 117.470 29.190 118.320 29.280 ;
      LAYER pwell ;
        RECT 103.750 29.030 104.170 29.040 ;
        RECT 146.690 28.420 148.000 29.280 ;
      LAYER nwell ;
        RECT 49.260 27.810 50.110 27.900 ;
      LAYER pwell ;
        RECT 2.170 26.190 3.070 27.720 ;
      LAYER nwell ;
        RECT 149.600 27.710 151.520 29.970 ;
      LAYER pwell ;
        RECT 238.970 29.170 239.870 30.700 ;
        RECT 248.810 30.120 250.120 30.980 ;
      LAYER nwell ;
        RECT 251.720 29.410 253.640 31.670 ;
        RECT 281.570 30.250 283.480 32.480 ;
      LAYER pwell ;
        RECT 340.020 32.390 340.920 33.330 ;
        RECT 340.010 32.130 340.920 32.390 ;
        RECT 285.210 30.950 286.520 31.810 ;
        RECT 340.010 31.230 340.910 32.130 ;
      LAYER nwell ;
        RECT 349.780 31.630 351.690 33.860 ;
        RECT 368.550 33.200 370.470 35.460 ;
      LAYER pwell ;
        RECT 353.420 32.330 354.730 33.190 ;
      LAYER nwell ;
        RECT 369.520 33.110 370.370 33.200 ;
        RECT 383.100 32.290 383.950 32.400 ;
        RECT 252.690 29.320 253.540 29.410 ;
      LAYER pwell ;
        RECT 238.970 29.160 239.390 29.170 ;
        RECT 281.910 28.550 283.220 29.410 ;
      LAYER nwell ;
        RECT 284.820 27.840 286.740 30.100 ;
      LAYER pwell ;
        RECT 340.280 28.980 341.180 30.510 ;
        RECT 350.120 29.930 351.430 30.790 ;
      LAYER nwell ;
        RECT 353.030 29.220 354.950 31.480 ;
        RECT 382.880 30.060 384.790 32.290 ;
      LAYER pwell ;
        RECT 386.520 30.760 387.830 31.620 ;
      LAYER nwell ;
        RECT 354.000 29.130 354.850 29.220 ;
      LAYER pwell ;
        RECT 340.280 28.970 340.700 28.980 ;
        RECT 383.220 28.360 384.530 29.220 ;
      LAYER nwell ;
        RECT 285.790 27.750 286.640 27.840 ;
        RECT 150.570 27.620 151.420 27.710 ;
      LAYER pwell ;
        RECT 2.170 26.180 2.590 26.190 ;
      LAYER nwell ;
        RECT 11.830 26.090 12.680 26.200 ;
      LAYER pwell ;
        RECT 2.050 23.620 2.950 24.560 ;
      LAYER nwell ;
        RECT 11.610 23.860 13.520 26.090 ;
      LAYER pwell ;
        RECT 103.480 26.000 104.380 27.530 ;
        RECT 238.700 26.130 239.600 27.660 ;
      LAYER nwell ;
        RECT 386.130 27.650 388.050 29.910 ;
        RECT 387.100 27.560 387.950 27.650 ;
      LAYER pwell ;
        RECT 238.700 26.120 239.120 26.130 ;
      LAYER nwell ;
        RECT 248.360 26.030 249.210 26.140 ;
      LAYER pwell ;
        RECT 103.480 25.990 103.900 26.000 ;
      LAYER nwell ;
        RECT 113.140 25.900 113.990 26.010 ;
      LAYER pwell ;
        RECT 15.250 24.560 16.560 25.420 ;
        RECT 2.040 23.360 2.950 23.620 ;
        RECT 2.040 22.460 2.940 23.360 ;
        RECT 2.010 21.380 2.910 22.320 ;
        RECT 11.950 22.160 13.260 23.020 ;
      LAYER nwell ;
        RECT 14.860 21.450 16.780 23.710 ;
        RECT 27.510 23.670 28.360 23.780 ;
      LAYER pwell ;
        RECT 2.000 21.120 2.910 21.380 ;
      LAYER nwell ;
        RECT 15.830 21.360 16.680 21.450 ;
        RECT 27.290 21.440 29.200 23.670 ;
      LAYER pwell ;
        RECT 103.360 23.430 104.260 24.370 ;
      LAYER nwell ;
        RECT 112.920 23.670 114.830 25.900 ;
      LAYER pwell ;
        RECT 116.560 24.370 117.870 25.230 ;
        RECT 103.350 23.170 104.260 23.430 ;
        RECT 30.930 22.140 32.240 23.000 ;
        RECT 103.350 22.270 104.250 23.170 ;
        RECT 2.000 20.220 2.900 21.120 ;
      LAYER nwell ;
        RECT 11.990 19.690 12.840 19.800 ;
      LAYER pwell ;
        RECT 27.630 19.740 28.940 20.600 ;
        RECT 2.010 18.220 2.910 19.160 ;
        RECT 2.000 17.960 2.910 18.220 ;
        RECT 2.000 17.060 2.900 17.960 ;
      LAYER nwell ;
        RECT 11.770 17.460 13.680 19.690 ;
        RECT 30.540 19.030 32.460 21.290 ;
      LAYER pwell ;
        RECT 103.320 21.190 104.220 22.130 ;
        RECT 113.260 21.970 114.570 22.830 ;
      LAYER nwell ;
        RECT 116.170 21.260 118.090 23.520 ;
        RECT 128.820 23.480 129.670 23.590 ;
      LAYER pwell ;
        RECT 238.580 23.560 239.480 24.500 ;
      LAYER nwell ;
        RECT 248.140 23.800 250.050 26.030 ;
      LAYER pwell ;
        RECT 340.010 25.940 340.910 27.470 ;
        RECT 340.010 25.930 340.430 25.940 ;
      LAYER nwell ;
        RECT 349.670 25.840 350.520 25.950 ;
      LAYER pwell ;
        RECT 251.780 24.500 253.090 25.360 ;
        RECT 103.310 20.930 104.220 21.190 ;
      LAYER nwell ;
        RECT 117.140 21.170 117.990 21.260 ;
        RECT 128.600 21.250 130.510 23.480 ;
      LAYER pwell ;
        RECT 238.570 23.300 239.480 23.560 ;
        RECT 132.240 21.950 133.550 22.810 ;
        RECT 238.570 22.400 239.470 23.300 ;
        RECT 238.540 21.320 239.440 22.260 ;
        RECT 248.480 22.100 249.790 22.960 ;
      LAYER nwell ;
        RECT 251.390 21.390 253.310 23.650 ;
        RECT 264.040 23.610 264.890 23.720 ;
      LAYER pwell ;
        RECT 103.310 20.030 104.210 20.930 ;
      LAYER nwell ;
        RECT 113.300 19.500 114.150 19.610 ;
      LAYER pwell ;
        RECT 128.940 19.550 130.250 20.410 ;
        RECT 15.410 18.160 16.720 19.020 ;
      LAYER nwell ;
        RECT 31.510 18.940 32.360 19.030 ;
      LAYER pwell ;
        RECT 103.320 18.030 104.220 18.970 ;
        RECT 103.310 17.770 104.220 18.030 ;
        RECT 2.270 14.810 3.170 16.340 ;
        RECT 12.110 15.760 13.420 16.620 ;
      LAYER nwell ;
        RECT 15.020 15.050 16.940 17.310 ;
      LAYER pwell ;
        RECT 103.310 16.870 104.210 17.770 ;
      LAYER nwell ;
        RECT 113.080 17.270 114.990 19.500 ;
        RECT 131.850 18.840 133.770 21.100 ;
      LAYER pwell ;
        RECT 238.530 21.060 239.440 21.320 ;
      LAYER nwell ;
        RECT 252.360 21.300 253.210 21.390 ;
        RECT 263.820 21.380 265.730 23.610 ;
      LAYER pwell ;
        RECT 339.890 23.370 340.790 24.310 ;
      LAYER nwell ;
        RECT 349.450 23.610 351.360 25.840 ;
      LAYER pwell ;
        RECT 353.090 24.310 354.400 25.170 ;
        RECT 339.880 23.110 340.790 23.370 ;
        RECT 267.460 22.080 268.770 22.940 ;
        RECT 339.880 22.210 340.780 23.110 ;
        RECT 238.530 20.160 239.430 21.060 ;
      LAYER nwell ;
        RECT 248.520 19.630 249.370 19.740 ;
      LAYER pwell ;
        RECT 264.160 19.680 265.470 20.540 ;
        RECT 116.720 17.970 118.030 18.830 ;
      LAYER nwell ;
        RECT 132.820 18.750 133.670 18.840 ;
      LAYER pwell ;
        RECT 238.540 18.160 239.440 19.100 ;
        RECT 238.530 17.900 239.440 18.160 ;
        RECT 238.530 17.000 239.430 17.900 ;
      LAYER nwell ;
        RECT 248.300 17.400 250.210 19.630 ;
        RECT 267.070 18.970 268.990 21.230 ;
      LAYER pwell ;
        RECT 339.850 21.130 340.750 22.070 ;
        RECT 349.790 21.910 351.100 22.770 ;
      LAYER nwell ;
        RECT 352.700 21.200 354.620 23.460 ;
        RECT 365.350 23.420 366.200 23.530 ;
      LAYER pwell ;
        RECT 339.840 20.870 340.750 21.130 ;
      LAYER nwell ;
        RECT 353.670 21.110 354.520 21.200 ;
        RECT 365.130 21.190 367.040 23.420 ;
      LAYER pwell ;
        RECT 368.770 21.890 370.080 22.750 ;
        RECT 339.840 19.970 340.740 20.870 ;
      LAYER nwell ;
        RECT 349.830 19.440 350.680 19.550 ;
      LAYER pwell ;
        RECT 365.470 19.490 366.780 20.350 ;
        RECT 251.940 18.100 253.250 18.960 ;
      LAYER nwell ;
        RECT 268.040 18.880 268.890 18.970 ;
      LAYER pwell ;
        RECT 339.850 17.970 340.750 18.910 ;
        RECT 339.840 17.710 340.750 17.970 ;
      LAYER nwell ;
        RECT 15.990 14.960 16.840 15.050 ;
      LAYER pwell ;
        RECT 2.270 14.800 2.690 14.810 ;
        RECT 103.580 14.620 104.480 16.150 ;
        RECT 113.420 15.570 114.730 16.430 ;
        RECT 238.800 14.750 239.700 16.280 ;
        RECT 248.640 15.700 249.950 16.560 ;
      LAYER nwell ;
        RECT 251.550 14.990 253.470 17.250 ;
      LAYER pwell ;
        RECT 339.840 16.810 340.740 17.710 ;
      LAYER nwell ;
        RECT 349.610 17.210 351.520 19.440 ;
        RECT 368.380 18.780 370.300 21.040 ;
      LAYER pwell ;
        RECT 353.250 17.910 354.560 18.770 ;
      LAYER nwell ;
        RECT 369.350 18.690 370.200 18.780 ;
        RECT 252.520 14.900 253.370 14.990 ;
      LAYER pwell ;
        RECT 238.800 14.740 239.220 14.750 ;
        RECT 103.580 14.610 104.000 14.620 ;
        RECT 340.110 14.560 341.010 16.090 ;
        RECT 349.950 15.510 351.260 16.370 ;
        RECT 340.110 14.550 340.530 14.560 ;
        RECT 1.390 11.050 2.920 11.530 ;
        RECT 1.390 10.630 2.930 11.050 ;
        RECT 237.920 10.990 239.450 11.470 ;
        RECT 102.970 10.380 104.500 10.860 ;
        RECT 237.920 10.570 239.460 10.990 ;
        RECT 102.970 9.960 104.510 10.380 ;
      LAYER li1 ;
        RECT 100.840 255.690 101.070 255.710 ;
        RECT 100.840 255.680 101.080 255.690 ;
        RECT 100.840 255.630 101.090 255.680 ;
        RECT 220.060 255.630 227.070 255.670 ;
        RECT 100.840 255.480 227.070 255.630 ;
        RECT 100.840 255.440 220.450 255.480 ;
        RECT 100.840 255.430 137.530 255.440 ;
        RECT 226.840 255.400 227.070 255.480 ;
        RECT 337.370 255.630 337.600 255.650 ;
        RECT 337.370 255.620 337.610 255.630 ;
        RECT 337.370 255.570 337.620 255.620 ;
        RECT 456.590 255.570 463.600 255.610 ;
        RECT 337.370 255.420 463.600 255.570 ;
        RECT 60.100 252.760 102.070 252.780 ;
        RECT 0.000 252.530 105.560 252.760 ;
        RECT 0.000 252.510 60.350 252.530 ;
        RECT 0.000 252.480 18.500 252.510 ;
        RECT 0.030 11.460 0.290 252.480 ;
        RECT 100.840 251.980 101.140 252.230 ;
        RECT 5.170 251.530 14.440 251.540 ;
        RECT 16.320 251.530 18.240 251.540 ;
        RECT 5.170 251.340 18.240 251.530 ;
        RECT 5.170 251.330 17.530 251.340 ;
        RECT 5.170 250.320 5.380 251.330 ;
        RECT 14.430 251.320 16.330 251.330 ;
        RECT 18.060 250.590 18.240 251.340 ;
        RECT 5.170 249.310 5.370 250.320 ;
        RECT 12.980 250.290 18.240 250.590 ;
        RECT 3.210 247.230 4.170 247.680 ;
        RECT 3.920 247.180 4.170 247.230 ;
        RECT 5.180 247.180 5.370 249.310 ;
        RECT 3.920 246.980 5.370 247.180 ;
        RECT 8.900 248.650 9.160 249.850 ;
        RECT 8.900 248.140 9.150 248.650 ;
        RECT 10.790 248.640 11.050 249.850 ;
        RECT 13.180 248.740 13.430 250.290 ;
        RECT 10.790 248.480 11.180 248.640 ;
        RECT 10.780 248.350 11.180 248.480 ;
        RECT 13.880 248.350 14.140 249.960 ;
        RECT 16.430 248.890 16.730 249.940 ;
        RECT 17.180 249.340 17.480 250.290 ;
        RECT 17.680 249.390 17.980 249.440 ;
        RECT 17.680 249.040 18.580 249.390 ;
        RECT 20.290 249.260 20.510 249.270 ;
        RECT 20.290 249.070 33.970 249.260 ;
        RECT 20.290 248.940 20.510 249.070 ;
        RECT 9.400 248.140 9.690 248.300 ;
        RECT 10.780 248.290 11.040 248.350 ;
        RECT 8.900 247.950 9.690 248.140 ;
        RECT 8.900 247.750 9.150 247.950 ;
        RECT 9.400 247.840 9.690 247.950 ;
        RECT 10.790 247.750 11.040 248.290 ;
        RECT 13.870 248.290 14.140 248.350 ;
        RECT 15.420 248.630 16.730 248.890 ;
        RECT 18.830 248.640 20.510 248.940 ;
        RECT 18.830 248.630 20.490 248.640 ;
        RECT 15.420 248.290 15.730 248.630 ;
        RECT 11.430 247.760 13.070 248.150 ;
        RECT 13.870 248.000 15.730 248.290 ;
        RECT 13.870 247.990 14.180 248.000 ;
        RECT 15.420 247.990 15.730 248.000 ;
        RECT 8.900 247.150 9.190 247.750 ;
        RECT 10.790 247.150 11.080 247.750 ;
        RECT 3.920 246.890 4.170 246.980 ;
        RECT 3.190 246.440 4.170 246.890 ;
        RECT 13.130 246.540 13.430 247.540 ;
        RECT 13.880 246.940 14.180 247.990 ;
        RECT 16.480 246.890 16.730 248.630 ;
        RECT 33.720 248.170 33.970 249.070 ;
        RECT 17.180 246.540 17.440 248.090 ;
        RECT 28.660 247.870 33.970 248.170 ;
        RECT 13.080 246.520 18.330 246.540 ;
        RECT 13.080 246.240 18.450 246.520 ;
        RECT 6.530 245.840 6.810 245.910 ;
        RECT 7.710 245.870 7.990 245.900 ;
        RECT 18.160 245.870 18.450 246.240 ;
        RECT 7.710 245.860 18.450 245.870 ;
        RECT 5.120 245.640 6.810 245.840 ;
        RECT 3.910 245.440 4.190 245.450 ;
        RECT 3.170 244.990 4.190 245.440 ;
        RECT 5.120 244.990 5.350 245.640 ;
        RECT 6.530 245.580 6.810 245.640 ;
        RECT 7.690 245.630 18.450 245.860 ;
        RECT 7.710 245.620 18.450 245.630 ;
        RECT 24.580 246.230 24.840 247.430 ;
        RECT 24.580 245.720 24.830 246.230 ;
        RECT 26.470 246.220 26.730 247.430 ;
        RECT 28.860 246.320 29.110 247.870 ;
        RECT 26.470 246.060 26.860 246.220 ;
        RECT 26.460 245.930 26.860 246.060 ;
        RECT 29.560 245.930 29.820 247.540 ;
        RECT 32.110 246.470 32.410 247.520 ;
        RECT 32.860 246.920 33.160 247.870 ;
        RECT 33.360 246.970 33.660 247.020 ;
        RECT 33.360 246.620 34.260 246.970 ;
        RECT 47.020 246.570 51.490 246.600 ;
        RECT 36.080 246.540 51.490 246.570 ;
        RECT 35.410 246.520 51.490 246.540 ;
        RECT 25.080 245.720 25.370 245.880 ;
        RECT 26.460 245.870 26.720 245.930 ;
        RECT 7.710 245.610 18.410 245.620 ;
        RECT 7.710 245.570 7.990 245.610 ;
        RECT 24.580 245.530 25.370 245.720 ;
        RECT 24.580 245.330 24.830 245.530 ;
        RECT 25.080 245.420 25.370 245.530 ;
        RECT 26.470 245.330 26.720 245.870 ;
        RECT 29.550 245.870 29.820 245.930 ;
        RECT 31.100 246.210 32.410 246.470 ;
        RECT 31.100 245.870 31.410 246.210 ;
        RECT 27.110 245.340 28.750 245.730 ;
        RECT 29.550 245.580 31.410 245.870 ;
        RECT 29.550 245.570 29.860 245.580 ;
        RECT 31.100 245.570 31.410 245.580 ;
        RECT 6.510 245.010 6.780 245.090 ;
        RECT 3.910 244.780 5.350 244.990 ;
        RECT 5.900 244.790 6.780 245.010 ;
        RECT 3.910 243.730 4.190 244.780 ;
        RECT 5.900 243.980 6.120 244.790 ;
        RECT 6.510 244.760 6.780 244.790 ;
        RECT 7.640 245.050 7.930 245.100 ;
        RECT 7.640 244.870 18.390 245.050 ;
        RECT 7.640 244.770 7.930 244.870 ;
        RECT 12.480 244.860 16.110 244.870 ;
        RECT 18.190 244.190 18.390 244.870 ;
        RECT 24.580 244.730 24.870 245.330 ;
        RECT 26.470 244.730 26.760 245.330 ;
        RECT 3.190 243.280 4.190 243.730 ;
        RECT 3.170 241.830 4.470 242.280 ;
        RECT 4.170 241.430 4.470 241.830 ;
        RECT 5.890 241.450 6.120 243.980 ;
        RECT 13.140 243.890 18.390 244.190 ;
        RECT 28.810 244.120 29.110 245.120 ;
        RECT 29.560 244.520 29.860 245.570 ;
        RECT 32.160 244.470 32.410 246.210 ;
        RECT 34.530 246.200 51.490 246.520 ;
        RECT 35.410 246.190 51.490 246.200 ;
        RECT 35.410 246.160 47.390 246.190 ;
        RECT 35.410 246.150 36.300 246.160 ;
        RECT 32.860 244.120 33.120 245.670 ;
        RECT 33.950 244.120 34.150 244.130 ;
        RECT 4.960 241.430 6.120 241.450 ;
        RECT 4.170 241.250 6.120 241.430 ;
        RECT 9.060 242.250 9.320 243.450 ;
        RECT 9.060 241.740 9.310 242.250 ;
        RECT 10.950 242.240 11.210 243.450 ;
        RECT 13.340 242.340 13.590 243.890 ;
        RECT 10.950 242.080 11.340 242.240 ;
        RECT 10.940 241.950 11.340 242.080 ;
        RECT 14.040 241.950 14.300 243.560 ;
        RECT 16.590 242.490 16.890 243.540 ;
        RECT 17.340 242.940 17.640 243.890 ;
        RECT 18.190 243.880 18.390 243.890 ;
        RECT 28.760 243.820 34.150 244.120 ;
        RECT 17.840 242.990 18.140 243.040 ;
        RECT 17.840 242.640 18.740 242.990 ;
        RECT 33.950 242.580 34.150 243.820 ;
        RECT 51.110 242.620 51.470 246.190 ;
        RECT 26.390 242.560 27.580 242.570 ;
        RECT 28.570 242.560 29.760 242.570 ;
        RECT 30.790 242.560 31.980 242.570 ;
        RECT 32.970 242.560 34.160 242.580 ;
        RECT 24.180 242.550 34.160 242.560 ;
        RECT 20.790 242.530 21.980 242.540 ;
        RECT 23.070 242.530 34.160 242.550 ;
        RECT 9.560 241.740 9.850 241.900 ;
        RECT 10.940 241.890 11.200 241.950 ;
        RECT 9.060 241.550 9.850 241.740 ;
        RECT 9.060 241.350 9.310 241.550 ;
        RECT 9.560 241.440 9.850 241.550 ;
        RECT 10.950 241.350 11.200 241.890 ;
        RECT 14.030 241.890 14.300 241.950 ;
        RECT 15.580 242.230 16.890 242.490 ;
        RECT 18.950 242.300 34.160 242.530 ;
        RECT 46.240 242.320 51.490 242.620 ;
        RECT 18.950 242.290 33.110 242.300 ;
        RECT 18.950 242.280 26.480 242.290 ;
        RECT 27.490 242.280 28.680 242.290 ;
        RECT 29.640 242.280 30.830 242.290 ;
        RECT 31.920 242.280 33.110 242.290 ;
        RECT 18.950 242.270 24.260 242.280 ;
        RECT 18.950 242.260 23.120 242.270 ;
        RECT 18.950 242.250 20.840 242.260 ;
        RECT 21.930 242.250 23.120 242.260 ;
        RECT 18.950 242.240 19.670 242.250 ;
        RECT 15.580 241.890 15.890 242.230 ;
        RECT 11.590 241.360 13.230 241.750 ;
        RECT 14.030 241.600 15.890 241.890 ;
        RECT 14.030 241.590 14.340 241.600 ;
        RECT 15.580 241.590 15.890 241.600 ;
        RECT 4.170 241.240 4.820 241.250 ;
        RECT 4.170 240.910 4.470 241.240 ;
        RECT 3.450 240.460 4.470 240.910 ;
        RECT 9.060 240.750 9.350 241.350 ;
        RECT 10.950 240.750 11.240 241.350 ;
        RECT 4.170 240.450 4.470 240.460 ;
        RECT 13.290 240.140 13.590 241.140 ;
        RECT 14.040 240.540 14.340 241.590 ;
        RECT 16.640 240.490 16.890 242.230 ;
        RECT 17.340 240.140 17.600 241.690 ;
        RECT 42.160 240.680 42.420 241.880 ;
        RECT 42.160 240.170 42.410 240.680 ;
        RECT 44.050 240.670 44.310 241.880 ;
        RECT 46.440 240.770 46.690 242.320 ;
        RECT 44.050 240.510 44.440 240.670 ;
        RECT 44.040 240.380 44.440 240.510 ;
        RECT 47.140 240.380 47.400 241.990 ;
        RECT 49.690 240.920 49.990 241.970 ;
        RECT 50.440 241.370 50.740 242.320 ;
        RECT 50.940 241.420 51.240 241.470 ;
        RECT 50.940 241.070 51.840 241.420 ;
        RECT 42.660 240.170 42.950 240.330 ;
        RECT 44.040 240.320 44.300 240.380 ;
        RECT 13.240 240.130 18.490 240.140 ;
        RECT 3.120 240.050 3.370 240.060 ;
        RECT 3.120 239.590 4.100 240.050 ;
        RECT 13.240 239.840 18.510 240.130 ;
        RECT 3.120 239.290 3.370 239.590 ;
        RECT 11.090 239.500 12.930 239.510 ;
        RECT 18.340 239.500 18.510 239.840 ;
        RECT 4.830 239.490 5.070 239.500 ;
        RECT 5.910 239.490 18.510 239.500 ;
        RECT 4.830 239.330 18.510 239.490 ;
        RECT 42.160 239.980 42.950 240.170 ;
        RECT 42.160 239.780 42.410 239.980 ;
        RECT 42.660 239.870 42.950 239.980 ;
        RECT 44.050 239.780 44.300 240.320 ;
        RECT 47.130 240.320 47.400 240.380 ;
        RECT 48.680 240.660 49.990 240.920 ;
        RECT 52.050 240.960 53.720 240.990 ;
        RECT 68.800 240.960 69.050 240.970 ;
        RECT 52.050 240.690 69.050 240.960 ;
        RECT 52.050 240.680 65.550 240.690 ;
        RECT 53.330 240.660 65.550 240.680 ;
        RECT 48.680 240.320 48.990 240.660 ;
        RECT 44.690 239.790 46.330 240.180 ;
        RECT 47.130 240.030 48.990 240.320 ;
        RECT 47.130 240.020 47.440 240.030 ;
        RECT 48.680 240.020 48.990 240.030 ;
        RECT 4.830 239.320 16.340 239.330 ;
        RECT 4.820 239.310 11.140 239.320 ;
        RECT 12.690 239.310 16.340 239.320 ;
        RECT 4.820 239.300 6.690 239.310 ;
        RECT 4.820 239.290 5.070 239.300 ;
        RECT 3.120 239.120 5.070 239.290 ;
        RECT 42.160 239.180 42.450 239.780 ;
        RECT 44.050 239.180 44.340 239.780 ;
        RECT 3.120 238.900 3.370 239.120 ;
        RECT 3.120 238.730 4.160 238.900 ;
        RECT 3.970 237.870 4.160 238.730 ;
        RECT 46.390 238.570 46.690 239.570 ;
        RECT 47.140 238.970 47.440 240.020 ;
        RECT 49.740 238.920 49.990 240.660 ;
        RECT 50.440 238.570 50.700 240.120 ;
        RECT 51.320 238.570 51.660 238.640 ;
        RECT 46.340 238.270 51.660 238.570 ;
        RECT 3.180 237.430 4.160 237.870 ;
        RECT 3.180 237.420 4.130 237.430 ;
        RECT 5.000 237.110 14.270 237.120 ;
        RECT 16.150 237.110 18.070 237.120 ;
        RECT 2.850 237.010 3.040 237.020 ;
        RECT 2.850 236.550 3.830 237.010 ;
        RECT 5.000 236.920 18.070 237.110 ;
        RECT 5.000 236.910 17.360 236.920 ;
        RECT 2.850 235.760 3.040 236.550 ;
        RECT 5.000 235.900 5.210 236.910 ;
        RECT 14.260 236.900 16.160 236.910 ;
        RECT 17.890 236.170 18.070 236.920 ;
        RECT 3.850 235.760 4.120 235.770 ;
        RECT 2.850 235.550 4.120 235.760 ;
        RECT 3.850 235.340 4.120 235.550 ;
        RECT 3.850 234.710 4.100 235.340 ;
        RECT 5.000 234.890 5.200 235.900 ;
        RECT 12.810 235.870 18.070 236.170 ;
        RECT 3.060 234.260 4.100 234.710 ;
        RECT 3.040 232.810 4.000 233.260 ;
        RECT 3.750 232.760 4.000 232.810 ;
        RECT 5.010 232.760 5.200 234.890 ;
        RECT 3.750 232.560 5.200 232.760 ;
        RECT 8.730 234.230 8.990 235.430 ;
        RECT 8.730 233.720 8.980 234.230 ;
        RECT 10.620 234.220 10.880 235.430 ;
        RECT 13.010 234.320 13.260 235.870 ;
        RECT 10.620 234.060 11.010 234.220 ;
        RECT 10.610 233.930 11.010 234.060 ;
        RECT 13.710 233.930 13.970 235.540 ;
        RECT 16.260 234.470 16.560 235.520 ;
        RECT 17.010 234.920 17.310 235.870 ;
        RECT 17.510 234.970 17.810 235.020 ;
        RECT 17.510 234.620 18.410 234.970 ;
        RECT 20.120 234.840 20.340 234.850 ;
        RECT 20.120 234.650 33.800 234.840 ;
        RECT 20.120 234.520 20.340 234.650 ;
        RECT 9.230 233.720 9.520 233.880 ;
        RECT 10.610 233.870 10.870 233.930 ;
        RECT 8.730 233.530 9.520 233.720 ;
        RECT 8.730 233.330 8.980 233.530 ;
        RECT 9.230 233.420 9.520 233.530 ;
        RECT 10.620 233.330 10.870 233.870 ;
        RECT 13.700 233.870 13.970 233.930 ;
        RECT 15.250 234.210 16.560 234.470 ;
        RECT 18.660 234.220 20.340 234.520 ;
        RECT 18.660 234.210 20.320 234.220 ;
        RECT 15.250 233.870 15.560 234.210 ;
        RECT 11.260 233.340 12.900 233.730 ;
        RECT 13.700 233.580 15.560 233.870 ;
        RECT 13.700 233.570 14.010 233.580 ;
        RECT 15.250 233.570 15.560 233.580 ;
        RECT 8.730 232.730 9.020 233.330 ;
        RECT 10.620 232.730 10.910 233.330 ;
        RECT 3.750 232.470 4.000 232.560 ;
        RECT 3.020 232.020 4.000 232.470 ;
        RECT 12.960 232.120 13.260 233.120 ;
        RECT 13.710 232.520 14.010 233.570 ;
        RECT 16.310 232.470 16.560 234.210 ;
        RECT 33.550 233.750 33.800 234.650 ;
        RECT 17.010 232.120 17.270 233.670 ;
        RECT 28.490 233.450 33.800 233.750 ;
        RECT 12.910 232.100 18.160 232.120 ;
        RECT 12.910 231.820 18.280 232.100 ;
        RECT 6.360 231.420 6.640 231.490 ;
        RECT 7.540 231.450 7.820 231.480 ;
        RECT 17.990 231.450 18.280 231.820 ;
        RECT 7.540 231.440 18.280 231.450 ;
        RECT 4.950 231.220 6.640 231.420 ;
        RECT 3.740 231.020 4.020 231.030 ;
        RECT 3.000 230.570 4.020 231.020 ;
        RECT 4.950 230.570 5.180 231.220 ;
        RECT 6.360 231.160 6.640 231.220 ;
        RECT 7.520 231.210 18.280 231.440 ;
        RECT 7.540 231.200 18.280 231.210 ;
        RECT 24.410 231.810 24.670 233.010 ;
        RECT 24.410 231.300 24.660 231.810 ;
        RECT 26.300 231.800 26.560 233.010 ;
        RECT 28.690 231.900 28.940 233.450 ;
        RECT 26.300 231.640 26.690 231.800 ;
        RECT 26.290 231.510 26.690 231.640 ;
        RECT 29.390 231.510 29.650 233.120 ;
        RECT 31.940 232.050 32.240 233.100 ;
        RECT 32.690 232.500 32.990 233.450 ;
        RECT 33.190 232.550 33.490 232.600 ;
        RECT 33.190 232.200 34.090 232.550 ;
        RECT 51.320 232.150 51.660 238.270 ;
        RECT 50.750 232.130 51.710 232.150 ;
        RECT 35.230 232.110 39.510 232.120 ;
        RECT 46.910 232.110 51.710 232.130 ;
        RECT 35.230 232.100 51.710 232.110 ;
        RECT 24.910 231.300 25.200 231.460 ;
        RECT 26.290 231.450 26.550 231.510 ;
        RECT 7.540 231.190 18.240 231.200 ;
        RECT 7.540 231.150 7.820 231.190 ;
        RECT 24.410 231.110 25.200 231.300 ;
        RECT 24.410 230.910 24.660 231.110 ;
        RECT 24.910 231.000 25.200 231.110 ;
        RECT 26.300 230.910 26.550 231.450 ;
        RECT 29.380 231.450 29.650 231.510 ;
        RECT 30.930 231.790 32.240 232.050 ;
        RECT 30.930 231.450 31.240 231.790 ;
        RECT 26.940 230.920 28.580 231.310 ;
        RECT 29.380 231.160 31.240 231.450 ;
        RECT 29.380 231.150 29.690 231.160 ;
        RECT 30.930 231.150 31.240 231.160 ;
        RECT 6.340 230.590 6.610 230.670 ;
        RECT 3.740 230.360 5.180 230.570 ;
        RECT 5.730 230.370 6.610 230.590 ;
        RECT 3.740 229.310 4.020 230.360 ;
        RECT 5.730 229.560 5.950 230.370 ;
        RECT 6.340 230.340 6.610 230.370 ;
        RECT 7.470 230.630 7.760 230.680 ;
        RECT 7.470 230.450 18.220 230.630 ;
        RECT 7.470 230.350 7.760 230.450 ;
        RECT 12.310 230.440 15.940 230.450 ;
        RECT 18.020 229.770 18.220 230.450 ;
        RECT 24.410 230.310 24.700 230.910 ;
        RECT 26.300 230.310 26.590 230.910 ;
        RECT 3.020 228.860 4.020 229.310 ;
        RECT 3.000 227.410 4.300 227.860 ;
        RECT 4.000 227.010 4.300 227.410 ;
        RECT 5.720 227.030 5.950 229.560 ;
        RECT 12.970 229.470 18.220 229.770 ;
        RECT 28.640 229.700 28.940 230.700 ;
        RECT 29.390 230.100 29.690 231.150 ;
        RECT 31.990 230.050 32.240 231.790 ;
        RECT 34.360 231.790 51.710 232.100 ;
        RECT 34.360 231.780 47.370 231.790 ;
        RECT 39.220 231.770 47.370 231.780 ;
        RECT 50.750 231.750 51.710 231.790 ;
        RECT 51.320 231.740 51.660 231.750 ;
        RECT 32.690 229.700 32.950 231.250 ;
        RECT 33.780 229.700 33.980 229.710 ;
        RECT 4.790 227.010 5.950 227.030 ;
        RECT 4.000 226.830 5.950 227.010 ;
        RECT 8.890 227.830 9.150 229.030 ;
        RECT 8.890 227.320 9.140 227.830 ;
        RECT 10.780 227.820 11.040 229.030 ;
        RECT 13.170 227.920 13.420 229.470 ;
        RECT 10.780 227.660 11.170 227.820 ;
        RECT 10.770 227.530 11.170 227.660 ;
        RECT 13.870 227.530 14.130 229.140 ;
        RECT 16.420 228.070 16.720 229.120 ;
        RECT 17.170 228.520 17.470 229.470 ;
        RECT 18.020 229.460 18.220 229.470 ;
        RECT 28.590 229.400 33.980 229.700 ;
        RECT 17.670 228.570 17.970 228.620 ;
        RECT 17.670 228.220 18.570 228.570 ;
        RECT 33.780 228.160 33.980 229.400 ;
        RECT 26.220 228.140 27.410 228.150 ;
        RECT 28.400 228.140 29.590 228.150 ;
        RECT 30.620 228.140 31.810 228.150 ;
        RECT 32.800 228.140 33.990 228.160 ;
        RECT 24.010 228.130 33.990 228.140 ;
        RECT 20.620 228.110 21.810 228.120 ;
        RECT 22.900 228.110 33.990 228.130 ;
        RECT 9.390 227.320 9.680 227.480 ;
        RECT 10.770 227.470 11.030 227.530 ;
        RECT 8.890 227.130 9.680 227.320 ;
        RECT 8.890 226.930 9.140 227.130 ;
        RECT 9.390 227.020 9.680 227.130 ;
        RECT 10.780 226.930 11.030 227.470 ;
        RECT 13.860 227.470 14.130 227.530 ;
        RECT 15.410 227.810 16.720 228.070 ;
        RECT 18.780 227.880 33.990 228.110 ;
        RECT 18.780 227.870 32.940 227.880 ;
        RECT 18.780 227.860 26.310 227.870 ;
        RECT 27.320 227.860 28.510 227.870 ;
        RECT 29.470 227.860 30.660 227.870 ;
        RECT 31.750 227.860 32.940 227.870 ;
        RECT 18.780 227.850 24.090 227.860 ;
        RECT 18.780 227.840 22.950 227.850 ;
        RECT 18.780 227.830 20.670 227.840 ;
        RECT 21.760 227.830 22.950 227.840 ;
        RECT 18.780 227.820 19.500 227.830 ;
        RECT 15.410 227.470 15.720 227.810 ;
        RECT 11.420 226.940 13.060 227.330 ;
        RECT 13.860 227.180 15.720 227.470 ;
        RECT 13.860 227.170 14.170 227.180 ;
        RECT 15.410 227.170 15.720 227.180 ;
        RECT 4.000 226.820 4.650 226.830 ;
        RECT 4.000 226.490 4.300 226.820 ;
        RECT 3.280 226.040 4.300 226.490 ;
        RECT 8.890 226.330 9.180 226.930 ;
        RECT 10.780 226.330 11.070 226.930 ;
        RECT 4.000 226.030 4.300 226.040 ;
        RECT 13.120 225.720 13.420 226.720 ;
        RECT 13.870 226.120 14.170 227.170 ;
        RECT 16.470 226.070 16.720 227.810 ;
        RECT 68.800 227.550 69.060 240.690 ;
        RECT 68.790 227.430 69.060 227.550 ;
        RECT 17.170 225.720 17.430 227.270 ;
        RECT 68.790 226.600 69.050 227.430 ;
        RECT 63.770 226.300 69.050 226.600 ;
        RECT 13.070 225.710 18.320 225.720 ;
        RECT 2.950 225.630 3.200 225.640 ;
        RECT 2.950 225.170 3.930 225.630 ;
        RECT 13.070 225.420 18.340 225.710 ;
        RECT 2.950 224.870 3.200 225.170 ;
        RECT 10.920 225.080 12.760 225.090 ;
        RECT 18.170 225.080 18.340 225.420 ;
        RECT 4.660 225.070 4.900 225.080 ;
        RECT 5.740 225.070 18.340 225.080 ;
        RECT 4.660 224.910 18.340 225.070 ;
        RECT 4.660 224.900 16.170 224.910 ;
        RECT 4.650 224.890 10.970 224.900 ;
        RECT 12.520 224.890 16.170 224.900 ;
        RECT 4.650 224.880 6.520 224.890 ;
        RECT 4.650 224.870 4.900 224.880 ;
        RECT 2.950 224.700 4.900 224.870 ;
        RECT 2.950 224.400 3.220 224.700 ;
        RECT 2.960 224.140 3.220 224.400 ;
        RECT 59.690 224.660 59.950 225.860 ;
        RECT 59.690 224.150 59.940 224.660 ;
        RECT 61.580 224.650 61.840 225.860 ;
        RECT 63.970 224.750 64.220 226.300 ;
        RECT 61.580 224.490 61.970 224.650 ;
        RECT 61.570 224.360 61.970 224.490 ;
        RECT 64.670 224.360 64.930 225.970 ;
        RECT 67.220 224.900 67.520 225.950 ;
        RECT 67.970 225.350 68.270 226.300 ;
        RECT 68.470 225.400 68.770 225.450 ;
        RECT 68.470 225.050 69.370 225.400 ;
        RECT 60.190 224.150 60.480 224.310 ;
        RECT 61.570 224.300 61.830 224.360 ;
        RECT 2.940 223.750 3.240 224.140 ;
        RECT 59.690 223.960 60.480 224.150 ;
        RECT 59.690 223.760 59.940 223.960 ;
        RECT 60.190 223.850 60.480 223.960 ;
        RECT 61.580 223.760 61.830 224.300 ;
        RECT 64.660 224.300 64.930 224.360 ;
        RECT 66.210 224.640 67.520 224.900 ;
        RECT 69.640 224.840 70.420 224.940 ;
        RECT 69.640 224.670 83.220 224.840 ;
        RECT 69.640 224.660 83.210 224.670 ;
        RECT 69.640 224.640 70.420 224.660 ;
        RECT 66.210 224.300 66.520 224.640 ;
        RECT 62.220 223.770 63.860 224.160 ;
        RECT 64.660 224.010 66.520 224.300 ;
        RECT 64.660 224.000 64.970 224.010 ;
        RECT 66.210 224.000 66.520 224.010 ;
        RECT 2.940 223.520 4.430 223.750 ;
        RECT 4.180 222.590 4.430 223.520 ;
        RECT 59.690 223.160 59.980 223.760 ;
        RECT 61.580 223.160 61.870 223.760 ;
        RECT 3.380 222.130 4.430 222.590 ;
        RECT 63.920 222.550 64.220 223.550 ;
        RECT 64.670 222.950 64.970 224.000 ;
        RECT 67.270 222.900 67.520 224.640 ;
        RECT 67.970 222.550 68.230 224.100 ;
        RECT 63.870 222.250 69.140 222.550 ;
        RECT 4.180 222.120 4.430 222.130 ;
        RECT 3.050 221.720 3.300 221.730 ;
        RECT 3.050 221.270 4.030 221.720 ;
        RECT 5.140 221.460 14.410 221.470 ;
        RECT 16.290 221.460 18.210 221.470 ;
        RECT 5.140 221.270 18.210 221.460 ;
        RECT 3.050 220.660 3.300 221.270 ;
        RECT 5.140 221.260 17.500 221.270 ;
        RECT 3.050 220.410 4.260 220.660 ;
        RECT 3.990 219.660 4.250 220.410 ;
        RECT 5.140 220.250 5.350 221.260 ;
        RECT 14.400 221.250 16.300 221.260 ;
        RECT 18.030 220.520 18.210 221.270 ;
        RECT 3.990 219.060 4.240 219.660 ;
        RECT 5.140 219.240 5.340 220.250 ;
        RECT 12.950 220.220 18.210 220.520 ;
        RECT 3.200 218.610 4.240 219.060 ;
        RECT 3.180 217.160 4.140 217.610 ;
        RECT 3.890 217.110 4.140 217.160 ;
        RECT 5.150 217.110 5.340 219.240 ;
        RECT 3.890 216.910 5.340 217.110 ;
        RECT 8.870 218.580 9.130 219.780 ;
        RECT 8.870 218.070 9.120 218.580 ;
        RECT 10.760 218.570 11.020 219.780 ;
        RECT 13.150 218.670 13.400 220.220 ;
        RECT 10.760 218.410 11.150 218.570 ;
        RECT 10.750 218.280 11.150 218.410 ;
        RECT 13.850 218.280 14.110 219.890 ;
        RECT 16.400 218.820 16.700 219.870 ;
        RECT 17.150 219.270 17.450 220.220 ;
        RECT 17.650 219.320 17.950 219.370 ;
        RECT 17.650 218.970 18.550 219.320 ;
        RECT 20.260 219.190 20.480 219.200 ;
        RECT 20.260 219.000 33.940 219.190 ;
        RECT 20.260 218.870 20.480 219.000 ;
        RECT 9.370 218.070 9.660 218.230 ;
        RECT 10.750 218.220 11.010 218.280 ;
        RECT 8.870 217.880 9.660 218.070 ;
        RECT 8.870 217.680 9.120 217.880 ;
        RECT 9.370 217.770 9.660 217.880 ;
        RECT 10.760 217.680 11.010 218.220 ;
        RECT 13.840 218.220 14.110 218.280 ;
        RECT 15.390 218.560 16.700 218.820 ;
        RECT 18.800 218.570 20.480 218.870 ;
        RECT 18.800 218.560 20.460 218.570 ;
        RECT 15.390 218.220 15.700 218.560 ;
        RECT 11.400 217.690 13.040 218.080 ;
        RECT 13.840 217.930 15.700 218.220 ;
        RECT 13.840 217.920 14.150 217.930 ;
        RECT 15.390 217.920 15.700 217.930 ;
        RECT 8.870 217.080 9.160 217.680 ;
        RECT 10.760 217.080 11.050 217.680 ;
        RECT 3.890 216.820 4.140 216.910 ;
        RECT 3.160 216.370 4.140 216.820 ;
        RECT 13.100 216.470 13.400 217.470 ;
        RECT 13.850 216.870 14.150 217.920 ;
        RECT 16.450 216.820 16.700 218.560 ;
        RECT 33.690 218.100 33.940 219.000 ;
        RECT 17.150 216.470 17.410 218.020 ;
        RECT 28.630 217.800 33.940 218.100 ;
        RECT 13.050 216.450 18.300 216.470 ;
        RECT 13.050 216.170 18.420 216.450 ;
        RECT 6.500 215.770 6.780 215.840 ;
        RECT 7.680 215.800 7.960 215.830 ;
        RECT 18.130 215.800 18.420 216.170 ;
        RECT 7.680 215.790 18.420 215.800 ;
        RECT 5.090 215.570 6.780 215.770 ;
        RECT 3.880 215.370 4.160 215.380 ;
        RECT 3.140 214.920 4.160 215.370 ;
        RECT 5.090 214.920 5.320 215.570 ;
        RECT 6.500 215.510 6.780 215.570 ;
        RECT 7.660 215.560 18.420 215.790 ;
        RECT 7.680 215.550 18.420 215.560 ;
        RECT 24.550 216.160 24.810 217.360 ;
        RECT 24.550 215.650 24.800 216.160 ;
        RECT 26.440 216.150 26.700 217.360 ;
        RECT 28.830 216.250 29.080 217.800 ;
        RECT 26.440 215.990 26.830 216.150 ;
        RECT 26.430 215.860 26.830 215.990 ;
        RECT 29.530 215.860 29.790 217.470 ;
        RECT 32.080 216.400 32.380 217.450 ;
        RECT 32.830 216.850 33.130 217.800 ;
        RECT 33.330 216.900 33.630 216.950 ;
        RECT 33.330 216.550 34.230 216.900 ;
        RECT 46.990 216.500 51.460 216.530 ;
        RECT 36.050 216.470 51.460 216.500 ;
        RECT 35.380 216.450 51.460 216.470 ;
        RECT 25.050 215.650 25.340 215.810 ;
        RECT 26.430 215.800 26.690 215.860 ;
        RECT 7.680 215.540 18.380 215.550 ;
        RECT 7.680 215.500 7.960 215.540 ;
        RECT 24.550 215.460 25.340 215.650 ;
        RECT 24.550 215.260 24.800 215.460 ;
        RECT 25.050 215.350 25.340 215.460 ;
        RECT 26.440 215.260 26.690 215.800 ;
        RECT 29.520 215.800 29.790 215.860 ;
        RECT 31.070 216.140 32.380 216.400 ;
        RECT 31.070 215.800 31.380 216.140 ;
        RECT 27.080 215.270 28.720 215.660 ;
        RECT 29.520 215.510 31.380 215.800 ;
        RECT 29.520 215.500 29.830 215.510 ;
        RECT 31.070 215.500 31.380 215.510 ;
        RECT 6.480 214.940 6.750 215.020 ;
        RECT 3.880 214.710 5.320 214.920 ;
        RECT 5.870 214.720 6.750 214.940 ;
        RECT 3.880 213.660 4.160 214.710 ;
        RECT 5.870 213.910 6.090 214.720 ;
        RECT 6.480 214.690 6.750 214.720 ;
        RECT 7.610 214.980 7.900 215.030 ;
        RECT 7.610 214.800 18.360 214.980 ;
        RECT 7.610 214.700 7.900 214.800 ;
        RECT 12.450 214.790 16.080 214.800 ;
        RECT 18.160 214.120 18.360 214.800 ;
        RECT 24.550 214.660 24.840 215.260 ;
        RECT 26.440 214.660 26.730 215.260 ;
        RECT 3.160 213.210 4.160 213.660 ;
        RECT 3.140 211.760 4.440 212.210 ;
        RECT 4.140 211.360 4.440 211.760 ;
        RECT 5.860 211.380 6.090 213.910 ;
        RECT 13.110 213.820 18.360 214.120 ;
        RECT 28.780 214.050 29.080 215.050 ;
        RECT 29.530 214.450 29.830 215.500 ;
        RECT 32.130 214.400 32.380 216.140 ;
        RECT 34.500 216.130 51.460 216.450 ;
        RECT 35.380 216.120 51.460 216.130 ;
        RECT 35.380 216.090 47.360 216.120 ;
        RECT 35.380 216.080 36.270 216.090 ;
        RECT 32.830 214.050 33.090 215.600 ;
        RECT 33.920 214.050 34.120 214.060 ;
        RECT 4.930 211.360 6.090 211.380 ;
        RECT 4.140 211.180 6.090 211.360 ;
        RECT 9.030 212.180 9.290 213.380 ;
        RECT 9.030 211.670 9.280 212.180 ;
        RECT 10.920 212.170 11.180 213.380 ;
        RECT 13.310 212.270 13.560 213.820 ;
        RECT 10.920 212.010 11.310 212.170 ;
        RECT 10.910 211.880 11.310 212.010 ;
        RECT 14.010 211.880 14.270 213.490 ;
        RECT 16.560 212.420 16.860 213.470 ;
        RECT 17.310 212.870 17.610 213.820 ;
        RECT 18.160 213.810 18.360 213.820 ;
        RECT 28.730 213.750 34.120 214.050 ;
        RECT 17.810 212.920 18.110 212.970 ;
        RECT 17.810 212.570 18.710 212.920 ;
        RECT 33.920 212.510 34.120 213.750 ;
        RECT 51.080 212.550 51.440 216.120 ;
        RECT 26.360 212.490 27.550 212.500 ;
        RECT 28.540 212.490 29.730 212.500 ;
        RECT 30.760 212.490 31.950 212.500 ;
        RECT 32.940 212.490 34.130 212.510 ;
        RECT 24.150 212.480 34.130 212.490 ;
        RECT 20.760 212.460 21.950 212.470 ;
        RECT 23.040 212.460 34.130 212.480 ;
        RECT 9.530 211.670 9.820 211.830 ;
        RECT 10.910 211.820 11.170 211.880 ;
        RECT 9.030 211.480 9.820 211.670 ;
        RECT 9.030 211.280 9.280 211.480 ;
        RECT 9.530 211.370 9.820 211.480 ;
        RECT 10.920 211.280 11.170 211.820 ;
        RECT 14.000 211.820 14.270 211.880 ;
        RECT 15.550 212.160 16.860 212.420 ;
        RECT 18.920 212.230 34.130 212.460 ;
        RECT 46.210 212.250 51.460 212.550 ;
        RECT 18.920 212.220 33.080 212.230 ;
        RECT 18.920 212.210 26.450 212.220 ;
        RECT 27.460 212.210 28.650 212.220 ;
        RECT 29.610 212.210 30.800 212.220 ;
        RECT 31.890 212.210 33.080 212.220 ;
        RECT 18.920 212.200 24.230 212.210 ;
        RECT 18.920 212.190 23.090 212.200 ;
        RECT 18.920 212.180 20.810 212.190 ;
        RECT 21.900 212.180 23.090 212.190 ;
        RECT 18.920 212.170 19.640 212.180 ;
        RECT 15.550 211.820 15.860 212.160 ;
        RECT 11.560 211.290 13.200 211.680 ;
        RECT 14.000 211.530 15.860 211.820 ;
        RECT 14.000 211.520 14.310 211.530 ;
        RECT 15.550 211.520 15.860 211.530 ;
        RECT 4.140 211.170 4.790 211.180 ;
        RECT 4.140 210.840 4.440 211.170 ;
        RECT 3.420 210.390 4.440 210.840 ;
        RECT 9.030 210.680 9.320 211.280 ;
        RECT 10.920 210.680 11.210 211.280 ;
        RECT 4.140 210.380 4.440 210.390 ;
        RECT 13.260 210.070 13.560 211.070 ;
        RECT 14.010 210.470 14.310 211.520 ;
        RECT 16.610 210.420 16.860 212.160 ;
        RECT 17.310 210.070 17.570 211.620 ;
        RECT 42.130 210.610 42.390 211.810 ;
        RECT 42.130 210.100 42.380 210.610 ;
        RECT 44.020 210.600 44.280 211.810 ;
        RECT 46.410 210.700 46.660 212.250 ;
        RECT 44.020 210.440 44.410 210.600 ;
        RECT 44.010 210.310 44.410 210.440 ;
        RECT 47.110 210.310 47.370 211.920 ;
        RECT 49.660 210.850 49.960 211.900 ;
        RECT 50.410 211.300 50.710 212.250 ;
        RECT 50.910 211.350 51.210 211.400 ;
        RECT 50.910 211.000 51.810 211.350 ;
        RECT 42.630 210.100 42.920 210.260 ;
        RECT 44.010 210.250 44.270 210.310 ;
        RECT 13.210 210.060 18.460 210.070 ;
        RECT 3.090 209.980 3.340 209.990 ;
        RECT 3.090 209.520 4.070 209.980 ;
        RECT 13.210 209.770 18.480 210.060 ;
        RECT 3.090 209.220 3.340 209.520 ;
        RECT 11.060 209.430 12.900 209.440 ;
        RECT 18.310 209.430 18.480 209.770 ;
        RECT 4.800 209.420 5.040 209.430 ;
        RECT 5.880 209.420 18.480 209.430 ;
        RECT 4.800 209.260 18.480 209.420 ;
        RECT 42.130 209.910 42.920 210.100 ;
        RECT 42.130 209.710 42.380 209.910 ;
        RECT 42.630 209.800 42.920 209.910 ;
        RECT 44.020 209.710 44.270 210.250 ;
        RECT 47.100 210.250 47.370 210.310 ;
        RECT 48.650 210.590 49.960 210.850 ;
        RECT 52.020 210.900 53.690 210.920 ;
        RECT 68.830 210.900 69.140 222.250 ;
        RECT 52.020 210.610 69.180 210.900 ;
        RECT 52.710 210.600 69.180 210.610 ;
        RECT 48.650 210.250 48.960 210.590 ;
        RECT 44.660 209.720 46.300 210.110 ;
        RECT 47.100 209.960 48.960 210.250 ;
        RECT 47.100 209.950 47.410 209.960 ;
        RECT 48.650 209.950 48.960 209.960 ;
        RECT 4.800 209.250 16.310 209.260 ;
        RECT 4.790 209.240 11.110 209.250 ;
        RECT 12.660 209.240 16.310 209.250 ;
        RECT 4.790 209.230 6.660 209.240 ;
        RECT 4.790 209.220 5.040 209.230 ;
        RECT 3.090 209.050 5.040 209.220 ;
        RECT 42.130 209.110 42.420 209.710 ;
        RECT 44.020 209.110 44.310 209.710 ;
        RECT 3.090 208.830 3.340 209.050 ;
        RECT 3.090 208.660 4.130 208.830 ;
        RECT 3.940 207.800 4.130 208.660 ;
        RECT 46.360 208.500 46.660 209.500 ;
        RECT 47.110 208.900 47.410 209.950 ;
        RECT 49.710 208.850 49.960 210.590 ;
        RECT 50.410 208.500 50.670 210.050 ;
        RECT 51.290 208.500 51.630 208.570 ;
        RECT 46.310 208.200 51.630 208.500 ;
        RECT 3.150 207.360 4.130 207.800 ;
        RECT 3.150 207.350 4.100 207.360 ;
        RECT 4.970 207.040 14.240 207.050 ;
        RECT 16.120 207.040 18.040 207.050 ;
        RECT 2.820 206.940 3.010 206.950 ;
        RECT 2.820 206.480 3.800 206.940 ;
        RECT 4.970 206.850 18.040 207.040 ;
        RECT 4.970 206.840 17.330 206.850 ;
        RECT 2.820 205.690 3.010 206.480 ;
        RECT 4.970 205.830 5.180 206.840 ;
        RECT 14.230 206.830 16.130 206.840 ;
        RECT 17.860 206.100 18.040 206.850 ;
        RECT 3.820 205.690 4.090 205.700 ;
        RECT 2.820 205.480 4.090 205.690 ;
        RECT 3.820 205.270 4.090 205.480 ;
        RECT 3.820 204.640 4.070 205.270 ;
        RECT 4.970 204.820 5.170 205.830 ;
        RECT 12.780 205.800 18.040 206.100 ;
        RECT 3.030 204.190 4.070 204.640 ;
        RECT 3.010 202.740 3.970 203.190 ;
        RECT 3.720 202.690 3.970 202.740 ;
        RECT 4.980 202.690 5.170 204.820 ;
        RECT 3.720 202.490 5.170 202.690 ;
        RECT 8.700 204.160 8.960 205.360 ;
        RECT 8.700 203.650 8.950 204.160 ;
        RECT 10.590 204.150 10.850 205.360 ;
        RECT 12.980 204.250 13.230 205.800 ;
        RECT 10.590 203.990 10.980 204.150 ;
        RECT 10.580 203.860 10.980 203.990 ;
        RECT 13.680 203.860 13.940 205.470 ;
        RECT 16.230 204.400 16.530 205.450 ;
        RECT 16.980 204.850 17.280 205.800 ;
        RECT 17.480 204.900 17.780 204.950 ;
        RECT 17.480 204.550 18.380 204.900 ;
        RECT 20.090 204.770 20.310 204.780 ;
        RECT 20.090 204.580 33.770 204.770 ;
        RECT 20.090 204.450 20.310 204.580 ;
        RECT 9.200 203.650 9.490 203.810 ;
        RECT 10.580 203.800 10.840 203.860 ;
        RECT 8.700 203.460 9.490 203.650 ;
        RECT 8.700 203.260 8.950 203.460 ;
        RECT 9.200 203.350 9.490 203.460 ;
        RECT 10.590 203.260 10.840 203.800 ;
        RECT 13.670 203.800 13.940 203.860 ;
        RECT 15.220 204.140 16.530 204.400 ;
        RECT 18.630 204.150 20.310 204.450 ;
        RECT 18.630 204.140 20.290 204.150 ;
        RECT 15.220 203.800 15.530 204.140 ;
        RECT 11.230 203.270 12.870 203.660 ;
        RECT 13.670 203.510 15.530 203.800 ;
        RECT 13.670 203.500 13.980 203.510 ;
        RECT 15.220 203.500 15.530 203.510 ;
        RECT 8.700 202.660 8.990 203.260 ;
        RECT 10.590 202.660 10.880 203.260 ;
        RECT 3.720 202.400 3.970 202.490 ;
        RECT 2.990 201.950 3.970 202.400 ;
        RECT 12.930 202.050 13.230 203.050 ;
        RECT 13.680 202.450 13.980 203.500 ;
        RECT 16.280 202.400 16.530 204.140 ;
        RECT 33.520 203.680 33.770 204.580 ;
        RECT 16.980 202.050 17.240 203.600 ;
        RECT 28.460 203.380 33.770 203.680 ;
        RECT 12.880 202.030 18.130 202.050 ;
        RECT 12.880 201.750 18.250 202.030 ;
        RECT 6.330 201.350 6.610 201.420 ;
        RECT 7.510 201.380 7.790 201.410 ;
        RECT 17.960 201.380 18.250 201.750 ;
        RECT 7.510 201.370 18.250 201.380 ;
        RECT 4.920 201.150 6.610 201.350 ;
        RECT 3.710 200.950 3.990 200.960 ;
        RECT 2.970 200.500 3.990 200.950 ;
        RECT 4.920 200.500 5.150 201.150 ;
        RECT 6.330 201.090 6.610 201.150 ;
        RECT 7.490 201.140 18.250 201.370 ;
        RECT 7.510 201.130 18.250 201.140 ;
        RECT 24.380 201.740 24.640 202.940 ;
        RECT 24.380 201.230 24.630 201.740 ;
        RECT 26.270 201.730 26.530 202.940 ;
        RECT 28.660 201.830 28.910 203.380 ;
        RECT 26.270 201.570 26.660 201.730 ;
        RECT 26.260 201.440 26.660 201.570 ;
        RECT 29.360 201.440 29.620 203.050 ;
        RECT 31.910 201.980 32.210 203.030 ;
        RECT 32.660 202.430 32.960 203.380 ;
        RECT 33.160 202.480 33.460 202.530 ;
        RECT 33.160 202.130 34.060 202.480 ;
        RECT 51.290 202.080 51.630 208.200 ;
        RECT 83.030 205.400 83.210 224.660 ;
        RECT 83.010 204.350 83.220 205.400 ;
        RECT 83.010 204.270 83.230 204.350 ;
        RECT 83.020 202.200 83.230 204.270 ;
        RECT 83.010 202.160 83.230 202.200 ;
        RECT 50.720 202.060 51.680 202.080 ;
        RECT 35.200 202.040 39.480 202.050 ;
        RECT 46.880 202.040 51.680 202.060 ;
        RECT 35.200 202.030 51.680 202.040 ;
        RECT 24.880 201.230 25.170 201.390 ;
        RECT 26.260 201.380 26.520 201.440 ;
        RECT 7.510 201.120 18.210 201.130 ;
        RECT 7.510 201.080 7.790 201.120 ;
        RECT 24.380 201.040 25.170 201.230 ;
        RECT 24.380 200.840 24.630 201.040 ;
        RECT 24.880 200.930 25.170 201.040 ;
        RECT 26.270 200.840 26.520 201.380 ;
        RECT 29.350 201.380 29.620 201.440 ;
        RECT 30.900 201.720 32.210 201.980 ;
        RECT 30.900 201.380 31.210 201.720 ;
        RECT 26.910 200.850 28.550 201.240 ;
        RECT 29.350 201.090 31.210 201.380 ;
        RECT 29.350 201.080 29.660 201.090 ;
        RECT 30.900 201.080 31.210 201.090 ;
        RECT 6.310 200.520 6.580 200.600 ;
        RECT 3.710 200.290 5.150 200.500 ;
        RECT 5.700 200.300 6.580 200.520 ;
        RECT 3.710 199.240 3.990 200.290 ;
        RECT 5.700 199.490 5.920 200.300 ;
        RECT 6.310 200.270 6.580 200.300 ;
        RECT 7.440 200.560 7.730 200.610 ;
        RECT 7.440 200.380 18.190 200.560 ;
        RECT 7.440 200.280 7.730 200.380 ;
        RECT 12.280 200.370 15.910 200.380 ;
        RECT 17.990 199.700 18.190 200.380 ;
        RECT 24.380 200.240 24.670 200.840 ;
        RECT 26.270 200.240 26.560 200.840 ;
        RECT 2.990 198.790 3.990 199.240 ;
        RECT 2.970 197.340 4.270 197.790 ;
        RECT 3.970 196.940 4.270 197.340 ;
        RECT 5.690 196.960 5.920 199.490 ;
        RECT 12.940 199.400 18.190 199.700 ;
        RECT 28.610 199.630 28.910 200.630 ;
        RECT 29.360 200.030 29.660 201.080 ;
        RECT 31.960 199.980 32.210 201.720 ;
        RECT 34.330 201.720 51.680 202.030 ;
        RECT 34.330 201.710 47.340 201.720 ;
        RECT 39.190 201.700 47.340 201.710 ;
        RECT 50.720 201.680 51.680 201.720 ;
        RECT 51.290 201.670 51.630 201.680 ;
        RECT 32.660 199.630 32.920 201.180 ;
        RECT 83.010 200.310 83.220 202.160 ;
        RECT 77.970 200.010 83.220 200.310 ;
        RECT 33.750 199.630 33.950 199.640 ;
        RECT 4.760 196.940 5.920 196.960 ;
        RECT 3.970 196.760 5.920 196.940 ;
        RECT 8.860 197.760 9.120 198.960 ;
        RECT 8.860 197.250 9.110 197.760 ;
        RECT 10.750 197.750 11.010 198.960 ;
        RECT 13.140 197.850 13.390 199.400 ;
        RECT 10.750 197.590 11.140 197.750 ;
        RECT 10.740 197.460 11.140 197.590 ;
        RECT 13.840 197.460 14.100 199.070 ;
        RECT 16.390 198.000 16.690 199.050 ;
        RECT 17.140 198.450 17.440 199.400 ;
        RECT 17.990 199.390 18.190 199.400 ;
        RECT 28.560 199.330 33.950 199.630 ;
        RECT 17.640 198.500 17.940 198.550 ;
        RECT 17.640 198.150 18.540 198.500 ;
        RECT 33.750 198.090 33.950 199.330 ;
        RECT 73.890 198.370 74.150 199.570 ;
        RECT 26.190 198.070 27.380 198.080 ;
        RECT 28.370 198.070 29.560 198.080 ;
        RECT 30.590 198.070 31.780 198.080 ;
        RECT 32.770 198.070 33.960 198.090 ;
        RECT 23.980 198.060 33.960 198.070 ;
        RECT 20.590 198.040 21.780 198.050 ;
        RECT 22.870 198.040 33.960 198.060 ;
        RECT 9.360 197.250 9.650 197.410 ;
        RECT 10.740 197.400 11.000 197.460 ;
        RECT 8.860 197.060 9.650 197.250 ;
        RECT 8.860 196.860 9.110 197.060 ;
        RECT 9.360 196.950 9.650 197.060 ;
        RECT 10.750 196.860 11.000 197.400 ;
        RECT 13.830 197.400 14.100 197.460 ;
        RECT 15.380 197.740 16.690 198.000 ;
        RECT 18.750 197.810 33.960 198.040 ;
        RECT 73.890 197.860 74.140 198.370 ;
        RECT 75.780 198.360 76.040 199.570 ;
        RECT 78.170 198.460 78.420 200.010 ;
        RECT 75.780 198.200 76.170 198.360 ;
        RECT 75.770 198.070 76.170 198.200 ;
        RECT 78.870 198.070 79.130 199.680 ;
        RECT 81.420 198.610 81.720 199.660 ;
        RECT 82.170 199.060 82.470 200.010 ;
        RECT 83.010 200.000 83.220 200.010 ;
        RECT 82.670 199.110 82.970 199.160 ;
        RECT 82.670 198.760 83.570 199.110 ;
        RECT 84.530 198.640 99.520 198.710 ;
        RECT 74.390 197.860 74.680 198.020 ;
        RECT 75.770 198.010 76.030 198.070 ;
        RECT 18.750 197.800 32.910 197.810 ;
        RECT 18.750 197.790 26.280 197.800 ;
        RECT 27.290 197.790 28.480 197.800 ;
        RECT 29.440 197.790 30.630 197.800 ;
        RECT 31.720 197.790 32.910 197.800 ;
        RECT 18.750 197.780 24.060 197.790 ;
        RECT 18.750 197.770 22.920 197.780 ;
        RECT 18.750 197.760 20.640 197.770 ;
        RECT 21.730 197.760 22.920 197.770 ;
        RECT 18.750 197.750 19.470 197.760 ;
        RECT 15.380 197.400 15.690 197.740 ;
        RECT 11.390 196.870 13.030 197.260 ;
        RECT 13.830 197.110 15.690 197.400 ;
        RECT 13.830 197.100 14.140 197.110 ;
        RECT 15.380 197.100 15.690 197.110 ;
        RECT 3.970 196.750 4.620 196.760 ;
        RECT 3.970 196.420 4.270 196.750 ;
        RECT 3.250 195.970 4.270 196.420 ;
        RECT 8.860 196.260 9.150 196.860 ;
        RECT 10.750 196.260 11.040 196.860 ;
        RECT 3.970 195.960 4.270 195.970 ;
        RECT 13.090 195.650 13.390 196.650 ;
        RECT 13.840 196.050 14.140 197.100 ;
        RECT 16.440 196.000 16.690 197.740 ;
        RECT 73.890 197.670 74.680 197.860 ;
        RECT 73.890 197.470 74.140 197.670 ;
        RECT 74.390 197.560 74.680 197.670 ;
        RECT 75.780 197.470 76.030 198.010 ;
        RECT 78.860 198.010 79.130 198.070 ;
        RECT 80.410 198.350 81.720 198.610 ;
        RECT 83.860 198.390 99.520 198.640 ;
        RECT 83.860 198.360 84.680 198.390 ;
        RECT 80.410 198.010 80.720 198.350 ;
        RECT 76.420 197.480 78.060 197.870 ;
        RECT 78.860 197.720 80.720 198.010 ;
        RECT 78.860 197.710 79.170 197.720 ;
        RECT 80.410 197.710 80.720 197.720 ;
        RECT 17.140 195.650 17.400 197.200 ;
        RECT 73.890 196.870 74.180 197.470 ;
        RECT 75.780 196.870 76.070 197.470 ;
        RECT 78.120 196.260 78.420 197.260 ;
        RECT 78.870 196.660 79.170 197.710 ;
        RECT 81.470 196.610 81.720 198.350 ;
        RECT 99.270 198.180 99.520 198.390 ;
        RECT 82.170 196.260 82.430 197.810 ;
        RECT 99.270 196.340 99.540 198.180 ;
        RECT 83.130 196.260 83.310 196.270 ;
        RECT 78.070 195.960 83.320 196.260 ;
        RECT 13.040 195.640 18.290 195.650 ;
        RECT 2.920 195.560 3.170 195.570 ;
        RECT 2.920 195.100 3.900 195.560 ;
        RECT 13.040 195.350 18.310 195.640 ;
        RECT 2.920 194.800 3.170 195.100 ;
        RECT 10.890 195.010 12.730 195.020 ;
        RECT 18.140 195.010 18.310 195.350 ;
        RECT 4.630 195.000 4.870 195.010 ;
        RECT 5.710 195.000 18.310 195.010 ;
        RECT 4.630 194.840 18.310 195.000 ;
        RECT 4.630 194.830 16.140 194.840 ;
        RECT 4.620 194.820 10.940 194.830 ;
        RECT 12.490 194.820 16.140 194.830 ;
        RECT 4.620 194.810 6.490 194.820 ;
        RECT 4.620 194.800 4.870 194.810 ;
        RECT 2.920 194.630 4.870 194.800 ;
        RECT 2.920 194.330 3.190 194.630 ;
        RECT 2.930 194.070 3.190 194.330 ;
        RECT 2.910 193.680 3.210 194.070 ;
        RECT 2.900 193.280 3.210 193.680 ;
        RECT 2.890 192.520 3.200 193.280 ;
        RECT 2.790 192.500 3.200 192.520 ;
        RECT 2.760 191.550 3.210 192.500 ;
        RECT 3.620 191.260 4.080 192.200 ;
        RECT 4.820 191.610 14.090 191.620 ;
        RECT 15.970 191.610 17.890 191.620 ;
        RECT 4.820 191.420 17.890 191.610 ;
        RECT 4.820 191.410 17.180 191.420 ;
        RECT 3.660 190.940 3.960 191.260 ;
        RECT 3.660 190.610 3.950 190.940 ;
        RECT 3.670 189.810 3.930 190.610 ;
        RECT 4.820 190.400 5.030 191.410 ;
        RECT 14.080 191.400 15.980 191.410 ;
        RECT 17.710 190.670 17.890 191.420 ;
        RECT 3.670 189.210 3.920 189.810 ;
        RECT 4.820 189.390 5.020 190.400 ;
        RECT 12.630 190.370 17.890 190.670 ;
        RECT 2.880 188.760 3.920 189.210 ;
        RECT 2.860 187.310 3.820 187.760 ;
        RECT 3.570 187.260 3.820 187.310 ;
        RECT 4.830 187.260 5.020 189.390 ;
        RECT 3.570 187.060 5.020 187.260 ;
        RECT 8.550 188.730 8.810 189.930 ;
        RECT 8.550 188.220 8.800 188.730 ;
        RECT 10.440 188.720 10.700 189.930 ;
        RECT 12.830 188.820 13.080 190.370 ;
        RECT 10.440 188.560 10.830 188.720 ;
        RECT 10.430 188.430 10.830 188.560 ;
        RECT 13.530 188.430 13.790 190.040 ;
        RECT 16.080 188.970 16.380 190.020 ;
        RECT 16.830 189.420 17.130 190.370 ;
        RECT 17.330 189.470 17.630 189.520 ;
        RECT 17.330 189.120 18.230 189.470 ;
        RECT 19.940 189.340 20.160 189.350 ;
        RECT 19.940 189.150 33.620 189.340 ;
        RECT 19.940 189.020 20.160 189.150 ;
        RECT 9.050 188.220 9.340 188.380 ;
        RECT 10.430 188.370 10.690 188.430 ;
        RECT 8.550 188.030 9.340 188.220 ;
        RECT 8.550 187.830 8.800 188.030 ;
        RECT 9.050 187.920 9.340 188.030 ;
        RECT 10.440 187.830 10.690 188.370 ;
        RECT 13.520 188.370 13.790 188.430 ;
        RECT 15.070 188.710 16.380 188.970 ;
        RECT 18.480 188.720 20.160 189.020 ;
        RECT 18.480 188.710 20.140 188.720 ;
        RECT 15.070 188.370 15.380 188.710 ;
        RECT 11.080 187.840 12.720 188.230 ;
        RECT 13.520 188.080 15.380 188.370 ;
        RECT 13.520 188.070 13.830 188.080 ;
        RECT 15.070 188.070 15.380 188.080 ;
        RECT 8.550 187.230 8.840 187.830 ;
        RECT 10.440 187.230 10.730 187.830 ;
        RECT 3.570 186.970 3.820 187.060 ;
        RECT 2.840 186.520 3.820 186.970 ;
        RECT 12.780 186.620 13.080 187.620 ;
        RECT 13.530 187.020 13.830 188.070 ;
        RECT 16.130 186.970 16.380 188.710 ;
        RECT 33.370 188.250 33.620 189.150 ;
        RECT 16.830 186.620 17.090 188.170 ;
        RECT 28.310 187.950 33.620 188.250 ;
        RECT 12.730 186.600 17.980 186.620 ;
        RECT 12.730 186.320 18.100 186.600 ;
        RECT 6.180 185.920 6.460 185.990 ;
        RECT 7.360 185.950 7.640 185.980 ;
        RECT 17.810 185.950 18.100 186.320 ;
        RECT 7.360 185.940 18.100 185.950 ;
        RECT 4.770 185.720 6.460 185.920 ;
        RECT 3.560 185.520 3.840 185.530 ;
        RECT 2.820 185.070 3.840 185.520 ;
        RECT 4.770 185.070 5.000 185.720 ;
        RECT 6.180 185.660 6.460 185.720 ;
        RECT 7.340 185.710 18.100 185.940 ;
        RECT 7.360 185.700 18.100 185.710 ;
        RECT 24.230 186.310 24.490 187.510 ;
        RECT 24.230 185.800 24.480 186.310 ;
        RECT 26.120 186.300 26.380 187.510 ;
        RECT 28.510 186.400 28.760 187.950 ;
        RECT 26.120 186.140 26.510 186.300 ;
        RECT 26.110 186.010 26.510 186.140 ;
        RECT 29.210 186.010 29.470 187.620 ;
        RECT 31.760 186.550 32.060 187.600 ;
        RECT 32.510 187.000 32.810 187.950 ;
        RECT 33.010 187.050 33.310 187.100 ;
        RECT 33.010 186.700 33.910 187.050 ;
        RECT 46.670 186.650 51.140 186.680 ;
        RECT 35.730 186.620 51.140 186.650 ;
        RECT 35.060 186.600 51.140 186.620 ;
        RECT 24.730 185.800 25.020 185.960 ;
        RECT 26.110 185.950 26.370 186.010 ;
        RECT 7.360 185.690 18.060 185.700 ;
        RECT 7.360 185.650 7.640 185.690 ;
        RECT 24.230 185.610 25.020 185.800 ;
        RECT 24.230 185.410 24.480 185.610 ;
        RECT 24.730 185.500 25.020 185.610 ;
        RECT 26.120 185.410 26.370 185.950 ;
        RECT 29.200 185.950 29.470 186.010 ;
        RECT 30.750 186.290 32.060 186.550 ;
        RECT 30.750 185.950 31.060 186.290 ;
        RECT 26.760 185.420 28.400 185.810 ;
        RECT 29.200 185.660 31.060 185.950 ;
        RECT 29.200 185.650 29.510 185.660 ;
        RECT 30.750 185.650 31.060 185.660 ;
        RECT 6.160 185.090 6.430 185.170 ;
        RECT 3.560 184.860 5.000 185.070 ;
        RECT 5.550 184.870 6.430 185.090 ;
        RECT 3.560 183.810 3.840 184.860 ;
        RECT 5.550 184.060 5.770 184.870 ;
        RECT 6.160 184.840 6.430 184.870 ;
        RECT 7.290 185.130 7.580 185.180 ;
        RECT 7.290 184.950 18.040 185.130 ;
        RECT 7.290 184.850 7.580 184.950 ;
        RECT 12.130 184.940 15.760 184.950 ;
        RECT 17.840 184.270 18.040 184.950 ;
        RECT 24.230 184.810 24.520 185.410 ;
        RECT 26.120 184.810 26.410 185.410 ;
        RECT 2.840 183.360 3.840 183.810 ;
        RECT 2.820 181.910 4.120 182.360 ;
        RECT 3.820 181.510 4.120 181.910 ;
        RECT 5.540 181.530 5.770 184.060 ;
        RECT 12.790 183.970 18.040 184.270 ;
        RECT 28.460 184.200 28.760 185.200 ;
        RECT 29.210 184.600 29.510 185.650 ;
        RECT 31.810 184.550 32.060 186.290 ;
        RECT 34.180 186.280 51.140 186.600 ;
        RECT 83.130 186.300 83.310 195.960 ;
        RECT 35.060 186.270 51.140 186.280 ;
        RECT 35.060 186.240 47.040 186.270 ;
        RECT 35.060 186.230 35.950 186.240 ;
        RECT 32.510 184.200 32.770 185.750 ;
        RECT 33.600 184.200 33.800 184.210 ;
        RECT 4.610 181.510 5.770 181.530 ;
        RECT 3.820 181.330 5.770 181.510 ;
        RECT 8.710 182.330 8.970 183.530 ;
        RECT 8.710 181.820 8.960 182.330 ;
        RECT 10.600 182.320 10.860 183.530 ;
        RECT 12.990 182.420 13.240 183.970 ;
        RECT 10.600 182.160 10.990 182.320 ;
        RECT 10.590 182.030 10.990 182.160 ;
        RECT 13.690 182.030 13.950 183.640 ;
        RECT 16.240 182.570 16.540 183.620 ;
        RECT 16.990 183.020 17.290 183.970 ;
        RECT 17.840 183.960 18.040 183.970 ;
        RECT 28.410 183.900 33.800 184.200 ;
        RECT 17.490 183.070 17.790 183.120 ;
        RECT 17.490 182.720 18.390 183.070 ;
        RECT 33.600 182.660 33.800 183.900 ;
        RECT 50.760 182.700 51.120 186.270 ;
        RECT 26.040 182.640 27.230 182.650 ;
        RECT 28.220 182.640 29.410 182.650 ;
        RECT 30.440 182.640 31.630 182.650 ;
        RECT 32.620 182.640 33.810 182.660 ;
        RECT 23.830 182.630 33.810 182.640 ;
        RECT 20.440 182.610 21.630 182.620 ;
        RECT 22.720 182.610 33.810 182.630 ;
        RECT 9.210 181.820 9.500 181.980 ;
        RECT 10.590 181.970 10.850 182.030 ;
        RECT 8.710 181.630 9.500 181.820 ;
        RECT 8.710 181.430 8.960 181.630 ;
        RECT 9.210 181.520 9.500 181.630 ;
        RECT 10.600 181.430 10.850 181.970 ;
        RECT 13.680 181.970 13.950 182.030 ;
        RECT 15.230 182.310 16.540 182.570 ;
        RECT 18.600 182.380 33.810 182.610 ;
        RECT 45.890 182.400 51.140 182.700 ;
        RECT 18.600 182.370 32.760 182.380 ;
        RECT 18.600 182.360 26.130 182.370 ;
        RECT 27.140 182.360 28.330 182.370 ;
        RECT 29.290 182.360 30.480 182.370 ;
        RECT 31.570 182.360 32.760 182.370 ;
        RECT 18.600 182.350 23.910 182.360 ;
        RECT 18.600 182.340 22.770 182.350 ;
        RECT 18.600 182.330 20.490 182.340 ;
        RECT 21.580 182.330 22.770 182.340 ;
        RECT 18.600 182.320 19.320 182.330 ;
        RECT 15.230 181.970 15.540 182.310 ;
        RECT 11.240 181.440 12.880 181.830 ;
        RECT 13.680 181.680 15.540 181.970 ;
        RECT 13.680 181.670 13.990 181.680 ;
        RECT 15.230 181.670 15.540 181.680 ;
        RECT 3.820 181.320 4.470 181.330 ;
        RECT 3.820 180.990 4.120 181.320 ;
        RECT 3.100 180.540 4.120 180.990 ;
        RECT 8.710 180.830 9.000 181.430 ;
        RECT 10.600 180.830 10.890 181.430 ;
        RECT 3.820 180.530 4.120 180.540 ;
        RECT 12.940 180.220 13.240 181.220 ;
        RECT 13.690 180.620 13.990 181.670 ;
        RECT 16.290 180.570 16.540 182.310 ;
        RECT 16.990 180.220 17.250 181.770 ;
        RECT 41.810 180.760 42.070 181.960 ;
        RECT 41.810 180.250 42.060 180.760 ;
        RECT 43.700 180.750 43.960 181.960 ;
        RECT 46.090 180.850 46.340 182.400 ;
        RECT 43.700 180.590 44.090 180.750 ;
        RECT 43.690 180.460 44.090 180.590 ;
        RECT 46.790 180.460 47.050 182.070 ;
        RECT 49.340 181.000 49.640 182.050 ;
        RECT 50.090 181.450 50.390 182.400 ;
        RECT 50.590 181.500 50.890 181.550 ;
        RECT 50.590 181.150 51.490 181.500 ;
        RECT 42.310 180.250 42.600 180.410 ;
        RECT 43.690 180.400 43.950 180.460 ;
        RECT 12.890 180.210 18.140 180.220 ;
        RECT 2.770 180.130 3.020 180.140 ;
        RECT 2.770 179.670 3.750 180.130 ;
        RECT 12.890 179.920 18.160 180.210 ;
        RECT 2.770 179.370 3.020 179.670 ;
        RECT 10.740 179.580 12.580 179.590 ;
        RECT 17.990 179.580 18.160 179.920 ;
        RECT 4.480 179.570 4.720 179.580 ;
        RECT 5.560 179.570 18.160 179.580 ;
        RECT 4.480 179.410 18.160 179.570 ;
        RECT 41.810 180.060 42.600 180.250 ;
        RECT 41.810 179.860 42.060 180.060 ;
        RECT 42.310 179.950 42.600 180.060 ;
        RECT 43.700 179.860 43.950 180.400 ;
        RECT 46.780 180.400 47.050 180.460 ;
        RECT 48.330 180.740 49.640 181.000 ;
        RECT 51.700 181.040 53.370 181.070 ;
        RECT 68.450 181.040 68.700 181.050 ;
        RECT 51.700 180.770 68.700 181.040 ;
        RECT 51.700 180.760 65.200 180.770 ;
        RECT 52.980 180.740 65.200 180.760 ;
        RECT 48.330 180.400 48.640 180.740 ;
        RECT 44.340 179.870 45.980 180.260 ;
        RECT 46.780 180.110 48.640 180.400 ;
        RECT 46.780 180.100 47.090 180.110 ;
        RECT 48.330 180.100 48.640 180.110 ;
        RECT 4.480 179.400 15.990 179.410 ;
        RECT 4.470 179.390 10.790 179.400 ;
        RECT 12.340 179.390 15.990 179.400 ;
        RECT 4.470 179.380 6.340 179.390 ;
        RECT 4.470 179.370 4.720 179.380 ;
        RECT 2.770 179.200 4.720 179.370 ;
        RECT 41.810 179.260 42.100 179.860 ;
        RECT 43.700 179.260 43.990 179.860 ;
        RECT 2.770 178.980 3.020 179.200 ;
        RECT 2.770 178.810 3.810 178.980 ;
        RECT 3.620 177.950 3.810 178.810 ;
        RECT 46.040 178.650 46.340 179.650 ;
        RECT 46.790 179.050 47.090 180.100 ;
        RECT 49.390 179.000 49.640 180.740 ;
        RECT 50.090 178.650 50.350 180.200 ;
        RECT 50.970 178.650 51.310 178.720 ;
        RECT 45.990 178.350 51.310 178.650 ;
        RECT 2.830 177.510 3.810 177.950 ;
        RECT 2.830 177.500 3.780 177.510 ;
        RECT 4.650 177.190 13.920 177.200 ;
        RECT 15.800 177.190 17.720 177.200 ;
        RECT 2.500 177.090 2.690 177.100 ;
        RECT 2.500 176.630 3.480 177.090 ;
        RECT 4.650 177.000 17.720 177.190 ;
        RECT 4.650 176.990 17.010 177.000 ;
        RECT 2.500 175.840 2.690 176.630 ;
        RECT 4.650 175.980 4.860 176.990 ;
        RECT 13.910 176.980 15.810 176.990 ;
        RECT 17.540 176.250 17.720 177.000 ;
        RECT 3.500 175.840 3.770 175.850 ;
        RECT 2.500 175.630 3.770 175.840 ;
        RECT 3.500 175.420 3.770 175.630 ;
        RECT 3.500 174.790 3.750 175.420 ;
        RECT 4.650 174.970 4.850 175.980 ;
        RECT 12.460 175.950 17.720 176.250 ;
        RECT 2.710 174.340 3.750 174.790 ;
        RECT 2.690 172.890 3.650 173.340 ;
        RECT 3.400 172.840 3.650 172.890 ;
        RECT 4.660 172.840 4.850 174.970 ;
        RECT 3.400 172.640 4.850 172.840 ;
        RECT 8.380 174.310 8.640 175.510 ;
        RECT 8.380 173.800 8.630 174.310 ;
        RECT 10.270 174.300 10.530 175.510 ;
        RECT 12.660 174.400 12.910 175.950 ;
        RECT 10.270 174.140 10.660 174.300 ;
        RECT 10.260 174.010 10.660 174.140 ;
        RECT 13.360 174.010 13.620 175.620 ;
        RECT 15.910 174.550 16.210 175.600 ;
        RECT 16.660 175.000 16.960 175.950 ;
        RECT 17.160 175.050 17.460 175.100 ;
        RECT 17.160 174.700 18.060 175.050 ;
        RECT 19.770 174.920 19.990 174.930 ;
        RECT 19.770 174.730 33.450 174.920 ;
        RECT 19.770 174.600 19.990 174.730 ;
        RECT 8.880 173.800 9.170 173.960 ;
        RECT 10.260 173.950 10.520 174.010 ;
        RECT 8.380 173.610 9.170 173.800 ;
        RECT 8.380 173.410 8.630 173.610 ;
        RECT 8.880 173.500 9.170 173.610 ;
        RECT 10.270 173.410 10.520 173.950 ;
        RECT 13.350 173.950 13.620 174.010 ;
        RECT 14.900 174.290 16.210 174.550 ;
        RECT 18.310 174.300 19.990 174.600 ;
        RECT 18.310 174.290 19.970 174.300 ;
        RECT 14.900 173.950 15.210 174.290 ;
        RECT 10.910 173.420 12.550 173.810 ;
        RECT 13.350 173.660 15.210 173.950 ;
        RECT 13.350 173.650 13.660 173.660 ;
        RECT 14.900 173.650 15.210 173.660 ;
        RECT 8.380 172.810 8.670 173.410 ;
        RECT 10.270 172.810 10.560 173.410 ;
        RECT 3.400 172.550 3.650 172.640 ;
        RECT 2.670 172.100 3.650 172.550 ;
        RECT 12.610 172.200 12.910 173.200 ;
        RECT 13.360 172.600 13.660 173.650 ;
        RECT 15.960 172.550 16.210 174.290 ;
        RECT 33.200 173.830 33.450 174.730 ;
        RECT 16.660 172.200 16.920 173.750 ;
        RECT 28.140 173.530 33.450 173.830 ;
        RECT 12.560 172.180 17.810 172.200 ;
        RECT 12.560 171.900 17.930 172.180 ;
        RECT 6.010 171.500 6.290 171.570 ;
        RECT 7.190 171.530 7.470 171.560 ;
        RECT 17.640 171.530 17.930 171.900 ;
        RECT 7.190 171.520 17.930 171.530 ;
        RECT 4.600 171.300 6.290 171.500 ;
        RECT 3.390 171.100 3.670 171.110 ;
        RECT 2.650 170.650 3.670 171.100 ;
        RECT 4.600 170.650 4.830 171.300 ;
        RECT 6.010 171.240 6.290 171.300 ;
        RECT 7.170 171.290 17.930 171.520 ;
        RECT 7.190 171.280 17.930 171.290 ;
        RECT 24.060 171.890 24.320 173.090 ;
        RECT 24.060 171.380 24.310 171.890 ;
        RECT 25.950 171.880 26.210 173.090 ;
        RECT 28.340 171.980 28.590 173.530 ;
        RECT 25.950 171.720 26.340 171.880 ;
        RECT 25.940 171.590 26.340 171.720 ;
        RECT 29.040 171.590 29.300 173.200 ;
        RECT 31.590 172.130 31.890 173.180 ;
        RECT 32.340 172.580 32.640 173.530 ;
        RECT 32.840 172.630 33.140 172.680 ;
        RECT 32.840 172.280 33.740 172.630 ;
        RECT 50.970 172.230 51.310 178.350 ;
        RECT 50.400 172.210 51.360 172.230 ;
        RECT 34.880 172.190 39.160 172.200 ;
        RECT 46.560 172.190 51.360 172.210 ;
        RECT 34.880 172.180 51.360 172.190 ;
        RECT 24.560 171.380 24.850 171.540 ;
        RECT 25.940 171.530 26.200 171.590 ;
        RECT 7.190 171.270 17.890 171.280 ;
        RECT 7.190 171.230 7.470 171.270 ;
        RECT 24.060 171.190 24.850 171.380 ;
        RECT 24.060 170.990 24.310 171.190 ;
        RECT 24.560 171.080 24.850 171.190 ;
        RECT 25.950 170.990 26.200 171.530 ;
        RECT 29.030 171.530 29.300 171.590 ;
        RECT 30.580 171.870 31.890 172.130 ;
        RECT 30.580 171.530 30.890 171.870 ;
        RECT 26.590 171.000 28.230 171.390 ;
        RECT 29.030 171.240 30.890 171.530 ;
        RECT 29.030 171.230 29.340 171.240 ;
        RECT 30.580 171.230 30.890 171.240 ;
        RECT 5.990 170.670 6.260 170.750 ;
        RECT 3.390 170.440 4.830 170.650 ;
        RECT 5.380 170.450 6.260 170.670 ;
        RECT 3.390 169.390 3.670 170.440 ;
        RECT 5.380 169.640 5.600 170.450 ;
        RECT 5.990 170.420 6.260 170.450 ;
        RECT 7.120 170.710 7.410 170.760 ;
        RECT 7.120 170.530 17.870 170.710 ;
        RECT 7.120 170.430 7.410 170.530 ;
        RECT 11.960 170.520 15.590 170.530 ;
        RECT 17.670 169.850 17.870 170.530 ;
        RECT 24.060 170.390 24.350 170.990 ;
        RECT 25.950 170.390 26.240 170.990 ;
        RECT 2.670 168.940 3.670 169.390 ;
        RECT 2.650 167.490 3.950 167.940 ;
        RECT 3.650 167.090 3.950 167.490 ;
        RECT 5.370 167.110 5.600 169.640 ;
        RECT 12.620 169.550 17.870 169.850 ;
        RECT 28.290 169.780 28.590 170.780 ;
        RECT 29.040 170.180 29.340 171.230 ;
        RECT 31.640 170.130 31.890 171.870 ;
        RECT 34.010 171.870 51.360 172.180 ;
        RECT 34.010 171.860 47.020 171.870 ;
        RECT 38.870 171.850 47.020 171.860 ;
        RECT 50.400 171.830 51.360 171.870 ;
        RECT 50.970 171.820 51.310 171.830 ;
        RECT 32.340 169.780 32.600 171.330 ;
        RECT 33.430 169.780 33.630 169.790 ;
        RECT 4.440 167.090 5.600 167.110 ;
        RECT 3.650 166.910 5.600 167.090 ;
        RECT 8.540 167.910 8.800 169.110 ;
        RECT 8.540 167.400 8.790 167.910 ;
        RECT 10.430 167.900 10.690 169.110 ;
        RECT 12.820 168.000 13.070 169.550 ;
        RECT 10.430 167.740 10.820 167.900 ;
        RECT 10.420 167.610 10.820 167.740 ;
        RECT 13.520 167.610 13.780 169.220 ;
        RECT 16.070 168.150 16.370 169.200 ;
        RECT 16.820 168.600 17.120 169.550 ;
        RECT 17.670 169.540 17.870 169.550 ;
        RECT 28.240 169.480 33.630 169.780 ;
        RECT 17.320 168.650 17.620 168.700 ;
        RECT 17.320 168.300 18.220 168.650 ;
        RECT 33.430 168.240 33.630 169.480 ;
        RECT 25.870 168.220 27.060 168.230 ;
        RECT 28.050 168.220 29.240 168.230 ;
        RECT 30.270 168.220 31.460 168.230 ;
        RECT 32.450 168.220 33.640 168.240 ;
        RECT 23.660 168.210 33.640 168.220 ;
        RECT 20.270 168.190 21.460 168.200 ;
        RECT 22.550 168.190 33.640 168.210 ;
        RECT 9.040 167.400 9.330 167.560 ;
        RECT 10.420 167.550 10.680 167.610 ;
        RECT 8.540 167.210 9.330 167.400 ;
        RECT 8.540 167.010 8.790 167.210 ;
        RECT 9.040 167.100 9.330 167.210 ;
        RECT 10.430 167.010 10.680 167.550 ;
        RECT 13.510 167.550 13.780 167.610 ;
        RECT 15.060 167.890 16.370 168.150 ;
        RECT 18.430 167.960 33.640 168.190 ;
        RECT 18.430 167.950 32.590 167.960 ;
        RECT 18.430 167.940 25.960 167.950 ;
        RECT 26.970 167.940 28.160 167.950 ;
        RECT 29.120 167.940 30.310 167.950 ;
        RECT 31.400 167.940 32.590 167.950 ;
        RECT 18.430 167.930 23.740 167.940 ;
        RECT 18.430 167.920 22.600 167.930 ;
        RECT 18.430 167.910 20.320 167.920 ;
        RECT 21.410 167.910 22.600 167.920 ;
        RECT 18.430 167.900 19.150 167.910 ;
        RECT 15.060 167.550 15.370 167.890 ;
        RECT 11.070 167.020 12.710 167.410 ;
        RECT 13.510 167.260 15.370 167.550 ;
        RECT 13.510 167.250 13.820 167.260 ;
        RECT 15.060 167.250 15.370 167.260 ;
        RECT 3.650 166.900 4.300 166.910 ;
        RECT 3.650 166.570 3.950 166.900 ;
        RECT 2.930 166.120 3.950 166.570 ;
        RECT 8.540 166.410 8.830 167.010 ;
        RECT 10.430 166.410 10.720 167.010 ;
        RECT 3.650 166.110 3.950 166.120 ;
        RECT 12.770 165.800 13.070 166.800 ;
        RECT 13.520 166.200 13.820 167.250 ;
        RECT 16.120 166.150 16.370 167.890 ;
        RECT 68.450 167.630 68.710 180.770 ;
        RECT 68.440 167.510 68.710 167.630 ;
        RECT 83.040 176.780 83.310 186.300 ;
        RECT 99.270 192.670 99.580 196.340 ;
        RECT 99.270 190.890 99.600 192.670 ;
        RECT 99.270 188.920 99.560 190.890 ;
        RECT 99.270 187.090 99.580 188.920 ;
        RECT 99.270 183.270 99.560 187.090 ;
        RECT 99.270 181.300 99.540 183.270 ;
        RECT 99.270 179.580 99.600 181.300 ;
        RECT 99.270 177.660 99.560 179.580 ;
        RECT 16.820 165.800 17.080 167.350 ;
        RECT 68.440 166.680 68.700 167.510 ;
        RECT 83.040 166.830 83.220 176.780 ;
        RECT 99.270 168.120 99.540 177.660 ;
        RECT 63.420 166.380 68.700 166.680 ;
        RECT 12.720 165.790 17.970 165.800 ;
        RECT 2.600 165.710 2.850 165.720 ;
        RECT 2.600 165.250 3.580 165.710 ;
        RECT 12.720 165.500 17.990 165.790 ;
        RECT 2.600 164.950 2.850 165.250 ;
        RECT 10.570 165.160 12.410 165.170 ;
        RECT 17.820 165.160 17.990 165.500 ;
        RECT 4.310 165.150 4.550 165.160 ;
        RECT 5.390 165.150 17.990 165.160 ;
        RECT 4.310 164.990 17.990 165.150 ;
        RECT 4.310 164.980 15.820 164.990 ;
        RECT 4.300 164.970 10.620 164.980 ;
        RECT 12.170 164.970 15.820 164.980 ;
        RECT 4.300 164.960 6.170 164.970 ;
        RECT 4.300 164.950 4.550 164.960 ;
        RECT 2.600 164.780 4.550 164.950 ;
        RECT 2.600 164.480 2.870 164.780 ;
        RECT 2.610 164.220 2.870 164.480 ;
        RECT 59.340 164.740 59.600 165.940 ;
        RECT 59.340 164.230 59.590 164.740 ;
        RECT 61.230 164.730 61.490 165.940 ;
        RECT 63.620 164.830 63.870 166.380 ;
        RECT 61.230 164.570 61.620 164.730 ;
        RECT 61.220 164.440 61.620 164.570 ;
        RECT 64.320 164.440 64.580 166.050 ;
        RECT 66.870 164.980 67.170 166.030 ;
        RECT 67.620 165.430 67.920 166.380 ;
        RECT 68.120 165.480 68.420 165.530 ;
        RECT 68.120 165.130 69.020 165.480 ;
        RECT 83.030 165.020 83.230 166.830 ;
        RECT 59.840 164.230 60.130 164.390 ;
        RECT 61.220 164.380 61.480 164.440 ;
        RECT 2.590 163.830 2.890 164.220 ;
        RECT 59.340 164.040 60.130 164.230 ;
        RECT 59.340 163.840 59.590 164.040 ;
        RECT 59.840 163.930 60.130 164.040 ;
        RECT 61.230 163.840 61.480 164.380 ;
        RECT 64.310 164.380 64.580 164.440 ;
        RECT 65.860 164.720 67.170 164.980 ;
        RECT 69.290 164.730 83.230 165.020 ;
        RECT 99.310 166.250 99.580 168.120 ;
        RECT 69.290 164.720 83.190 164.730 ;
        RECT 65.860 164.380 66.170 164.720 ;
        RECT 61.870 163.850 63.510 164.240 ;
        RECT 64.310 164.090 66.170 164.380 ;
        RECT 64.310 164.080 64.620 164.090 ;
        RECT 65.860 164.080 66.170 164.090 ;
        RECT 2.590 163.600 4.080 163.830 ;
        RECT 3.830 162.670 4.080 163.600 ;
        RECT 59.340 163.240 59.630 163.840 ;
        RECT 61.230 163.240 61.520 163.840 ;
        RECT 3.030 162.210 4.080 162.670 ;
        RECT 63.570 162.630 63.870 163.630 ;
        RECT 64.320 163.030 64.620 164.080 ;
        RECT 66.920 162.980 67.170 164.720 ;
        RECT 69.880 164.710 83.190 164.720 ;
        RECT 67.620 162.630 67.880 164.180 ;
        RECT 63.520 162.330 68.790 162.630 ;
        RECT 3.830 162.200 4.080 162.210 ;
        RECT 2.700 161.800 2.950 161.810 ;
        RECT 2.700 161.350 3.680 161.800 ;
        RECT 4.790 161.540 14.060 161.550 ;
        RECT 15.940 161.540 17.860 161.550 ;
        RECT 4.790 161.350 17.860 161.540 ;
        RECT 2.700 160.740 2.950 161.350 ;
        RECT 4.790 161.340 17.150 161.350 ;
        RECT 2.700 160.490 3.910 160.740 ;
        RECT 3.640 159.740 3.900 160.490 ;
        RECT 4.790 160.330 5.000 161.340 ;
        RECT 14.050 161.330 15.950 161.340 ;
        RECT 17.680 160.600 17.860 161.350 ;
        RECT 3.640 159.140 3.890 159.740 ;
        RECT 4.790 159.320 4.990 160.330 ;
        RECT 12.600 160.300 17.860 160.600 ;
        RECT 2.850 158.690 3.890 159.140 ;
        RECT 2.830 157.240 3.790 157.690 ;
        RECT 3.540 157.190 3.790 157.240 ;
        RECT 4.800 157.190 4.990 159.320 ;
        RECT 3.540 156.990 4.990 157.190 ;
        RECT 8.520 158.660 8.780 159.860 ;
        RECT 8.520 158.150 8.770 158.660 ;
        RECT 10.410 158.650 10.670 159.860 ;
        RECT 12.800 158.750 13.050 160.300 ;
        RECT 10.410 158.490 10.800 158.650 ;
        RECT 10.400 158.360 10.800 158.490 ;
        RECT 13.500 158.360 13.760 159.970 ;
        RECT 16.050 158.900 16.350 159.950 ;
        RECT 16.800 159.350 17.100 160.300 ;
        RECT 17.300 159.400 17.600 159.450 ;
        RECT 17.300 159.050 18.200 159.400 ;
        RECT 19.910 159.270 20.130 159.280 ;
        RECT 19.910 159.080 33.590 159.270 ;
        RECT 19.910 158.950 20.130 159.080 ;
        RECT 9.020 158.150 9.310 158.310 ;
        RECT 10.400 158.300 10.660 158.360 ;
        RECT 8.520 157.960 9.310 158.150 ;
        RECT 8.520 157.760 8.770 157.960 ;
        RECT 9.020 157.850 9.310 157.960 ;
        RECT 10.410 157.760 10.660 158.300 ;
        RECT 13.490 158.300 13.760 158.360 ;
        RECT 15.040 158.640 16.350 158.900 ;
        RECT 18.450 158.650 20.130 158.950 ;
        RECT 18.450 158.640 20.110 158.650 ;
        RECT 15.040 158.300 15.350 158.640 ;
        RECT 11.050 157.770 12.690 158.160 ;
        RECT 13.490 158.010 15.350 158.300 ;
        RECT 13.490 158.000 13.800 158.010 ;
        RECT 15.040 158.000 15.350 158.010 ;
        RECT 8.520 157.160 8.810 157.760 ;
        RECT 10.410 157.160 10.700 157.760 ;
        RECT 3.540 156.900 3.790 156.990 ;
        RECT 2.810 156.450 3.790 156.900 ;
        RECT 12.750 156.550 13.050 157.550 ;
        RECT 13.500 156.950 13.800 158.000 ;
        RECT 16.100 156.900 16.350 158.640 ;
        RECT 33.340 158.180 33.590 159.080 ;
        RECT 16.800 156.550 17.060 158.100 ;
        RECT 28.280 157.880 33.590 158.180 ;
        RECT 12.700 156.530 17.950 156.550 ;
        RECT 12.700 156.250 18.070 156.530 ;
        RECT 6.150 155.850 6.430 155.920 ;
        RECT 7.330 155.880 7.610 155.910 ;
        RECT 17.780 155.880 18.070 156.250 ;
        RECT 7.330 155.870 18.070 155.880 ;
        RECT 4.740 155.650 6.430 155.850 ;
        RECT 3.530 155.450 3.810 155.460 ;
        RECT 2.790 155.000 3.810 155.450 ;
        RECT 4.740 155.000 4.970 155.650 ;
        RECT 6.150 155.590 6.430 155.650 ;
        RECT 7.310 155.640 18.070 155.870 ;
        RECT 7.330 155.630 18.070 155.640 ;
        RECT 24.200 156.240 24.460 157.440 ;
        RECT 24.200 155.730 24.450 156.240 ;
        RECT 26.090 156.230 26.350 157.440 ;
        RECT 28.480 156.330 28.730 157.880 ;
        RECT 26.090 156.070 26.480 156.230 ;
        RECT 26.080 155.940 26.480 156.070 ;
        RECT 29.180 155.940 29.440 157.550 ;
        RECT 31.730 156.480 32.030 157.530 ;
        RECT 32.480 156.930 32.780 157.880 ;
        RECT 32.980 156.980 33.280 157.030 ;
        RECT 32.980 156.630 33.880 156.980 ;
        RECT 46.640 156.580 51.110 156.610 ;
        RECT 35.700 156.550 51.110 156.580 ;
        RECT 35.030 156.530 51.110 156.550 ;
        RECT 24.700 155.730 24.990 155.890 ;
        RECT 26.080 155.880 26.340 155.940 ;
        RECT 7.330 155.620 18.030 155.630 ;
        RECT 7.330 155.580 7.610 155.620 ;
        RECT 24.200 155.540 24.990 155.730 ;
        RECT 24.200 155.340 24.450 155.540 ;
        RECT 24.700 155.430 24.990 155.540 ;
        RECT 26.090 155.340 26.340 155.880 ;
        RECT 29.170 155.880 29.440 155.940 ;
        RECT 30.720 156.220 32.030 156.480 ;
        RECT 30.720 155.880 31.030 156.220 ;
        RECT 26.730 155.350 28.370 155.740 ;
        RECT 29.170 155.590 31.030 155.880 ;
        RECT 29.170 155.580 29.480 155.590 ;
        RECT 30.720 155.580 31.030 155.590 ;
        RECT 6.130 155.020 6.400 155.100 ;
        RECT 3.530 154.790 4.970 155.000 ;
        RECT 5.520 154.800 6.400 155.020 ;
        RECT 3.530 153.740 3.810 154.790 ;
        RECT 5.520 153.990 5.740 154.800 ;
        RECT 6.130 154.770 6.400 154.800 ;
        RECT 7.260 155.060 7.550 155.110 ;
        RECT 7.260 154.880 18.010 155.060 ;
        RECT 7.260 154.780 7.550 154.880 ;
        RECT 12.100 154.870 15.730 154.880 ;
        RECT 17.810 154.200 18.010 154.880 ;
        RECT 24.200 154.740 24.490 155.340 ;
        RECT 26.090 154.740 26.380 155.340 ;
        RECT 2.810 153.290 3.810 153.740 ;
        RECT 2.790 151.840 4.090 152.290 ;
        RECT 3.790 151.440 4.090 151.840 ;
        RECT 5.510 151.460 5.740 153.990 ;
        RECT 12.760 153.900 18.010 154.200 ;
        RECT 28.430 154.130 28.730 155.130 ;
        RECT 29.180 154.530 29.480 155.580 ;
        RECT 31.780 154.480 32.030 156.220 ;
        RECT 34.150 156.210 51.110 156.530 ;
        RECT 35.030 156.200 51.110 156.210 ;
        RECT 35.030 156.170 47.010 156.200 ;
        RECT 35.030 156.160 35.920 156.170 ;
        RECT 32.480 154.130 32.740 155.680 ;
        RECT 33.570 154.130 33.770 154.140 ;
        RECT 4.580 151.440 5.740 151.460 ;
        RECT 3.790 151.260 5.740 151.440 ;
        RECT 8.680 152.260 8.940 153.460 ;
        RECT 8.680 151.750 8.930 152.260 ;
        RECT 10.570 152.250 10.830 153.460 ;
        RECT 12.960 152.350 13.210 153.900 ;
        RECT 10.570 152.090 10.960 152.250 ;
        RECT 10.560 151.960 10.960 152.090 ;
        RECT 13.660 151.960 13.920 153.570 ;
        RECT 16.210 152.500 16.510 153.550 ;
        RECT 16.960 152.950 17.260 153.900 ;
        RECT 17.810 153.890 18.010 153.900 ;
        RECT 28.380 153.830 33.770 154.130 ;
        RECT 17.460 153.000 17.760 153.050 ;
        RECT 17.460 152.650 18.360 153.000 ;
        RECT 33.570 152.590 33.770 153.830 ;
        RECT 50.730 152.630 51.090 156.200 ;
        RECT 26.010 152.570 27.200 152.580 ;
        RECT 28.190 152.570 29.380 152.580 ;
        RECT 30.410 152.570 31.600 152.580 ;
        RECT 32.590 152.570 33.780 152.590 ;
        RECT 23.800 152.560 33.780 152.570 ;
        RECT 20.410 152.540 21.600 152.550 ;
        RECT 22.690 152.540 33.780 152.560 ;
        RECT 9.180 151.750 9.470 151.910 ;
        RECT 10.560 151.900 10.820 151.960 ;
        RECT 8.680 151.560 9.470 151.750 ;
        RECT 8.680 151.360 8.930 151.560 ;
        RECT 9.180 151.450 9.470 151.560 ;
        RECT 10.570 151.360 10.820 151.900 ;
        RECT 13.650 151.900 13.920 151.960 ;
        RECT 15.200 152.240 16.510 152.500 ;
        RECT 18.570 152.310 33.780 152.540 ;
        RECT 45.860 152.330 51.110 152.630 ;
        RECT 18.570 152.300 32.730 152.310 ;
        RECT 18.570 152.290 26.100 152.300 ;
        RECT 27.110 152.290 28.300 152.300 ;
        RECT 29.260 152.290 30.450 152.300 ;
        RECT 31.540 152.290 32.730 152.300 ;
        RECT 18.570 152.280 23.880 152.290 ;
        RECT 18.570 152.270 22.740 152.280 ;
        RECT 18.570 152.260 20.460 152.270 ;
        RECT 21.550 152.260 22.740 152.270 ;
        RECT 18.570 152.250 19.290 152.260 ;
        RECT 15.200 151.900 15.510 152.240 ;
        RECT 11.210 151.370 12.850 151.760 ;
        RECT 13.650 151.610 15.510 151.900 ;
        RECT 13.650 151.600 13.960 151.610 ;
        RECT 15.200 151.600 15.510 151.610 ;
        RECT 3.790 151.250 4.440 151.260 ;
        RECT 3.790 150.920 4.090 151.250 ;
        RECT 3.070 150.470 4.090 150.920 ;
        RECT 8.680 150.760 8.970 151.360 ;
        RECT 10.570 150.760 10.860 151.360 ;
        RECT 3.790 150.460 4.090 150.470 ;
        RECT 12.910 150.150 13.210 151.150 ;
        RECT 13.660 150.550 13.960 151.600 ;
        RECT 16.260 150.500 16.510 152.240 ;
        RECT 16.960 150.150 17.220 151.700 ;
        RECT 41.780 150.690 42.040 151.890 ;
        RECT 41.780 150.180 42.030 150.690 ;
        RECT 43.670 150.680 43.930 151.890 ;
        RECT 46.060 150.780 46.310 152.330 ;
        RECT 43.670 150.520 44.060 150.680 ;
        RECT 43.660 150.390 44.060 150.520 ;
        RECT 46.760 150.390 47.020 152.000 ;
        RECT 49.310 150.930 49.610 151.980 ;
        RECT 50.060 151.380 50.360 152.330 ;
        RECT 50.560 151.430 50.860 151.480 ;
        RECT 50.560 151.080 51.460 151.430 ;
        RECT 42.280 150.180 42.570 150.340 ;
        RECT 43.660 150.330 43.920 150.390 ;
        RECT 12.860 150.140 18.110 150.150 ;
        RECT 2.740 150.060 2.990 150.070 ;
        RECT 2.740 149.600 3.720 150.060 ;
        RECT 12.860 149.850 18.130 150.140 ;
        RECT 2.740 149.300 2.990 149.600 ;
        RECT 10.710 149.510 12.550 149.520 ;
        RECT 17.960 149.510 18.130 149.850 ;
        RECT 4.450 149.500 4.690 149.510 ;
        RECT 5.530 149.500 18.130 149.510 ;
        RECT 4.450 149.340 18.130 149.500 ;
        RECT 41.780 149.990 42.570 150.180 ;
        RECT 41.780 149.790 42.030 149.990 ;
        RECT 42.280 149.880 42.570 149.990 ;
        RECT 43.670 149.790 43.920 150.330 ;
        RECT 46.750 150.330 47.020 150.390 ;
        RECT 48.300 150.670 49.610 150.930 ;
        RECT 51.670 150.980 53.340 151.000 ;
        RECT 68.480 150.980 68.790 162.330 ;
        RECT 99.310 160.610 99.560 166.250 ;
        RECT 100.850 166.180 101.080 251.980 ;
        RECT 105.310 251.410 105.550 252.530 ;
        RECT 105.300 251.190 105.580 251.410 ;
        RECT 106.480 251.340 115.750 251.350 ;
        RECT 117.630 251.340 119.550 251.350 ;
        RECT 105.300 251.010 105.590 251.190 ;
        RECT 105.310 250.740 105.590 251.010 ;
        RECT 106.480 251.150 119.550 251.340 ;
        RECT 106.480 251.140 118.840 251.150 ;
        RECT 105.310 250.510 105.610 250.740 ;
        RECT 105.320 250.340 105.610 250.510 ;
        RECT 105.330 249.540 105.590 250.340 ;
        RECT 106.480 250.130 106.690 251.140 ;
        RECT 115.740 251.130 117.640 251.140 ;
        RECT 119.370 250.400 119.550 251.150 ;
        RECT 105.330 248.940 105.580 249.540 ;
        RECT 106.480 249.120 106.680 250.130 ;
        RECT 114.290 250.100 119.550 250.400 ;
        RECT 104.540 248.490 105.580 248.940 ;
        RECT 104.520 247.040 105.480 247.490 ;
        RECT 105.230 246.990 105.480 247.040 ;
        RECT 106.490 246.990 106.680 249.120 ;
        RECT 105.230 246.790 106.680 246.990 ;
        RECT 110.210 248.460 110.470 249.660 ;
        RECT 110.210 247.950 110.460 248.460 ;
        RECT 112.100 248.450 112.360 249.660 ;
        RECT 114.490 248.550 114.740 250.100 ;
        RECT 112.100 248.290 112.490 248.450 ;
        RECT 112.090 248.160 112.490 248.290 ;
        RECT 115.190 248.160 115.450 249.770 ;
        RECT 117.740 248.700 118.040 249.750 ;
        RECT 118.490 249.150 118.790 250.100 ;
        RECT 118.990 249.200 119.290 249.250 ;
        RECT 118.990 248.850 119.890 249.200 ;
        RECT 121.600 249.070 121.820 249.080 ;
        RECT 121.600 248.880 135.280 249.070 ;
        RECT 121.600 248.750 121.820 248.880 ;
        RECT 110.710 247.950 111.000 248.110 ;
        RECT 112.090 248.100 112.350 248.160 ;
        RECT 110.210 247.760 111.000 247.950 ;
        RECT 110.210 247.560 110.460 247.760 ;
        RECT 110.710 247.650 111.000 247.760 ;
        RECT 112.100 247.560 112.350 248.100 ;
        RECT 115.180 248.100 115.450 248.160 ;
        RECT 116.730 248.440 118.040 248.700 ;
        RECT 120.140 248.450 121.820 248.750 ;
        RECT 120.140 248.440 121.800 248.450 ;
        RECT 116.730 248.100 117.040 248.440 ;
        RECT 112.740 247.570 114.380 247.960 ;
        RECT 115.180 247.810 117.040 248.100 ;
        RECT 115.180 247.800 115.490 247.810 ;
        RECT 116.730 247.800 117.040 247.810 ;
        RECT 110.210 246.960 110.500 247.560 ;
        RECT 112.100 246.960 112.390 247.560 ;
        RECT 105.230 246.700 105.480 246.790 ;
        RECT 104.500 246.250 105.480 246.700 ;
        RECT 114.440 246.350 114.740 247.350 ;
        RECT 115.190 246.750 115.490 247.800 ;
        RECT 117.790 246.700 118.040 248.440 ;
        RECT 135.030 247.980 135.280 248.880 ;
        RECT 118.490 246.350 118.750 247.900 ;
        RECT 129.970 247.680 135.280 247.980 ;
        RECT 114.390 246.330 119.640 246.350 ;
        RECT 114.390 246.050 119.760 246.330 ;
        RECT 107.840 245.650 108.120 245.720 ;
        RECT 109.020 245.680 109.300 245.710 ;
        RECT 119.470 245.680 119.760 246.050 ;
        RECT 109.020 245.670 119.760 245.680 ;
        RECT 106.430 245.450 108.120 245.650 ;
        RECT 105.220 245.250 105.500 245.260 ;
        RECT 104.480 244.800 105.500 245.250 ;
        RECT 106.430 244.800 106.660 245.450 ;
        RECT 107.840 245.390 108.120 245.450 ;
        RECT 109.000 245.440 119.760 245.670 ;
        RECT 109.020 245.430 119.760 245.440 ;
        RECT 125.890 246.040 126.150 247.240 ;
        RECT 125.890 245.530 126.140 246.040 ;
        RECT 127.780 246.030 128.040 247.240 ;
        RECT 130.170 246.130 130.420 247.680 ;
        RECT 127.780 245.870 128.170 246.030 ;
        RECT 127.770 245.740 128.170 245.870 ;
        RECT 130.870 245.740 131.130 247.350 ;
        RECT 133.420 246.280 133.720 247.330 ;
        RECT 134.170 246.730 134.470 247.680 ;
        RECT 134.670 246.780 134.970 246.830 ;
        RECT 134.670 246.430 135.570 246.780 ;
        RECT 148.330 246.380 152.800 246.410 ;
        RECT 137.390 246.350 152.800 246.380 ;
        RECT 136.720 246.330 152.800 246.350 ;
        RECT 126.390 245.530 126.680 245.690 ;
        RECT 127.770 245.680 128.030 245.740 ;
        RECT 109.020 245.420 119.720 245.430 ;
        RECT 109.020 245.380 109.300 245.420 ;
        RECT 125.890 245.340 126.680 245.530 ;
        RECT 125.890 245.140 126.140 245.340 ;
        RECT 126.390 245.230 126.680 245.340 ;
        RECT 127.780 245.140 128.030 245.680 ;
        RECT 130.860 245.680 131.130 245.740 ;
        RECT 132.410 246.020 133.720 246.280 ;
        RECT 132.410 245.680 132.720 246.020 ;
        RECT 128.420 245.150 130.060 245.540 ;
        RECT 130.860 245.390 132.720 245.680 ;
        RECT 130.860 245.380 131.170 245.390 ;
        RECT 132.410 245.380 132.720 245.390 ;
        RECT 107.820 244.820 108.090 244.900 ;
        RECT 105.220 244.590 106.660 244.800 ;
        RECT 107.210 244.600 108.090 244.820 ;
        RECT 105.220 243.540 105.500 244.590 ;
        RECT 107.210 243.790 107.430 244.600 ;
        RECT 107.820 244.570 108.090 244.600 ;
        RECT 108.950 244.860 109.240 244.910 ;
        RECT 108.950 244.680 119.700 244.860 ;
        RECT 108.950 244.580 109.240 244.680 ;
        RECT 113.790 244.670 117.420 244.680 ;
        RECT 119.500 244.000 119.700 244.680 ;
        RECT 125.890 244.540 126.180 245.140 ;
        RECT 127.780 244.540 128.070 245.140 ;
        RECT 104.500 243.090 105.500 243.540 ;
        RECT 104.480 241.640 105.780 242.090 ;
        RECT 105.480 241.240 105.780 241.640 ;
        RECT 107.200 241.260 107.430 243.790 ;
        RECT 114.450 243.700 119.700 244.000 ;
        RECT 130.120 243.930 130.420 244.930 ;
        RECT 130.870 244.330 131.170 245.380 ;
        RECT 133.470 244.280 133.720 246.020 ;
        RECT 135.840 246.010 152.800 246.330 ;
        RECT 136.720 246.000 152.800 246.010 ;
        RECT 136.720 245.970 148.700 246.000 ;
        RECT 136.720 245.960 137.610 245.970 ;
        RECT 134.170 243.930 134.430 245.480 ;
        RECT 135.260 243.930 135.460 243.940 ;
        RECT 106.270 241.240 107.430 241.260 ;
        RECT 105.480 241.060 107.430 241.240 ;
        RECT 110.370 242.060 110.630 243.260 ;
        RECT 110.370 241.550 110.620 242.060 ;
        RECT 112.260 242.050 112.520 243.260 ;
        RECT 114.650 242.150 114.900 243.700 ;
        RECT 112.260 241.890 112.650 242.050 ;
        RECT 112.250 241.760 112.650 241.890 ;
        RECT 115.350 241.760 115.610 243.370 ;
        RECT 117.900 242.300 118.200 243.350 ;
        RECT 118.650 242.750 118.950 243.700 ;
        RECT 119.500 243.690 119.700 243.700 ;
        RECT 130.070 243.630 135.460 243.930 ;
        RECT 119.150 242.800 119.450 242.850 ;
        RECT 119.150 242.450 120.050 242.800 ;
        RECT 135.260 242.390 135.460 243.630 ;
        RECT 152.420 242.430 152.780 246.000 ;
        RECT 226.840 242.980 227.090 255.400 ;
        RECT 337.370 255.380 456.980 255.420 ;
        RECT 337.370 255.370 374.060 255.380 ;
        RECT 463.370 255.340 463.600 255.420 ;
        RECT 296.630 252.700 338.600 252.720 ;
        RECT 236.530 252.470 342.090 252.700 ;
        RECT 236.530 252.450 296.880 252.470 ;
        RECT 236.530 252.420 255.030 252.450 ;
        RECT 127.700 242.370 128.890 242.380 ;
        RECT 129.880 242.370 131.070 242.380 ;
        RECT 132.100 242.370 133.290 242.380 ;
        RECT 134.280 242.370 135.470 242.390 ;
        RECT 125.490 242.360 135.470 242.370 ;
        RECT 122.100 242.340 123.290 242.350 ;
        RECT 124.380 242.340 135.470 242.360 ;
        RECT 110.870 241.550 111.160 241.710 ;
        RECT 112.250 241.700 112.510 241.760 ;
        RECT 110.370 241.360 111.160 241.550 ;
        RECT 110.370 241.160 110.620 241.360 ;
        RECT 110.870 241.250 111.160 241.360 ;
        RECT 112.260 241.160 112.510 241.700 ;
        RECT 115.340 241.700 115.610 241.760 ;
        RECT 116.890 242.040 118.200 242.300 ;
        RECT 120.260 242.110 135.470 242.340 ;
        RECT 147.550 242.130 152.800 242.430 ;
        RECT 120.260 242.100 134.420 242.110 ;
        RECT 120.260 242.090 127.790 242.100 ;
        RECT 128.800 242.090 129.990 242.100 ;
        RECT 130.950 242.090 132.140 242.100 ;
        RECT 133.230 242.090 134.420 242.100 ;
        RECT 120.260 242.080 125.570 242.090 ;
        RECT 120.260 242.070 124.430 242.080 ;
        RECT 120.260 242.060 122.150 242.070 ;
        RECT 123.240 242.060 124.430 242.070 ;
        RECT 120.260 242.050 120.980 242.060 ;
        RECT 116.890 241.700 117.200 242.040 ;
        RECT 112.900 241.170 114.540 241.560 ;
        RECT 115.340 241.410 117.200 241.700 ;
        RECT 115.340 241.400 115.650 241.410 ;
        RECT 116.890 241.400 117.200 241.410 ;
        RECT 105.480 241.050 106.130 241.060 ;
        RECT 105.480 240.720 105.780 241.050 ;
        RECT 104.760 240.270 105.780 240.720 ;
        RECT 110.370 240.560 110.660 241.160 ;
        RECT 112.260 240.560 112.550 241.160 ;
        RECT 105.480 240.260 105.780 240.270 ;
        RECT 114.600 239.950 114.900 240.950 ;
        RECT 115.350 240.350 115.650 241.400 ;
        RECT 117.950 240.300 118.200 242.040 ;
        RECT 118.650 239.950 118.910 241.500 ;
        RECT 143.470 240.490 143.730 241.690 ;
        RECT 143.470 239.980 143.720 240.490 ;
        RECT 145.360 240.480 145.620 241.690 ;
        RECT 147.750 240.580 148.000 242.130 ;
        RECT 145.360 240.320 145.750 240.480 ;
        RECT 145.350 240.190 145.750 240.320 ;
        RECT 148.450 240.190 148.710 241.800 ;
        RECT 151.000 240.730 151.300 241.780 ;
        RECT 151.750 241.180 152.050 242.130 ;
        RECT 152.250 241.230 152.550 241.280 ;
        RECT 152.250 240.880 153.150 241.230 ;
        RECT 143.970 239.980 144.260 240.140 ;
        RECT 145.350 240.130 145.610 240.190 ;
        RECT 114.550 239.940 119.800 239.950 ;
        RECT 104.430 239.860 104.680 239.870 ;
        RECT 104.430 239.400 105.410 239.860 ;
        RECT 114.550 239.650 119.820 239.940 ;
        RECT 104.430 239.100 104.680 239.400 ;
        RECT 112.400 239.310 114.240 239.320 ;
        RECT 119.650 239.310 119.820 239.650 ;
        RECT 106.140 239.300 106.380 239.310 ;
        RECT 107.220 239.300 119.820 239.310 ;
        RECT 106.140 239.140 119.820 239.300 ;
        RECT 143.470 239.790 144.260 239.980 ;
        RECT 143.470 239.590 143.720 239.790 ;
        RECT 143.970 239.680 144.260 239.790 ;
        RECT 145.360 239.590 145.610 240.130 ;
        RECT 148.440 240.130 148.710 240.190 ;
        RECT 149.990 240.470 151.300 240.730 ;
        RECT 153.360 240.770 155.030 240.800 ;
        RECT 170.110 240.770 170.360 240.780 ;
        RECT 153.360 240.500 170.360 240.770 ;
        RECT 153.360 240.490 166.860 240.500 ;
        RECT 154.640 240.470 166.860 240.490 ;
        RECT 149.990 240.130 150.300 240.470 ;
        RECT 146.000 239.600 147.640 239.990 ;
        RECT 148.440 239.840 150.300 240.130 ;
        RECT 148.440 239.830 148.750 239.840 ;
        RECT 149.990 239.830 150.300 239.840 ;
        RECT 106.140 239.130 117.650 239.140 ;
        RECT 106.130 239.120 112.450 239.130 ;
        RECT 114.000 239.120 117.650 239.130 ;
        RECT 106.130 239.110 108.000 239.120 ;
        RECT 106.130 239.100 106.380 239.110 ;
        RECT 104.430 238.930 106.380 239.100 ;
        RECT 143.470 238.990 143.760 239.590 ;
        RECT 145.360 238.990 145.650 239.590 ;
        RECT 104.430 238.710 104.680 238.930 ;
        RECT 104.430 238.540 105.470 238.710 ;
        RECT 105.280 237.680 105.470 238.540 ;
        RECT 147.700 238.380 148.000 239.380 ;
        RECT 148.450 238.780 148.750 239.830 ;
        RECT 151.050 238.730 151.300 240.470 ;
        RECT 151.750 238.380 152.010 239.930 ;
        RECT 152.630 238.380 152.970 238.450 ;
        RECT 147.650 238.080 152.970 238.380 ;
        RECT 104.490 237.240 105.470 237.680 ;
        RECT 104.490 237.230 105.440 237.240 ;
        RECT 106.310 236.920 115.580 236.930 ;
        RECT 117.460 236.920 119.380 236.930 ;
        RECT 104.160 236.820 104.350 236.830 ;
        RECT 104.160 236.360 105.140 236.820 ;
        RECT 106.310 236.730 119.380 236.920 ;
        RECT 106.310 236.720 118.670 236.730 ;
        RECT 104.160 235.570 104.350 236.360 ;
        RECT 106.310 235.710 106.520 236.720 ;
        RECT 115.570 236.710 117.470 236.720 ;
        RECT 119.200 235.980 119.380 236.730 ;
        RECT 105.160 235.570 105.430 235.580 ;
        RECT 104.160 235.360 105.430 235.570 ;
        RECT 105.160 235.150 105.430 235.360 ;
        RECT 105.160 234.520 105.410 235.150 ;
        RECT 106.310 234.700 106.510 235.710 ;
        RECT 114.120 235.680 119.380 235.980 ;
        RECT 104.370 234.070 105.410 234.520 ;
        RECT 104.350 232.620 105.310 233.070 ;
        RECT 105.060 232.570 105.310 232.620 ;
        RECT 106.320 232.570 106.510 234.700 ;
        RECT 105.060 232.370 106.510 232.570 ;
        RECT 110.040 234.040 110.300 235.240 ;
        RECT 110.040 233.530 110.290 234.040 ;
        RECT 111.930 234.030 112.190 235.240 ;
        RECT 114.320 234.130 114.570 235.680 ;
        RECT 111.930 233.870 112.320 234.030 ;
        RECT 111.920 233.740 112.320 233.870 ;
        RECT 115.020 233.740 115.280 235.350 ;
        RECT 117.570 234.280 117.870 235.330 ;
        RECT 118.320 234.730 118.620 235.680 ;
        RECT 118.820 234.780 119.120 234.830 ;
        RECT 118.820 234.430 119.720 234.780 ;
        RECT 121.430 234.650 121.650 234.660 ;
        RECT 121.430 234.460 135.110 234.650 ;
        RECT 121.430 234.330 121.650 234.460 ;
        RECT 110.540 233.530 110.830 233.690 ;
        RECT 111.920 233.680 112.180 233.740 ;
        RECT 110.040 233.340 110.830 233.530 ;
        RECT 110.040 233.140 110.290 233.340 ;
        RECT 110.540 233.230 110.830 233.340 ;
        RECT 111.930 233.140 112.180 233.680 ;
        RECT 115.010 233.680 115.280 233.740 ;
        RECT 116.560 234.020 117.870 234.280 ;
        RECT 119.970 234.030 121.650 234.330 ;
        RECT 119.970 234.020 121.630 234.030 ;
        RECT 116.560 233.680 116.870 234.020 ;
        RECT 112.570 233.150 114.210 233.540 ;
        RECT 115.010 233.390 116.870 233.680 ;
        RECT 115.010 233.380 115.320 233.390 ;
        RECT 116.560 233.380 116.870 233.390 ;
        RECT 110.040 232.540 110.330 233.140 ;
        RECT 111.930 232.540 112.220 233.140 ;
        RECT 105.060 232.280 105.310 232.370 ;
        RECT 104.330 231.830 105.310 232.280 ;
        RECT 114.270 231.930 114.570 232.930 ;
        RECT 115.020 232.330 115.320 233.380 ;
        RECT 117.620 232.280 117.870 234.020 ;
        RECT 134.860 233.560 135.110 234.460 ;
        RECT 118.320 231.930 118.580 233.480 ;
        RECT 129.800 233.260 135.110 233.560 ;
        RECT 114.220 231.910 119.470 231.930 ;
        RECT 114.220 231.630 119.590 231.910 ;
        RECT 107.670 231.230 107.950 231.300 ;
        RECT 108.850 231.260 109.130 231.290 ;
        RECT 119.300 231.260 119.590 231.630 ;
        RECT 108.850 231.250 119.590 231.260 ;
        RECT 106.260 231.030 107.950 231.230 ;
        RECT 105.050 230.830 105.330 230.840 ;
        RECT 104.310 230.380 105.330 230.830 ;
        RECT 106.260 230.380 106.490 231.030 ;
        RECT 107.670 230.970 107.950 231.030 ;
        RECT 108.830 231.020 119.590 231.250 ;
        RECT 108.850 231.010 119.590 231.020 ;
        RECT 125.720 231.620 125.980 232.820 ;
        RECT 125.720 231.110 125.970 231.620 ;
        RECT 127.610 231.610 127.870 232.820 ;
        RECT 130.000 231.710 130.250 233.260 ;
        RECT 127.610 231.450 128.000 231.610 ;
        RECT 127.600 231.320 128.000 231.450 ;
        RECT 130.700 231.320 130.960 232.930 ;
        RECT 133.250 231.860 133.550 232.910 ;
        RECT 134.000 232.310 134.300 233.260 ;
        RECT 134.500 232.360 134.800 232.410 ;
        RECT 134.500 232.010 135.400 232.360 ;
        RECT 152.630 231.960 152.970 238.080 ;
        RECT 152.060 231.940 153.020 231.960 ;
        RECT 136.540 231.920 140.820 231.930 ;
        RECT 148.220 231.920 153.020 231.940 ;
        RECT 136.540 231.910 153.020 231.920 ;
        RECT 126.220 231.110 126.510 231.270 ;
        RECT 127.600 231.260 127.860 231.320 ;
        RECT 108.850 231.000 119.550 231.010 ;
        RECT 108.850 230.960 109.130 231.000 ;
        RECT 125.720 230.920 126.510 231.110 ;
        RECT 125.720 230.720 125.970 230.920 ;
        RECT 126.220 230.810 126.510 230.920 ;
        RECT 127.610 230.720 127.860 231.260 ;
        RECT 130.690 231.260 130.960 231.320 ;
        RECT 132.240 231.600 133.550 231.860 ;
        RECT 132.240 231.260 132.550 231.600 ;
        RECT 128.250 230.730 129.890 231.120 ;
        RECT 130.690 230.970 132.550 231.260 ;
        RECT 130.690 230.960 131.000 230.970 ;
        RECT 132.240 230.960 132.550 230.970 ;
        RECT 107.650 230.400 107.920 230.480 ;
        RECT 105.050 230.170 106.490 230.380 ;
        RECT 107.040 230.180 107.920 230.400 ;
        RECT 105.050 229.120 105.330 230.170 ;
        RECT 107.040 229.370 107.260 230.180 ;
        RECT 107.650 230.150 107.920 230.180 ;
        RECT 108.780 230.440 109.070 230.490 ;
        RECT 108.780 230.260 119.530 230.440 ;
        RECT 108.780 230.160 109.070 230.260 ;
        RECT 113.620 230.250 117.250 230.260 ;
        RECT 119.330 229.580 119.530 230.260 ;
        RECT 125.720 230.120 126.010 230.720 ;
        RECT 127.610 230.120 127.900 230.720 ;
        RECT 104.330 228.670 105.330 229.120 ;
        RECT 104.310 227.220 105.610 227.670 ;
        RECT 105.310 226.820 105.610 227.220 ;
        RECT 107.030 226.840 107.260 229.370 ;
        RECT 114.280 229.280 119.530 229.580 ;
        RECT 129.950 229.510 130.250 230.510 ;
        RECT 130.700 229.910 131.000 230.960 ;
        RECT 133.300 229.860 133.550 231.600 ;
        RECT 135.670 231.600 153.020 231.910 ;
        RECT 135.670 231.590 148.680 231.600 ;
        RECT 140.530 231.580 148.680 231.590 ;
        RECT 152.060 231.560 153.020 231.600 ;
        RECT 152.630 231.550 152.970 231.560 ;
        RECT 134.000 229.510 134.260 231.060 ;
        RECT 135.090 229.510 135.290 229.520 ;
        RECT 106.100 226.820 107.260 226.840 ;
        RECT 105.310 226.640 107.260 226.820 ;
        RECT 110.200 227.640 110.460 228.840 ;
        RECT 110.200 227.130 110.450 227.640 ;
        RECT 112.090 227.630 112.350 228.840 ;
        RECT 114.480 227.730 114.730 229.280 ;
        RECT 112.090 227.470 112.480 227.630 ;
        RECT 112.080 227.340 112.480 227.470 ;
        RECT 115.180 227.340 115.440 228.950 ;
        RECT 117.730 227.880 118.030 228.930 ;
        RECT 118.480 228.330 118.780 229.280 ;
        RECT 119.330 229.270 119.530 229.280 ;
        RECT 129.900 229.210 135.290 229.510 ;
        RECT 118.980 228.380 119.280 228.430 ;
        RECT 118.980 228.030 119.880 228.380 ;
        RECT 135.090 227.970 135.290 229.210 ;
        RECT 127.530 227.950 128.720 227.960 ;
        RECT 129.710 227.950 130.900 227.960 ;
        RECT 131.930 227.950 133.120 227.960 ;
        RECT 134.110 227.950 135.300 227.970 ;
        RECT 125.320 227.940 135.300 227.950 ;
        RECT 121.930 227.920 123.120 227.930 ;
        RECT 124.210 227.920 135.300 227.940 ;
        RECT 110.700 227.130 110.990 227.290 ;
        RECT 112.080 227.280 112.340 227.340 ;
        RECT 110.200 226.940 110.990 227.130 ;
        RECT 110.200 226.740 110.450 226.940 ;
        RECT 110.700 226.830 110.990 226.940 ;
        RECT 112.090 226.740 112.340 227.280 ;
        RECT 115.170 227.280 115.440 227.340 ;
        RECT 116.720 227.620 118.030 227.880 ;
        RECT 120.090 227.690 135.300 227.920 ;
        RECT 120.090 227.680 134.250 227.690 ;
        RECT 120.090 227.670 127.620 227.680 ;
        RECT 128.630 227.670 129.820 227.680 ;
        RECT 130.780 227.670 131.970 227.680 ;
        RECT 133.060 227.670 134.250 227.680 ;
        RECT 120.090 227.660 125.400 227.670 ;
        RECT 120.090 227.650 124.260 227.660 ;
        RECT 120.090 227.640 121.980 227.650 ;
        RECT 123.070 227.640 124.260 227.650 ;
        RECT 120.090 227.630 120.810 227.640 ;
        RECT 116.720 227.280 117.030 227.620 ;
        RECT 112.730 226.750 114.370 227.140 ;
        RECT 115.170 226.990 117.030 227.280 ;
        RECT 115.170 226.980 115.480 226.990 ;
        RECT 116.720 226.980 117.030 226.990 ;
        RECT 105.310 226.630 105.960 226.640 ;
        RECT 105.310 226.300 105.610 226.630 ;
        RECT 104.590 225.850 105.610 226.300 ;
        RECT 110.200 226.140 110.490 226.740 ;
        RECT 112.090 226.140 112.380 226.740 ;
        RECT 105.310 225.840 105.610 225.850 ;
        RECT 114.430 225.530 114.730 226.530 ;
        RECT 115.180 225.930 115.480 226.980 ;
        RECT 117.780 225.880 118.030 227.620 ;
        RECT 170.110 227.360 170.370 240.500 ;
        RECT 170.100 227.240 170.370 227.360 ;
        RECT 118.480 225.530 118.740 227.080 ;
        RECT 170.100 226.410 170.360 227.240 ;
        RECT 165.080 226.110 170.360 226.410 ;
        RECT 114.380 225.520 119.630 225.530 ;
        RECT 104.260 225.440 104.510 225.450 ;
        RECT 104.260 224.980 105.240 225.440 ;
        RECT 114.380 225.230 119.650 225.520 ;
        RECT 104.260 224.680 104.510 224.980 ;
        RECT 112.230 224.890 114.070 224.900 ;
        RECT 119.480 224.890 119.650 225.230 ;
        RECT 105.970 224.880 106.210 224.890 ;
        RECT 107.050 224.880 119.650 224.890 ;
        RECT 105.970 224.720 119.650 224.880 ;
        RECT 105.970 224.710 117.480 224.720 ;
        RECT 105.960 224.700 112.280 224.710 ;
        RECT 113.830 224.700 117.480 224.710 ;
        RECT 105.960 224.690 107.830 224.700 ;
        RECT 105.960 224.680 106.210 224.690 ;
        RECT 104.260 224.510 106.210 224.680 ;
        RECT 104.260 224.210 104.530 224.510 ;
        RECT 104.270 223.950 104.530 224.210 ;
        RECT 161.000 224.470 161.260 225.670 ;
        RECT 161.000 223.960 161.250 224.470 ;
        RECT 162.890 224.460 163.150 225.670 ;
        RECT 165.280 224.560 165.530 226.110 ;
        RECT 162.890 224.300 163.280 224.460 ;
        RECT 162.880 224.170 163.280 224.300 ;
        RECT 165.980 224.170 166.240 225.780 ;
        RECT 168.530 224.710 168.830 225.760 ;
        RECT 169.280 225.160 169.580 226.110 ;
        RECT 169.780 225.210 170.080 225.260 ;
        RECT 169.780 224.860 170.680 225.210 ;
        RECT 161.500 223.960 161.790 224.120 ;
        RECT 162.880 224.110 163.140 224.170 ;
        RECT 104.250 223.560 104.550 223.950 ;
        RECT 161.000 223.770 161.790 223.960 ;
        RECT 161.000 223.570 161.250 223.770 ;
        RECT 161.500 223.660 161.790 223.770 ;
        RECT 162.890 223.570 163.140 224.110 ;
        RECT 165.970 224.110 166.240 224.170 ;
        RECT 167.520 224.450 168.830 224.710 ;
        RECT 170.950 224.650 171.730 224.750 ;
        RECT 170.950 224.480 184.530 224.650 ;
        RECT 170.950 224.470 184.520 224.480 ;
        RECT 170.950 224.450 171.730 224.470 ;
        RECT 167.520 224.110 167.830 224.450 ;
        RECT 163.530 223.580 165.170 223.970 ;
        RECT 165.970 223.820 167.830 224.110 ;
        RECT 165.970 223.810 166.280 223.820 ;
        RECT 167.520 223.810 167.830 223.820 ;
        RECT 104.250 223.330 105.740 223.560 ;
        RECT 105.490 222.400 105.740 223.330 ;
        RECT 161.000 222.970 161.290 223.570 ;
        RECT 162.890 222.970 163.180 223.570 ;
        RECT 104.690 221.940 105.740 222.400 ;
        RECT 165.230 222.360 165.530 223.360 ;
        RECT 165.980 222.760 166.280 223.810 ;
        RECT 168.580 222.710 168.830 224.450 ;
        RECT 169.280 222.360 169.540 223.910 ;
        RECT 165.180 222.060 170.450 222.360 ;
        RECT 105.490 221.930 105.740 221.940 ;
        RECT 104.360 221.530 104.610 221.540 ;
        RECT 104.360 221.080 105.340 221.530 ;
        RECT 106.450 221.270 115.720 221.280 ;
        RECT 117.600 221.270 119.520 221.280 ;
        RECT 106.450 221.080 119.520 221.270 ;
        RECT 104.360 220.470 104.610 221.080 ;
        RECT 106.450 221.070 118.810 221.080 ;
        RECT 104.360 220.220 105.570 220.470 ;
        RECT 105.300 219.470 105.560 220.220 ;
        RECT 106.450 220.060 106.660 221.070 ;
        RECT 115.710 221.060 117.610 221.070 ;
        RECT 119.340 220.330 119.520 221.080 ;
        RECT 105.300 218.870 105.550 219.470 ;
        RECT 106.450 219.050 106.650 220.060 ;
        RECT 114.260 220.030 119.520 220.330 ;
        RECT 104.510 218.420 105.550 218.870 ;
        RECT 104.490 216.970 105.450 217.420 ;
        RECT 105.200 216.920 105.450 216.970 ;
        RECT 106.460 216.920 106.650 219.050 ;
        RECT 105.200 216.720 106.650 216.920 ;
        RECT 110.180 218.390 110.440 219.590 ;
        RECT 110.180 217.880 110.430 218.390 ;
        RECT 112.070 218.380 112.330 219.590 ;
        RECT 114.460 218.480 114.710 220.030 ;
        RECT 112.070 218.220 112.460 218.380 ;
        RECT 112.060 218.090 112.460 218.220 ;
        RECT 115.160 218.090 115.420 219.700 ;
        RECT 117.710 218.630 118.010 219.680 ;
        RECT 118.460 219.080 118.760 220.030 ;
        RECT 118.960 219.130 119.260 219.180 ;
        RECT 118.960 218.780 119.860 219.130 ;
        RECT 121.570 219.000 121.790 219.010 ;
        RECT 121.570 218.810 135.250 219.000 ;
        RECT 121.570 218.680 121.790 218.810 ;
        RECT 110.680 217.880 110.970 218.040 ;
        RECT 112.060 218.030 112.320 218.090 ;
        RECT 110.180 217.690 110.970 217.880 ;
        RECT 110.180 217.490 110.430 217.690 ;
        RECT 110.680 217.580 110.970 217.690 ;
        RECT 112.070 217.490 112.320 218.030 ;
        RECT 115.150 218.030 115.420 218.090 ;
        RECT 116.700 218.370 118.010 218.630 ;
        RECT 120.110 218.380 121.790 218.680 ;
        RECT 120.110 218.370 121.770 218.380 ;
        RECT 116.700 218.030 117.010 218.370 ;
        RECT 112.710 217.500 114.350 217.890 ;
        RECT 115.150 217.740 117.010 218.030 ;
        RECT 115.150 217.730 115.460 217.740 ;
        RECT 116.700 217.730 117.010 217.740 ;
        RECT 110.180 216.890 110.470 217.490 ;
        RECT 112.070 216.890 112.360 217.490 ;
        RECT 105.200 216.630 105.450 216.720 ;
        RECT 104.470 216.180 105.450 216.630 ;
        RECT 114.410 216.280 114.710 217.280 ;
        RECT 115.160 216.680 115.460 217.730 ;
        RECT 117.760 216.630 118.010 218.370 ;
        RECT 135.000 217.910 135.250 218.810 ;
        RECT 118.460 216.280 118.720 217.830 ;
        RECT 129.940 217.610 135.250 217.910 ;
        RECT 114.360 216.260 119.610 216.280 ;
        RECT 114.360 215.980 119.730 216.260 ;
        RECT 107.810 215.580 108.090 215.650 ;
        RECT 108.990 215.610 109.270 215.640 ;
        RECT 119.440 215.610 119.730 215.980 ;
        RECT 108.990 215.600 119.730 215.610 ;
        RECT 106.400 215.380 108.090 215.580 ;
        RECT 105.190 215.180 105.470 215.190 ;
        RECT 104.450 214.730 105.470 215.180 ;
        RECT 106.400 214.730 106.630 215.380 ;
        RECT 107.810 215.320 108.090 215.380 ;
        RECT 108.970 215.370 119.730 215.600 ;
        RECT 108.990 215.360 119.730 215.370 ;
        RECT 125.860 215.970 126.120 217.170 ;
        RECT 125.860 215.460 126.110 215.970 ;
        RECT 127.750 215.960 128.010 217.170 ;
        RECT 130.140 216.060 130.390 217.610 ;
        RECT 127.750 215.800 128.140 215.960 ;
        RECT 127.740 215.670 128.140 215.800 ;
        RECT 130.840 215.670 131.100 217.280 ;
        RECT 133.390 216.210 133.690 217.260 ;
        RECT 134.140 216.660 134.440 217.610 ;
        RECT 134.640 216.710 134.940 216.760 ;
        RECT 134.640 216.360 135.540 216.710 ;
        RECT 148.300 216.310 152.770 216.340 ;
        RECT 137.360 216.280 152.770 216.310 ;
        RECT 136.690 216.260 152.770 216.280 ;
        RECT 126.360 215.460 126.650 215.620 ;
        RECT 127.740 215.610 128.000 215.670 ;
        RECT 108.990 215.350 119.690 215.360 ;
        RECT 108.990 215.310 109.270 215.350 ;
        RECT 125.860 215.270 126.650 215.460 ;
        RECT 125.860 215.070 126.110 215.270 ;
        RECT 126.360 215.160 126.650 215.270 ;
        RECT 127.750 215.070 128.000 215.610 ;
        RECT 130.830 215.610 131.100 215.670 ;
        RECT 132.380 215.950 133.690 216.210 ;
        RECT 132.380 215.610 132.690 215.950 ;
        RECT 128.390 215.080 130.030 215.470 ;
        RECT 130.830 215.320 132.690 215.610 ;
        RECT 130.830 215.310 131.140 215.320 ;
        RECT 132.380 215.310 132.690 215.320 ;
        RECT 107.790 214.750 108.060 214.830 ;
        RECT 105.190 214.520 106.630 214.730 ;
        RECT 107.180 214.530 108.060 214.750 ;
        RECT 105.190 213.470 105.470 214.520 ;
        RECT 107.180 213.720 107.400 214.530 ;
        RECT 107.790 214.500 108.060 214.530 ;
        RECT 108.920 214.790 109.210 214.840 ;
        RECT 108.920 214.610 119.670 214.790 ;
        RECT 108.920 214.510 109.210 214.610 ;
        RECT 113.760 214.600 117.390 214.610 ;
        RECT 119.470 213.930 119.670 214.610 ;
        RECT 125.860 214.470 126.150 215.070 ;
        RECT 127.750 214.470 128.040 215.070 ;
        RECT 104.470 213.020 105.470 213.470 ;
        RECT 104.450 211.570 105.750 212.020 ;
        RECT 105.450 211.170 105.750 211.570 ;
        RECT 107.170 211.190 107.400 213.720 ;
        RECT 114.420 213.630 119.670 213.930 ;
        RECT 130.090 213.860 130.390 214.860 ;
        RECT 130.840 214.260 131.140 215.310 ;
        RECT 133.440 214.210 133.690 215.950 ;
        RECT 135.810 215.940 152.770 216.260 ;
        RECT 136.690 215.930 152.770 215.940 ;
        RECT 136.690 215.900 148.670 215.930 ;
        RECT 136.690 215.890 137.580 215.900 ;
        RECT 134.140 213.860 134.400 215.410 ;
        RECT 135.230 213.860 135.430 213.870 ;
        RECT 106.240 211.170 107.400 211.190 ;
        RECT 105.450 210.990 107.400 211.170 ;
        RECT 110.340 211.990 110.600 213.190 ;
        RECT 110.340 211.480 110.590 211.990 ;
        RECT 112.230 211.980 112.490 213.190 ;
        RECT 114.620 212.080 114.870 213.630 ;
        RECT 112.230 211.820 112.620 211.980 ;
        RECT 112.220 211.690 112.620 211.820 ;
        RECT 115.320 211.690 115.580 213.300 ;
        RECT 117.870 212.230 118.170 213.280 ;
        RECT 118.620 212.680 118.920 213.630 ;
        RECT 119.470 213.620 119.670 213.630 ;
        RECT 130.040 213.560 135.430 213.860 ;
        RECT 119.120 212.730 119.420 212.780 ;
        RECT 119.120 212.380 120.020 212.730 ;
        RECT 135.230 212.320 135.430 213.560 ;
        RECT 152.390 212.360 152.750 215.930 ;
        RECT 127.670 212.300 128.860 212.310 ;
        RECT 129.850 212.300 131.040 212.310 ;
        RECT 132.070 212.300 133.260 212.310 ;
        RECT 134.250 212.300 135.440 212.320 ;
        RECT 125.460 212.290 135.440 212.300 ;
        RECT 122.070 212.270 123.260 212.280 ;
        RECT 124.350 212.270 135.440 212.290 ;
        RECT 110.840 211.480 111.130 211.640 ;
        RECT 112.220 211.630 112.480 211.690 ;
        RECT 110.340 211.290 111.130 211.480 ;
        RECT 110.340 211.090 110.590 211.290 ;
        RECT 110.840 211.180 111.130 211.290 ;
        RECT 112.230 211.090 112.480 211.630 ;
        RECT 115.310 211.630 115.580 211.690 ;
        RECT 116.860 211.970 118.170 212.230 ;
        RECT 120.230 212.040 135.440 212.270 ;
        RECT 147.520 212.060 152.770 212.360 ;
        RECT 120.230 212.030 134.390 212.040 ;
        RECT 120.230 212.020 127.760 212.030 ;
        RECT 128.770 212.020 129.960 212.030 ;
        RECT 130.920 212.020 132.110 212.030 ;
        RECT 133.200 212.020 134.390 212.030 ;
        RECT 120.230 212.010 125.540 212.020 ;
        RECT 120.230 212.000 124.400 212.010 ;
        RECT 120.230 211.990 122.120 212.000 ;
        RECT 123.210 211.990 124.400 212.000 ;
        RECT 120.230 211.980 120.950 211.990 ;
        RECT 116.860 211.630 117.170 211.970 ;
        RECT 112.870 211.100 114.510 211.490 ;
        RECT 115.310 211.340 117.170 211.630 ;
        RECT 115.310 211.330 115.620 211.340 ;
        RECT 116.860 211.330 117.170 211.340 ;
        RECT 105.450 210.980 106.100 210.990 ;
        RECT 105.450 210.650 105.750 210.980 ;
        RECT 104.730 210.200 105.750 210.650 ;
        RECT 110.340 210.490 110.630 211.090 ;
        RECT 112.230 210.490 112.520 211.090 ;
        RECT 105.450 210.190 105.750 210.200 ;
        RECT 114.570 209.880 114.870 210.880 ;
        RECT 115.320 210.280 115.620 211.330 ;
        RECT 117.920 210.230 118.170 211.970 ;
        RECT 118.620 209.880 118.880 211.430 ;
        RECT 143.440 210.420 143.700 211.620 ;
        RECT 143.440 209.910 143.690 210.420 ;
        RECT 145.330 210.410 145.590 211.620 ;
        RECT 147.720 210.510 147.970 212.060 ;
        RECT 145.330 210.250 145.720 210.410 ;
        RECT 145.320 210.120 145.720 210.250 ;
        RECT 148.420 210.120 148.680 211.730 ;
        RECT 150.970 210.660 151.270 211.710 ;
        RECT 151.720 211.110 152.020 212.060 ;
        RECT 152.220 211.160 152.520 211.210 ;
        RECT 152.220 210.810 153.120 211.160 ;
        RECT 143.940 209.910 144.230 210.070 ;
        RECT 145.320 210.060 145.580 210.120 ;
        RECT 114.520 209.870 119.770 209.880 ;
        RECT 104.400 209.790 104.650 209.800 ;
        RECT 104.400 209.330 105.380 209.790 ;
        RECT 114.520 209.580 119.790 209.870 ;
        RECT 104.400 209.030 104.650 209.330 ;
        RECT 112.370 209.240 114.210 209.250 ;
        RECT 119.620 209.240 119.790 209.580 ;
        RECT 106.110 209.230 106.350 209.240 ;
        RECT 107.190 209.230 119.790 209.240 ;
        RECT 106.110 209.070 119.790 209.230 ;
        RECT 143.440 209.720 144.230 209.910 ;
        RECT 143.440 209.520 143.690 209.720 ;
        RECT 143.940 209.610 144.230 209.720 ;
        RECT 145.330 209.520 145.580 210.060 ;
        RECT 148.410 210.060 148.680 210.120 ;
        RECT 149.960 210.400 151.270 210.660 ;
        RECT 153.330 210.710 155.000 210.730 ;
        RECT 170.140 210.710 170.450 222.060 ;
        RECT 153.330 210.420 170.490 210.710 ;
        RECT 154.020 210.410 170.490 210.420 ;
        RECT 149.960 210.060 150.270 210.400 ;
        RECT 145.970 209.530 147.610 209.920 ;
        RECT 148.410 209.770 150.270 210.060 ;
        RECT 148.410 209.760 148.720 209.770 ;
        RECT 149.960 209.760 150.270 209.770 ;
        RECT 106.110 209.060 117.620 209.070 ;
        RECT 106.100 209.050 112.420 209.060 ;
        RECT 113.970 209.050 117.620 209.060 ;
        RECT 106.100 209.040 107.970 209.050 ;
        RECT 106.100 209.030 106.350 209.040 ;
        RECT 104.400 208.860 106.350 209.030 ;
        RECT 143.440 208.920 143.730 209.520 ;
        RECT 145.330 208.920 145.620 209.520 ;
        RECT 104.400 208.640 104.650 208.860 ;
        RECT 104.400 208.470 105.440 208.640 ;
        RECT 105.250 207.610 105.440 208.470 ;
        RECT 147.670 208.310 147.970 209.310 ;
        RECT 148.420 208.710 148.720 209.760 ;
        RECT 151.020 208.660 151.270 210.400 ;
        RECT 151.720 208.310 151.980 209.860 ;
        RECT 152.600 208.310 152.940 208.380 ;
        RECT 147.620 208.010 152.940 208.310 ;
        RECT 104.460 207.170 105.440 207.610 ;
        RECT 104.460 207.160 105.410 207.170 ;
        RECT 106.280 206.850 115.550 206.860 ;
        RECT 117.430 206.850 119.350 206.860 ;
        RECT 104.130 206.750 104.320 206.760 ;
        RECT 104.130 206.290 105.110 206.750 ;
        RECT 106.280 206.660 119.350 206.850 ;
        RECT 106.280 206.650 118.640 206.660 ;
        RECT 104.130 205.500 104.320 206.290 ;
        RECT 106.280 205.640 106.490 206.650 ;
        RECT 115.540 206.640 117.440 206.650 ;
        RECT 119.170 205.910 119.350 206.660 ;
        RECT 105.130 205.500 105.400 205.510 ;
        RECT 104.130 205.290 105.400 205.500 ;
        RECT 105.130 205.080 105.400 205.290 ;
        RECT 105.130 204.450 105.380 205.080 ;
        RECT 106.280 204.630 106.480 205.640 ;
        RECT 114.090 205.610 119.350 205.910 ;
        RECT 104.340 204.000 105.380 204.450 ;
        RECT 104.320 202.550 105.280 203.000 ;
        RECT 105.030 202.500 105.280 202.550 ;
        RECT 106.290 202.500 106.480 204.630 ;
        RECT 105.030 202.300 106.480 202.500 ;
        RECT 110.010 203.970 110.270 205.170 ;
        RECT 110.010 203.460 110.260 203.970 ;
        RECT 111.900 203.960 112.160 205.170 ;
        RECT 114.290 204.060 114.540 205.610 ;
        RECT 111.900 203.800 112.290 203.960 ;
        RECT 111.890 203.670 112.290 203.800 ;
        RECT 114.990 203.670 115.250 205.280 ;
        RECT 117.540 204.210 117.840 205.260 ;
        RECT 118.290 204.660 118.590 205.610 ;
        RECT 118.790 204.710 119.090 204.760 ;
        RECT 118.790 204.360 119.690 204.710 ;
        RECT 121.400 204.580 121.620 204.590 ;
        RECT 121.400 204.390 135.080 204.580 ;
        RECT 121.400 204.260 121.620 204.390 ;
        RECT 110.510 203.460 110.800 203.620 ;
        RECT 111.890 203.610 112.150 203.670 ;
        RECT 110.010 203.270 110.800 203.460 ;
        RECT 110.010 203.070 110.260 203.270 ;
        RECT 110.510 203.160 110.800 203.270 ;
        RECT 111.900 203.070 112.150 203.610 ;
        RECT 114.980 203.610 115.250 203.670 ;
        RECT 116.530 203.950 117.840 204.210 ;
        RECT 119.940 203.960 121.620 204.260 ;
        RECT 119.940 203.950 121.600 203.960 ;
        RECT 116.530 203.610 116.840 203.950 ;
        RECT 112.540 203.080 114.180 203.470 ;
        RECT 114.980 203.320 116.840 203.610 ;
        RECT 114.980 203.310 115.290 203.320 ;
        RECT 116.530 203.310 116.840 203.320 ;
        RECT 110.010 202.470 110.300 203.070 ;
        RECT 111.900 202.470 112.190 203.070 ;
        RECT 105.030 202.210 105.280 202.300 ;
        RECT 104.300 201.760 105.280 202.210 ;
        RECT 114.240 201.860 114.540 202.860 ;
        RECT 114.990 202.260 115.290 203.310 ;
        RECT 117.590 202.210 117.840 203.950 ;
        RECT 134.830 203.490 135.080 204.390 ;
        RECT 118.290 201.860 118.550 203.410 ;
        RECT 129.770 203.190 135.080 203.490 ;
        RECT 114.190 201.840 119.440 201.860 ;
        RECT 114.190 201.560 119.560 201.840 ;
        RECT 107.640 201.160 107.920 201.230 ;
        RECT 108.820 201.190 109.100 201.220 ;
        RECT 119.270 201.190 119.560 201.560 ;
        RECT 108.820 201.180 119.560 201.190 ;
        RECT 106.230 200.960 107.920 201.160 ;
        RECT 105.020 200.760 105.300 200.770 ;
        RECT 104.280 200.310 105.300 200.760 ;
        RECT 106.230 200.310 106.460 200.960 ;
        RECT 107.640 200.900 107.920 200.960 ;
        RECT 108.800 200.950 119.560 201.180 ;
        RECT 108.820 200.940 119.560 200.950 ;
        RECT 125.690 201.550 125.950 202.750 ;
        RECT 125.690 201.040 125.940 201.550 ;
        RECT 127.580 201.540 127.840 202.750 ;
        RECT 129.970 201.640 130.220 203.190 ;
        RECT 127.580 201.380 127.970 201.540 ;
        RECT 127.570 201.250 127.970 201.380 ;
        RECT 130.670 201.250 130.930 202.860 ;
        RECT 133.220 201.790 133.520 202.840 ;
        RECT 133.970 202.240 134.270 203.190 ;
        RECT 134.470 202.290 134.770 202.340 ;
        RECT 134.470 201.940 135.370 202.290 ;
        RECT 152.600 201.890 152.940 208.010 ;
        RECT 184.340 205.210 184.520 224.470 ;
        RECT 184.320 204.160 184.530 205.210 ;
        RECT 184.320 204.080 184.540 204.160 ;
        RECT 184.330 202.010 184.540 204.080 ;
        RECT 184.320 201.970 184.540 202.010 ;
        RECT 152.030 201.870 152.990 201.890 ;
        RECT 136.510 201.850 140.790 201.860 ;
        RECT 148.190 201.850 152.990 201.870 ;
        RECT 136.510 201.840 152.990 201.850 ;
        RECT 126.190 201.040 126.480 201.200 ;
        RECT 127.570 201.190 127.830 201.250 ;
        RECT 108.820 200.930 119.520 200.940 ;
        RECT 108.820 200.890 109.100 200.930 ;
        RECT 125.690 200.850 126.480 201.040 ;
        RECT 125.690 200.650 125.940 200.850 ;
        RECT 126.190 200.740 126.480 200.850 ;
        RECT 127.580 200.650 127.830 201.190 ;
        RECT 130.660 201.190 130.930 201.250 ;
        RECT 132.210 201.530 133.520 201.790 ;
        RECT 132.210 201.190 132.520 201.530 ;
        RECT 128.220 200.660 129.860 201.050 ;
        RECT 130.660 200.900 132.520 201.190 ;
        RECT 130.660 200.890 130.970 200.900 ;
        RECT 132.210 200.890 132.520 200.900 ;
        RECT 107.620 200.330 107.890 200.410 ;
        RECT 105.020 200.100 106.460 200.310 ;
        RECT 107.010 200.110 107.890 200.330 ;
        RECT 105.020 199.050 105.300 200.100 ;
        RECT 107.010 199.300 107.230 200.110 ;
        RECT 107.620 200.080 107.890 200.110 ;
        RECT 108.750 200.370 109.040 200.420 ;
        RECT 108.750 200.190 119.500 200.370 ;
        RECT 108.750 200.090 109.040 200.190 ;
        RECT 113.590 200.180 117.220 200.190 ;
        RECT 119.300 199.510 119.500 200.190 ;
        RECT 125.690 200.050 125.980 200.650 ;
        RECT 127.580 200.050 127.870 200.650 ;
        RECT 104.300 198.600 105.300 199.050 ;
        RECT 104.280 197.150 105.580 197.600 ;
        RECT 105.280 196.750 105.580 197.150 ;
        RECT 107.000 196.770 107.230 199.300 ;
        RECT 114.250 199.210 119.500 199.510 ;
        RECT 129.920 199.440 130.220 200.440 ;
        RECT 130.670 199.840 130.970 200.890 ;
        RECT 133.270 199.790 133.520 201.530 ;
        RECT 135.640 201.530 152.990 201.840 ;
        RECT 135.640 201.520 148.650 201.530 ;
        RECT 140.500 201.510 148.650 201.520 ;
        RECT 152.030 201.490 152.990 201.530 ;
        RECT 152.600 201.480 152.940 201.490 ;
        RECT 133.970 199.440 134.230 200.990 ;
        RECT 184.320 200.120 184.530 201.970 ;
        RECT 179.280 199.820 184.530 200.120 ;
        RECT 135.060 199.440 135.260 199.450 ;
        RECT 106.070 196.750 107.230 196.770 ;
        RECT 105.280 196.570 107.230 196.750 ;
        RECT 110.170 197.570 110.430 198.770 ;
        RECT 110.170 197.060 110.420 197.570 ;
        RECT 112.060 197.560 112.320 198.770 ;
        RECT 114.450 197.660 114.700 199.210 ;
        RECT 112.060 197.400 112.450 197.560 ;
        RECT 112.050 197.270 112.450 197.400 ;
        RECT 115.150 197.270 115.410 198.880 ;
        RECT 117.700 197.810 118.000 198.860 ;
        RECT 118.450 198.260 118.750 199.210 ;
        RECT 119.300 199.200 119.500 199.210 ;
        RECT 129.870 199.140 135.260 199.440 ;
        RECT 118.950 198.310 119.250 198.360 ;
        RECT 118.950 197.960 119.850 198.310 ;
        RECT 135.060 197.900 135.260 199.140 ;
        RECT 175.200 198.180 175.460 199.380 ;
        RECT 127.500 197.880 128.690 197.890 ;
        RECT 129.680 197.880 130.870 197.890 ;
        RECT 131.900 197.880 133.090 197.890 ;
        RECT 134.080 197.880 135.270 197.900 ;
        RECT 125.290 197.870 135.270 197.880 ;
        RECT 121.900 197.850 123.090 197.860 ;
        RECT 124.180 197.850 135.270 197.870 ;
        RECT 110.670 197.060 110.960 197.220 ;
        RECT 112.050 197.210 112.310 197.270 ;
        RECT 110.170 196.870 110.960 197.060 ;
        RECT 110.170 196.670 110.420 196.870 ;
        RECT 110.670 196.760 110.960 196.870 ;
        RECT 112.060 196.670 112.310 197.210 ;
        RECT 115.140 197.210 115.410 197.270 ;
        RECT 116.690 197.550 118.000 197.810 ;
        RECT 120.060 197.620 135.270 197.850 ;
        RECT 175.200 197.670 175.450 198.180 ;
        RECT 177.090 198.170 177.350 199.380 ;
        RECT 179.480 198.270 179.730 199.820 ;
        RECT 177.090 198.010 177.480 198.170 ;
        RECT 177.080 197.880 177.480 198.010 ;
        RECT 180.180 197.880 180.440 199.490 ;
        RECT 182.730 198.420 183.030 199.470 ;
        RECT 183.480 198.870 183.780 199.820 ;
        RECT 184.320 199.810 184.530 199.820 ;
        RECT 183.980 198.920 184.280 198.970 ;
        RECT 183.980 198.570 184.880 198.920 ;
        RECT 185.840 198.450 200.830 198.520 ;
        RECT 175.700 197.670 175.990 197.830 ;
        RECT 177.080 197.820 177.340 197.880 ;
        RECT 120.060 197.610 134.220 197.620 ;
        RECT 120.060 197.600 127.590 197.610 ;
        RECT 128.600 197.600 129.790 197.610 ;
        RECT 130.750 197.600 131.940 197.610 ;
        RECT 133.030 197.600 134.220 197.610 ;
        RECT 120.060 197.590 125.370 197.600 ;
        RECT 120.060 197.580 124.230 197.590 ;
        RECT 120.060 197.570 121.950 197.580 ;
        RECT 123.040 197.570 124.230 197.580 ;
        RECT 120.060 197.560 120.780 197.570 ;
        RECT 116.690 197.210 117.000 197.550 ;
        RECT 112.700 196.680 114.340 197.070 ;
        RECT 115.140 196.920 117.000 197.210 ;
        RECT 115.140 196.910 115.450 196.920 ;
        RECT 116.690 196.910 117.000 196.920 ;
        RECT 105.280 196.560 105.930 196.570 ;
        RECT 105.280 196.230 105.580 196.560 ;
        RECT 104.560 195.780 105.580 196.230 ;
        RECT 110.170 196.070 110.460 196.670 ;
        RECT 112.060 196.070 112.350 196.670 ;
        RECT 105.280 195.770 105.580 195.780 ;
        RECT 114.400 195.460 114.700 196.460 ;
        RECT 115.150 195.860 115.450 196.910 ;
        RECT 117.750 195.810 118.000 197.550 ;
        RECT 175.200 197.480 175.990 197.670 ;
        RECT 175.200 197.280 175.450 197.480 ;
        RECT 175.700 197.370 175.990 197.480 ;
        RECT 177.090 197.280 177.340 197.820 ;
        RECT 180.170 197.820 180.440 197.880 ;
        RECT 181.720 198.160 183.030 198.420 ;
        RECT 185.170 198.200 200.830 198.450 ;
        RECT 185.170 198.170 185.990 198.200 ;
        RECT 181.720 197.820 182.030 198.160 ;
        RECT 177.730 197.290 179.370 197.680 ;
        RECT 180.170 197.530 182.030 197.820 ;
        RECT 180.170 197.520 180.480 197.530 ;
        RECT 181.720 197.520 182.030 197.530 ;
        RECT 118.450 195.460 118.710 197.010 ;
        RECT 175.200 196.680 175.490 197.280 ;
        RECT 177.090 196.680 177.380 197.280 ;
        RECT 179.430 196.070 179.730 197.070 ;
        RECT 180.180 196.470 180.480 197.520 ;
        RECT 182.780 196.420 183.030 198.160 ;
        RECT 200.580 197.990 200.830 198.200 ;
        RECT 183.480 196.070 183.740 197.620 ;
        RECT 200.580 196.150 200.850 197.990 ;
        RECT 184.440 196.070 184.620 196.080 ;
        RECT 179.380 195.770 184.630 196.070 ;
        RECT 114.350 195.450 119.600 195.460 ;
        RECT 104.230 195.370 104.480 195.380 ;
        RECT 104.230 194.910 105.210 195.370 ;
        RECT 114.350 195.160 119.620 195.450 ;
        RECT 104.230 194.610 104.480 194.910 ;
        RECT 112.200 194.820 114.040 194.830 ;
        RECT 119.450 194.820 119.620 195.160 ;
        RECT 105.940 194.810 106.180 194.820 ;
        RECT 107.020 194.810 119.620 194.820 ;
        RECT 105.940 194.650 119.620 194.810 ;
        RECT 105.940 194.640 117.450 194.650 ;
        RECT 105.930 194.630 112.250 194.640 ;
        RECT 113.800 194.630 117.450 194.640 ;
        RECT 105.930 194.620 107.800 194.630 ;
        RECT 105.930 194.610 106.180 194.620 ;
        RECT 104.230 194.440 106.180 194.610 ;
        RECT 104.230 194.140 104.500 194.440 ;
        RECT 104.240 193.880 104.500 194.140 ;
        RECT 104.220 193.490 104.520 193.880 ;
        RECT 104.210 193.090 104.520 193.490 ;
        RECT 104.200 192.330 104.510 193.090 ;
        RECT 104.100 192.310 104.510 192.330 ;
        RECT 104.070 191.360 104.520 192.310 ;
        RECT 104.930 191.070 105.390 192.010 ;
        RECT 106.130 191.420 115.400 191.430 ;
        RECT 117.280 191.420 119.200 191.430 ;
        RECT 106.130 191.230 119.200 191.420 ;
        RECT 106.130 191.220 118.490 191.230 ;
        RECT 104.970 190.750 105.270 191.070 ;
        RECT 104.970 190.420 105.260 190.750 ;
        RECT 104.980 189.620 105.240 190.420 ;
        RECT 106.130 190.210 106.340 191.220 ;
        RECT 115.390 191.210 117.290 191.220 ;
        RECT 119.020 190.480 119.200 191.230 ;
        RECT 104.980 189.020 105.230 189.620 ;
        RECT 106.130 189.200 106.330 190.210 ;
        RECT 113.940 190.180 119.200 190.480 ;
        RECT 104.190 188.570 105.230 189.020 ;
        RECT 104.170 187.120 105.130 187.570 ;
        RECT 104.880 187.070 105.130 187.120 ;
        RECT 106.140 187.070 106.330 189.200 ;
        RECT 104.880 186.870 106.330 187.070 ;
        RECT 109.860 188.540 110.120 189.740 ;
        RECT 109.860 188.030 110.110 188.540 ;
        RECT 111.750 188.530 112.010 189.740 ;
        RECT 114.140 188.630 114.390 190.180 ;
        RECT 111.750 188.370 112.140 188.530 ;
        RECT 111.740 188.240 112.140 188.370 ;
        RECT 114.840 188.240 115.100 189.850 ;
        RECT 117.390 188.780 117.690 189.830 ;
        RECT 118.140 189.230 118.440 190.180 ;
        RECT 118.640 189.280 118.940 189.330 ;
        RECT 118.640 188.930 119.540 189.280 ;
        RECT 121.250 189.150 121.470 189.160 ;
        RECT 121.250 188.960 134.930 189.150 ;
        RECT 121.250 188.830 121.470 188.960 ;
        RECT 110.360 188.030 110.650 188.190 ;
        RECT 111.740 188.180 112.000 188.240 ;
        RECT 109.860 187.840 110.650 188.030 ;
        RECT 109.860 187.640 110.110 187.840 ;
        RECT 110.360 187.730 110.650 187.840 ;
        RECT 111.750 187.640 112.000 188.180 ;
        RECT 114.830 188.180 115.100 188.240 ;
        RECT 116.380 188.520 117.690 188.780 ;
        RECT 119.790 188.530 121.470 188.830 ;
        RECT 119.790 188.520 121.450 188.530 ;
        RECT 116.380 188.180 116.690 188.520 ;
        RECT 112.390 187.650 114.030 188.040 ;
        RECT 114.830 187.890 116.690 188.180 ;
        RECT 114.830 187.880 115.140 187.890 ;
        RECT 116.380 187.880 116.690 187.890 ;
        RECT 109.860 187.040 110.150 187.640 ;
        RECT 111.750 187.040 112.040 187.640 ;
        RECT 104.880 186.780 105.130 186.870 ;
        RECT 104.150 186.330 105.130 186.780 ;
        RECT 114.090 186.430 114.390 187.430 ;
        RECT 114.840 186.830 115.140 187.880 ;
        RECT 117.440 186.780 117.690 188.520 ;
        RECT 134.680 188.060 134.930 188.960 ;
        RECT 118.140 186.430 118.400 187.980 ;
        RECT 129.620 187.760 134.930 188.060 ;
        RECT 114.040 186.410 119.290 186.430 ;
        RECT 114.040 186.130 119.410 186.410 ;
        RECT 107.490 185.730 107.770 185.800 ;
        RECT 108.670 185.760 108.950 185.790 ;
        RECT 119.120 185.760 119.410 186.130 ;
        RECT 108.670 185.750 119.410 185.760 ;
        RECT 106.080 185.530 107.770 185.730 ;
        RECT 104.870 185.330 105.150 185.340 ;
        RECT 104.130 184.880 105.150 185.330 ;
        RECT 106.080 184.880 106.310 185.530 ;
        RECT 107.490 185.470 107.770 185.530 ;
        RECT 108.650 185.520 119.410 185.750 ;
        RECT 108.670 185.510 119.410 185.520 ;
        RECT 125.540 186.120 125.800 187.320 ;
        RECT 125.540 185.610 125.790 186.120 ;
        RECT 127.430 186.110 127.690 187.320 ;
        RECT 129.820 186.210 130.070 187.760 ;
        RECT 127.430 185.950 127.820 186.110 ;
        RECT 127.420 185.820 127.820 185.950 ;
        RECT 130.520 185.820 130.780 187.430 ;
        RECT 133.070 186.360 133.370 187.410 ;
        RECT 133.820 186.810 134.120 187.760 ;
        RECT 134.320 186.860 134.620 186.910 ;
        RECT 134.320 186.510 135.220 186.860 ;
        RECT 147.980 186.460 152.450 186.490 ;
        RECT 137.040 186.430 152.450 186.460 ;
        RECT 136.370 186.410 152.450 186.430 ;
        RECT 126.040 185.610 126.330 185.770 ;
        RECT 127.420 185.760 127.680 185.820 ;
        RECT 108.670 185.500 119.370 185.510 ;
        RECT 108.670 185.460 108.950 185.500 ;
        RECT 125.540 185.420 126.330 185.610 ;
        RECT 125.540 185.220 125.790 185.420 ;
        RECT 126.040 185.310 126.330 185.420 ;
        RECT 127.430 185.220 127.680 185.760 ;
        RECT 130.510 185.760 130.780 185.820 ;
        RECT 132.060 186.100 133.370 186.360 ;
        RECT 132.060 185.760 132.370 186.100 ;
        RECT 128.070 185.230 129.710 185.620 ;
        RECT 130.510 185.470 132.370 185.760 ;
        RECT 130.510 185.460 130.820 185.470 ;
        RECT 132.060 185.460 132.370 185.470 ;
        RECT 107.470 184.900 107.740 184.980 ;
        RECT 104.870 184.670 106.310 184.880 ;
        RECT 106.860 184.680 107.740 184.900 ;
        RECT 104.870 183.620 105.150 184.670 ;
        RECT 106.860 183.870 107.080 184.680 ;
        RECT 107.470 184.650 107.740 184.680 ;
        RECT 108.600 184.940 108.890 184.990 ;
        RECT 108.600 184.760 119.350 184.940 ;
        RECT 108.600 184.660 108.890 184.760 ;
        RECT 113.440 184.750 117.070 184.760 ;
        RECT 119.150 184.080 119.350 184.760 ;
        RECT 125.540 184.620 125.830 185.220 ;
        RECT 127.430 184.620 127.720 185.220 ;
        RECT 104.150 183.170 105.150 183.620 ;
        RECT 104.130 181.720 105.430 182.170 ;
        RECT 105.130 181.320 105.430 181.720 ;
        RECT 106.850 181.340 107.080 183.870 ;
        RECT 114.100 183.780 119.350 184.080 ;
        RECT 129.770 184.010 130.070 185.010 ;
        RECT 130.520 184.410 130.820 185.460 ;
        RECT 133.120 184.360 133.370 186.100 ;
        RECT 135.490 186.090 152.450 186.410 ;
        RECT 184.440 186.110 184.620 195.770 ;
        RECT 136.370 186.080 152.450 186.090 ;
        RECT 136.370 186.050 148.350 186.080 ;
        RECT 136.370 186.040 137.260 186.050 ;
        RECT 133.820 184.010 134.080 185.560 ;
        RECT 134.910 184.010 135.110 184.020 ;
        RECT 105.920 181.320 107.080 181.340 ;
        RECT 105.130 181.140 107.080 181.320 ;
        RECT 110.020 182.140 110.280 183.340 ;
        RECT 110.020 181.630 110.270 182.140 ;
        RECT 111.910 182.130 112.170 183.340 ;
        RECT 114.300 182.230 114.550 183.780 ;
        RECT 111.910 181.970 112.300 182.130 ;
        RECT 111.900 181.840 112.300 181.970 ;
        RECT 115.000 181.840 115.260 183.450 ;
        RECT 117.550 182.380 117.850 183.430 ;
        RECT 118.300 182.830 118.600 183.780 ;
        RECT 119.150 183.770 119.350 183.780 ;
        RECT 129.720 183.710 135.110 184.010 ;
        RECT 118.800 182.880 119.100 182.930 ;
        RECT 118.800 182.530 119.700 182.880 ;
        RECT 134.910 182.470 135.110 183.710 ;
        RECT 152.070 182.510 152.430 186.080 ;
        RECT 127.350 182.450 128.540 182.460 ;
        RECT 129.530 182.450 130.720 182.460 ;
        RECT 131.750 182.450 132.940 182.460 ;
        RECT 133.930 182.450 135.120 182.470 ;
        RECT 125.140 182.440 135.120 182.450 ;
        RECT 121.750 182.420 122.940 182.430 ;
        RECT 124.030 182.420 135.120 182.440 ;
        RECT 110.520 181.630 110.810 181.790 ;
        RECT 111.900 181.780 112.160 181.840 ;
        RECT 110.020 181.440 110.810 181.630 ;
        RECT 110.020 181.240 110.270 181.440 ;
        RECT 110.520 181.330 110.810 181.440 ;
        RECT 111.910 181.240 112.160 181.780 ;
        RECT 114.990 181.780 115.260 181.840 ;
        RECT 116.540 182.120 117.850 182.380 ;
        RECT 119.910 182.190 135.120 182.420 ;
        RECT 147.200 182.210 152.450 182.510 ;
        RECT 119.910 182.180 134.070 182.190 ;
        RECT 119.910 182.170 127.440 182.180 ;
        RECT 128.450 182.170 129.640 182.180 ;
        RECT 130.600 182.170 131.790 182.180 ;
        RECT 132.880 182.170 134.070 182.180 ;
        RECT 119.910 182.160 125.220 182.170 ;
        RECT 119.910 182.150 124.080 182.160 ;
        RECT 119.910 182.140 121.800 182.150 ;
        RECT 122.890 182.140 124.080 182.150 ;
        RECT 119.910 182.130 120.630 182.140 ;
        RECT 116.540 181.780 116.850 182.120 ;
        RECT 112.550 181.250 114.190 181.640 ;
        RECT 114.990 181.490 116.850 181.780 ;
        RECT 114.990 181.480 115.300 181.490 ;
        RECT 116.540 181.480 116.850 181.490 ;
        RECT 105.130 181.130 105.780 181.140 ;
        RECT 105.130 180.800 105.430 181.130 ;
        RECT 104.410 180.350 105.430 180.800 ;
        RECT 110.020 180.640 110.310 181.240 ;
        RECT 111.910 180.640 112.200 181.240 ;
        RECT 105.130 180.340 105.430 180.350 ;
        RECT 114.250 180.030 114.550 181.030 ;
        RECT 115.000 180.430 115.300 181.480 ;
        RECT 117.600 180.380 117.850 182.120 ;
        RECT 118.300 180.030 118.560 181.580 ;
        RECT 143.120 180.570 143.380 181.770 ;
        RECT 143.120 180.060 143.370 180.570 ;
        RECT 145.010 180.560 145.270 181.770 ;
        RECT 147.400 180.660 147.650 182.210 ;
        RECT 145.010 180.400 145.400 180.560 ;
        RECT 145.000 180.270 145.400 180.400 ;
        RECT 148.100 180.270 148.360 181.880 ;
        RECT 150.650 180.810 150.950 181.860 ;
        RECT 151.400 181.260 151.700 182.210 ;
        RECT 151.900 181.310 152.200 181.360 ;
        RECT 151.900 180.960 152.800 181.310 ;
        RECT 143.620 180.060 143.910 180.220 ;
        RECT 145.000 180.210 145.260 180.270 ;
        RECT 114.200 180.020 119.450 180.030 ;
        RECT 104.080 179.940 104.330 179.950 ;
        RECT 104.080 179.480 105.060 179.940 ;
        RECT 114.200 179.730 119.470 180.020 ;
        RECT 104.080 179.180 104.330 179.480 ;
        RECT 112.050 179.390 113.890 179.400 ;
        RECT 119.300 179.390 119.470 179.730 ;
        RECT 105.790 179.380 106.030 179.390 ;
        RECT 106.870 179.380 119.470 179.390 ;
        RECT 105.790 179.220 119.470 179.380 ;
        RECT 143.120 179.870 143.910 180.060 ;
        RECT 143.120 179.670 143.370 179.870 ;
        RECT 143.620 179.760 143.910 179.870 ;
        RECT 145.010 179.670 145.260 180.210 ;
        RECT 148.090 180.210 148.360 180.270 ;
        RECT 149.640 180.550 150.950 180.810 ;
        RECT 153.010 180.850 154.680 180.880 ;
        RECT 169.760 180.850 170.010 180.860 ;
        RECT 153.010 180.580 170.010 180.850 ;
        RECT 153.010 180.570 166.510 180.580 ;
        RECT 154.290 180.550 166.510 180.570 ;
        RECT 149.640 180.210 149.950 180.550 ;
        RECT 145.650 179.680 147.290 180.070 ;
        RECT 148.090 179.920 149.950 180.210 ;
        RECT 148.090 179.910 148.400 179.920 ;
        RECT 149.640 179.910 149.950 179.920 ;
        RECT 105.790 179.210 117.300 179.220 ;
        RECT 105.780 179.200 112.100 179.210 ;
        RECT 113.650 179.200 117.300 179.210 ;
        RECT 105.780 179.190 107.650 179.200 ;
        RECT 105.780 179.180 106.030 179.190 ;
        RECT 104.080 179.010 106.030 179.180 ;
        RECT 143.120 179.070 143.410 179.670 ;
        RECT 145.010 179.070 145.300 179.670 ;
        RECT 104.080 178.790 104.330 179.010 ;
        RECT 104.080 178.620 105.120 178.790 ;
        RECT 104.930 177.760 105.120 178.620 ;
        RECT 147.350 178.460 147.650 179.460 ;
        RECT 148.100 178.860 148.400 179.910 ;
        RECT 150.700 178.810 150.950 180.550 ;
        RECT 151.400 178.460 151.660 180.010 ;
        RECT 152.280 178.460 152.620 178.530 ;
        RECT 147.300 178.160 152.620 178.460 ;
        RECT 104.140 177.320 105.120 177.760 ;
        RECT 104.140 177.310 105.090 177.320 ;
        RECT 105.960 177.000 115.230 177.010 ;
        RECT 117.110 177.000 119.030 177.010 ;
        RECT 103.810 176.900 104.000 176.910 ;
        RECT 103.810 176.440 104.790 176.900 ;
        RECT 105.960 176.810 119.030 177.000 ;
        RECT 105.960 176.800 118.320 176.810 ;
        RECT 103.810 175.650 104.000 176.440 ;
        RECT 105.960 175.790 106.170 176.800 ;
        RECT 115.220 176.790 117.120 176.800 ;
        RECT 118.850 176.060 119.030 176.810 ;
        RECT 104.810 175.650 105.080 175.660 ;
        RECT 103.810 175.440 105.080 175.650 ;
        RECT 104.810 175.230 105.080 175.440 ;
        RECT 104.810 174.600 105.060 175.230 ;
        RECT 105.960 174.780 106.160 175.790 ;
        RECT 113.770 175.760 119.030 176.060 ;
        RECT 104.020 174.150 105.060 174.600 ;
        RECT 104.000 172.700 104.960 173.150 ;
        RECT 104.710 172.650 104.960 172.700 ;
        RECT 105.970 172.650 106.160 174.780 ;
        RECT 104.710 172.450 106.160 172.650 ;
        RECT 109.690 174.120 109.950 175.320 ;
        RECT 109.690 173.610 109.940 174.120 ;
        RECT 111.580 174.110 111.840 175.320 ;
        RECT 113.970 174.210 114.220 175.760 ;
        RECT 111.580 173.950 111.970 174.110 ;
        RECT 111.570 173.820 111.970 173.950 ;
        RECT 114.670 173.820 114.930 175.430 ;
        RECT 117.220 174.360 117.520 175.410 ;
        RECT 117.970 174.810 118.270 175.760 ;
        RECT 118.470 174.860 118.770 174.910 ;
        RECT 118.470 174.510 119.370 174.860 ;
        RECT 121.080 174.730 121.300 174.740 ;
        RECT 121.080 174.540 134.760 174.730 ;
        RECT 121.080 174.410 121.300 174.540 ;
        RECT 110.190 173.610 110.480 173.770 ;
        RECT 111.570 173.760 111.830 173.820 ;
        RECT 109.690 173.420 110.480 173.610 ;
        RECT 109.690 173.220 109.940 173.420 ;
        RECT 110.190 173.310 110.480 173.420 ;
        RECT 111.580 173.220 111.830 173.760 ;
        RECT 114.660 173.760 114.930 173.820 ;
        RECT 116.210 174.100 117.520 174.360 ;
        RECT 119.620 174.110 121.300 174.410 ;
        RECT 119.620 174.100 121.280 174.110 ;
        RECT 116.210 173.760 116.520 174.100 ;
        RECT 112.220 173.230 113.860 173.620 ;
        RECT 114.660 173.470 116.520 173.760 ;
        RECT 114.660 173.460 114.970 173.470 ;
        RECT 116.210 173.460 116.520 173.470 ;
        RECT 109.690 172.620 109.980 173.220 ;
        RECT 111.580 172.620 111.870 173.220 ;
        RECT 104.710 172.360 104.960 172.450 ;
        RECT 103.980 171.910 104.960 172.360 ;
        RECT 113.920 172.010 114.220 173.010 ;
        RECT 114.670 172.410 114.970 173.460 ;
        RECT 117.270 172.360 117.520 174.100 ;
        RECT 134.510 173.640 134.760 174.540 ;
        RECT 117.970 172.010 118.230 173.560 ;
        RECT 129.450 173.340 134.760 173.640 ;
        RECT 113.870 171.990 119.120 172.010 ;
        RECT 113.870 171.710 119.240 171.990 ;
        RECT 107.320 171.310 107.600 171.380 ;
        RECT 108.500 171.340 108.780 171.370 ;
        RECT 118.950 171.340 119.240 171.710 ;
        RECT 108.500 171.330 119.240 171.340 ;
        RECT 105.910 171.110 107.600 171.310 ;
        RECT 104.700 170.910 104.980 170.920 ;
        RECT 103.960 170.460 104.980 170.910 ;
        RECT 105.910 170.460 106.140 171.110 ;
        RECT 107.320 171.050 107.600 171.110 ;
        RECT 108.480 171.100 119.240 171.330 ;
        RECT 108.500 171.090 119.240 171.100 ;
        RECT 125.370 171.700 125.630 172.900 ;
        RECT 125.370 171.190 125.620 171.700 ;
        RECT 127.260 171.690 127.520 172.900 ;
        RECT 129.650 171.790 129.900 173.340 ;
        RECT 127.260 171.530 127.650 171.690 ;
        RECT 127.250 171.400 127.650 171.530 ;
        RECT 130.350 171.400 130.610 173.010 ;
        RECT 132.900 171.940 133.200 172.990 ;
        RECT 133.650 172.390 133.950 173.340 ;
        RECT 134.150 172.440 134.450 172.490 ;
        RECT 134.150 172.090 135.050 172.440 ;
        RECT 152.280 172.040 152.620 178.160 ;
        RECT 151.710 172.020 152.670 172.040 ;
        RECT 136.190 172.000 140.470 172.010 ;
        RECT 147.870 172.000 152.670 172.020 ;
        RECT 136.190 171.990 152.670 172.000 ;
        RECT 125.870 171.190 126.160 171.350 ;
        RECT 127.250 171.340 127.510 171.400 ;
        RECT 108.500 171.080 119.200 171.090 ;
        RECT 108.500 171.040 108.780 171.080 ;
        RECT 125.370 171.000 126.160 171.190 ;
        RECT 125.370 170.800 125.620 171.000 ;
        RECT 125.870 170.890 126.160 171.000 ;
        RECT 127.260 170.800 127.510 171.340 ;
        RECT 130.340 171.340 130.610 171.400 ;
        RECT 131.890 171.680 133.200 171.940 ;
        RECT 131.890 171.340 132.200 171.680 ;
        RECT 127.900 170.810 129.540 171.200 ;
        RECT 130.340 171.050 132.200 171.340 ;
        RECT 130.340 171.040 130.650 171.050 ;
        RECT 131.890 171.040 132.200 171.050 ;
        RECT 107.300 170.480 107.570 170.560 ;
        RECT 104.700 170.250 106.140 170.460 ;
        RECT 106.690 170.260 107.570 170.480 ;
        RECT 104.700 169.200 104.980 170.250 ;
        RECT 106.690 169.450 106.910 170.260 ;
        RECT 107.300 170.230 107.570 170.260 ;
        RECT 108.430 170.520 108.720 170.570 ;
        RECT 108.430 170.340 119.180 170.520 ;
        RECT 108.430 170.240 108.720 170.340 ;
        RECT 113.270 170.330 116.900 170.340 ;
        RECT 118.980 169.660 119.180 170.340 ;
        RECT 125.370 170.200 125.660 170.800 ;
        RECT 127.260 170.200 127.550 170.800 ;
        RECT 103.980 168.750 104.980 169.200 ;
        RECT 103.960 167.300 105.260 167.750 ;
        RECT 104.960 166.900 105.260 167.300 ;
        RECT 106.680 166.920 106.910 169.450 ;
        RECT 113.930 169.360 119.180 169.660 ;
        RECT 129.600 169.590 129.900 170.590 ;
        RECT 130.350 169.990 130.650 171.040 ;
        RECT 132.950 169.940 133.200 171.680 ;
        RECT 135.320 171.680 152.670 171.990 ;
        RECT 135.320 171.670 148.330 171.680 ;
        RECT 140.180 171.660 148.330 171.670 ;
        RECT 151.710 171.640 152.670 171.680 ;
        RECT 152.280 171.630 152.620 171.640 ;
        RECT 133.650 169.590 133.910 171.140 ;
        RECT 134.740 169.590 134.940 169.600 ;
        RECT 105.750 166.900 106.910 166.920 ;
        RECT 104.960 166.720 106.910 166.900 ;
        RECT 109.850 167.720 110.110 168.920 ;
        RECT 109.850 167.210 110.100 167.720 ;
        RECT 111.740 167.710 112.000 168.920 ;
        RECT 114.130 167.810 114.380 169.360 ;
        RECT 111.740 167.550 112.130 167.710 ;
        RECT 111.730 167.420 112.130 167.550 ;
        RECT 114.830 167.420 115.090 169.030 ;
        RECT 117.380 167.960 117.680 169.010 ;
        RECT 118.130 168.410 118.430 169.360 ;
        RECT 118.980 169.350 119.180 169.360 ;
        RECT 129.550 169.290 134.940 169.590 ;
        RECT 118.630 168.460 118.930 168.510 ;
        RECT 118.630 168.110 119.530 168.460 ;
        RECT 134.740 168.050 134.940 169.290 ;
        RECT 127.180 168.030 128.370 168.040 ;
        RECT 129.360 168.030 130.550 168.040 ;
        RECT 131.580 168.030 132.770 168.040 ;
        RECT 133.760 168.030 134.950 168.050 ;
        RECT 124.970 168.020 134.950 168.030 ;
        RECT 121.580 168.000 122.770 168.010 ;
        RECT 123.860 168.000 134.950 168.020 ;
        RECT 110.350 167.210 110.640 167.370 ;
        RECT 111.730 167.360 111.990 167.420 ;
        RECT 109.850 167.020 110.640 167.210 ;
        RECT 109.850 166.820 110.100 167.020 ;
        RECT 110.350 166.910 110.640 167.020 ;
        RECT 111.740 166.820 111.990 167.360 ;
        RECT 114.820 167.360 115.090 167.420 ;
        RECT 116.370 167.700 117.680 167.960 ;
        RECT 119.740 167.770 134.950 168.000 ;
        RECT 119.740 167.760 133.900 167.770 ;
        RECT 119.740 167.750 127.270 167.760 ;
        RECT 128.280 167.750 129.470 167.760 ;
        RECT 130.430 167.750 131.620 167.760 ;
        RECT 132.710 167.750 133.900 167.760 ;
        RECT 119.740 167.740 125.050 167.750 ;
        RECT 119.740 167.730 123.910 167.740 ;
        RECT 119.740 167.720 121.630 167.730 ;
        RECT 122.720 167.720 123.910 167.730 ;
        RECT 119.740 167.710 120.460 167.720 ;
        RECT 116.370 167.360 116.680 167.700 ;
        RECT 112.380 166.830 114.020 167.220 ;
        RECT 114.820 167.070 116.680 167.360 ;
        RECT 114.820 167.060 115.130 167.070 ;
        RECT 116.370 167.060 116.680 167.070 ;
        RECT 104.960 166.710 105.610 166.720 ;
        RECT 104.960 166.380 105.260 166.710 ;
        RECT 100.850 166.000 101.110 166.180 ;
        RECT 99.310 158.640 99.540 160.610 ;
        RECT 99.310 156.750 99.560 158.640 ;
        RECT 99.310 154.950 99.580 156.750 ;
        RECT 51.670 150.690 68.830 150.980 ;
        RECT 52.360 150.680 68.830 150.690 ;
        RECT 48.300 150.330 48.610 150.670 ;
        RECT 44.310 149.800 45.950 150.190 ;
        RECT 46.750 150.040 48.610 150.330 ;
        RECT 46.750 150.030 47.060 150.040 ;
        RECT 48.300 150.030 48.610 150.040 ;
        RECT 4.450 149.330 15.960 149.340 ;
        RECT 4.440 149.320 10.760 149.330 ;
        RECT 12.310 149.320 15.960 149.330 ;
        RECT 4.440 149.310 6.310 149.320 ;
        RECT 4.440 149.300 4.690 149.310 ;
        RECT 2.740 149.130 4.690 149.300 ;
        RECT 41.780 149.190 42.070 149.790 ;
        RECT 43.670 149.190 43.960 149.790 ;
        RECT 2.740 148.910 2.990 149.130 ;
        RECT 2.740 148.740 3.780 148.910 ;
        RECT 3.590 147.880 3.780 148.740 ;
        RECT 46.010 148.580 46.310 149.580 ;
        RECT 46.760 148.980 47.060 150.030 ;
        RECT 49.360 148.930 49.610 150.670 ;
        RECT 50.060 148.580 50.320 150.130 ;
        RECT 99.310 149.710 99.600 154.950 ;
        RECT 50.940 148.580 51.280 148.650 ;
        RECT 45.960 148.280 51.280 148.580 ;
        RECT 2.800 147.440 3.780 147.880 ;
        RECT 2.800 147.430 3.750 147.440 ;
        RECT 4.620 147.120 13.890 147.130 ;
        RECT 15.770 147.120 17.690 147.130 ;
        RECT 2.470 147.020 2.660 147.030 ;
        RECT 2.470 146.560 3.450 147.020 ;
        RECT 4.620 146.930 17.690 147.120 ;
        RECT 4.620 146.920 16.980 146.930 ;
        RECT 2.470 145.770 2.660 146.560 ;
        RECT 4.620 145.910 4.830 146.920 ;
        RECT 13.880 146.910 15.780 146.920 ;
        RECT 17.510 146.180 17.690 146.930 ;
        RECT 3.470 145.770 3.740 145.780 ;
        RECT 2.470 145.560 3.740 145.770 ;
        RECT 3.470 145.350 3.740 145.560 ;
        RECT 3.470 144.720 3.720 145.350 ;
        RECT 4.620 144.900 4.820 145.910 ;
        RECT 12.430 145.880 17.690 146.180 ;
        RECT 2.680 144.270 3.720 144.720 ;
        RECT 2.660 142.820 3.620 143.270 ;
        RECT 3.370 142.770 3.620 142.820 ;
        RECT 4.630 142.770 4.820 144.900 ;
        RECT 3.370 142.570 4.820 142.770 ;
        RECT 8.350 144.240 8.610 145.440 ;
        RECT 8.350 143.730 8.600 144.240 ;
        RECT 10.240 144.230 10.500 145.440 ;
        RECT 12.630 144.330 12.880 145.880 ;
        RECT 10.240 144.070 10.630 144.230 ;
        RECT 10.230 143.940 10.630 144.070 ;
        RECT 13.330 143.940 13.590 145.550 ;
        RECT 15.880 144.480 16.180 145.530 ;
        RECT 16.630 144.930 16.930 145.880 ;
        RECT 17.130 144.980 17.430 145.030 ;
        RECT 17.130 144.630 18.030 144.980 ;
        RECT 19.740 144.850 19.960 144.860 ;
        RECT 19.740 144.660 33.420 144.850 ;
        RECT 19.740 144.530 19.960 144.660 ;
        RECT 8.850 143.730 9.140 143.890 ;
        RECT 10.230 143.880 10.490 143.940 ;
        RECT 8.350 143.540 9.140 143.730 ;
        RECT 8.350 143.340 8.600 143.540 ;
        RECT 8.850 143.430 9.140 143.540 ;
        RECT 10.240 143.340 10.490 143.880 ;
        RECT 13.320 143.880 13.590 143.940 ;
        RECT 14.870 144.220 16.180 144.480 ;
        RECT 18.280 144.230 19.960 144.530 ;
        RECT 18.280 144.220 19.940 144.230 ;
        RECT 14.870 143.880 15.180 144.220 ;
        RECT 10.880 143.350 12.520 143.740 ;
        RECT 13.320 143.590 15.180 143.880 ;
        RECT 13.320 143.580 13.630 143.590 ;
        RECT 14.870 143.580 15.180 143.590 ;
        RECT 8.350 142.740 8.640 143.340 ;
        RECT 10.240 142.740 10.530 143.340 ;
        RECT 3.370 142.480 3.620 142.570 ;
        RECT 2.640 142.030 3.620 142.480 ;
        RECT 12.580 142.130 12.880 143.130 ;
        RECT 13.330 142.530 13.630 143.580 ;
        RECT 15.930 142.480 16.180 144.220 ;
        RECT 33.170 143.760 33.420 144.660 ;
        RECT 16.630 142.130 16.890 143.680 ;
        RECT 28.110 143.460 33.420 143.760 ;
        RECT 12.530 142.110 17.780 142.130 ;
        RECT 12.530 141.830 17.900 142.110 ;
        RECT 5.980 141.430 6.260 141.500 ;
        RECT 7.160 141.460 7.440 141.490 ;
        RECT 17.610 141.460 17.900 141.830 ;
        RECT 7.160 141.450 17.900 141.460 ;
        RECT 4.570 141.230 6.260 141.430 ;
        RECT 3.360 141.030 3.640 141.040 ;
        RECT 2.620 140.580 3.640 141.030 ;
        RECT 4.570 140.580 4.800 141.230 ;
        RECT 5.980 141.170 6.260 141.230 ;
        RECT 7.140 141.220 17.900 141.450 ;
        RECT 7.160 141.210 17.900 141.220 ;
        RECT 24.030 141.820 24.290 143.020 ;
        RECT 24.030 141.310 24.280 141.820 ;
        RECT 25.920 141.810 26.180 143.020 ;
        RECT 28.310 141.910 28.560 143.460 ;
        RECT 25.920 141.650 26.310 141.810 ;
        RECT 25.910 141.520 26.310 141.650 ;
        RECT 29.010 141.520 29.270 143.130 ;
        RECT 31.560 142.060 31.860 143.110 ;
        RECT 32.310 142.510 32.610 143.460 ;
        RECT 32.810 142.560 33.110 142.610 ;
        RECT 32.810 142.210 33.710 142.560 ;
        RECT 50.940 142.160 51.280 148.280 ;
        RECT 99.310 147.740 99.540 149.710 ;
        RECT 100.870 149.200 101.110 166.000 ;
        RECT 104.240 165.930 105.260 166.380 ;
        RECT 109.850 166.220 110.140 166.820 ;
        RECT 111.740 166.220 112.030 166.820 ;
        RECT 104.960 165.920 105.260 165.930 ;
        RECT 114.080 165.610 114.380 166.610 ;
        RECT 114.830 166.010 115.130 167.060 ;
        RECT 117.430 165.960 117.680 167.700 ;
        RECT 169.760 167.440 170.020 180.580 ;
        RECT 169.750 167.320 170.020 167.440 ;
        RECT 184.350 176.590 184.620 186.110 ;
        RECT 200.580 192.480 200.890 196.150 ;
        RECT 200.580 190.700 200.910 192.480 ;
        RECT 200.580 188.730 200.870 190.700 ;
        RECT 200.580 186.900 200.890 188.730 ;
        RECT 200.580 183.080 200.870 186.900 ;
        RECT 200.580 181.110 200.850 183.080 ;
        RECT 200.580 179.390 200.910 181.110 ;
        RECT 200.580 177.470 200.870 179.390 ;
        RECT 118.130 165.610 118.390 167.160 ;
        RECT 169.750 166.490 170.010 167.320 ;
        RECT 184.350 166.640 184.530 176.590 ;
        RECT 200.580 167.930 200.850 177.470 ;
        RECT 164.730 166.190 170.010 166.490 ;
        RECT 114.030 165.600 119.280 165.610 ;
        RECT 103.910 165.520 104.160 165.530 ;
        RECT 103.910 165.060 104.890 165.520 ;
        RECT 114.030 165.310 119.300 165.600 ;
        RECT 103.910 164.760 104.160 165.060 ;
        RECT 111.880 164.970 113.720 164.980 ;
        RECT 119.130 164.970 119.300 165.310 ;
        RECT 105.620 164.960 105.860 164.970 ;
        RECT 106.700 164.960 119.300 164.970 ;
        RECT 105.620 164.800 119.300 164.960 ;
        RECT 105.620 164.790 117.130 164.800 ;
        RECT 105.610 164.780 111.930 164.790 ;
        RECT 113.480 164.780 117.130 164.790 ;
        RECT 105.610 164.770 107.480 164.780 ;
        RECT 105.610 164.760 105.860 164.770 ;
        RECT 103.910 164.590 105.860 164.760 ;
        RECT 103.910 164.290 104.180 164.590 ;
        RECT 103.920 164.030 104.180 164.290 ;
        RECT 160.650 164.550 160.910 165.750 ;
        RECT 160.650 164.040 160.900 164.550 ;
        RECT 162.540 164.540 162.800 165.750 ;
        RECT 164.930 164.640 165.180 166.190 ;
        RECT 162.540 164.380 162.930 164.540 ;
        RECT 162.530 164.250 162.930 164.380 ;
        RECT 165.630 164.250 165.890 165.860 ;
        RECT 168.180 164.790 168.480 165.840 ;
        RECT 168.930 165.240 169.230 166.190 ;
        RECT 169.430 165.290 169.730 165.340 ;
        RECT 169.430 164.940 170.330 165.290 ;
        RECT 184.340 164.830 184.540 166.640 ;
        RECT 161.150 164.040 161.440 164.200 ;
        RECT 162.530 164.190 162.790 164.250 ;
        RECT 103.900 163.640 104.200 164.030 ;
        RECT 160.650 163.850 161.440 164.040 ;
        RECT 160.650 163.650 160.900 163.850 ;
        RECT 161.150 163.740 161.440 163.850 ;
        RECT 162.540 163.650 162.790 164.190 ;
        RECT 165.620 164.190 165.890 164.250 ;
        RECT 167.170 164.530 168.480 164.790 ;
        RECT 170.600 164.540 184.540 164.830 ;
        RECT 200.620 166.060 200.890 167.930 ;
        RECT 170.600 164.530 184.500 164.540 ;
        RECT 167.170 164.190 167.480 164.530 ;
        RECT 163.180 163.660 164.820 164.050 ;
        RECT 165.620 163.900 167.480 164.190 ;
        RECT 165.620 163.890 165.930 163.900 ;
        RECT 167.170 163.890 167.480 163.900 ;
        RECT 103.900 163.410 105.390 163.640 ;
        RECT 105.140 162.480 105.390 163.410 ;
        RECT 160.650 163.050 160.940 163.650 ;
        RECT 162.540 163.050 162.830 163.650 ;
        RECT 104.340 162.020 105.390 162.480 ;
        RECT 164.880 162.440 165.180 163.440 ;
        RECT 165.630 162.840 165.930 163.890 ;
        RECT 168.230 162.790 168.480 164.530 ;
        RECT 171.190 164.520 184.500 164.530 ;
        RECT 168.930 162.440 169.190 163.990 ;
        RECT 164.830 162.140 170.100 162.440 ;
        RECT 105.140 162.010 105.390 162.020 ;
        RECT 104.010 161.610 104.260 161.620 ;
        RECT 104.010 161.160 104.990 161.610 ;
        RECT 106.100 161.350 115.370 161.360 ;
        RECT 117.250 161.350 119.170 161.360 ;
        RECT 106.100 161.160 119.170 161.350 ;
        RECT 104.010 160.550 104.260 161.160 ;
        RECT 106.100 161.150 118.460 161.160 ;
        RECT 104.010 160.300 105.220 160.550 ;
        RECT 104.950 159.550 105.210 160.300 ;
        RECT 106.100 160.140 106.310 161.150 ;
        RECT 115.360 161.140 117.260 161.150 ;
        RECT 118.990 160.410 119.170 161.160 ;
        RECT 104.950 158.950 105.200 159.550 ;
        RECT 106.100 159.130 106.300 160.140 ;
        RECT 113.910 160.110 119.170 160.410 ;
        RECT 104.160 158.500 105.200 158.950 ;
        RECT 104.140 157.050 105.100 157.500 ;
        RECT 104.850 157.000 105.100 157.050 ;
        RECT 106.110 157.000 106.300 159.130 ;
        RECT 104.850 156.800 106.300 157.000 ;
        RECT 109.830 158.470 110.090 159.670 ;
        RECT 109.830 157.960 110.080 158.470 ;
        RECT 111.720 158.460 111.980 159.670 ;
        RECT 114.110 158.560 114.360 160.110 ;
        RECT 111.720 158.300 112.110 158.460 ;
        RECT 111.710 158.170 112.110 158.300 ;
        RECT 114.810 158.170 115.070 159.780 ;
        RECT 117.360 158.710 117.660 159.760 ;
        RECT 118.110 159.160 118.410 160.110 ;
        RECT 118.610 159.210 118.910 159.260 ;
        RECT 118.610 158.860 119.510 159.210 ;
        RECT 121.220 159.080 121.440 159.090 ;
        RECT 121.220 158.890 134.900 159.080 ;
        RECT 121.220 158.760 121.440 158.890 ;
        RECT 110.330 157.960 110.620 158.120 ;
        RECT 111.710 158.110 111.970 158.170 ;
        RECT 109.830 157.770 110.620 157.960 ;
        RECT 109.830 157.570 110.080 157.770 ;
        RECT 110.330 157.660 110.620 157.770 ;
        RECT 111.720 157.570 111.970 158.110 ;
        RECT 114.800 158.110 115.070 158.170 ;
        RECT 116.350 158.450 117.660 158.710 ;
        RECT 119.760 158.460 121.440 158.760 ;
        RECT 119.760 158.450 121.420 158.460 ;
        RECT 116.350 158.110 116.660 158.450 ;
        RECT 112.360 157.580 114.000 157.970 ;
        RECT 114.800 157.820 116.660 158.110 ;
        RECT 114.800 157.810 115.110 157.820 ;
        RECT 116.350 157.810 116.660 157.820 ;
        RECT 109.830 156.970 110.120 157.570 ;
        RECT 111.720 156.970 112.010 157.570 ;
        RECT 104.850 156.710 105.100 156.800 ;
        RECT 104.120 156.260 105.100 156.710 ;
        RECT 114.060 156.360 114.360 157.360 ;
        RECT 114.810 156.760 115.110 157.810 ;
        RECT 117.410 156.710 117.660 158.450 ;
        RECT 134.650 157.990 134.900 158.890 ;
        RECT 118.110 156.360 118.370 157.910 ;
        RECT 129.590 157.690 134.900 157.990 ;
        RECT 114.010 156.340 119.260 156.360 ;
        RECT 114.010 156.060 119.380 156.340 ;
        RECT 107.460 155.660 107.740 155.730 ;
        RECT 108.640 155.690 108.920 155.720 ;
        RECT 119.090 155.690 119.380 156.060 ;
        RECT 108.640 155.680 119.380 155.690 ;
        RECT 106.050 155.460 107.740 155.660 ;
        RECT 104.840 155.260 105.120 155.270 ;
        RECT 104.100 154.810 105.120 155.260 ;
        RECT 106.050 154.810 106.280 155.460 ;
        RECT 107.460 155.400 107.740 155.460 ;
        RECT 108.620 155.450 119.380 155.680 ;
        RECT 108.640 155.440 119.380 155.450 ;
        RECT 125.510 156.050 125.770 157.250 ;
        RECT 125.510 155.540 125.760 156.050 ;
        RECT 127.400 156.040 127.660 157.250 ;
        RECT 129.790 156.140 130.040 157.690 ;
        RECT 127.400 155.880 127.790 156.040 ;
        RECT 127.390 155.750 127.790 155.880 ;
        RECT 130.490 155.750 130.750 157.360 ;
        RECT 133.040 156.290 133.340 157.340 ;
        RECT 133.790 156.740 134.090 157.690 ;
        RECT 134.290 156.790 134.590 156.840 ;
        RECT 134.290 156.440 135.190 156.790 ;
        RECT 147.950 156.390 152.420 156.420 ;
        RECT 137.010 156.360 152.420 156.390 ;
        RECT 136.340 156.340 152.420 156.360 ;
        RECT 126.010 155.540 126.300 155.700 ;
        RECT 127.390 155.690 127.650 155.750 ;
        RECT 108.640 155.430 119.340 155.440 ;
        RECT 108.640 155.390 108.920 155.430 ;
        RECT 125.510 155.350 126.300 155.540 ;
        RECT 125.510 155.150 125.760 155.350 ;
        RECT 126.010 155.240 126.300 155.350 ;
        RECT 127.400 155.150 127.650 155.690 ;
        RECT 130.480 155.690 130.750 155.750 ;
        RECT 132.030 156.030 133.340 156.290 ;
        RECT 132.030 155.690 132.340 156.030 ;
        RECT 128.040 155.160 129.680 155.550 ;
        RECT 130.480 155.400 132.340 155.690 ;
        RECT 130.480 155.390 130.790 155.400 ;
        RECT 132.030 155.390 132.340 155.400 ;
        RECT 107.440 154.830 107.710 154.910 ;
        RECT 104.840 154.600 106.280 154.810 ;
        RECT 106.830 154.610 107.710 154.830 ;
        RECT 104.840 153.550 105.120 154.600 ;
        RECT 106.830 153.800 107.050 154.610 ;
        RECT 107.440 154.580 107.710 154.610 ;
        RECT 108.570 154.870 108.860 154.920 ;
        RECT 108.570 154.690 119.320 154.870 ;
        RECT 108.570 154.590 108.860 154.690 ;
        RECT 113.410 154.680 117.040 154.690 ;
        RECT 119.120 154.010 119.320 154.690 ;
        RECT 125.510 154.550 125.800 155.150 ;
        RECT 127.400 154.550 127.690 155.150 ;
        RECT 104.120 153.100 105.120 153.550 ;
        RECT 104.100 151.650 105.400 152.100 ;
        RECT 105.100 151.250 105.400 151.650 ;
        RECT 106.820 151.270 107.050 153.800 ;
        RECT 114.070 153.710 119.320 154.010 ;
        RECT 129.740 153.940 130.040 154.940 ;
        RECT 130.490 154.340 130.790 155.390 ;
        RECT 133.090 154.290 133.340 156.030 ;
        RECT 135.460 156.020 152.420 156.340 ;
        RECT 136.340 156.010 152.420 156.020 ;
        RECT 136.340 155.980 148.320 156.010 ;
        RECT 136.340 155.970 137.230 155.980 ;
        RECT 133.790 153.940 134.050 155.490 ;
        RECT 134.880 153.940 135.080 153.950 ;
        RECT 105.890 151.250 107.050 151.270 ;
        RECT 105.100 151.070 107.050 151.250 ;
        RECT 109.990 152.070 110.250 153.270 ;
        RECT 109.990 151.560 110.240 152.070 ;
        RECT 111.880 152.060 112.140 153.270 ;
        RECT 114.270 152.160 114.520 153.710 ;
        RECT 111.880 151.900 112.270 152.060 ;
        RECT 111.870 151.770 112.270 151.900 ;
        RECT 114.970 151.770 115.230 153.380 ;
        RECT 117.520 152.310 117.820 153.360 ;
        RECT 118.270 152.760 118.570 153.710 ;
        RECT 119.120 153.700 119.320 153.710 ;
        RECT 129.690 153.640 135.080 153.940 ;
        RECT 118.770 152.810 119.070 152.860 ;
        RECT 118.770 152.460 119.670 152.810 ;
        RECT 134.880 152.400 135.080 153.640 ;
        RECT 152.040 152.440 152.400 156.010 ;
        RECT 127.320 152.380 128.510 152.390 ;
        RECT 129.500 152.380 130.690 152.390 ;
        RECT 131.720 152.380 132.910 152.390 ;
        RECT 133.900 152.380 135.090 152.400 ;
        RECT 125.110 152.370 135.090 152.380 ;
        RECT 121.720 152.350 122.910 152.360 ;
        RECT 124.000 152.350 135.090 152.370 ;
        RECT 110.490 151.560 110.780 151.720 ;
        RECT 111.870 151.710 112.130 151.770 ;
        RECT 109.990 151.370 110.780 151.560 ;
        RECT 109.990 151.170 110.240 151.370 ;
        RECT 110.490 151.260 110.780 151.370 ;
        RECT 111.880 151.170 112.130 151.710 ;
        RECT 114.960 151.710 115.230 151.770 ;
        RECT 116.510 152.050 117.820 152.310 ;
        RECT 119.880 152.120 135.090 152.350 ;
        RECT 147.170 152.140 152.420 152.440 ;
        RECT 119.880 152.110 134.040 152.120 ;
        RECT 119.880 152.100 127.410 152.110 ;
        RECT 128.420 152.100 129.610 152.110 ;
        RECT 130.570 152.100 131.760 152.110 ;
        RECT 132.850 152.100 134.040 152.110 ;
        RECT 119.880 152.090 125.190 152.100 ;
        RECT 119.880 152.080 124.050 152.090 ;
        RECT 119.880 152.070 121.770 152.080 ;
        RECT 122.860 152.070 124.050 152.080 ;
        RECT 119.880 152.060 120.600 152.070 ;
        RECT 116.510 151.710 116.820 152.050 ;
        RECT 112.520 151.180 114.160 151.570 ;
        RECT 114.960 151.420 116.820 151.710 ;
        RECT 114.960 151.410 115.270 151.420 ;
        RECT 116.510 151.410 116.820 151.420 ;
        RECT 105.100 151.060 105.750 151.070 ;
        RECT 105.100 150.730 105.400 151.060 ;
        RECT 104.380 150.280 105.400 150.730 ;
        RECT 109.990 150.570 110.280 151.170 ;
        RECT 111.880 150.570 112.170 151.170 ;
        RECT 105.100 150.270 105.400 150.280 ;
        RECT 114.220 149.960 114.520 150.960 ;
        RECT 114.970 150.360 115.270 151.410 ;
        RECT 117.570 150.310 117.820 152.050 ;
        RECT 118.270 149.960 118.530 151.510 ;
        RECT 143.090 150.500 143.350 151.700 ;
        RECT 143.090 149.990 143.340 150.500 ;
        RECT 144.980 150.490 145.240 151.700 ;
        RECT 147.370 150.590 147.620 152.140 ;
        RECT 144.980 150.330 145.370 150.490 ;
        RECT 144.970 150.200 145.370 150.330 ;
        RECT 148.070 150.200 148.330 151.810 ;
        RECT 150.620 150.740 150.920 151.790 ;
        RECT 151.370 151.190 151.670 152.140 ;
        RECT 151.870 151.240 152.170 151.290 ;
        RECT 151.870 150.890 152.770 151.240 ;
        RECT 143.590 149.990 143.880 150.150 ;
        RECT 144.970 150.140 145.230 150.200 ;
        RECT 114.170 149.950 119.420 149.960 ;
        RECT 100.840 148.990 101.110 149.200 ;
        RECT 104.050 149.870 104.300 149.880 ;
        RECT 104.050 149.410 105.030 149.870 ;
        RECT 114.170 149.660 119.440 149.950 ;
        RECT 104.050 149.110 104.300 149.410 ;
        RECT 112.020 149.320 113.860 149.330 ;
        RECT 119.270 149.320 119.440 149.660 ;
        RECT 105.760 149.310 106.000 149.320 ;
        RECT 106.840 149.310 119.440 149.320 ;
        RECT 105.760 149.150 119.440 149.310 ;
        RECT 143.090 149.800 143.880 149.990 ;
        RECT 143.090 149.600 143.340 149.800 ;
        RECT 143.590 149.690 143.880 149.800 ;
        RECT 144.980 149.600 145.230 150.140 ;
        RECT 148.060 150.140 148.330 150.200 ;
        RECT 149.610 150.480 150.920 150.740 ;
        RECT 152.980 150.790 154.650 150.810 ;
        RECT 169.790 150.790 170.100 162.140 ;
        RECT 200.620 160.420 200.870 166.060 ;
        RECT 200.620 158.450 200.850 160.420 ;
        RECT 200.620 156.560 200.870 158.450 ;
        RECT 200.620 154.760 200.890 156.560 ;
        RECT 152.980 150.500 170.140 150.790 ;
        RECT 153.670 150.490 170.140 150.500 ;
        RECT 149.610 150.140 149.920 150.480 ;
        RECT 145.620 149.610 147.260 150.000 ;
        RECT 148.060 149.850 149.920 150.140 ;
        RECT 148.060 149.840 148.370 149.850 ;
        RECT 149.610 149.840 149.920 149.850 ;
        RECT 105.760 149.140 117.270 149.150 ;
        RECT 105.750 149.130 112.070 149.140 ;
        RECT 113.620 149.130 117.270 149.140 ;
        RECT 105.750 149.120 107.620 149.130 ;
        RECT 105.750 149.110 106.000 149.120 ;
        RECT 99.310 144.150 99.580 147.740 ;
        RECT 100.840 145.760 101.080 148.990 ;
        RECT 104.050 148.940 106.000 149.110 ;
        RECT 143.090 149.000 143.380 149.600 ;
        RECT 144.980 149.000 145.270 149.600 ;
        RECT 104.050 148.720 104.300 148.940 ;
        RECT 104.050 148.550 105.090 148.720 ;
        RECT 104.900 147.690 105.090 148.550 ;
        RECT 147.320 148.390 147.620 149.390 ;
        RECT 148.070 148.790 148.370 149.840 ;
        RECT 150.670 148.740 150.920 150.480 ;
        RECT 151.370 148.390 151.630 149.940 ;
        RECT 200.620 149.520 200.910 154.760 ;
        RECT 152.250 148.390 152.590 148.460 ;
        RECT 147.270 148.090 152.590 148.390 ;
        RECT 104.110 147.250 105.090 147.690 ;
        RECT 104.110 147.240 105.060 147.250 ;
        RECT 105.930 146.930 115.200 146.940 ;
        RECT 117.080 146.930 119.000 146.940 ;
        RECT 103.780 146.830 103.970 146.840 ;
        RECT 103.780 146.370 104.760 146.830 ;
        RECT 105.930 146.740 119.000 146.930 ;
        RECT 105.930 146.730 118.290 146.740 ;
        RECT 100.840 145.590 101.090 145.760 ;
        RECT 99.310 142.330 99.560 144.150 ;
        RECT 50.370 142.140 51.330 142.160 ;
        RECT 34.850 142.120 39.130 142.130 ;
        RECT 46.530 142.120 51.330 142.140 ;
        RECT 34.850 142.110 51.330 142.120 ;
        RECT 24.530 141.310 24.820 141.470 ;
        RECT 25.910 141.460 26.170 141.520 ;
        RECT 7.160 141.200 17.860 141.210 ;
        RECT 7.160 141.160 7.440 141.200 ;
        RECT 24.030 141.120 24.820 141.310 ;
        RECT 24.030 140.920 24.280 141.120 ;
        RECT 24.530 141.010 24.820 141.120 ;
        RECT 25.920 140.920 26.170 141.460 ;
        RECT 29.000 141.460 29.270 141.520 ;
        RECT 30.550 141.800 31.860 142.060 ;
        RECT 30.550 141.460 30.860 141.800 ;
        RECT 26.560 140.930 28.200 141.320 ;
        RECT 29.000 141.170 30.860 141.460 ;
        RECT 29.000 141.160 29.310 141.170 ;
        RECT 30.550 141.160 30.860 141.170 ;
        RECT 5.960 140.600 6.230 140.680 ;
        RECT 3.360 140.370 4.800 140.580 ;
        RECT 5.350 140.380 6.230 140.600 ;
        RECT 3.360 139.320 3.640 140.370 ;
        RECT 5.350 139.570 5.570 140.380 ;
        RECT 5.960 140.350 6.230 140.380 ;
        RECT 7.090 140.640 7.380 140.690 ;
        RECT 7.090 140.460 17.840 140.640 ;
        RECT 7.090 140.360 7.380 140.460 ;
        RECT 11.930 140.450 15.560 140.460 ;
        RECT 17.640 139.780 17.840 140.460 ;
        RECT 24.030 140.320 24.320 140.920 ;
        RECT 25.920 140.320 26.210 140.920 ;
        RECT 2.640 138.870 3.640 139.320 ;
        RECT 2.620 137.420 3.920 137.870 ;
        RECT 3.620 137.020 3.920 137.420 ;
        RECT 5.340 137.040 5.570 139.570 ;
        RECT 12.590 139.480 17.840 139.780 ;
        RECT 28.260 139.710 28.560 140.710 ;
        RECT 29.010 140.110 29.310 141.160 ;
        RECT 31.610 140.060 31.860 141.800 ;
        RECT 33.980 141.800 51.330 142.110 ;
        RECT 33.980 141.790 46.990 141.800 ;
        RECT 38.840 141.780 46.990 141.790 ;
        RECT 50.370 141.760 51.330 141.800 ;
        RECT 50.940 141.750 51.280 141.760 ;
        RECT 32.310 139.710 32.570 141.260 ;
        RECT 33.400 139.710 33.600 139.720 ;
        RECT 4.410 137.020 5.570 137.040 ;
        RECT 3.620 136.840 5.570 137.020 ;
        RECT 8.510 137.840 8.770 139.040 ;
        RECT 8.510 137.330 8.760 137.840 ;
        RECT 10.400 137.830 10.660 139.040 ;
        RECT 12.790 137.930 13.040 139.480 ;
        RECT 10.400 137.670 10.790 137.830 ;
        RECT 10.390 137.540 10.790 137.670 ;
        RECT 13.490 137.540 13.750 139.150 ;
        RECT 16.040 138.080 16.340 139.130 ;
        RECT 16.790 138.530 17.090 139.480 ;
        RECT 17.640 139.470 17.840 139.480 ;
        RECT 28.210 139.410 33.600 139.710 ;
        RECT 17.290 138.580 17.590 138.630 ;
        RECT 17.290 138.230 18.190 138.580 ;
        RECT 33.400 138.170 33.600 139.410 ;
        RECT 99.310 138.870 99.540 142.330 ;
        RECT 100.850 142.300 101.090 145.590 ;
        RECT 103.780 145.580 103.970 146.370 ;
        RECT 105.930 145.720 106.140 146.730 ;
        RECT 115.190 146.720 117.090 146.730 ;
        RECT 118.820 145.990 119.000 146.740 ;
        RECT 104.780 145.580 105.050 145.590 ;
        RECT 103.780 145.370 105.050 145.580 ;
        RECT 104.780 145.160 105.050 145.370 ;
        RECT 104.780 144.530 105.030 145.160 ;
        RECT 105.930 144.710 106.130 145.720 ;
        RECT 113.740 145.690 119.000 145.990 ;
        RECT 103.990 144.080 105.030 144.530 ;
        RECT 103.970 142.630 104.930 143.080 ;
        RECT 104.680 142.580 104.930 142.630 ;
        RECT 105.940 142.580 106.130 144.710 ;
        RECT 104.680 142.380 106.130 142.580 ;
        RECT 109.660 144.050 109.920 145.250 ;
        RECT 109.660 143.540 109.910 144.050 ;
        RECT 111.550 144.040 111.810 145.250 ;
        RECT 113.940 144.140 114.190 145.690 ;
        RECT 111.550 143.880 111.940 144.040 ;
        RECT 111.540 143.750 111.940 143.880 ;
        RECT 114.640 143.750 114.900 145.360 ;
        RECT 117.190 144.290 117.490 145.340 ;
        RECT 117.940 144.740 118.240 145.690 ;
        RECT 118.440 144.790 118.740 144.840 ;
        RECT 118.440 144.440 119.340 144.790 ;
        RECT 121.050 144.660 121.270 144.670 ;
        RECT 121.050 144.470 134.730 144.660 ;
        RECT 121.050 144.340 121.270 144.470 ;
        RECT 110.160 143.540 110.450 143.700 ;
        RECT 111.540 143.690 111.800 143.750 ;
        RECT 109.660 143.350 110.450 143.540 ;
        RECT 109.660 143.150 109.910 143.350 ;
        RECT 110.160 143.240 110.450 143.350 ;
        RECT 111.550 143.150 111.800 143.690 ;
        RECT 114.630 143.690 114.900 143.750 ;
        RECT 116.180 144.030 117.490 144.290 ;
        RECT 119.590 144.040 121.270 144.340 ;
        RECT 119.590 144.030 121.250 144.040 ;
        RECT 116.180 143.690 116.490 144.030 ;
        RECT 112.190 143.160 113.830 143.550 ;
        RECT 114.630 143.400 116.490 143.690 ;
        RECT 114.630 143.390 114.940 143.400 ;
        RECT 116.180 143.390 116.490 143.400 ;
        RECT 109.660 142.550 109.950 143.150 ;
        RECT 111.550 142.550 111.840 143.150 ;
        RECT 100.850 142.150 101.110 142.300 ;
        RECT 104.680 142.290 104.930 142.380 ;
        RECT 99.270 138.460 99.540 138.870 ;
        RECT 25.840 138.150 27.030 138.160 ;
        RECT 28.020 138.150 29.210 138.160 ;
        RECT 30.240 138.150 31.430 138.160 ;
        RECT 32.420 138.150 33.610 138.170 ;
        RECT 23.630 138.140 33.610 138.150 ;
        RECT 20.240 138.120 21.430 138.130 ;
        RECT 22.520 138.120 33.610 138.140 ;
        RECT 9.010 137.330 9.300 137.490 ;
        RECT 10.390 137.480 10.650 137.540 ;
        RECT 8.510 137.140 9.300 137.330 ;
        RECT 8.510 136.940 8.760 137.140 ;
        RECT 9.010 137.030 9.300 137.140 ;
        RECT 10.400 136.940 10.650 137.480 ;
        RECT 13.480 137.480 13.750 137.540 ;
        RECT 15.030 137.820 16.340 138.080 ;
        RECT 18.400 137.890 33.610 138.120 ;
        RECT 18.400 137.880 32.560 137.890 ;
        RECT 18.400 137.870 25.930 137.880 ;
        RECT 26.940 137.870 28.130 137.880 ;
        RECT 29.090 137.870 30.280 137.880 ;
        RECT 31.370 137.870 32.560 137.880 ;
        RECT 18.400 137.860 23.710 137.870 ;
        RECT 18.400 137.850 22.570 137.860 ;
        RECT 18.400 137.840 20.290 137.850 ;
        RECT 21.380 137.840 22.570 137.850 ;
        RECT 18.400 137.830 19.120 137.840 ;
        RECT 15.030 137.480 15.340 137.820 ;
        RECT 11.040 136.950 12.680 137.340 ;
        RECT 13.480 137.190 15.340 137.480 ;
        RECT 13.480 137.180 13.790 137.190 ;
        RECT 15.030 137.180 15.340 137.190 ;
        RECT 3.620 136.830 4.270 136.840 ;
        RECT 3.620 136.500 3.920 136.830 ;
        RECT 2.900 136.050 3.920 136.500 ;
        RECT 8.510 136.340 8.800 136.940 ;
        RECT 10.400 136.340 10.690 136.940 ;
        RECT 3.620 136.040 3.920 136.050 ;
        RECT 12.740 135.730 13.040 136.730 ;
        RECT 13.490 136.130 13.790 137.180 ;
        RECT 16.090 136.080 16.340 137.820 ;
        RECT 16.790 135.730 17.050 137.280 ;
        RECT 99.270 137.170 99.520 138.460 ;
        RECT 94.300 136.870 99.550 137.170 ;
        RECT 12.690 135.720 17.940 135.730 ;
        RECT 2.570 135.640 2.820 135.650 ;
        RECT 2.570 135.180 3.550 135.640 ;
        RECT 12.690 135.430 17.960 135.720 ;
        RECT 2.570 134.880 2.820 135.180 ;
        RECT 10.540 135.090 12.380 135.100 ;
        RECT 17.790 135.090 17.960 135.430 ;
        RECT 4.280 135.080 4.520 135.090 ;
        RECT 5.360 135.080 17.960 135.090 ;
        RECT 4.280 134.920 17.960 135.080 ;
        RECT 90.220 135.230 90.480 136.430 ;
        RECT 4.280 134.910 15.790 134.920 ;
        RECT 4.270 134.900 10.590 134.910 ;
        RECT 12.140 134.900 15.790 134.910 ;
        RECT 4.270 134.890 6.140 134.900 ;
        RECT 4.270 134.880 4.520 134.890 ;
        RECT 2.570 134.710 4.520 134.880 ;
        RECT 90.220 134.720 90.470 135.230 ;
        RECT 92.110 135.220 92.370 136.430 ;
        RECT 94.500 135.320 94.750 136.870 ;
        RECT 92.110 135.060 92.500 135.220 ;
        RECT 92.100 134.930 92.500 135.060 ;
        RECT 95.200 134.930 95.460 136.540 ;
        RECT 97.750 135.470 98.050 136.520 ;
        RECT 98.500 135.920 98.800 136.870 ;
        RECT 99.000 135.970 99.300 136.020 ;
        RECT 99.000 135.620 99.900 135.970 ;
        RECT 100.870 135.520 101.110 142.150 ;
        RECT 103.950 141.840 104.930 142.290 ;
        RECT 113.890 141.940 114.190 142.940 ;
        RECT 114.640 142.340 114.940 143.390 ;
        RECT 117.240 142.290 117.490 144.030 ;
        RECT 134.480 143.570 134.730 144.470 ;
        RECT 117.940 141.940 118.200 143.490 ;
        RECT 129.420 143.270 134.730 143.570 ;
        RECT 113.840 141.920 119.090 141.940 ;
        RECT 113.840 141.640 119.210 141.920 ;
        RECT 107.290 141.240 107.570 141.310 ;
        RECT 108.470 141.270 108.750 141.300 ;
        RECT 118.920 141.270 119.210 141.640 ;
        RECT 108.470 141.260 119.210 141.270 ;
        RECT 105.880 141.040 107.570 141.240 ;
        RECT 104.670 140.840 104.950 140.850 ;
        RECT 103.930 140.390 104.950 140.840 ;
        RECT 105.880 140.390 106.110 141.040 ;
        RECT 107.290 140.980 107.570 141.040 ;
        RECT 108.450 141.030 119.210 141.260 ;
        RECT 108.470 141.020 119.210 141.030 ;
        RECT 125.340 141.630 125.600 142.830 ;
        RECT 125.340 141.120 125.590 141.630 ;
        RECT 127.230 141.620 127.490 142.830 ;
        RECT 129.620 141.720 129.870 143.270 ;
        RECT 127.230 141.460 127.620 141.620 ;
        RECT 127.220 141.330 127.620 141.460 ;
        RECT 130.320 141.330 130.580 142.940 ;
        RECT 132.870 141.870 133.170 142.920 ;
        RECT 133.620 142.320 133.920 143.270 ;
        RECT 134.120 142.370 134.420 142.420 ;
        RECT 134.120 142.020 135.020 142.370 ;
        RECT 152.250 141.970 152.590 148.090 ;
        RECT 200.620 147.550 200.850 149.520 ;
        RECT 200.620 143.960 200.890 147.550 ;
        RECT 200.620 142.140 200.870 143.960 ;
        RECT 226.840 143.480 227.110 242.980 ;
        RECT 226.840 143.300 227.160 143.480 ;
        RECT 151.680 141.950 152.640 141.970 ;
        RECT 136.160 141.930 140.440 141.940 ;
        RECT 147.840 141.930 152.640 141.950 ;
        RECT 136.160 141.920 152.640 141.930 ;
        RECT 125.840 141.120 126.130 141.280 ;
        RECT 127.220 141.270 127.480 141.330 ;
        RECT 108.470 141.010 119.170 141.020 ;
        RECT 108.470 140.970 108.750 141.010 ;
        RECT 125.340 140.930 126.130 141.120 ;
        RECT 125.340 140.730 125.590 140.930 ;
        RECT 125.840 140.820 126.130 140.930 ;
        RECT 127.230 140.730 127.480 141.270 ;
        RECT 130.310 141.270 130.580 141.330 ;
        RECT 131.860 141.610 133.170 141.870 ;
        RECT 131.860 141.270 132.170 141.610 ;
        RECT 127.870 140.740 129.510 141.130 ;
        RECT 130.310 140.980 132.170 141.270 ;
        RECT 130.310 140.970 130.620 140.980 ;
        RECT 131.860 140.970 132.170 140.980 ;
        RECT 107.270 140.410 107.540 140.490 ;
        RECT 104.670 140.180 106.110 140.390 ;
        RECT 106.660 140.190 107.540 140.410 ;
        RECT 104.670 139.130 104.950 140.180 ;
        RECT 106.660 139.380 106.880 140.190 ;
        RECT 107.270 140.160 107.540 140.190 ;
        RECT 108.400 140.450 108.690 140.500 ;
        RECT 108.400 140.270 119.150 140.450 ;
        RECT 108.400 140.170 108.690 140.270 ;
        RECT 113.240 140.260 116.870 140.270 ;
        RECT 118.950 139.590 119.150 140.270 ;
        RECT 125.340 140.130 125.630 140.730 ;
        RECT 127.230 140.130 127.520 140.730 ;
        RECT 103.950 138.680 104.950 139.130 ;
        RECT 103.930 137.230 105.230 137.680 ;
        RECT 104.930 136.830 105.230 137.230 ;
        RECT 106.650 136.850 106.880 139.380 ;
        RECT 113.900 139.290 119.150 139.590 ;
        RECT 129.570 139.520 129.870 140.520 ;
        RECT 130.320 139.920 130.620 140.970 ;
        RECT 132.920 139.870 133.170 141.610 ;
        RECT 135.290 141.610 152.640 141.920 ;
        RECT 135.290 141.600 148.300 141.610 ;
        RECT 140.150 141.590 148.300 141.600 ;
        RECT 151.680 141.570 152.640 141.610 ;
        RECT 152.250 141.560 152.590 141.570 ;
        RECT 133.620 139.520 133.880 141.070 ;
        RECT 134.710 139.520 134.910 139.530 ;
        RECT 105.720 136.830 106.880 136.850 ;
        RECT 104.930 136.650 106.880 136.830 ;
        RECT 109.820 137.650 110.080 138.850 ;
        RECT 109.820 137.140 110.070 137.650 ;
        RECT 111.710 137.640 111.970 138.850 ;
        RECT 114.100 137.740 114.350 139.290 ;
        RECT 111.710 137.480 112.100 137.640 ;
        RECT 111.700 137.350 112.100 137.480 ;
        RECT 114.800 137.350 115.060 138.960 ;
        RECT 117.350 137.890 117.650 138.940 ;
        RECT 118.100 138.340 118.400 139.290 ;
        RECT 118.950 139.280 119.150 139.290 ;
        RECT 129.520 139.220 134.910 139.520 ;
        RECT 118.600 138.390 118.900 138.440 ;
        RECT 118.600 138.040 119.500 138.390 ;
        RECT 134.710 137.980 134.910 139.220 ;
        RECT 200.620 138.680 200.850 142.140 ;
        RECT 226.860 140.800 227.160 143.300 ;
        RECT 226.870 139.310 227.140 140.800 ;
        RECT 221.890 139.010 227.140 139.310 ;
        RECT 200.580 138.270 200.850 138.680 ;
        RECT 127.150 137.960 128.340 137.970 ;
        RECT 129.330 137.960 130.520 137.970 ;
        RECT 131.550 137.960 132.740 137.970 ;
        RECT 133.730 137.960 134.920 137.980 ;
        RECT 124.940 137.950 134.920 137.960 ;
        RECT 121.550 137.930 122.740 137.940 ;
        RECT 123.830 137.930 134.920 137.950 ;
        RECT 110.320 137.140 110.610 137.300 ;
        RECT 111.700 137.290 111.960 137.350 ;
        RECT 109.820 136.950 110.610 137.140 ;
        RECT 109.820 136.750 110.070 136.950 ;
        RECT 110.320 136.840 110.610 136.950 ;
        RECT 111.710 136.750 111.960 137.290 ;
        RECT 114.790 137.290 115.060 137.350 ;
        RECT 116.340 137.630 117.650 137.890 ;
        RECT 119.710 137.700 134.920 137.930 ;
        RECT 119.710 137.690 133.870 137.700 ;
        RECT 119.710 137.680 127.240 137.690 ;
        RECT 128.250 137.680 129.440 137.690 ;
        RECT 130.400 137.680 131.590 137.690 ;
        RECT 132.680 137.680 133.870 137.690 ;
        RECT 119.710 137.670 125.020 137.680 ;
        RECT 119.710 137.660 123.880 137.670 ;
        RECT 119.710 137.650 121.600 137.660 ;
        RECT 122.690 137.650 123.880 137.660 ;
        RECT 119.710 137.640 120.430 137.650 ;
        RECT 116.340 137.290 116.650 137.630 ;
        RECT 112.350 136.760 113.990 137.150 ;
        RECT 114.790 137.000 116.650 137.290 ;
        RECT 114.790 136.990 115.100 137.000 ;
        RECT 116.340 136.990 116.650 137.000 ;
        RECT 104.930 136.640 105.580 136.650 ;
        RECT 104.930 136.310 105.230 136.640 ;
        RECT 104.210 135.860 105.230 136.310 ;
        RECT 109.820 136.150 110.110 136.750 ;
        RECT 111.710 136.150 112.000 136.750 ;
        RECT 104.930 135.850 105.230 135.860 ;
        RECT 114.050 135.540 114.350 136.540 ;
        RECT 114.800 135.940 115.100 136.990 ;
        RECT 117.400 135.890 117.650 137.630 ;
        RECT 118.100 135.540 118.360 137.090 ;
        RECT 200.580 136.980 200.830 138.270 ;
        RECT 217.810 137.370 218.070 138.570 ;
        RECT 195.610 136.680 200.860 136.980 ;
        RECT 217.810 136.860 218.060 137.370 ;
        RECT 219.700 137.360 219.960 138.570 ;
        RECT 222.090 137.460 222.340 139.010 ;
        RECT 226.090 138.060 226.390 139.010 ;
        RECT 226.590 138.110 226.890 138.160 ;
        RECT 226.590 137.760 227.490 138.110 ;
        RECT 219.700 137.200 220.090 137.360 ;
        RECT 219.690 137.070 220.090 137.200 ;
        RECT 218.310 136.860 218.600 137.020 ;
        RECT 219.690 137.010 219.950 137.070 ;
        RECT 90.720 134.720 91.010 134.880 ;
        RECT 92.100 134.870 92.360 134.930 ;
        RECT 2.570 134.410 2.840 134.710 ;
        RECT 2.580 134.150 2.840 134.410 ;
        RECT 90.220 134.530 91.010 134.720 ;
        RECT 90.220 134.330 90.470 134.530 ;
        RECT 90.720 134.420 91.010 134.530 ;
        RECT 92.110 134.330 92.360 134.870 ;
        RECT 95.190 134.870 95.460 134.930 ;
        RECT 96.740 135.210 98.050 135.470 ;
        RECT 100.230 135.210 101.110 135.520 ;
        RECT 114.000 135.530 119.250 135.540 ;
        RECT 103.880 135.450 104.130 135.460 ;
        RECT 96.740 134.870 97.050 135.210 ;
        RECT 92.750 134.340 94.390 134.730 ;
        RECT 95.190 134.580 97.050 134.870 ;
        RECT 95.190 134.570 95.500 134.580 ;
        RECT 96.740 134.570 97.050 134.580 ;
        RECT 2.560 133.760 2.860 134.150 ;
        RECT 2.550 133.360 2.860 133.760 ;
        RECT 90.220 133.730 90.510 134.330 ;
        RECT 92.110 133.730 92.400 134.330 ;
        RECT 2.550 133.030 2.840 133.360 ;
        RECT 94.450 133.120 94.750 134.120 ;
        RECT 95.200 133.520 95.500 134.570 ;
        RECT 97.800 133.470 98.050 135.210 ;
        RECT 103.880 134.990 104.860 135.450 ;
        RECT 114.000 135.240 119.270 135.530 ;
        RECT 103.880 134.690 104.130 134.990 ;
        RECT 111.850 134.900 113.690 134.910 ;
        RECT 119.100 134.900 119.270 135.240 ;
        RECT 105.590 134.890 105.830 134.900 ;
        RECT 106.670 134.890 119.270 134.900 ;
        RECT 105.590 134.730 119.270 134.890 ;
        RECT 191.530 135.040 191.790 136.240 ;
        RECT 105.590 134.720 117.100 134.730 ;
        RECT 105.580 134.710 111.900 134.720 ;
        RECT 113.450 134.710 117.100 134.720 ;
        RECT 105.580 134.700 107.450 134.710 ;
        RECT 105.580 134.690 105.830 134.700 ;
        RECT 98.500 133.120 98.760 134.670 ;
        RECT 103.880 134.520 105.830 134.690 ;
        RECT 191.530 134.530 191.780 135.040 ;
        RECT 193.420 135.030 193.680 136.240 ;
        RECT 195.810 135.130 196.060 136.680 ;
        RECT 193.420 134.870 193.810 135.030 ;
        RECT 193.410 134.740 193.810 134.870 ;
        RECT 196.510 134.740 196.770 136.350 ;
        RECT 199.060 135.280 199.360 136.330 ;
        RECT 199.810 135.730 200.110 136.680 ;
        RECT 217.810 136.670 218.600 136.860 ;
        RECT 217.810 136.470 218.060 136.670 ;
        RECT 218.310 136.560 218.600 136.670 ;
        RECT 219.700 136.470 219.950 137.010 ;
        RECT 220.340 136.480 221.980 136.870 ;
        RECT 217.810 135.870 218.100 136.470 ;
        RECT 219.700 135.870 219.990 136.470 ;
        RECT 200.310 135.780 200.610 135.830 ;
        RECT 200.310 135.430 201.210 135.780 ;
        RECT 209.280 135.330 213.110 135.350 ;
        RECT 192.030 134.530 192.320 134.690 ;
        RECT 193.410 134.680 193.670 134.740 ;
        RECT 103.880 134.220 104.150 134.520 ;
        RECT 103.890 133.960 104.150 134.220 ;
        RECT 191.530 134.340 192.320 134.530 ;
        RECT 191.530 134.140 191.780 134.340 ;
        RECT 192.030 134.230 192.320 134.340 ;
        RECT 193.420 134.140 193.670 134.680 ;
        RECT 196.500 134.680 196.770 134.740 ;
        RECT 198.050 135.020 199.360 135.280 ;
        RECT 201.540 135.050 213.120 135.330 ;
        RECT 222.040 135.260 222.340 136.260 ;
        RECT 226.090 135.260 226.350 136.810 ;
        RECT 227.140 135.260 227.340 135.290 ;
        RECT 201.540 135.030 209.730 135.050 ;
        RECT 201.540 135.020 202.370 135.030 ;
        RECT 198.050 134.680 198.360 135.020 ;
        RECT 194.060 134.150 195.700 134.540 ;
        RECT 196.500 134.390 198.360 134.680 ;
        RECT 196.500 134.380 196.810 134.390 ;
        RECT 198.050 134.380 198.360 134.390 ;
        RECT 103.870 133.570 104.170 133.960 ;
        RECT 103.860 133.170 104.170 133.570 ;
        RECT 191.530 133.540 191.820 134.140 ;
        RECT 193.420 133.540 193.710 134.140 ;
        RECT 99.590 133.120 100.140 133.140 ;
        RECT 2.530 132.370 2.880 133.030 ;
        RECT 94.400 132.830 100.140 133.120 ;
        RECT 103.860 132.840 104.150 133.170 ;
        RECT 195.760 132.930 196.060 133.930 ;
        RECT 196.510 133.330 196.810 134.380 ;
        RECT 199.110 133.280 199.360 135.020 ;
        RECT 199.810 132.930 200.070 134.480 ;
        RECT 212.920 133.090 213.120 135.050 ;
        RECT 221.990 134.960 227.340 135.260 ;
        RECT 227.140 133.110 227.340 134.960 ;
        RECT 220.680 133.090 227.370 133.110 ;
        RECT 200.900 132.930 201.450 132.950 ;
        RECT 94.400 132.820 99.650 132.830 ;
        RECT 1.260 132.030 2.880 132.370 ;
        RECT 1.260 131.180 1.710 132.030 ;
        RECT 2.530 132.020 2.880 132.030 ;
        RECT 2.120 131.000 2.580 131.830 ;
        RECT 4.670 131.290 13.940 131.300 ;
        RECT 15.820 131.290 17.740 131.300 ;
        RECT 3.500 131.000 3.780 131.140 ;
        RECT 2.120 130.890 3.780 131.000 ;
        RECT 2.130 130.690 3.780 130.890 ;
        RECT 4.670 131.100 17.740 131.290 ;
        RECT 4.670 131.090 17.030 131.100 ;
        RECT 2.130 130.680 3.800 130.690 ;
        RECT 3.500 130.460 3.800 130.680 ;
        RECT 3.510 130.290 3.800 130.460 ;
        RECT 3.520 129.490 3.780 130.290 ;
        RECT 4.670 130.080 4.880 131.090 ;
        RECT 13.930 131.080 15.830 131.090 ;
        RECT 17.560 130.350 17.740 131.100 ;
        RECT 3.520 128.890 3.770 129.490 ;
        RECT 4.670 129.070 4.870 130.080 ;
        RECT 12.480 130.050 17.740 130.350 ;
        RECT 2.730 128.440 3.770 128.890 ;
        RECT 2.710 126.990 3.670 127.440 ;
        RECT 3.420 126.940 3.670 126.990 ;
        RECT 4.680 126.940 4.870 129.070 ;
        RECT 3.420 126.740 4.870 126.940 ;
        RECT 8.400 128.410 8.660 129.610 ;
        RECT 8.400 127.900 8.650 128.410 ;
        RECT 10.290 128.400 10.550 129.610 ;
        RECT 12.680 128.500 12.930 130.050 ;
        RECT 10.290 128.240 10.680 128.400 ;
        RECT 10.280 128.110 10.680 128.240 ;
        RECT 13.380 128.110 13.640 129.720 ;
        RECT 15.930 128.650 16.230 129.700 ;
        RECT 16.680 129.100 16.980 130.050 ;
        RECT 17.180 129.150 17.480 129.200 ;
        RECT 17.180 128.800 18.080 129.150 ;
        RECT 19.790 129.020 20.010 129.030 ;
        RECT 19.790 128.830 33.470 129.020 ;
        RECT 19.790 128.700 20.010 128.830 ;
        RECT 8.900 127.900 9.190 128.060 ;
        RECT 10.280 128.050 10.540 128.110 ;
        RECT 8.400 127.710 9.190 127.900 ;
        RECT 8.400 127.510 8.650 127.710 ;
        RECT 8.900 127.600 9.190 127.710 ;
        RECT 10.290 127.510 10.540 128.050 ;
        RECT 13.370 128.050 13.640 128.110 ;
        RECT 14.920 128.390 16.230 128.650 ;
        RECT 18.330 128.400 20.010 128.700 ;
        RECT 18.330 128.390 19.990 128.400 ;
        RECT 14.920 128.050 15.230 128.390 ;
        RECT 10.930 127.520 12.570 127.910 ;
        RECT 13.370 127.760 15.230 128.050 ;
        RECT 13.370 127.750 13.680 127.760 ;
        RECT 14.920 127.750 15.230 127.760 ;
        RECT 8.400 126.910 8.690 127.510 ;
        RECT 10.290 126.910 10.580 127.510 ;
        RECT 3.420 126.650 3.670 126.740 ;
        RECT 2.690 126.200 3.670 126.650 ;
        RECT 12.630 126.300 12.930 127.300 ;
        RECT 13.380 126.700 13.680 127.750 ;
        RECT 15.980 126.650 16.230 128.390 ;
        RECT 33.220 127.930 33.470 128.830 ;
        RECT 16.680 126.300 16.940 127.850 ;
        RECT 28.160 127.630 33.470 127.930 ;
        RECT 12.580 126.280 17.830 126.300 ;
        RECT 12.580 126.000 17.950 126.280 ;
        RECT 6.030 125.600 6.310 125.670 ;
        RECT 7.210 125.630 7.490 125.660 ;
        RECT 17.660 125.630 17.950 126.000 ;
        RECT 7.210 125.620 17.950 125.630 ;
        RECT 4.620 125.400 6.310 125.600 ;
        RECT 3.410 125.200 3.690 125.210 ;
        RECT 2.670 124.750 3.690 125.200 ;
        RECT 4.620 124.750 4.850 125.400 ;
        RECT 6.030 125.340 6.310 125.400 ;
        RECT 7.190 125.390 17.950 125.620 ;
        RECT 7.210 125.380 17.950 125.390 ;
        RECT 24.080 125.990 24.340 127.190 ;
        RECT 24.080 125.480 24.330 125.990 ;
        RECT 25.970 125.980 26.230 127.190 ;
        RECT 28.360 126.080 28.610 127.630 ;
        RECT 25.970 125.820 26.360 125.980 ;
        RECT 25.960 125.690 26.360 125.820 ;
        RECT 29.060 125.690 29.320 127.300 ;
        RECT 31.610 126.230 31.910 127.280 ;
        RECT 32.360 126.680 32.660 127.630 ;
        RECT 32.860 126.730 33.160 126.780 ;
        RECT 32.860 126.380 33.760 126.730 ;
        RECT 46.520 126.330 50.990 126.360 ;
        RECT 35.580 126.300 50.990 126.330 ;
        RECT 34.910 126.280 50.990 126.300 ;
        RECT 24.580 125.480 24.870 125.640 ;
        RECT 25.960 125.630 26.220 125.690 ;
        RECT 7.210 125.370 17.910 125.380 ;
        RECT 7.210 125.330 7.490 125.370 ;
        RECT 24.080 125.290 24.870 125.480 ;
        RECT 24.080 125.090 24.330 125.290 ;
        RECT 24.580 125.180 24.870 125.290 ;
        RECT 25.970 125.090 26.220 125.630 ;
        RECT 29.050 125.630 29.320 125.690 ;
        RECT 30.600 125.970 31.910 126.230 ;
        RECT 30.600 125.630 30.910 125.970 ;
        RECT 26.610 125.100 28.250 125.490 ;
        RECT 29.050 125.340 30.910 125.630 ;
        RECT 29.050 125.330 29.360 125.340 ;
        RECT 30.600 125.330 30.910 125.340 ;
        RECT 6.010 124.770 6.280 124.850 ;
        RECT 3.410 124.540 4.850 124.750 ;
        RECT 5.400 124.550 6.280 124.770 ;
        RECT 3.410 123.490 3.690 124.540 ;
        RECT 5.400 123.740 5.620 124.550 ;
        RECT 6.010 124.520 6.280 124.550 ;
        RECT 7.140 124.810 7.430 124.860 ;
        RECT 7.140 124.630 17.890 124.810 ;
        RECT 7.140 124.530 7.430 124.630 ;
        RECT 11.980 124.620 15.610 124.630 ;
        RECT 17.690 123.950 17.890 124.630 ;
        RECT 24.080 124.490 24.370 125.090 ;
        RECT 25.970 124.490 26.260 125.090 ;
        RECT 2.690 123.040 3.690 123.490 ;
        RECT 2.670 121.590 3.970 122.040 ;
        RECT 3.670 121.190 3.970 121.590 ;
        RECT 5.390 121.210 5.620 123.740 ;
        RECT 12.640 123.650 17.890 123.950 ;
        RECT 28.310 123.880 28.610 124.880 ;
        RECT 29.060 124.280 29.360 125.330 ;
        RECT 31.660 124.230 31.910 125.970 ;
        RECT 34.030 125.960 50.990 126.280 ;
        RECT 34.910 125.950 50.990 125.960 ;
        RECT 34.910 125.920 46.890 125.950 ;
        RECT 34.910 125.910 35.800 125.920 ;
        RECT 32.360 123.880 32.620 125.430 ;
        RECT 33.450 123.880 33.650 123.890 ;
        RECT 4.460 121.190 5.620 121.210 ;
        RECT 3.670 121.010 5.620 121.190 ;
        RECT 8.560 122.010 8.820 123.210 ;
        RECT 8.560 121.500 8.810 122.010 ;
        RECT 10.450 122.000 10.710 123.210 ;
        RECT 12.840 122.100 13.090 123.650 ;
        RECT 10.450 121.840 10.840 122.000 ;
        RECT 10.440 121.710 10.840 121.840 ;
        RECT 13.540 121.710 13.800 123.320 ;
        RECT 16.090 122.250 16.390 123.300 ;
        RECT 16.840 122.700 17.140 123.650 ;
        RECT 17.690 123.640 17.890 123.650 ;
        RECT 28.260 123.580 33.650 123.880 ;
        RECT 17.340 122.750 17.640 122.800 ;
        RECT 17.340 122.400 18.240 122.750 ;
        RECT 33.450 122.340 33.650 123.580 ;
        RECT 50.610 122.380 50.970 125.950 ;
        RECT 25.890 122.320 27.080 122.330 ;
        RECT 28.070 122.320 29.260 122.330 ;
        RECT 30.290 122.320 31.480 122.330 ;
        RECT 32.470 122.320 33.660 122.340 ;
        RECT 23.680 122.310 33.660 122.320 ;
        RECT 20.290 122.290 21.480 122.300 ;
        RECT 22.570 122.290 33.660 122.310 ;
        RECT 9.060 121.500 9.350 121.660 ;
        RECT 10.440 121.650 10.700 121.710 ;
        RECT 8.560 121.310 9.350 121.500 ;
        RECT 8.560 121.110 8.810 121.310 ;
        RECT 9.060 121.200 9.350 121.310 ;
        RECT 10.450 121.110 10.700 121.650 ;
        RECT 13.530 121.650 13.800 121.710 ;
        RECT 15.080 121.990 16.390 122.250 ;
        RECT 18.450 122.060 33.660 122.290 ;
        RECT 45.740 122.080 50.990 122.380 ;
        RECT 18.450 122.050 32.610 122.060 ;
        RECT 18.450 122.040 25.980 122.050 ;
        RECT 26.990 122.040 28.180 122.050 ;
        RECT 29.140 122.040 30.330 122.050 ;
        RECT 31.420 122.040 32.610 122.050 ;
        RECT 18.450 122.030 23.760 122.040 ;
        RECT 18.450 122.020 22.620 122.030 ;
        RECT 18.450 122.010 20.340 122.020 ;
        RECT 21.430 122.010 22.620 122.020 ;
        RECT 18.450 122.000 19.170 122.010 ;
        RECT 15.080 121.650 15.390 121.990 ;
        RECT 11.090 121.120 12.730 121.510 ;
        RECT 13.530 121.360 15.390 121.650 ;
        RECT 13.530 121.350 13.840 121.360 ;
        RECT 15.080 121.350 15.390 121.360 ;
        RECT 3.670 121.000 4.320 121.010 ;
        RECT 3.670 120.670 3.970 121.000 ;
        RECT 2.950 120.220 3.970 120.670 ;
        RECT 8.560 120.510 8.850 121.110 ;
        RECT 10.450 120.510 10.740 121.110 ;
        RECT 3.670 120.210 3.970 120.220 ;
        RECT 12.790 119.900 13.090 120.900 ;
        RECT 13.540 120.300 13.840 121.350 ;
        RECT 16.140 120.250 16.390 121.990 ;
        RECT 16.840 119.900 17.100 121.450 ;
        RECT 41.660 120.440 41.920 121.640 ;
        RECT 41.660 119.930 41.910 120.440 ;
        RECT 43.550 120.430 43.810 121.640 ;
        RECT 45.940 120.530 46.190 122.080 ;
        RECT 43.550 120.270 43.940 120.430 ;
        RECT 43.540 120.140 43.940 120.270 ;
        RECT 46.640 120.140 46.900 121.750 ;
        RECT 49.190 120.680 49.490 121.730 ;
        RECT 49.940 121.130 50.240 122.080 ;
        RECT 50.440 121.180 50.740 121.230 ;
        RECT 50.440 120.830 51.340 121.180 ;
        RECT 42.160 119.930 42.450 120.090 ;
        RECT 43.540 120.080 43.800 120.140 ;
        RECT 12.740 119.890 17.990 119.900 ;
        RECT 2.620 119.810 2.870 119.820 ;
        RECT 2.620 119.350 3.600 119.810 ;
        RECT 12.740 119.600 18.010 119.890 ;
        RECT 2.620 119.050 2.870 119.350 ;
        RECT 10.590 119.260 12.430 119.270 ;
        RECT 17.840 119.260 18.010 119.600 ;
        RECT 4.330 119.250 4.570 119.260 ;
        RECT 5.410 119.250 18.010 119.260 ;
        RECT 4.330 119.090 18.010 119.250 ;
        RECT 41.660 119.740 42.450 119.930 ;
        RECT 41.660 119.540 41.910 119.740 ;
        RECT 42.160 119.630 42.450 119.740 ;
        RECT 43.550 119.540 43.800 120.080 ;
        RECT 46.630 120.080 46.900 120.140 ;
        RECT 48.180 120.420 49.490 120.680 ;
        RECT 51.550 120.720 53.220 120.750 ;
        RECT 68.300 120.720 68.550 120.730 ;
        RECT 51.550 120.450 68.550 120.720 ;
        RECT 51.550 120.440 65.050 120.450 ;
        RECT 52.830 120.420 65.050 120.440 ;
        RECT 48.180 120.080 48.490 120.420 ;
        RECT 44.190 119.550 45.830 119.940 ;
        RECT 46.630 119.790 48.490 120.080 ;
        RECT 46.630 119.780 46.940 119.790 ;
        RECT 48.180 119.780 48.490 119.790 ;
        RECT 4.330 119.080 15.840 119.090 ;
        RECT 4.320 119.070 10.640 119.080 ;
        RECT 12.190 119.070 15.840 119.080 ;
        RECT 4.320 119.060 6.190 119.070 ;
        RECT 4.320 119.050 4.570 119.060 ;
        RECT 2.620 118.880 4.570 119.050 ;
        RECT 41.660 118.940 41.950 119.540 ;
        RECT 43.550 118.940 43.840 119.540 ;
        RECT 2.620 118.660 2.870 118.880 ;
        RECT 2.620 118.490 3.660 118.660 ;
        RECT 3.470 117.630 3.660 118.490 ;
        RECT 45.890 118.330 46.190 119.330 ;
        RECT 46.640 118.730 46.940 119.780 ;
        RECT 49.240 118.680 49.490 120.420 ;
        RECT 49.940 118.330 50.200 119.880 ;
        RECT 50.820 118.330 51.160 118.400 ;
        RECT 45.840 118.030 51.160 118.330 ;
        RECT 2.680 117.190 3.660 117.630 ;
        RECT 2.680 117.180 3.630 117.190 ;
        RECT 4.500 116.870 13.770 116.880 ;
        RECT 15.650 116.870 17.570 116.880 ;
        RECT 2.350 116.770 2.540 116.780 ;
        RECT 2.350 116.310 3.330 116.770 ;
        RECT 4.500 116.680 17.570 116.870 ;
        RECT 4.500 116.670 16.860 116.680 ;
        RECT 2.350 115.520 2.540 116.310 ;
        RECT 4.500 115.660 4.710 116.670 ;
        RECT 13.760 116.660 15.660 116.670 ;
        RECT 17.390 115.930 17.570 116.680 ;
        RECT 3.350 115.520 3.620 115.530 ;
        RECT 2.350 115.310 3.620 115.520 ;
        RECT 3.350 115.100 3.620 115.310 ;
        RECT 3.350 114.470 3.600 115.100 ;
        RECT 4.500 114.650 4.700 115.660 ;
        RECT 12.310 115.630 17.570 115.930 ;
        RECT 2.560 114.020 3.600 114.470 ;
        RECT 2.540 112.570 3.500 113.020 ;
        RECT 3.250 112.520 3.500 112.570 ;
        RECT 4.510 112.520 4.700 114.650 ;
        RECT 3.250 112.320 4.700 112.520 ;
        RECT 8.230 113.990 8.490 115.190 ;
        RECT 8.230 113.480 8.480 113.990 ;
        RECT 10.120 113.980 10.380 115.190 ;
        RECT 12.510 114.080 12.760 115.630 ;
        RECT 10.120 113.820 10.510 113.980 ;
        RECT 10.110 113.690 10.510 113.820 ;
        RECT 13.210 113.690 13.470 115.300 ;
        RECT 15.760 114.230 16.060 115.280 ;
        RECT 16.510 114.680 16.810 115.630 ;
        RECT 17.010 114.730 17.310 114.780 ;
        RECT 17.010 114.380 17.910 114.730 ;
        RECT 19.620 114.600 19.840 114.610 ;
        RECT 19.620 114.410 33.300 114.600 ;
        RECT 19.620 114.280 19.840 114.410 ;
        RECT 8.730 113.480 9.020 113.640 ;
        RECT 10.110 113.630 10.370 113.690 ;
        RECT 8.230 113.290 9.020 113.480 ;
        RECT 8.230 113.090 8.480 113.290 ;
        RECT 8.730 113.180 9.020 113.290 ;
        RECT 10.120 113.090 10.370 113.630 ;
        RECT 13.200 113.630 13.470 113.690 ;
        RECT 14.750 113.970 16.060 114.230 ;
        RECT 18.160 113.980 19.840 114.280 ;
        RECT 18.160 113.970 19.820 113.980 ;
        RECT 14.750 113.630 15.060 113.970 ;
        RECT 10.760 113.100 12.400 113.490 ;
        RECT 13.200 113.340 15.060 113.630 ;
        RECT 13.200 113.330 13.510 113.340 ;
        RECT 14.750 113.330 15.060 113.340 ;
        RECT 8.230 112.490 8.520 113.090 ;
        RECT 10.120 112.490 10.410 113.090 ;
        RECT 3.250 112.230 3.500 112.320 ;
        RECT 2.520 111.780 3.500 112.230 ;
        RECT 12.460 111.880 12.760 112.880 ;
        RECT 13.210 112.280 13.510 113.330 ;
        RECT 15.810 112.230 16.060 113.970 ;
        RECT 33.050 113.510 33.300 114.410 ;
        RECT 16.510 111.880 16.770 113.430 ;
        RECT 27.990 113.210 33.300 113.510 ;
        RECT 12.410 111.860 17.660 111.880 ;
        RECT 12.410 111.580 17.780 111.860 ;
        RECT 5.860 111.180 6.140 111.250 ;
        RECT 7.040 111.210 7.320 111.240 ;
        RECT 17.490 111.210 17.780 111.580 ;
        RECT 7.040 111.200 17.780 111.210 ;
        RECT 4.450 110.980 6.140 111.180 ;
        RECT 3.240 110.780 3.520 110.790 ;
        RECT 2.500 110.330 3.520 110.780 ;
        RECT 4.450 110.330 4.680 110.980 ;
        RECT 5.860 110.920 6.140 110.980 ;
        RECT 7.020 110.970 17.780 111.200 ;
        RECT 7.040 110.960 17.780 110.970 ;
        RECT 23.910 111.570 24.170 112.770 ;
        RECT 23.910 111.060 24.160 111.570 ;
        RECT 25.800 111.560 26.060 112.770 ;
        RECT 28.190 111.660 28.440 113.210 ;
        RECT 25.800 111.400 26.190 111.560 ;
        RECT 25.790 111.270 26.190 111.400 ;
        RECT 28.890 111.270 29.150 112.880 ;
        RECT 31.440 111.810 31.740 112.860 ;
        RECT 32.190 112.260 32.490 113.210 ;
        RECT 32.690 112.310 32.990 112.360 ;
        RECT 32.690 111.960 33.590 112.310 ;
        RECT 50.820 111.910 51.160 118.030 ;
        RECT 50.250 111.890 51.210 111.910 ;
        RECT 34.730 111.870 39.010 111.880 ;
        RECT 46.410 111.870 51.210 111.890 ;
        RECT 34.730 111.860 51.210 111.870 ;
        RECT 24.410 111.060 24.700 111.220 ;
        RECT 25.790 111.210 26.050 111.270 ;
        RECT 7.040 110.950 17.740 110.960 ;
        RECT 7.040 110.910 7.320 110.950 ;
        RECT 23.910 110.870 24.700 111.060 ;
        RECT 23.910 110.670 24.160 110.870 ;
        RECT 24.410 110.760 24.700 110.870 ;
        RECT 25.800 110.670 26.050 111.210 ;
        RECT 28.880 111.210 29.150 111.270 ;
        RECT 30.430 111.550 31.740 111.810 ;
        RECT 30.430 111.210 30.740 111.550 ;
        RECT 26.440 110.680 28.080 111.070 ;
        RECT 28.880 110.920 30.740 111.210 ;
        RECT 28.880 110.910 29.190 110.920 ;
        RECT 30.430 110.910 30.740 110.920 ;
        RECT 5.840 110.350 6.110 110.430 ;
        RECT 3.240 110.120 4.680 110.330 ;
        RECT 5.230 110.130 6.110 110.350 ;
        RECT 3.240 109.070 3.520 110.120 ;
        RECT 5.230 109.320 5.450 110.130 ;
        RECT 5.840 110.100 6.110 110.130 ;
        RECT 6.970 110.390 7.260 110.440 ;
        RECT 6.970 110.210 17.720 110.390 ;
        RECT 6.970 110.110 7.260 110.210 ;
        RECT 11.810 110.200 15.440 110.210 ;
        RECT 17.520 109.530 17.720 110.210 ;
        RECT 23.910 110.070 24.200 110.670 ;
        RECT 25.800 110.070 26.090 110.670 ;
        RECT 2.520 108.620 3.520 109.070 ;
        RECT 2.500 107.170 3.800 107.620 ;
        RECT 3.500 106.770 3.800 107.170 ;
        RECT 5.220 106.790 5.450 109.320 ;
        RECT 12.470 109.230 17.720 109.530 ;
        RECT 28.140 109.460 28.440 110.460 ;
        RECT 28.890 109.860 29.190 110.910 ;
        RECT 31.490 109.810 31.740 111.550 ;
        RECT 33.860 111.550 51.210 111.860 ;
        RECT 33.860 111.540 46.870 111.550 ;
        RECT 38.720 111.530 46.870 111.540 ;
        RECT 50.250 111.510 51.210 111.550 ;
        RECT 50.820 111.500 51.160 111.510 ;
        RECT 32.190 109.460 32.450 111.010 ;
        RECT 33.280 109.460 33.480 109.470 ;
        RECT 4.290 106.770 5.450 106.790 ;
        RECT 3.500 106.590 5.450 106.770 ;
        RECT 8.390 107.590 8.650 108.790 ;
        RECT 8.390 107.080 8.640 107.590 ;
        RECT 10.280 107.580 10.540 108.790 ;
        RECT 12.670 107.680 12.920 109.230 ;
        RECT 10.280 107.420 10.670 107.580 ;
        RECT 10.270 107.290 10.670 107.420 ;
        RECT 13.370 107.290 13.630 108.900 ;
        RECT 15.920 107.830 16.220 108.880 ;
        RECT 16.670 108.280 16.970 109.230 ;
        RECT 17.520 109.220 17.720 109.230 ;
        RECT 28.090 109.160 33.480 109.460 ;
        RECT 17.170 108.330 17.470 108.380 ;
        RECT 17.170 107.980 18.070 108.330 ;
        RECT 33.280 107.920 33.480 109.160 ;
        RECT 25.720 107.900 26.910 107.910 ;
        RECT 27.900 107.900 29.090 107.910 ;
        RECT 30.120 107.900 31.310 107.910 ;
        RECT 32.300 107.900 33.490 107.920 ;
        RECT 23.510 107.890 33.490 107.900 ;
        RECT 20.120 107.870 21.310 107.880 ;
        RECT 22.400 107.870 33.490 107.890 ;
        RECT 8.890 107.080 9.180 107.240 ;
        RECT 10.270 107.230 10.530 107.290 ;
        RECT 8.390 106.890 9.180 107.080 ;
        RECT 8.390 106.690 8.640 106.890 ;
        RECT 8.890 106.780 9.180 106.890 ;
        RECT 10.280 106.690 10.530 107.230 ;
        RECT 13.360 107.230 13.630 107.290 ;
        RECT 14.910 107.570 16.220 107.830 ;
        RECT 18.280 107.640 33.490 107.870 ;
        RECT 18.280 107.630 32.440 107.640 ;
        RECT 18.280 107.620 25.810 107.630 ;
        RECT 26.820 107.620 28.010 107.630 ;
        RECT 28.970 107.620 30.160 107.630 ;
        RECT 31.250 107.620 32.440 107.630 ;
        RECT 18.280 107.610 23.590 107.620 ;
        RECT 18.280 107.600 22.450 107.610 ;
        RECT 18.280 107.590 20.170 107.600 ;
        RECT 21.260 107.590 22.450 107.600 ;
        RECT 18.280 107.580 19.000 107.590 ;
        RECT 14.910 107.230 15.220 107.570 ;
        RECT 10.920 106.700 12.560 107.090 ;
        RECT 13.360 106.940 15.220 107.230 ;
        RECT 13.360 106.930 13.670 106.940 ;
        RECT 14.910 106.930 15.220 106.940 ;
        RECT 3.500 106.580 4.150 106.590 ;
        RECT 3.500 106.250 3.800 106.580 ;
        RECT 2.780 105.800 3.800 106.250 ;
        RECT 8.390 106.090 8.680 106.690 ;
        RECT 10.280 106.090 10.570 106.690 ;
        RECT 3.500 105.790 3.800 105.800 ;
        RECT 12.620 105.480 12.920 106.480 ;
        RECT 13.370 105.880 13.670 106.930 ;
        RECT 15.970 105.830 16.220 107.570 ;
        RECT 68.300 107.310 68.560 120.450 ;
        RECT 68.290 107.190 68.560 107.310 ;
        RECT 16.670 105.480 16.930 107.030 ;
        RECT 68.290 106.360 68.550 107.190 ;
        RECT 63.270 106.060 68.550 106.360 ;
        RECT 12.570 105.470 17.820 105.480 ;
        RECT 2.450 105.390 2.700 105.400 ;
        RECT 2.450 104.930 3.430 105.390 ;
        RECT 12.570 105.180 17.840 105.470 ;
        RECT 2.450 104.630 2.700 104.930 ;
        RECT 10.420 104.840 12.260 104.850 ;
        RECT 17.670 104.840 17.840 105.180 ;
        RECT 4.160 104.830 4.400 104.840 ;
        RECT 5.240 104.830 17.840 104.840 ;
        RECT 4.160 104.670 17.840 104.830 ;
        RECT 4.160 104.660 15.670 104.670 ;
        RECT 4.150 104.650 10.470 104.660 ;
        RECT 12.020 104.650 15.670 104.660 ;
        RECT 4.150 104.640 6.020 104.650 ;
        RECT 4.150 104.630 4.400 104.640 ;
        RECT 2.450 104.460 4.400 104.630 ;
        RECT 2.450 104.160 2.720 104.460 ;
        RECT 2.460 103.900 2.720 104.160 ;
        RECT 59.190 104.420 59.450 105.620 ;
        RECT 59.190 103.910 59.440 104.420 ;
        RECT 61.080 104.410 61.340 105.620 ;
        RECT 63.470 104.510 63.720 106.060 ;
        RECT 61.080 104.250 61.470 104.410 ;
        RECT 61.070 104.120 61.470 104.250 ;
        RECT 64.170 104.120 64.430 105.730 ;
        RECT 66.720 104.660 67.020 105.710 ;
        RECT 67.470 105.110 67.770 106.060 ;
        RECT 67.970 105.160 68.270 105.210 ;
        RECT 67.970 104.810 68.870 105.160 ;
        RECT 59.690 103.910 59.980 104.070 ;
        RECT 61.070 104.060 61.330 104.120 ;
        RECT 2.440 103.510 2.740 103.900 ;
        RECT 59.190 103.720 59.980 103.910 ;
        RECT 59.190 103.520 59.440 103.720 ;
        RECT 59.690 103.610 59.980 103.720 ;
        RECT 61.080 103.520 61.330 104.060 ;
        RECT 64.160 104.060 64.430 104.120 ;
        RECT 65.710 104.400 67.020 104.660 ;
        RECT 69.140 104.600 69.920 104.700 ;
        RECT 69.140 104.430 82.720 104.600 ;
        RECT 69.140 104.420 82.710 104.430 ;
        RECT 69.140 104.400 69.920 104.420 ;
        RECT 65.710 104.060 66.020 104.400 ;
        RECT 61.720 103.530 63.360 103.920 ;
        RECT 64.160 103.770 66.020 104.060 ;
        RECT 64.160 103.760 64.470 103.770 ;
        RECT 65.710 103.760 66.020 103.770 ;
        RECT 2.440 103.280 3.930 103.510 ;
        RECT 3.680 102.350 3.930 103.280 ;
        RECT 59.190 102.920 59.480 103.520 ;
        RECT 61.080 102.920 61.370 103.520 ;
        RECT 2.880 101.890 3.930 102.350 ;
        RECT 63.420 102.310 63.720 103.310 ;
        RECT 64.170 102.710 64.470 103.760 ;
        RECT 66.770 102.660 67.020 104.400 ;
        RECT 67.470 102.310 67.730 103.860 ;
        RECT 63.370 102.010 68.640 102.310 ;
        RECT 3.680 101.880 3.930 101.890 ;
        RECT 2.550 101.480 2.800 101.490 ;
        RECT 2.550 101.030 3.530 101.480 ;
        RECT 4.640 101.220 13.910 101.230 ;
        RECT 15.790 101.220 17.710 101.230 ;
        RECT 4.640 101.030 17.710 101.220 ;
        RECT 2.550 100.420 2.800 101.030 ;
        RECT 4.640 101.020 17.000 101.030 ;
        RECT 2.550 100.170 3.760 100.420 ;
        RECT 3.490 99.420 3.750 100.170 ;
        RECT 4.640 100.010 4.850 101.020 ;
        RECT 13.900 101.010 15.800 101.020 ;
        RECT 17.530 100.280 17.710 101.030 ;
        RECT 3.490 98.820 3.740 99.420 ;
        RECT 4.640 99.000 4.840 100.010 ;
        RECT 12.450 99.980 17.710 100.280 ;
        RECT 2.700 98.370 3.740 98.820 ;
        RECT 2.680 96.920 3.640 97.370 ;
        RECT 3.390 96.870 3.640 96.920 ;
        RECT 4.650 96.870 4.840 99.000 ;
        RECT 3.390 96.670 4.840 96.870 ;
        RECT 8.370 98.340 8.630 99.540 ;
        RECT 8.370 97.830 8.620 98.340 ;
        RECT 10.260 98.330 10.520 99.540 ;
        RECT 12.650 98.430 12.900 99.980 ;
        RECT 10.260 98.170 10.650 98.330 ;
        RECT 10.250 98.040 10.650 98.170 ;
        RECT 13.350 98.040 13.610 99.650 ;
        RECT 15.900 98.580 16.200 99.630 ;
        RECT 16.650 99.030 16.950 99.980 ;
        RECT 17.150 99.080 17.450 99.130 ;
        RECT 17.150 98.730 18.050 99.080 ;
        RECT 19.760 98.950 19.980 98.960 ;
        RECT 19.760 98.760 33.440 98.950 ;
        RECT 19.760 98.630 19.980 98.760 ;
        RECT 8.870 97.830 9.160 97.990 ;
        RECT 10.250 97.980 10.510 98.040 ;
        RECT 8.370 97.640 9.160 97.830 ;
        RECT 8.370 97.440 8.620 97.640 ;
        RECT 8.870 97.530 9.160 97.640 ;
        RECT 10.260 97.440 10.510 97.980 ;
        RECT 13.340 97.980 13.610 98.040 ;
        RECT 14.890 98.320 16.200 98.580 ;
        RECT 18.300 98.330 19.980 98.630 ;
        RECT 18.300 98.320 19.960 98.330 ;
        RECT 14.890 97.980 15.200 98.320 ;
        RECT 10.900 97.450 12.540 97.840 ;
        RECT 13.340 97.690 15.200 97.980 ;
        RECT 13.340 97.680 13.650 97.690 ;
        RECT 14.890 97.680 15.200 97.690 ;
        RECT 8.370 96.840 8.660 97.440 ;
        RECT 10.260 96.840 10.550 97.440 ;
        RECT 3.390 96.580 3.640 96.670 ;
        RECT 2.660 96.130 3.640 96.580 ;
        RECT 12.600 96.230 12.900 97.230 ;
        RECT 13.350 96.630 13.650 97.680 ;
        RECT 15.950 96.580 16.200 98.320 ;
        RECT 33.190 97.860 33.440 98.760 ;
        RECT 16.650 96.230 16.910 97.780 ;
        RECT 28.130 97.560 33.440 97.860 ;
        RECT 12.550 96.210 17.800 96.230 ;
        RECT 12.550 95.930 17.920 96.210 ;
        RECT 6.000 95.530 6.280 95.600 ;
        RECT 7.180 95.560 7.460 95.590 ;
        RECT 17.630 95.560 17.920 95.930 ;
        RECT 7.180 95.550 17.920 95.560 ;
        RECT 4.590 95.330 6.280 95.530 ;
        RECT 3.380 95.130 3.660 95.140 ;
        RECT 2.640 94.680 3.660 95.130 ;
        RECT 4.590 94.680 4.820 95.330 ;
        RECT 6.000 95.270 6.280 95.330 ;
        RECT 7.160 95.320 17.920 95.550 ;
        RECT 7.180 95.310 17.920 95.320 ;
        RECT 24.050 95.920 24.310 97.120 ;
        RECT 24.050 95.410 24.300 95.920 ;
        RECT 25.940 95.910 26.200 97.120 ;
        RECT 28.330 96.010 28.580 97.560 ;
        RECT 25.940 95.750 26.330 95.910 ;
        RECT 25.930 95.620 26.330 95.750 ;
        RECT 29.030 95.620 29.290 97.230 ;
        RECT 31.580 96.160 31.880 97.210 ;
        RECT 32.330 96.610 32.630 97.560 ;
        RECT 32.830 96.660 33.130 96.710 ;
        RECT 32.830 96.310 33.730 96.660 ;
        RECT 46.490 96.260 50.960 96.290 ;
        RECT 35.550 96.230 50.960 96.260 ;
        RECT 34.880 96.210 50.960 96.230 ;
        RECT 24.550 95.410 24.840 95.570 ;
        RECT 25.930 95.560 26.190 95.620 ;
        RECT 7.180 95.300 17.880 95.310 ;
        RECT 7.180 95.260 7.460 95.300 ;
        RECT 24.050 95.220 24.840 95.410 ;
        RECT 24.050 95.020 24.300 95.220 ;
        RECT 24.550 95.110 24.840 95.220 ;
        RECT 25.940 95.020 26.190 95.560 ;
        RECT 29.020 95.560 29.290 95.620 ;
        RECT 30.570 95.900 31.880 96.160 ;
        RECT 30.570 95.560 30.880 95.900 ;
        RECT 26.580 95.030 28.220 95.420 ;
        RECT 29.020 95.270 30.880 95.560 ;
        RECT 29.020 95.260 29.330 95.270 ;
        RECT 30.570 95.260 30.880 95.270 ;
        RECT 5.980 94.700 6.250 94.780 ;
        RECT 3.380 94.470 4.820 94.680 ;
        RECT 5.370 94.480 6.250 94.700 ;
        RECT 3.380 93.420 3.660 94.470 ;
        RECT 5.370 93.670 5.590 94.480 ;
        RECT 5.980 94.450 6.250 94.480 ;
        RECT 7.110 94.740 7.400 94.790 ;
        RECT 7.110 94.560 17.860 94.740 ;
        RECT 7.110 94.460 7.400 94.560 ;
        RECT 11.950 94.550 15.580 94.560 ;
        RECT 17.660 93.880 17.860 94.560 ;
        RECT 24.050 94.420 24.340 95.020 ;
        RECT 25.940 94.420 26.230 95.020 ;
        RECT 2.660 92.970 3.660 93.420 ;
        RECT 2.640 91.520 3.940 91.970 ;
        RECT 3.640 91.120 3.940 91.520 ;
        RECT 5.360 91.140 5.590 93.670 ;
        RECT 12.610 93.580 17.860 93.880 ;
        RECT 28.280 93.810 28.580 94.810 ;
        RECT 29.030 94.210 29.330 95.260 ;
        RECT 31.630 94.160 31.880 95.900 ;
        RECT 34.000 95.890 50.960 96.210 ;
        RECT 34.880 95.880 50.960 95.890 ;
        RECT 34.880 95.850 46.860 95.880 ;
        RECT 34.880 95.840 35.770 95.850 ;
        RECT 32.330 93.810 32.590 95.360 ;
        RECT 33.420 93.810 33.620 93.820 ;
        RECT 4.430 91.120 5.590 91.140 ;
        RECT 3.640 90.940 5.590 91.120 ;
        RECT 8.530 91.940 8.790 93.140 ;
        RECT 8.530 91.430 8.780 91.940 ;
        RECT 10.420 91.930 10.680 93.140 ;
        RECT 12.810 92.030 13.060 93.580 ;
        RECT 10.420 91.770 10.810 91.930 ;
        RECT 10.410 91.640 10.810 91.770 ;
        RECT 13.510 91.640 13.770 93.250 ;
        RECT 16.060 92.180 16.360 93.230 ;
        RECT 16.810 92.630 17.110 93.580 ;
        RECT 17.660 93.570 17.860 93.580 ;
        RECT 28.230 93.510 33.620 93.810 ;
        RECT 17.310 92.680 17.610 92.730 ;
        RECT 17.310 92.330 18.210 92.680 ;
        RECT 33.420 92.270 33.620 93.510 ;
        RECT 50.580 92.310 50.940 95.880 ;
        RECT 25.860 92.250 27.050 92.260 ;
        RECT 28.040 92.250 29.230 92.260 ;
        RECT 30.260 92.250 31.450 92.260 ;
        RECT 32.440 92.250 33.630 92.270 ;
        RECT 23.650 92.240 33.630 92.250 ;
        RECT 20.260 92.220 21.450 92.230 ;
        RECT 22.540 92.220 33.630 92.240 ;
        RECT 9.030 91.430 9.320 91.590 ;
        RECT 10.410 91.580 10.670 91.640 ;
        RECT 8.530 91.240 9.320 91.430 ;
        RECT 8.530 91.040 8.780 91.240 ;
        RECT 9.030 91.130 9.320 91.240 ;
        RECT 10.420 91.040 10.670 91.580 ;
        RECT 13.500 91.580 13.770 91.640 ;
        RECT 15.050 91.920 16.360 92.180 ;
        RECT 18.420 91.990 33.630 92.220 ;
        RECT 45.710 92.010 50.960 92.310 ;
        RECT 18.420 91.980 32.580 91.990 ;
        RECT 18.420 91.970 25.950 91.980 ;
        RECT 26.960 91.970 28.150 91.980 ;
        RECT 29.110 91.970 30.300 91.980 ;
        RECT 31.390 91.970 32.580 91.980 ;
        RECT 18.420 91.960 23.730 91.970 ;
        RECT 18.420 91.950 22.590 91.960 ;
        RECT 18.420 91.940 20.310 91.950 ;
        RECT 21.400 91.940 22.590 91.950 ;
        RECT 18.420 91.930 19.140 91.940 ;
        RECT 15.050 91.580 15.360 91.920 ;
        RECT 11.060 91.050 12.700 91.440 ;
        RECT 13.500 91.290 15.360 91.580 ;
        RECT 13.500 91.280 13.810 91.290 ;
        RECT 15.050 91.280 15.360 91.290 ;
        RECT 3.640 90.930 4.290 90.940 ;
        RECT 3.640 90.600 3.940 90.930 ;
        RECT 2.920 90.150 3.940 90.600 ;
        RECT 8.530 90.440 8.820 91.040 ;
        RECT 10.420 90.440 10.710 91.040 ;
        RECT 3.640 90.140 3.940 90.150 ;
        RECT 12.760 89.830 13.060 90.830 ;
        RECT 13.510 90.230 13.810 91.280 ;
        RECT 16.110 90.180 16.360 91.920 ;
        RECT 16.810 89.830 17.070 91.380 ;
        RECT 41.630 90.370 41.890 91.570 ;
        RECT 41.630 89.860 41.880 90.370 ;
        RECT 43.520 90.360 43.780 91.570 ;
        RECT 45.910 90.460 46.160 92.010 ;
        RECT 43.520 90.200 43.910 90.360 ;
        RECT 43.510 90.070 43.910 90.200 ;
        RECT 46.610 90.070 46.870 91.680 ;
        RECT 49.160 90.610 49.460 91.660 ;
        RECT 49.910 91.060 50.210 92.010 ;
        RECT 50.410 91.110 50.710 91.160 ;
        RECT 50.410 90.760 51.310 91.110 ;
        RECT 42.130 89.860 42.420 90.020 ;
        RECT 43.510 90.010 43.770 90.070 ;
        RECT 12.710 89.820 17.960 89.830 ;
        RECT 2.590 89.740 2.840 89.750 ;
        RECT 2.590 89.280 3.570 89.740 ;
        RECT 12.710 89.530 17.980 89.820 ;
        RECT 2.590 88.980 2.840 89.280 ;
        RECT 10.560 89.190 12.400 89.200 ;
        RECT 17.810 89.190 17.980 89.530 ;
        RECT 4.300 89.180 4.540 89.190 ;
        RECT 5.380 89.180 17.980 89.190 ;
        RECT 4.300 89.020 17.980 89.180 ;
        RECT 41.630 89.670 42.420 89.860 ;
        RECT 41.630 89.470 41.880 89.670 ;
        RECT 42.130 89.560 42.420 89.670 ;
        RECT 43.520 89.470 43.770 90.010 ;
        RECT 46.600 90.010 46.870 90.070 ;
        RECT 48.150 90.350 49.460 90.610 ;
        RECT 51.520 90.660 53.190 90.680 ;
        RECT 68.330 90.660 68.640 102.010 ;
        RECT 51.520 90.370 68.680 90.660 ;
        RECT 52.210 90.360 68.680 90.370 ;
        RECT 48.150 90.010 48.460 90.350 ;
        RECT 44.160 89.480 45.800 89.870 ;
        RECT 46.600 89.720 48.460 90.010 ;
        RECT 46.600 89.710 46.910 89.720 ;
        RECT 48.150 89.710 48.460 89.720 ;
        RECT 4.300 89.010 15.810 89.020 ;
        RECT 4.290 89.000 10.610 89.010 ;
        RECT 12.160 89.000 15.810 89.010 ;
        RECT 4.290 88.990 6.160 89.000 ;
        RECT 4.290 88.980 4.540 88.990 ;
        RECT 2.590 88.810 4.540 88.980 ;
        RECT 41.630 88.870 41.920 89.470 ;
        RECT 43.520 88.870 43.810 89.470 ;
        RECT 2.590 88.590 2.840 88.810 ;
        RECT 2.590 88.420 3.630 88.590 ;
        RECT 3.440 87.560 3.630 88.420 ;
        RECT 45.860 88.260 46.160 89.260 ;
        RECT 46.610 88.660 46.910 89.710 ;
        RECT 49.210 88.610 49.460 90.350 ;
        RECT 49.910 88.260 50.170 89.810 ;
        RECT 50.790 88.260 51.130 88.330 ;
        RECT 45.810 87.960 51.130 88.260 ;
        RECT 2.650 87.120 3.630 87.560 ;
        RECT 2.650 87.110 3.600 87.120 ;
        RECT 4.470 86.800 13.740 86.810 ;
        RECT 15.620 86.800 17.540 86.810 ;
        RECT 2.320 86.700 2.510 86.710 ;
        RECT 2.320 86.240 3.300 86.700 ;
        RECT 4.470 86.610 17.540 86.800 ;
        RECT 4.470 86.600 16.830 86.610 ;
        RECT 2.320 85.450 2.510 86.240 ;
        RECT 4.470 85.590 4.680 86.600 ;
        RECT 13.730 86.590 15.630 86.600 ;
        RECT 17.360 85.860 17.540 86.610 ;
        RECT 3.320 85.450 3.590 85.460 ;
        RECT 2.320 85.240 3.590 85.450 ;
        RECT 3.320 85.030 3.590 85.240 ;
        RECT 3.320 84.400 3.570 85.030 ;
        RECT 4.470 84.580 4.670 85.590 ;
        RECT 12.280 85.560 17.540 85.860 ;
        RECT 2.530 83.950 3.570 84.400 ;
        RECT 2.510 82.500 3.470 82.950 ;
        RECT 3.220 82.450 3.470 82.500 ;
        RECT 4.480 82.450 4.670 84.580 ;
        RECT 3.220 82.250 4.670 82.450 ;
        RECT 8.200 83.920 8.460 85.120 ;
        RECT 8.200 83.410 8.450 83.920 ;
        RECT 10.090 83.910 10.350 85.120 ;
        RECT 12.480 84.010 12.730 85.560 ;
        RECT 10.090 83.750 10.480 83.910 ;
        RECT 10.080 83.620 10.480 83.750 ;
        RECT 13.180 83.620 13.440 85.230 ;
        RECT 15.730 84.160 16.030 85.210 ;
        RECT 16.480 84.610 16.780 85.560 ;
        RECT 16.980 84.660 17.280 84.710 ;
        RECT 16.980 84.310 17.880 84.660 ;
        RECT 19.590 84.530 19.810 84.540 ;
        RECT 19.590 84.340 33.270 84.530 ;
        RECT 19.590 84.210 19.810 84.340 ;
        RECT 8.700 83.410 8.990 83.570 ;
        RECT 10.080 83.560 10.340 83.620 ;
        RECT 8.200 83.220 8.990 83.410 ;
        RECT 8.200 83.020 8.450 83.220 ;
        RECT 8.700 83.110 8.990 83.220 ;
        RECT 10.090 83.020 10.340 83.560 ;
        RECT 13.170 83.560 13.440 83.620 ;
        RECT 14.720 83.900 16.030 84.160 ;
        RECT 18.130 83.910 19.810 84.210 ;
        RECT 18.130 83.900 19.790 83.910 ;
        RECT 14.720 83.560 15.030 83.900 ;
        RECT 10.730 83.030 12.370 83.420 ;
        RECT 13.170 83.270 15.030 83.560 ;
        RECT 13.170 83.260 13.480 83.270 ;
        RECT 14.720 83.260 15.030 83.270 ;
        RECT 8.200 82.420 8.490 83.020 ;
        RECT 10.090 82.420 10.380 83.020 ;
        RECT 3.220 82.160 3.470 82.250 ;
        RECT 2.490 81.710 3.470 82.160 ;
        RECT 12.430 81.810 12.730 82.810 ;
        RECT 13.180 82.210 13.480 83.260 ;
        RECT 15.780 82.160 16.030 83.900 ;
        RECT 33.020 83.440 33.270 84.340 ;
        RECT 16.480 81.810 16.740 83.360 ;
        RECT 27.960 83.140 33.270 83.440 ;
        RECT 12.380 81.790 17.630 81.810 ;
        RECT 12.380 81.510 17.750 81.790 ;
        RECT 5.830 81.110 6.110 81.180 ;
        RECT 7.010 81.140 7.290 81.170 ;
        RECT 17.460 81.140 17.750 81.510 ;
        RECT 7.010 81.130 17.750 81.140 ;
        RECT 4.420 80.910 6.110 81.110 ;
        RECT 3.210 80.710 3.490 80.720 ;
        RECT 2.470 80.260 3.490 80.710 ;
        RECT 4.420 80.260 4.650 80.910 ;
        RECT 5.830 80.850 6.110 80.910 ;
        RECT 6.990 80.900 17.750 81.130 ;
        RECT 7.010 80.890 17.750 80.900 ;
        RECT 23.880 81.500 24.140 82.700 ;
        RECT 23.880 80.990 24.130 81.500 ;
        RECT 25.770 81.490 26.030 82.700 ;
        RECT 28.160 81.590 28.410 83.140 ;
        RECT 25.770 81.330 26.160 81.490 ;
        RECT 25.760 81.200 26.160 81.330 ;
        RECT 28.860 81.200 29.120 82.810 ;
        RECT 31.410 81.740 31.710 82.790 ;
        RECT 32.160 82.190 32.460 83.140 ;
        RECT 32.660 82.240 32.960 82.290 ;
        RECT 32.660 81.890 33.560 82.240 ;
        RECT 50.790 81.840 51.130 87.960 ;
        RECT 82.530 85.160 82.710 104.420 ;
        RECT 82.510 84.110 82.720 85.160 ;
        RECT 82.510 84.030 82.730 84.110 ;
        RECT 82.520 81.960 82.730 84.030 ;
        RECT 82.510 81.920 82.730 81.960 ;
        RECT 50.220 81.820 51.180 81.840 ;
        RECT 34.700 81.800 38.980 81.810 ;
        RECT 46.380 81.800 51.180 81.820 ;
        RECT 34.700 81.790 51.180 81.800 ;
        RECT 24.380 80.990 24.670 81.150 ;
        RECT 25.760 81.140 26.020 81.200 ;
        RECT 7.010 80.880 17.710 80.890 ;
        RECT 7.010 80.840 7.290 80.880 ;
        RECT 23.880 80.800 24.670 80.990 ;
        RECT 23.880 80.600 24.130 80.800 ;
        RECT 24.380 80.690 24.670 80.800 ;
        RECT 25.770 80.600 26.020 81.140 ;
        RECT 28.850 81.140 29.120 81.200 ;
        RECT 30.400 81.480 31.710 81.740 ;
        RECT 30.400 81.140 30.710 81.480 ;
        RECT 26.410 80.610 28.050 81.000 ;
        RECT 28.850 80.850 30.710 81.140 ;
        RECT 28.850 80.840 29.160 80.850 ;
        RECT 30.400 80.840 30.710 80.850 ;
        RECT 5.810 80.280 6.080 80.360 ;
        RECT 3.210 80.050 4.650 80.260 ;
        RECT 5.200 80.060 6.080 80.280 ;
        RECT 3.210 79.000 3.490 80.050 ;
        RECT 5.200 79.250 5.420 80.060 ;
        RECT 5.810 80.030 6.080 80.060 ;
        RECT 6.940 80.320 7.230 80.370 ;
        RECT 6.940 80.140 17.690 80.320 ;
        RECT 6.940 80.040 7.230 80.140 ;
        RECT 11.780 80.130 15.410 80.140 ;
        RECT 17.490 79.460 17.690 80.140 ;
        RECT 23.880 80.000 24.170 80.600 ;
        RECT 25.770 80.000 26.060 80.600 ;
        RECT 2.490 78.550 3.490 79.000 ;
        RECT 2.470 77.100 3.770 77.550 ;
        RECT 3.470 76.700 3.770 77.100 ;
        RECT 5.190 76.720 5.420 79.250 ;
        RECT 12.440 79.160 17.690 79.460 ;
        RECT 28.110 79.390 28.410 80.390 ;
        RECT 28.860 79.790 29.160 80.840 ;
        RECT 31.460 79.740 31.710 81.480 ;
        RECT 33.830 81.480 51.180 81.790 ;
        RECT 33.830 81.470 46.840 81.480 ;
        RECT 38.690 81.460 46.840 81.470 ;
        RECT 50.220 81.440 51.180 81.480 ;
        RECT 50.790 81.430 51.130 81.440 ;
        RECT 32.160 79.390 32.420 80.940 ;
        RECT 82.510 80.070 82.720 81.920 ;
        RECT 77.470 79.770 82.720 80.070 ;
        RECT 33.250 79.390 33.450 79.400 ;
        RECT 4.260 76.700 5.420 76.720 ;
        RECT 3.470 76.520 5.420 76.700 ;
        RECT 8.360 77.520 8.620 78.720 ;
        RECT 8.360 77.010 8.610 77.520 ;
        RECT 10.250 77.510 10.510 78.720 ;
        RECT 12.640 77.610 12.890 79.160 ;
        RECT 10.250 77.350 10.640 77.510 ;
        RECT 10.240 77.220 10.640 77.350 ;
        RECT 13.340 77.220 13.600 78.830 ;
        RECT 15.890 77.760 16.190 78.810 ;
        RECT 16.640 78.210 16.940 79.160 ;
        RECT 17.490 79.150 17.690 79.160 ;
        RECT 28.060 79.090 33.450 79.390 ;
        RECT 17.140 78.260 17.440 78.310 ;
        RECT 17.140 77.910 18.040 78.260 ;
        RECT 33.250 77.850 33.450 79.090 ;
        RECT 73.390 78.130 73.650 79.330 ;
        RECT 25.690 77.830 26.880 77.840 ;
        RECT 27.870 77.830 29.060 77.840 ;
        RECT 30.090 77.830 31.280 77.840 ;
        RECT 32.270 77.830 33.460 77.850 ;
        RECT 23.480 77.820 33.460 77.830 ;
        RECT 20.090 77.800 21.280 77.810 ;
        RECT 22.370 77.800 33.460 77.820 ;
        RECT 8.860 77.010 9.150 77.170 ;
        RECT 10.240 77.160 10.500 77.220 ;
        RECT 8.360 76.820 9.150 77.010 ;
        RECT 8.360 76.620 8.610 76.820 ;
        RECT 8.860 76.710 9.150 76.820 ;
        RECT 10.250 76.620 10.500 77.160 ;
        RECT 13.330 77.160 13.600 77.220 ;
        RECT 14.880 77.500 16.190 77.760 ;
        RECT 18.250 77.570 33.460 77.800 ;
        RECT 73.390 77.620 73.640 78.130 ;
        RECT 75.280 78.120 75.540 79.330 ;
        RECT 77.670 78.220 77.920 79.770 ;
        RECT 75.280 77.960 75.670 78.120 ;
        RECT 75.270 77.830 75.670 77.960 ;
        RECT 78.370 77.830 78.630 79.440 ;
        RECT 80.920 78.370 81.220 79.420 ;
        RECT 81.670 78.820 81.970 79.770 ;
        RECT 82.510 79.760 82.720 79.770 ;
        RECT 82.170 78.870 82.470 78.920 ;
        RECT 82.170 78.520 83.070 78.870 ;
        RECT 99.840 78.490 100.140 132.830 ;
        RECT 103.840 132.180 104.190 132.840 ;
        RECT 195.710 132.640 201.450 132.930 ;
        RECT 212.920 132.890 227.370 133.090 ;
        RECT 212.920 132.880 224.720 132.890 ;
        RECT 212.920 132.860 220.880 132.880 ;
        RECT 195.710 132.630 200.960 132.640 ;
        RECT 102.570 131.840 104.190 132.180 ;
        RECT 102.570 130.990 103.020 131.840 ;
        RECT 103.840 131.830 104.190 131.840 ;
        RECT 103.430 130.810 103.890 131.640 ;
        RECT 105.980 131.100 115.250 131.110 ;
        RECT 117.130 131.100 119.050 131.110 ;
        RECT 104.810 130.810 105.090 130.950 ;
        RECT 103.430 130.700 105.090 130.810 ;
        RECT 103.440 130.500 105.090 130.700 ;
        RECT 105.980 130.910 119.050 131.100 ;
        RECT 105.980 130.900 118.340 130.910 ;
        RECT 103.440 130.490 105.110 130.500 ;
        RECT 104.810 130.270 105.110 130.490 ;
        RECT 104.820 130.100 105.110 130.270 ;
        RECT 104.830 129.300 105.090 130.100 ;
        RECT 105.980 129.890 106.190 130.900 ;
        RECT 115.240 130.890 117.140 130.900 ;
        RECT 118.870 130.160 119.050 130.910 ;
        RECT 104.830 128.700 105.080 129.300 ;
        RECT 105.980 128.880 106.180 129.890 ;
        RECT 113.790 129.860 119.050 130.160 ;
        RECT 104.040 128.250 105.080 128.700 ;
        RECT 104.020 126.800 104.980 127.250 ;
        RECT 104.730 126.750 104.980 126.800 ;
        RECT 105.990 126.750 106.180 128.880 ;
        RECT 104.730 126.550 106.180 126.750 ;
        RECT 109.710 128.220 109.970 129.420 ;
        RECT 109.710 127.710 109.960 128.220 ;
        RECT 111.600 128.210 111.860 129.420 ;
        RECT 113.990 128.310 114.240 129.860 ;
        RECT 111.600 128.050 111.990 128.210 ;
        RECT 111.590 127.920 111.990 128.050 ;
        RECT 114.690 127.920 114.950 129.530 ;
        RECT 117.240 128.460 117.540 129.510 ;
        RECT 117.990 128.910 118.290 129.860 ;
        RECT 118.490 128.960 118.790 129.010 ;
        RECT 118.490 128.610 119.390 128.960 ;
        RECT 121.100 128.830 121.320 128.840 ;
        RECT 121.100 128.640 134.780 128.830 ;
        RECT 121.100 128.510 121.320 128.640 ;
        RECT 110.210 127.710 110.500 127.870 ;
        RECT 111.590 127.860 111.850 127.920 ;
        RECT 109.710 127.520 110.500 127.710 ;
        RECT 109.710 127.320 109.960 127.520 ;
        RECT 110.210 127.410 110.500 127.520 ;
        RECT 111.600 127.320 111.850 127.860 ;
        RECT 114.680 127.860 114.950 127.920 ;
        RECT 116.230 128.200 117.540 128.460 ;
        RECT 119.640 128.210 121.320 128.510 ;
        RECT 119.640 128.200 121.300 128.210 ;
        RECT 116.230 127.860 116.540 128.200 ;
        RECT 112.240 127.330 113.880 127.720 ;
        RECT 114.680 127.570 116.540 127.860 ;
        RECT 114.680 127.560 114.990 127.570 ;
        RECT 116.230 127.560 116.540 127.570 ;
        RECT 109.710 126.720 110.000 127.320 ;
        RECT 111.600 126.720 111.890 127.320 ;
        RECT 104.730 126.460 104.980 126.550 ;
        RECT 104.000 126.010 104.980 126.460 ;
        RECT 113.940 126.110 114.240 127.110 ;
        RECT 114.690 126.510 114.990 127.560 ;
        RECT 117.290 126.460 117.540 128.200 ;
        RECT 134.530 127.740 134.780 128.640 ;
        RECT 117.990 126.110 118.250 127.660 ;
        RECT 129.470 127.440 134.780 127.740 ;
        RECT 113.890 126.090 119.140 126.110 ;
        RECT 113.890 125.810 119.260 126.090 ;
        RECT 107.340 125.410 107.620 125.480 ;
        RECT 108.520 125.440 108.800 125.470 ;
        RECT 118.970 125.440 119.260 125.810 ;
        RECT 108.520 125.430 119.260 125.440 ;
        RECT 105.930 125.210 107.620 125.410 ;
        RECT 104.720 125.010 105.000 125.020 ;
        RECT 103.980 124.560 105.000 125.010 ;
        RECT 105.930 124.560 106.160 125.210 ;
        RECT 107.340 125.150 107.620 125.210 ;
        RECT 108.500 125.200 119.260 125.430 ;
        RECT 108.520 125.190 119.260 125.200 ;
        RECT 125.390 125.800 125.650 127.000 ;
        RECT 125.390 125.290 125.640 125.800 ;
        RECT 127.280 125.790 127.540 127.000 ;
        RECT 129.670 125.890 129.920 127.440 ;
        RECT 127.280 125.630 127.670 125.790 ;
        RECT 127.270 125.500 127.670 125.630 ;
        RECT 130.370 125.500 130.630 127.110 ;
        RECT 132.920 126.040 133.220 127.090 ;
        RECT 133.670 126.490 133.970 127.440 ;
        RECT 134.170 126.540 134.470 126.590 ;
        RECT 134.170 126.190 135.070 126.540 ;
        RECT 147.830 126.140 152.300 126.170 ;
        RECT 136.890 126.110 152.300 126.140 ;
        RECT 136.220 126.090 152.300 126.110 ;
        RECT 125.890 125.290 126.180 125.450 ;
        RECT 127.270 125.440 127.530 125.500 ;
        RECT 108.520 125.180 119.220 125.190 ;
        RECT 108.520 125.140 108.800 125.180 ;
        RECT 125.390 125.100 126.180 125.290 ;
        RECT 125.390 124.900 125.640 125.100 ;
        RECT 125.890 124.990 126.180 125.100 ;
        RECT 127.280 124.900 127.530 125.440 ;
        RECT 130.360 125.440 130.630 125.500 ;
        RECT 131.910 125.780 133.220 126.040 ;
        RECT 131.910 125.440 132.220 125.780 ;
        RECT 127.920 124.910 129.560 125.300 ;
        RECT 130.360 125.150 132.220 125.440 ;
        RECT 130.360 125.140 130.670 125.150 ;
        RECT 131.910 125.140 132.220 125.150 ;
        RECT 107.320 124.580 107.590 124.660 ;
        RECT 104.720 124.350 106.160 124.560 ;
        RECT 106.710 124.360 107.590 124.580 ;
        RECT 104.720 123.300 105.000 124.350 ;
        RECT 106.710 123.550 106.930 124.360 ;
        RECT 107.320 124.330 107.590 124.360 ;
        RECT 108.450 124.620 108.740 124.670 ;
        RECT 108.450 124.440 119.200 124.620 ;
        RECT 108.450 124.340 108.740 124.440 ;
        RECT 113.290 124.430 116.920 124.440 ;
        RECT 119.000 123.760 119.200 124.440 ;
        RECT 125.390 124.300 125.680 124.900 ;
        RECT 127.280 124.300 127.570 124.900 ;
        RECT 104.000 122.850 105.000 123.300 ;
        RECT 103.980 121.400 105.280 121.850 ;
        RECT 104.980 121.000 105.280 121.400 ;
        RECT 106.700 121.020 106.930 123.550 ;
        RECT 113.950 123.460 119.200 123.760 ;
        RECT 129.620 123.690 129.920 124.690 ;
        RECT 130.370 124.090 130.670 125.140 ;
        RECT 132.970 124.040 133.220 125.780 ;
        RECT 135.340 125.770 152.300 126.090 ;
        RECT 136.220 125.760 152.300 125.770 ;
        RECT 136.220 125.730 148.200 125.760 ;
        RECT 136.220 125.720 137.110 125.730 ;
        RECT 133.670 123.690 133.930 125.240 ;
        RECT 134.760 123.690 134.960 123.700 ;
        RECT 105.770 121.000 106.930 121.020 ;
        RECT 104.980 120.820 106.930 121.000 ;
        RECT 109.870 121.820 110.130 123.020 ;
        RECT 109.870 121.310 110.120 121.820 ;
        RECT 111.760 121.810 112.020 123.020 ;
        RECT 114.150 121.910 114.400 123.460 ;
        RECT 111.760 121.650 112.150 121.810 ;
        RECT 111.750 121.520 112.150 121.650 ;
        RECT 114.850 121.520 115.110 123.130 ;
        RECT 117.400 122.060 117.700 123.110 ;
        RECT 118.150 122.510 118.450 123.460 ;
        RECT 119.000 123.450 119.200 123.460 ;
        RECT 129.570 123.390 134.960 123.690 ;
        RECT 118.650 122.560 118.950 122.610 ;
        RECT 118.650 122.210 119.550 122.560 ;
        RECT 134.760 122.150 134.960 123.390 ;
        RECT 151.920 122.190 152.280 125.760 ;
        RECT 127.200 122.130 128.390 122.140 ;
        RECT 129.380 122.130 130.570 122.140 ;
        RECT 131.600 122.130 132.790 122.140 ;
        RECT 133.780 122.130 134.970 122.150 ;
        RECT 124.990 122.120 134.970 122.130 ;
        RECT 121.600 122.100 122.790 122.110 ;
        RECT 123.880 122.100 134.970 122.120 ;
        RECT 110.370 121.310 110.660 121.470 ;
        RECT 111.750 121.460 112.010 121.520 ;
        RECT 109.870 121.120 110.660 121.310 ;
        RECT 109.870 120.920 110.120 121.120 ;
        RECT 110.370 121.010 110.660 121.120 ;
        RECT 111.760 120.920 112.010 121.460 ;
        RECT 114.840 121.460 115.110 121.520 ;
        RECT 116.390 121.800 117.700 122.060 ;
        RECT 119.760 121.870 134.970 122.100 ;
        RECT 147.050 121.890 152.300 122.190 ;
        RECT 119.760 121.860 133.920 121.870 ;
        RECT 119.760 121.850 127.290 121.860 ;
        RECT 128.300 121.850 129.490 121.860 ;
        RECT 130.450 121.850 131.640 121.860 ;
        RECT 132.730 121.850 133.920 121.860 ;
        RECT 119.760 121.840 125.070 121.850 ;
        RECT 119.760 121.830 123.930 121.840 ;
        RECT 119.760 121.820 121.650 121.830 ;
        RECT 122.740 121.820 123.930 121.830 ;
        RECT 119.760 121.810 120.480 121.820 ;
        RECT 116.390 121.460 116.700 121.800 ;
        RECT 112.400 120.930 114.040 121.320 ;
        RECT 114.840 121.170 116.700 121.460 ;
        RECT 114.840 121.160 115.150 121.170 ;
        RECT 116.390 121.160 116.700 121.170 ;
        RECT 104.980 120.810 105.630 120.820 ;
        RECT 104.980 120.480 105.280 120.810 ;
        RECT 104.260 120.030 105.280 120.480 ;
        RECT 109.870 120.320 110.160 120.920 ;
        RECT 111.760 120.320 112.050 120.920 ;
        RECT 104.980 120.020 105.280 120.030 ;
        RECT 114.100 119.710 114.400 120.710 ;
        RECT 114.850 120.110 115.150 121.160 ;
        RECT 117.450 120.060 117.700 121.800 ;
        RECT 118.150 119.710 118.410 121.260 ;
        RECT 142.970 120.250 143.230 121.450 ;
        RECT 142.970 119.740 143.220 120.250 ;
        RECT 144.860 120.240 145.120 121.450 ;
        RECT 147.250 120.340 147.500 121.890 ;
        RECT 144.860 120.080 145.250 120.240 ;
        RECT 144.850 119.950 145.250 120.080 ;
        RECT 147.950 119.950 148.210 121.560 ;
        RECT 150.500 120.490 150.800 121.540 ;
        RECT 151.250 120.940 151.550 121.890 ;
        RECT 151.750 120.990 152.050 121.040 ;
        RECT 151.750 120.640 152.650 120.990 ;
        RECT 143.470 119.740 143.760 119.900 ;
        RECT 144.850 119.890 145.110 119.950 ;
        RECT 114.050 119.700 119.300 119.710 ;
        RECT 103.930 119.620 104.180 119.630 ;
        RECT 103.930 119.160 104.910 119.620 ;
        RECT 114.050 119.410 119.320 119.700 ;
        RECT 103.930 118.860 104.180 119.160 ;
        RECT 111.900 119.070 113.740 119.080 ;
        RECT 119.150 119.070 119.320 119.410 ;
        RECT 105.640 119.060 105.880 119.070 ;
        RECT 106.720 119.060 119.320 119.070 ;
        RECT 105.640 118.900 119.320 119.060 ;
        RECT 142.970 119.550 143.760 119.740 ;
        RECT 142.970 119.350 143.220 119.550 ;
        RECT 143.470 119.440 143.760 119.550 ;
        RECT 144.860 119.350 145.110 119.890 ;
        RECT 147.940 119.890 148.210 119.950 ;
        RECT 149.490 120.230 150.800 120.490 ;
        RECT 152.860 120.530 154.530 120.560 ;
        RECT 169.610 120.530 169.860 120.540 ;
        RECT 152.860 120.260 169.860 120.530 ;
        RECT 152.860 120.250 166.360 120.260 ;
        RECT 154.140 120.230 166.360 120.250 ;
        RECT 149.490 119.890 149.800 120.230 ;
        RECT 145.500 119.360 147.140 119.750 ;
        RECT 147.940 119.600 149.800 119.890 ;
        RECT 147.940 119.590 148.250 119.600 ;
        RECT 149.490 119.590 149.800 119.600 ;
        RECT 105.640 118.890 117.150 118.900 ;
        RECT 105.630 118.880 111.950 118.890 ;
        RECT 113.500 118.880 117.150 118.890 ;
        RECT 105.630 118.870 107.500 118.880 ;
        RECT 105.630 118.860 105.880 118.870 ;
        RECT 103.930 118.690 105.880 118.860 ;
        RECT 142.970 118.750 143.260 119.350 ;
        RECT 144.860 118.750 145.150 119.350 ;
        RECT 103.930 118.470 104.180 118.690 ;
        RECT 103.930 118.300 104.970 118.470 ;
        RECT 104.780 117.440 104.970 118.300 ;
        RECT 147.200 118.140 147.500 119.140 ;
        RECT 147.950 118.540 148.250 119.590 ;
        RECT 150.550 118.490 150.800 120.230 ;
        RECT 151.250 118.140 151.510 119.690 ;
        RECT 152.130 118.140 152.470 118.210 ;
        RECT 147.150 117.840 152.470 118.140 ;
        RECT 103.990 117.000 104.970 117.440 ;
        RECT 103.990 116.990 104.940 117.000 ;
        RECT 105.810 116.680 115.080 116.690 ;
        RECT 116.960 116.680 118.880 116.690 ;
        RECT 103.660 116.580 103.850 116.590 ;
        RECT 103.660 116.120 104.640 116.580 ;
        RECT 105.810 116.490 118.880 116.680 ;
        RECT 105.810 116.480 118.170 116.490 ;
        RECT 103.660 115.330 103.850 116.120 ;
        RECT 105.810 115.470 106.020 116.480 ;
        RECT 115.070 116.470 116.970 116.480 ;
        RECT 118.700 115.740 118.880 116.490 ;
        RECT 104.660 115.330 104.930 115.340 ;
        RECT 103.660 115.120 104.930 115.330 ;
        RECT 104.660 114.910 104.930 115.120 ;
        RECT 104.660 114.280 104.910 114.910 ;
        RECT 105.810 114.460 106.010 115.470 ;
        RECT 113.620 115.440 118.880 115.740 ;
        RECT 103.870 113.830 104.910 114.280 ;
        RECT 103.850 112.380 104.810 112.830 ;
        RECT 104.560 112.330 104.810 112.380 ;
        RECT 105.820 112.330 106.010 114.460 ;
        RECT 104.560 112.130 106.010 112.330 ;
        RECT 109.540 113.800 109.800 115.000 ;
        RECT 109.540 113.290 109.790 113.800 ;
        RECT 111.430 113.790 111.690 115.000 ;
        RECT 113.820 113.890 114.070 115.440 ;
        RECT 111.430 113.630 111.820 113.790 ;
        RECT 111.420 113.500 111.820 113.630 ;
        RECT 114.520 113.500 114.780 115.110 ;
        RECT 117.070 114.040 117.370 115.090 ;
        RECT 117.820 114.490 118.120 115.440 ;
        RECT 118.320 114.540 118.620 114.590 ;
        RECT 118.320 114.190 119.220 114.540 ;
        RECT 120.930 114.410 121.150 114.420 ;
        RECT 120.930 114.220 134.610 114.410 ;
        RECT 120.930 114.090 121.150 114.220 ;
        RECT 110.040 113.290 110.330 113.450 ;
        RECT 111.420 113.440 111.680 113.500 ;
        RECT 109.540 113.100 110.330 113.290 ;
        RECT 109.540 112.900 109.790 113.100 ;
        RECT 110.040 112.990 110.330 113.100 ;
        RECT 111.430 112.900 111.680 113.440 ;
        RECT 114.510 113.440 114.780 113.500 ;
        RECT 116.060 113.780 117.370 114.040 ;
        RECT 119.470 113.790 121.150 114.090 ;
        RECT 119.470 113.780 121.130 113.790 ;
        RECT 116.060 113.440 116.370 113.780 ;
        RECT 112.070 112.910 113.710 113.300 ;
        RECT 114.510 113.150 116.370 113.440 ;
        RECT 114.510 113.140 114.820 113.150 ;
        RECT 116.060 113.140 116.370 113.150 ;
        RECT 109.540 112.300 109.830 112.900 ;
        RECT 111.430 112.300 111.720 112.900 ;
        RECT 104.560 112.040 104.810 112.130 ;
        RECT 103.830 111.590 104.810 112.040 ;
        RECT 113.770 111.690 114.070 112.690 ;
        RECT 114.520 112.090 114.820 113.140 ;
        RECT 117.120 112.040 117.370 113.780 ;
        RECT 134.360 113.320 134.610 114.220 ;
        RECT 117.820 111.690 118.080 113.240 ;
        RECT 129.300 113.020 134.610 113.320 ;
        RECT 113.720 111.670 118.970 111.690 ;
        RECT 113.720 111.390 119.090 111.670 ;
        RECT 107.170 110.990 107.450 111.060 ;
        RECT 108.350 111.020 108.630 111.050 ;
        RECT 118.800 111.020 119.090 111.390 ;
        RECT 108.350 111.010 119.090 111.020 ;
        RECT 105.760 110.790 107.450 110.990 ;
        RECT 104.550 110.590 104.830 110.600 ;
        RECT 103.810 110.140 104.830 110.590 ;
        RECT 105.760 110.140 105.990 110.790 ;
        RECT 107.170 110.730 107.450 110.790 ;
        RECT 108.330 110.780 119.090 111.010 ;
        RECT 108.350 110.770 119.090 110.780 ;
        RECT 125.220 111.380 125.480 112.580 ;
        RECT 125.220 110.870 125.470 111.380 ;
        RECT 127.110 111.370 127.370 112.580 ;
        RECT 129.500 111.470 129.750 113.020 ;
        RECT 127.110 111.210 127.500 111.370 ;
        RECT 127.100 111.080 127.500 111.210 ;
        RECT 130.200 111.080 130.460 112.690 ;
        RECT 132.750 111.620 133.050 112.670 ;
        RECT 133.500 112.070 133.800 113.020 ;
        RECT 134.000 112.120 134.300 112.170 ;
        RECT 134.000 111.770 134.900 112.120 ;
        RECT 152.130 111.720 152.470 117.840 ;
        RECT 151.560 111.700 152.520 111.720 ;
        RECT 136.040 111.680 140.320 111.690 ;
        RECT 147.720 111.680 152.520 111.700 ;
        RECT 136.040 111.670 152.520 111.680 ;
        RECT 125.720 110.870 126.010 111.030 ;
        RECT 127.100 111.020 127.360 111.080 ;
        RECT 108.350 110.760 119.050 110.770 ;
        RECT 108.350 110.720 108.630 110.760 ;
        RECT 125.220 110.680 126.010 110.870 ;
        RECT 125.220 110.480 125.470 110.680 ;
        RECT 125.720 110.570 126.010 110.680 ;
        RECT 127.110 110.480 127.360 111.020 ;
        RECT 130.190 111.020 130.460 111.080 ;
        RECT 131.740 111.360 133.050 111.620 ;
        RECT 131.740 111.020 132.050 111.360 ;
        RECT 127.750 110.490 129.390 110.880 ;
        RECT 130.190 110.730 132.050 111.020 ;
        RECT 130.190 110.720 130.500 110.730 ;
        RECT 131.740 110.720 132.050 110.730 ;
        RECT 107.150 110.160 107.420 110.240 ;
        RECT 104.550 109.930 105.990 110.140 ;
        RECT 106.540 109.940 107.420 110.160 ;
        RECT 104.550 108.880 104.830 109.930 ;
        RECT 106.540 109.130 106.760 109.940 ;
        RECT 107.150 109.910 107.420 109.940 ;
        RECT 108.280 110.200 108.570 110.250 ;
        RECT 108.280 110.020 119.030 110.200 ;
        RECT 108.280 109.920 108.570 110.020 ;
        RECT 113.120 110.010 116.750 110.020 ;
        RECT 118.830 109.340 119.030 110.020 ;
        RECT 125.220 109.880 125.510 110.480 ;
        RECT 127.110 109.880 127.400 110.480 ;
        RECT 103.830 108.430 104.830 108.880 ;
        RECT 103.810 106.980 105.110 107.430 ;
        RECT 104.810 106.580 105.110 106.980 ;
        RECT 106.530 106.600 106.760 109.130 ;
        RECT 113.780 109.040 119.030 109.340 ;
        RECT 129.450 109.270 129.750 110.270 ;
        RECT 130.200 109.670 130.500 110.720 ;
        RECT 132.800 109.620 133.050 111.360 ;
        RECT 135.170 111.360 152.520 111.670 ;
        RECT 135.170 111.350 148.180 111.360 ;
        RECT 140.030 111.340 148.180 111.350 ;
        RECT 151.560 111.320 152.520 111.360 ;
        RECT 152.130 111.310 152.470 111.320 ;
        RECT 133.500 109.270 133.760 110.820 ;
        RECT 134.590 109.270 134.790 109.280 ;
        RECT 105.600 106.580 106.760 106.600 ;
        RECT 104.810 106.400 106.760 106.580 ;
        RECT 109.700 107.400 109.960 108.600 ;
        RECT 109.700 106.890 109.950 107.400 ;
        RECT 111.590 107.390 111.850 108.600 ;
        RECT 113.980 107.490 114.230 109.040 ;
        RECT 111.590 107.230 111.980 107.390 ;
        RECT 111.580 107.100 111.980 107.230 ;
        RECT 114.680 107.100 114.940 108.710 ;
        RECT 117.230 107.640 117.530 108.690 ;
        RECT 117.980 108.090 118.280 109.040 ;
        RECT 118.830 109.030 119.030 109.040 ;
        RECT 129.400 108.970 134.790 109.270 ;
        RECT 118.480 108.140 118.780 108.190 ;
        RECT 118.480 107.790 119.380 108.140 ;
        RECT 134.590 107.730 134.790 108.970 ;
        RECT 127.030 107.710 128.220 107.720 ;
        RECT 129.210 107.710 130.400 107.720 ;
        RECT 131.430 107.710 132.620 107.720 ;
        RECT 133.610 107.710 134.800 107.730 ;
        RECT 124.820 107.700 134.800 107.710 ;
        RECT 121.430 107.680 122.620 107.690 ;
        RECT 123.710 107.680 134.800 107.700 ;
        RECT 110.200 106.890 110.490 107.050 ;
        RECT 111.580 107.040 111.840 107.100 ;
        RECT 109.700 106.700 110.490 106.890 ;
        RECT 109.700 106.500 109.950 106.700 ;
        RECT 110.200 106.590 110.490 106.700 ;
        RECT 111.590 106.500 111.840 107.040 ;
        RECT 114.670 107.040 114.940 107.100 ;
        RECT 116.220 107.380 117.530 107.640 ;
        RECT 119.590 107.450 134.800 107.680 ;
        RECT 119.590 107.440 133.750 107.450 ;
        RECT 119.590 107.430 127.120 107.440 ;
        RECT 128.130 107.430 129.320 107.440 ;
        RECT 130.280 107.430 131.470 107.440 ;
        RECT 132.560 107.430 133.750 107.440 ;
        RECT 119.590 107.420 124.900 107.430 ;
        RECT 119.590 107.410 123.760 107.420 ;
        RECT 119.590 107.400 121.480 107.410 ;
        RECT 122.570 107.400 123.760 107.410 ;
        RECT 119.590 107.390 120.310 107.400 ;
        RECT 116.220 107.040 116.530 107.380 ;
        RECT 112.230 106.510 113.870 106.900 ;
        RECT 114.670 106.750 116.530 107.040 ;
        RECT 114.670 106.740 114.980 106.750 ;
        RECT 116.220 106.740 116.530 106.750 ;
        RECT 104.810 106.390 105.460 106.400 ;
        RECT 104.810 106.060 105.110 106.390 ;
        RECT 104.090 105.610 105.110 106.060 ;
        RECT 109.700 105.900 109.990 106.500 ;
        RECT 111.590 105.900 111.880 106.500 ;
        RECT 104.810 105.600 105.110 105.610 ;
        RECT 113.930 105.290 114.230 106.290 ;
        RECT 114.680 105.690 114.980 106.740 ;
        RECT 117.280 105.640 117.530 107.380 ;
        RECT 169.610 107.120 169.870 120.260 ;
        RECT 169.600 107.000 169.870 107.120 ;
        RECT 117.980 105.290 118.240 106.840 ;
        RECT 169.600 106.170 169.860 107.000 ;
        RECT 164.580 105.870 169.860 106.170 ;
        RECT 113.880 105.280 119.130 105.290 ;
        RECT 103.760 105.200 104.010 105.210 ;
        RECT 103.760 104.740 104.740 105.200 ;
        RECT 113.880 104.990 119.150 105.280 ;
        RECT 103.760 104.440 104.010 104.740 ;
        RECT 111.730 104.650 113.570 104.660 ;
        RECT 118.980 104.650 119.150 104.990 ;
        RECT 105.470 104.640 105.710 104.650 ;
        RECT 106.550 104.640 119.150 104.650 ;
        RECT 105.470 104.480 119.150 104.640 ;
        RECT 105.470 104.470 116.980 104.480 ;
        RECT 105.460 104.460 111.780 104.470 ;
        RECT 113.330 104.460 116.980 104.470 ;
        RECT 105.460 104.450 107.330 104.460 ;
        RECT 105.460 104.440 105.710 104.450 ;
        RECT 103.760 104.270 105.710 104.440 ;
        RECT 103.760 103.970 104.030 104.270 ;
        RECT 103.770 103.710 104.030 103.970 ;
        RECT 160.500 104.230 160.760 105.430 ;
        RECT 160.500 103.720 160.750 104.230 ;
        RECT 162.390 104.220 162.650 105.430 ;
        RECT 164.780 104.320 165.030 105.870 ;
        RECT 162.390 104.060 162.780 104.220 ;
        RECT 162.380 103.930 162.780 104.060 ;
        RECT 165.480 103.930 165.740 105.540 ;
        RECT 168.030 104.470 168.330 105.520 ;
        RECT 168.780 104.920 169.080 105.870 ;
        RECT 169.280 104.970 169.580 105.020 ;
        RECT 169.280 104.620 170.180 104.970 ;
        RECT 161.000 103.720 161.290 103.880 ;
        RECT 162.380 103.870 162.640 103.930 ;
        RECT 103.750 103.320 104.050 103.710 ;
        RECT 160.500 103.530 161.290 103.720 ;
        RECT 160.500 103.330 160.750 103.530 ;
        RECT 161.000 103.420 161.290 103.530 ;
        RECT 162.390 103.330 162.640 103.870 ;
        RECT 165.470 103.870 165.740 103.930 ;
        RECT 167.020 104.210 168.330 104.470 ;
        RECT 170.450 104.410 171.230 104.510 ;
        RECT 170.450 104.240 184.030 104.410 ;
        RECT 170.450 104.230 184.020 104.240 ;
        RECT 170.450 104.210 171.230 104.230 ;
        RECT 167.020 103.870 167.330 104.210 ;
        RECT 163.030 103.340 164.670 103.730 ;
        RECT 165.470 103.580 167.330 103.870 ;
        RECT 165.470 103.570 165.780 103.580 ;
        RECT 167.020 103.570 167.330 103.580 ;
        RECT 103.750 103.090 105.240 103.320 ;
        RECT 104.990 102.160 105.240 103.090 ;
        RECT 160.500 102.730 160.790 103.330 ;
        RECT 162.390 102.730 162.680 103.330 ;
        RECT 104.190 101.700 105.240 102.160 ;
        RECT 164.730 102.120 165.030 103.120 ;
        RECT 165.480 102.520 165.780 103.570 ;
        RECT 168.080 102.470 168.330 104.210 ;
        RECT 168.780 102.120 169.040 103.670 ;
        RECT 164.680 101.820 169.950 102.120 ;
        RECT 104.990 101.690 105.240 101.700 ;
        RECT 103.860 101.290 104.110 101.300 ;
        RECT 103.860 100.840 104.840 101.290 ;
        RECT 105.950 101.030 115.220 101.040 ;
        RECT 117.100 101.030 119.020 101.040 ;
        RECT 105.950 100.840 119.020 101.030 ;
        RECT 103.860 100.230 104.110 100.840 ;
        RECT 105.950 100.830 118.310 100.840 ;
        RECT 103.860 99.980 105.070 100.230 ;
        RECT 104.800 99.230 105.060 99.980 ;
        RECT 105.950 99.820 106.160 100.830 ;
        RECT 115.210 100.820 117.110 100.830 ;
        RECT 118.840 100.090 119.020 100.840 ;
        RECT 104.800 98.630 105.050 99.230 ;
        RECT 105.950 98.810 106.150 99.820 ;
        RECT 113.760 99.790 119.020 100.090 ;
        RECT 104.010 98.180 105.050 98.630 ;
        RECT 103.990 96.730 104.950 97.180 ;
        RECT 104.700 96.680 104.950 96.730 ;
        RECT 105.960 96.680 106.150 98.810 ;
        RECT 104.700 96.480 106.150 96.680 ;
        RECT 109.680 98.150 109.940 99.350 ;
        RECT 109.680 97.640 109.930 98.150 ;
        RECT 111.570 98.140 111.830 99.350 ;
        RECT 113.960 98.240 114.210 99.790 ;
        RECT 111.570 97.980 111.960 98.140 ;
        RECT 111.560 97.850 111.960 97.980 ;
        RECT 114.660 97.850 114.920 99.460 ;
        RECT 117.210 98.390 117.510 99.440 ;
        RECT 117.960 98.840 118.260 99.790 ;
        RECT 118.460 98.890 118.760 98.940 ;
        RECT 118.460 98.540 119.360 98.890 ;
        RECT 121.070 98.760 121.290 98.770 ;
        RECT 121.070 98.570 134.750 98.760 ;
        RECT 121.070 98.440 121.290 98.570 ;
        RECT 110.180 97.640 110.470 97.800 ;
        RECT 111.560 97.790 111.820 97.850 ;
        RECT 109.680 97.450 110.470 97.640 ;
        RECT 109.680 97.250 109.930 97.450 ;
        RECT 110.180 97.340 110.470 97.450 ;
        RECT 111.570 97.250 111.820 97.790 ;
        RECT 114.650 97.790 114.920 97.850 ;
        RECT 116.200 98.130 117.510 98.390 ;
        RECT 119.610 98.140 121.290 98.440 ;
        RECT 119.610 98.130 121.270 98.140 ;
        RECT 116.200 97.790 116.510 98.130 ;
        RECT 112.210 97.260 113.850 97.650 ;
        RECT 114.650 97.500 116.510 97.790 ;
        RECT 114.650 97.490 114.960 97.500 ;
        RECT 116.200 97.490 116.510 97.500 ;
        RECT 109.680 96.650 109.970 97.250 ;
        RECT 111.570 96.650 111.860 97.250 ;
        RECT 104.700 96.390 104.950 96.480 ;
        RECT 103.970 95.940 104.950 96.390 ;
        RECT 113.910 96.040 114.210 97.040 ;
        RECT 114.660 96.440 114.960 97.490 ;
        RECT 117.260 96.390 117.510 98.130 ;
        RECT 134.500 97.670 134.750 98.570 ;
        RECT 117.960 96.040 118.220 97.590 ;
        RECT 129.440 97.370 134.750 97.670 ;
        RECT 113.860 96.020 119.110 96.040 ;
        RECT 113.860 95.740 119.230 96.020 ;
        RECT 107.310 95.340 107.590 95.410 ;
        RECT 108.490 95.370 108.770 95.400 ;
        RECT 118.940 95.370 119.230 95.740 ;
        RECT 108.490 95.360 119.230 95.370 ;
        RECT 105.900 95.140 107.590 95.340 ;
        RECT 104.690 94.940 104.970 94.950 ;
        RECT 103.950 94.490 104.970 94.940 ;
        RECT 105.900 94.490 106.130 95.140 ;
        RECT 107.310 95.080 107.590 95.140 ;
        RECT 108.470 95.130 119.230 95.360 ;
        RECT 108.490 95.120 119.230 95.130 ;
        RECT 125.360 95.730 125.620 96.930 ;
        RECT 125.360 95.220 125.610 95.730 ;
        RECT 127.250 95.720 127.510 96.930 ;
        RECT 129.640 95.820 129.890 97.370 ;
        RECT 127.250 95.560 127.640 95.720 ;
        RECT 127.240 95.430 127.640 95.560 ;
        RECT 130.340 95.430 130.600 97.040 ;
        RECT 132.890 95.970 133.190 97.020 ;
        RECT 133.640 96.420 133.940 97.370 ;
        RECT 134.140 96.470 134.440 96.520 ;
        RECT 134.140 96.120 135.040 96.470 ;
        RECT 147.800 96.070 152.270 96.100 ;
        RECT 136.860 96.040 152.270 96.070 ;
        RECT 136.190 96.020 152.270 96.040 ;
        RECT 125.860 95.220 126.150 95.380 ;
        RECT 127.240 95.370 127.500 95.430 ;
        RECT 108.490 95.110 119.190 95.120 ;
        RECT 108.490 95.070 108.770 95.110 ;
        RECT 125.360 95.030 126.150 95.220 ;
        RECT 125.360 94.830 125.610 95.030 ;
        RECT 125.860 94.920 126.150 95.030 ;
        RECT 127.250 94.830 127.500 95.370 ;
        RECT 130.330 95.370 130.600 95.430 ;
        RECT 131.880 95.710 133.190 95.970 ;
        RECT 131.880 95.370 132.190 95.710 ;
        RECT 127.890 94.840 129.530 95.230 ;
        RECT 130.330 95.080 132.190 95.370 ;
        RECT 130.330 95.070 130.640 95.080 ;
        RECT 131.880 95.070 132.190 95.080 ;
        RECT 107.290 94.510 107.560 94.590 ;
        RECT 104.690 94.280 106.130 94.490 ;
        RECT 106.680 94.290 107.560 94.510 ;
        RECT 104.690 93.230 104.970 94.280 ;
        RECT 106.680 93.480 106.900 94.290 ;
        RECT 107.290 94.260 107.560 94.290 ;
        RECT 108.420 94.550 108.710 94.600 ;
        RECT 108.420 94.370 119.170 94.550 ;
        RECT 108.420 94.270 108.710 94.370 ;
        RECT 113.260 94.360 116.890 94.370 ;
        RECT 118.970 93.690 119.170 94.370 ;
        RECT 125.360 94.230 125.650 94.830 ;
        RECT 127.250 94.230 127.540 94.830 ;
        RECT 103.970 92.780 104.970 93.230 ;
        RECT 103.950 91.330 105.250 91.780 ;
        RECT 104.950 90.930 105.250 91.330 ;
        RECT 106.670 90.950 106.900 93.480 ;
        RECT 113.920 93.390 119.170 93.690 ;
        RECT 129.590 93.620 129.890 94.620 ;
        RECT 130.340 94.020 130.640 95.070 ;
        RECT 132.940 93.970 133.190 95.710 ;
        RECT 135.310 95.700 152.270 96.020 ;
        RECT 136.190 95.690 152.270 95.700 ;
        RECT 136.190 95.660 148.170 95.690 ;
        RECT 136.190 95.650 137.080 95.660 ;
        RECT 133.640 93.620 133.900 95.170 ;
        RECT 134.730 93.620 134.930 93.630 ;
        RECT 105.740 90.930 106.900 90.950 ;
        RECT 104.950 90.750 106.900 90.930 ;
        RECT 109.840 91.750 110.100 92.950 ;
        RECT 109.840 91.240 110.090 91.750 ;
        RECT 111.730 91.740 111.990 92.950 ;
        RECT 114.120 91.840 114.370 93.390 ;
        RECT 111.730 91.580 112.120 91.740 ;
        RECT 111.720 91.450 112.120 91.580 ;
        RECT 114.820 91.450 115.080 93.060 ;
        RECT 117.370 91.990 117.670 93.040 ;
        RECT 118.120 92.440 118.420 93.390 ;
        RECT 118.970 93.380 119.170 93.390 ;
        RECT 129.540 93.320 134.930 93.620 ;
        RECT 118.620 92.490 118.920 92.540 ;
        RECT 118.620 92.140 119.520 92.490 ;
        RECT 134.730 92.080 134.930 93.320 ;
        RECT 151.890 92.120 152.250 95.690 ;
        RECT 127.170 92.060 128.360 92.070 ;
        RECT 129.350 92.060 130.540 92.070 ;
        RECT 131.570 92.060 132.760 92.070 ;
        RECT 133.750 92.060 134.940 92.080 ;
        RECT 124.960 92.050 134.940 92.060 ;
        RECT 121.570 92.030 122.760 92.040 ;
        RECT 123.850 92.030 134.940 92.050 ;
        RECT 110.340 91.240 110.630 91.400 ;
        RECT 111.720 91.390 111.980 91.450 ;
        RECT 109.840 91.050 110.630 91.240 ;
        RECT 109.840 90.850 110.090 91.050 ;
        RECT 110.340 90.940 110.630 91.050 ;
        RECT 111.730 90.850 111.980 91.390 ;
        RECT 114.810 91.390 115.080 91.450 ;
        RECT 116.360 91.730 117.670 91.990 ;
        RECT 119.730 91.800 134.940 92.030 ;
        RECT 147.020 91.820 152.270 92.120 ;
        RECT 119.730 91.790 133.890 91.800 ;
        RECT 119.730 91.780 127.260 91.790 ;
        RECT 128.270 91.780 129.460 91.790 ;
        RECT 130.420 91.780 131.610 91.790 ;
        RECT 132.700 91.780 133.890 91.790 ;
        RECT 119.730 91.770 125.040 91.780 ;
        RECT 119.730 91.760 123.900 91.770 ;
        RECT 119.730 91.750 121.620 91.760 ;
        RECT 122.710 91.750 123.900 91.760 ;
        RECT 119.730 91.740 120.450 91.750 ;
        RECT 116.360 91.390 116.670 91.730 ;
        RECT 112.370 90.860 114.010 91.250 ;
        RECT 114.810 91.100 116.670 91.390 ;
        RECT 114.810 91.090 115.120 91.100 ;
        RECT 116.360 91.090 116.670 91.100 ;
        RECT 104.950 90.740 105.600 90.750 ;
        RECT 104.950 90.410 105.250 90.740 ;
        RECT 104.230 89.960 105.250 90.410 ;
        RECT 109.840 90.250 110.130 90.850 ;
        RECT 111.730 90.250 112.020 90.850 ;
        RECT 104.950 89.950 105.250 89.960 ;
        RECT 114.070 89.640 114.370 90.640 ;
        RECT 114.820 90.040 115.120 91.090 ;
        RECT 117.420 89.990 117.670 91.730 ;
        RECT 118.120 89.640 118.380 91.190 ;
        RECT 142.940 90.180 143.200 91.380 ;
        RECT 142.940 89.670 143.190 90.180 ;
        RECT 144.830 90.170 145.090 91.380 ;
        RECT 147.220 90.270 147.470 91.820 ;
        RECT 144.830 90.010 145.220 90.170 ;
        RECT 144.820 89.880 145.220 90.010 ;
        RECT 147.920 89.880 148.180 91.490 ;
        RECT 150.470 90.420 150.770 91.470 ;
        RECT 151.220 90.870 151.520 91.820 ;
        RECT 151.720 90.920 152.020 90.970 ;
        RECT 151.720 90.570 152.620 90.920 ;
        RECT 143.440 89.670 143.730 89.830 ;
        RECT 144.820 89.820 145.080 89.880 ;
        RECT 114.020 89.630 119.270 89.640 ;
        RECT 103.900 89.550 104.150 89.560 ;
        RECT 103.900 89.090 104.880 89.550 ;
        RECT 114.020 89.340 119.290 89.630 ;
        RECT 103.900 88.790 104.150 89.090 ;
        RECT 111.870 89.000 113.710 89.010 ;
        RECT 119.120 89.000 119.290 89.340 ;
        RECT 105.610 88.990 105.850 89.000 ;
        RECT 106.690 88.990 119.290 89.000 ;
        RECT 105.610 88.830 119.290 88.990 ;
        RECT 142.940 89.480 143.730 89.670 ;
        RECT 142.940 89.280 143.190 89.480 ;
        RECT 143.440 89.370 143.730 89.480 ;
        RECT 144.830 89.280 145.080 89.820 ;
        RECT 147.910 89.820 148.180 89.880 ;
        RECT 149.460 90.160 150.770 90.420 ;
        RECT 152.830 90.470 154.500 90.490 ;
        RECT 169.640 90.470 169.950 101.820 ;
        RECT 152.830 90.180 169.990 90.470 ;
        RECT 153.520 90.170 169.990 90.180 ;
        RECT 149.460 89.820 149.770 90.160 ;
        RECT 145.470 89.290 147.110 89.680 ;
        RECT 147.910 89.530 149.770 89.820 ;
        RECT 147.910 89.520 148.220 89.530 ;
        RECT 149.460 89.520 149.770 89.530 ;
        RECT 105.610 88.820 117.120 88.830 ;
        RECT 105.600 88.810 111.920 88.820 ;
        RECT 113.470 88.810 117.120 88.820 ;
        RECT 105.600 88.800 107.470 88.810 ;
        RECT 105.600 88.790 105.850 88.800 ;
        RECT 103.900 88.620 105.850 88.790 ;
        RECT 142.940 88.680 143.230 89.280 ;
        RECT 144.830 88.680 145.120 89.280 ;
        RECT 103.900 88.400 104.150 88.620 ;
        RECT 103.900 88.230 104.940 88.400 ;
        RECT 104.750 87.370 104.940 88.230 ;
        RECT 147.170 88.070 147.470 89.070 ;
        RECT 147.920 88.470 148.220 89.520 ;
        RECT 150.520 88.420 150.770 90.160 ;
        RECT 151.220 88.070 151.480 89.620 ;
        RECT 152.100 88.070 152.440 88.140 ;
        RECT 147.120 87.770 152.440 88.070 ;
        RECT 103.960 86.930 104.940 87.370 ;
        RECT 103.960 86.920 104.910 86.930 ;
        RECT 105.780 86.610 115.050 86.620 ;
        RECT 116.930 86.610 118.850 86.620 ;
        RECT 103.630 86.510 103.820 86.520 ;
        RECT 103.630 86.050 104.610 86.510 ;
        RECT 105.780 86.420 118.850 86.610 ;
        RECT 105.780 86.410 118.140 86.420 ;
        RECT 103.630 85.260 103.820 86.050 ;
        RECT 105.780 85.400 105.990 86.410 ;
        RECT 115.040 86.400 116.940 86.410 ;
        RECT 118.670 85.670 118.850 86.420 ;
        RECT 104.630 85.260 104.900 85.270 ;
        RECT 103.630 85.050 104.900 85.260 ;
        RECT 104.630 84.840 104.900 85.050 ;
        RECT 104.630 84.210 104.880 84.840 ;
        RECT 105.780 84.390 105.980 85.400 ;
        RECT 113.590 85.370 118.850 85.670 ;
        RECT 103.840 83.760 104.880 84.210 ;
        RECT 103.820 82.310 104.780 82.760 ;
        RECT 104.530 82.260 104.780 82.310 ;
        RECT 105.790 82.260 105.980 84.390 ;
        RECT 104.530 82.060 105.980 82.260 ;
        RECT 109.510 83.730 109.770 84.930 ;
        RECT 109.510 83.220 109.760 83.730 ;
        RECT 111.400 83.720 111.660 84.930 ;
        RECT 113.790 83.820 114.040 85.370 ;
        RECT 111.400 83.560 111.790 83.720 ;
        RECT 111.390 83.430 111.790 83.560 ;
        RECT 114.490 83.430 114.750 85.040 ;
        RECT 117.040 83.970 117.340 85.020 ;
        RECT 117.790 84.420 118.090 85.370 ;
        RECT 118.290 84.470 118.590 84.520 ;
        RECT 118.290 84.120 119.190 84.470 ;
        RECT 120.900 84.340 121.120 84.350 ;
        RECT 120.900 84.150 134.580 84.340 ;
        RECT 120.900 84.020 121.120 84.150 ;
        RECT 110.010 83.220 110.300 83.380 ;
        RECT 111.390 83.370 111.650 83.430 ;
        RECT 109.510 83.030 110.300 83.220 ;
        RECT 109.510 82.830 109.760 83.030 ;
        RECT 110.010 82.920 110.300 83.030 ;
        RECT 111.400 82.830 111.650 83.370 ;
        RECT 114.480 83.370 114.750 83.430 ;
        RECT 116.030 83.710 117.340 83.970 ;
        RECT 119.440 83.720 121.120 84.020 ;
        RECT 119.440 83.710 121.100 83.720 ;
        RECT 116.030 83.370 116.340 83.710 ;
        RECT 112.040 82.840 113.680 83.230 ;
        RECT 114.480 83.080 116.340 83.370 ;
        RECT 114.480 83.070 114.790 83.080 ;
        RECT 116.030 83.070 116.340 83.080 ;
        RECT 109.510 82.230 109.800 82.830 ;
        RECT 111.400 82.230 111.690 82.830 ;
        RECT 104.530 81.970 104.780 82.060 ;
        RECT 103.800 81.520 104.780 81.970 ;
        RECT 113.740 81.620 114.040 82.620 ;
        RECT 114.490 82.020 114.790 83.070 ;
        RECT 117.090 81.970 117.340 83.710 ;
        RECT 134.330 83.250 134.580 84.150 ;
        RECT 117.790 81.620 118.050 83.170 ;
        RECT 129.270 82.950 134.580 83.250 ;
        RECT 113.690 81.600 118.940 81.620 ;
        RECT 113.690 81.320 119.060 81.600 ;
        RECT 107.140 80.920 107.420 80.990 ;
        RECT 108.320 80.950 108.600 80.980 ;
        RECT 118.770 80.950 119.060 81.320 ;
        RECT 108.320 80.940 119.060 80.950 ;
        RECT 105.730 80.720 107.420 80.920 ;
        RECT 104.520 80.520 104.800 80.530 ;
        RECT 103.780 80.070 104.800 80.520 ;
        RECT 105.730 80.070 105.960 80.720 ;
        RECT 107.140 80.660 107.420 80.720 ;
        RECT 108.300 80.710 119.060 80.940 ;
        RECT 108.320 80.700 119.060 80.710 ;
        RECT 125.190 81.310 125.450 82.510 ;
        RECT 125.190 80.800 125.440 81.310 ;
        RECT 127.080 81.300 127.340 82.510 ;
        RECT 129.470 81.400 129.720 82.950 ;
        RECT 127.080 81.140 127.470 81.300 ;
        RECT 127.070 81.010 127.470 81.140 ;
        RECT 130.170 81.010 130.430 82.620 ;
        RECT 132.720 81.550 133.020 82.600 ;
        RECT 133.470 82.000 133.770 82.950 ;
        RECT 133.970 82.050 134.270 82.100 ;
        RECT 133.970 81.700 134.870 82.050 ;
        RECT 152.100 81.650 152.440 87.770 ;
        RECT 183.840 84.970 184.020 104.230 ;
        RECT 183.820 83.920 184.030 84.970 ;
        RECT 183.820 83.840 184.040 83.920 ;
        RECT 183.830 81.770 184.040 83.840 ;
        RECT 183.820 81.730 184.040 81.770 ;
        RECT 151.530 81.630 152.490 81.650 ;
        RECT 136.010 81.610 140.290 81.620 ;
        RECT 147.690 81.610 152.490 81.630 ;
        RECT 136.010 81.600 152.490 81.610 ;
        RECT 125.690 80.800 125.980 80.960 ;
        RECT 127.070 80.950 127.330 81.010 ;
        RECT 108.320 80.690 119.020 80.700 ;
        RECT 108.320 80.650 108.600 80.690 ;
        RECT 125.190 80.610 125.980 80.800 ;
        RECT 125.190 80.410 125.440 80.610 ;
        RECT 125.690 80.500 125.980 80.610 ;
        RECT 127.080 80.410 127.330 80.950 ;
        RECT 130.160 80.950 130.430 81.010 ;
        RECT 131.710 81.290 133.020 81.550 ;
        RECT 131.710 80.950 132.020 81.290 ;
        RECT 127.720 80.420 129.360 80.810 ;
        RECT 130.160 80.660 132.020 80.950 ;
        RECT 130.160 80.650 130.470 80.660 ;
        RECT 131.710 80.650 132.020 80.660 ;
        RECT 107.120 80.090 107.390 80.170 ;
        RECT 104.520 79.860 105.960 80.070 ;
        RECT 106.510 79.870 107.390 80.090 ;
        RECT 104.520 78.810 104.800 79.860 ;
        RECT 106.510 79.060 106.730 79.870 ;
        RECT 107.120 79.840 107.390 79.870 ;
        RECT 108.250 80.130 108.540 80.180 ;
        RECT 108.250 79.950 119.000 80.130 ;
        RECT 108.250 79.850 108.540 79.950 ;
        RECT 113.090 79.940 116.720 79.950 ;
        RECT 118.800 79.270 119.000 79.950 ;
        RECT 125.190 79.810 125.480 80.410 ;
        RECT 127.080 79.810 127.370 80.410 ;
        RECT 84.080 78.400 100.140 78.490 ;
        RECT 73.890 77.620 74.180 77.780 ;
        RECT 75.270 77.770 75.530 77.830 ;
        RECT 18.250 77.560 32.410 77.570 ;
        RECT 18.250 77.550 25.780 77.560 ;
        RECT 26.790 77.550 27.980 77.560 ;
        RECT 28.940 77.550 30.130 77.560 ;
        RECT 31.220 77.550 32.410 77.560 ;
        RECT 18.250 77.540 23.560 77.550 ;
        RECT 18.250 77.530 22.420 77.540 ;
        RECT 18.250 77.520 20.140 77.530 ;
        RECT 21.230 77.520 22.420 77.530 ;
        RECT 18.250 77.510 18.970 77.520 ;
        RECT 14.880 77.160 15.190 77.500 ;
        RECT 10.890 76.630 12.530 77.020 ;
        RECT 13.330 76.870 15.190 77.160 ;
        RECT 13.330 76.860 13.640 76.870 ;
        RECT 14.880 76.860 15.190 76.870 ;
        RECT 3.470 76.510 4.120 76.520 ;
        RECT 3.470 76.180 3.770 76.510 ;
        RECT 2.750 75.730 3.770 76.180 ;
        RECT 8.360 76.020 8.650 76.620 ;
        RECT 10.250 76.020 10.540 76.620 ;
        RECT 3.470 75.720 3.770 75.730 ;
        RECT 12.590 75.410 12.890 76.410 ;
        RECT 13.340 75.810 13.640 76.860 ;
        RECT 15.940 75.760 16.190 77.500 ;
        RECT 73.390 77.430 74.180 77.620 ;
        RECT 73.390 77.230 73.640 77.430 ;
        RECT 73.890 77.320 74.180 77.430 ;
        RECT 75.280 77.230 75.530 77.770 ;
        RECT 78.360 77.770 78.630 77.830 ;
        RECT 79.910 78.110 81.220 78.370 ;
        RECT 83.360 78.120 100.140 78.400 ;
        RECT 103.800 78.360 104.800 78.810 ;
        RECT 79.910 77.770 80.220 78.110 ;
        RECT 75.920 77.240 77.560 77.630 ;
        RECT 78.360 77.480 80.220 77.770 ;
        RECT 78.360 77.470 78.670 77.480 ;
        RECT 79.910 77.470 80.220 77.480 ;
        RECT 16.640 75.410 16.900 76.960 ;
        RECT 73.390 76.630 73.680 77.230 ;
        RECT 75.280 76.630 75.570 77.230 ;
        RECT 77.620 76.020 77.920 77.020 ;
        RECT 78.370 76.420 78.670 77.470 ;
        RECT 80.970 76.370 81.220 78.110 ;
        RECT 84.080 78.070 100.140 78.120 ;
        RECT 84.080 78.060 99.810 78.070 ;
        RECT 81.670 76.020 81.930 77.570 ;
        RECT 103.780 76.910 105.080 77.360 ;
        RECT 104.780 76.510 105.080 76.910 ;
        RECT 106.500 76.530 106.730 79.060 ;
        RECT 113.750 78.970 119.000 79.270 ;
        RECT 129.420 79.200 129.720 80.200 ;
        RECT 130.170 79.600 130.470 80.650 ;
        RECT 132.770 79.550 133.020 81.290 ;
        RECT 135.140 81.290 152.490 81.600 ;
        RECT 135.140 81.280 148.150 81.290 ;
        RECT 140.000 81.270 148.150 81.280 ;
        RECT 151.530 81.250 152.490 81.290 ;
        RECT 152.100 81.240 152.440 81.250 ;
        RECT 133.470 79.200 133.730 80.750 ;
        RECT 183.820 79.880 184.030 81.730 ;
        RECT 178.780 79.580 184.030 79.880 ;
        RECT 134.560 79.200 134.760 79.210 ;
        RECT 105.570 76.510 106.730 76.530 ;
        RECT 104.780 76.330 106.730 76.510 ;
        RECT 109.670 77.330 109.930 78.530 ;
        RECT 109.670 76.820 109.920 77.330 ;
        RECT 111.560 77.320 111.820 78.530 ;
        RECT 113.950 77.420 114.200 78.970 ;
        RECT 111.560 77.160 111.950 77.320 ;
        RECT 111.550 77.030 111.950 77.160 ;
        RECT 114.650 77.030 114.910 78.640 ;
        RECT 117.200 77.570 117.500 78.620 ;
        RECT 117.950 78.020 118.250 78.970 ;
        RECT 118.800 78.960 119.000 78.970 ;
        RECT 129.370 78.900 134.760 79.200 ;
        RECT 118.450 78.070 118.750 78.120 ;
        RECT 118.450 77.720 119.350 78.070 ;
        RECT 134.560 77.660 134.760 78.900 ;
        RECT 174.700 77.940 174.960 79.140 ;
        RECT 127.000 77.640 128.190 77.650 ;
        RECT 129.180 77.640 130.370 77.650 ;
        RECT 131.400 77.640 132.590 77.650 ;
        RECT 133.580 77.640 134.770 77.660 ;
        RECT 124.790 77.630 134.770 77.640 ;
        RECT 121.400 77.610 122.590 77.620 ;
        RECT 123.680 77.610 134.770 77.630 ;
        RECT 110.170 76.820 110.460 76.980 ;
        RECT 111.550 76.970 111.810 77.030 ;
        RECT 109.670 76.630 110.460 76.820 ;
        RECT 109.670 76.430 109.920 76.630 ;
        RECT 110.170 76.520 110.460 76.630 ;
        RECT 111.560 76.430 111.810 76.970 ;
        RECT 114.640 76.970 114.910 77.030 ;
        RECT 116.190 77.310 117.500 77.570 ;
        RECT 119.560 77.380 134.770 77.610 ;
        RECT 174.700 77.430 174.950 77.940 ;
        RECT 176.590 77.930 176.850 79.140 ;
        RECT 178.980 78.030 179.230 79.580 ;
        RECT 176.590 77.770 176.980 77.930 ;
        RECT 176.580 77.640 176.980 77.770 ;
        RECT 179.680 77.640 179.940 79.250 ;
        RECT 182.230 78.180 182.530 79.230 ;
        RECT 182.980 78.630 183.280 79.580 ;
        RECT 183.820 79.570 184.030 79.580 ;
        RECT 183.480 78.680 183.780 78.730 ;
        RECT 183.480 78.330 184.380 78.680 ;
        RECT 201.150 78.300 201.450 132.640 ;
        RECT 185.390 78.210 201.450 78.300 ;
        RECT 175.200 77.430 175.490 77.590 ;
        RECT 176.580 77.580 176.840 77.640 ;
        RECT 119.560 77.370 133.720 77.380 ;
        RECT 119.560 77.360 127.090 77.370 ;
        RECT 128.100 77.360 129.290 77.370 ;
        RECT 130.250 77.360 131.440 77.370 ;
        RECT 132.530 77.360 133.720 77.370 ;
        RECT 119.560 77.350 124.870 77.360 ;
        RECT 119.560 77.340 123.730 77.350 ;
        RECT 119.560 77.330 121.450 77.340 ;
        RECT 122.540 77.330 123.730 77.340 ;
        RECT 119.560 77.320 120.280 77.330 ;
        RECT 116.190 76.970 116.500 77.310 ;
        RECT 112.200 76.440 113.840 76.830 ;
        RECT 114.640 76.680 116.500 76.970 ;
        RECT 114.640 76.670 114.950 76.680 ;
        RECT 116.190 76.670 116.500 76.680 ;
        RECT 104.780 76.320 105.430 76.330 ;
        RECT 82.630 76.020 82.810 76.030 ;
        RECT 77.570 75.720 82.820 76.020 ;
        RECT 104.780 75.990 105.080 76.320 ;
        RECT 12.540 75.400 17.790 75.410 ;
        RECT 2.420 75.320 2.670 75.330 ;
        RECT 2.420 74.860 3.400 75.320 ;
        RECT 12.540 75.110 17.810 75.400 ;
        RECT 2.420 74.560 2.670 74.860 ;
        RECT 10.390 74.770 12.230 74.780 ;
        RECT 17.640 74.770 17.810 75.110 ;
        RECT 4.130 74.760 4.370 74.770 ;
        RECT 5.210 74.760 17.810 74.770 ;
        RECT 4.130 74.600 17.810 74.760 ;
        RECT 4.130 74.590 15.640 74.600 ;
        RECT 4.120 74.580 10.440 74.590 ;
        RECT 11.990 74.580 15.640 74.590 ;
        RECT 4.120 74.570 5.990 74.580 ;
        RECT 4.120 74.560 4.370 74.570 ;
        RECT 2.420 74.390 4.370 74.560 ;
        RECT 2.420 74.090 2.690 74.390 ;
        RECT 2.430 73.830 2.690 74.090 ;
        RECT 2.410 73.440 2.710 73.830 ;
        RECT 2.400 73.040 2.710 73.440 ;
        RECT 2.390 72.280 2.700 73.040 ;
        RECT 2.290 72.260 2.700 72.280 ;
        RECT 2.260 71.310 2.710 72.260 ;
        RECT 3.120 71.020 3.580 71.960 ;
        RECT 4.320 71.370 13.590 71.380 ;
        RECT 15.470 71.370 17.390 71.380 ;
        RECT 4.320 71.180 17.390 71.370 ;
        RECT 4.320 71.170 16.680 71.180 ;
        RECT 3.160 70.700 3.460 71.020 ;
        RECT 3.160 70.370 3.450 70.700 ;
        RECT 3.170 69.570 3.430 70.370 ;
        RECT 4.320 70.160 4.530 71.170 ;
        RECT 13.580 71.160 15.480 71.170 ;
        RECT 17.210 70.430 17.390 71.180 ;
        RECT 3.170 68.970 3.420 69.570 ;
        RECT 4.320 69.150 4.520 70.160 ;
        RECT 12.130 70.130 17.390 70.430 ;
        RECT 2.380 68.520 3.420 68.970 ;
        RECT 2.360 67.070 3.320 67.520 ;
        RECT 3.070 67.020 3.320 67.070 ;
        RECT 4.330 67.020 4.520 69.150 ;
        RECT 3.070 66.820 4.520 67.020 ;
        RECT 8.050 68.490 8.310 69.690 ;
        RECT 8.050 67.980 8.300 68.490 ;
        RECT 9.940 68.480 10.200 69.690 ;
        RECT 12.330 68.580 12.580 70.130 ;
        RECT 9.940 68.320 10.330 68.480 ;
        RECT 9.930 68.190 10.330 68.320 ;
        RECT 13.030 68.190 13.290 69.800 ;
        RECT 15.580 68.730 15.880 69.780 ;
        RECT 16.330 69.180 16.630 70.130 ;
        RECT 16.830 69.230 17.130 69.280 ;
        RECT 16.830 68.880 17.730 69.230 ;
        RECT 19.440 69.100 19.660 69.110 ;
        RECT 19.440 68.910 33.120 69.100 ;
        RECT 19.440 68.780 19.660 68.910 ;
        RECT 8.550 67.980 8.840 68.140 ;
        RECT 9.930 68.130 10.190 68.190 ;
        RECT 8.050 67.790 8.840 67.980 ;
        RECT 8.050 67.590 8.300 67.790 ;
        RECT 8.550 67.680 8.840 67.790 ;
        RECT 9.940 67.590 10.190 68.130 ;
        RECT 13.020 68.130 13.290 68.190 ;
        RECT 14.570 68.470 15.880 68.730 ;
        RECT 17.980 68.480 19.660 68.780 ;
        RECT 17.980 68.470 19.640 68.480 ;
        RECT 14.570 68.130 14.880 68.470 ;
        RECT 10.580 67.600 12.220 67.990 ;
        RECT 13.020 67.840 14.880 68.130 ;
        RECT 13.020 67.830 13.330 67.840 ;
        RECT 14.570 67.830 14.880 67.840 ;
        RECT 8.050 66.990 8.340 67.590 ;
        RECT 9.940 66.990 10.230 67.590 ;
        RECT 3.070 66.730 3.320 66.820 ;
        RECT 2.340 66.280 3.320 66.730 ;
        RECT 12.280 66.380 12.580 67.380 ;
        RECT 13.030 66.780 13.330 67.830 ;
        RECT 15.630 66.730 15.880 68.470 ;
        RECT 32.870 68.010 33.120 68.910 ;
        RECT 16.330 66.380 16.590 67.930 ;
        RECT 27.810 67.710 33.120 68.010 ;
        RECT 12.230 66.360 17.480 66.380 ;
        RECT 12.230 66.080 17.600 66.360 ;
        RECT 5.680 65.680 5.960 65.750 ;
        RECT 6.860 65.710 7.140 65.740 ;
        RECT 17.310 65.710 17.600 66.080 ;
        RECT 6.860 65.700 17.600 65.710 ;
        RECT 4.270 65.480 5.960 65.680 ;
        RECT 3.060 65.280 3.340 65.290 ;
        RECT 2.320 64.830 3.340 65.280 ;
        RECT 4.270 64.830 4.500 65.480 ;
        RECT 5.680 65.420 5.960 65.480 ;
        RECT 6.840 65.470 17.600 65.700 ;
        RECT 6.860 65.460 17.600 65.470 ;
        RECT 23.730 66.070 23.990 67.270 ;
        RECT 23.730 65.560 23.980 66.070 ;
        RECT 25.620 66.060 25.880 67.270 ;
        RECT 28.010 66.160 28.260 67.710 ;
        RECT 25.620 65.900 26.010 66.060 ;
        RECT 25.610 65.770 26.010 65.900 ;
        RECT 28.710 65.770 28.970 67.380 ;
        RECT 31.260 66.310 31.560 67.360 ;
        RECT 32.010 66.760 32.310 67.710 ;
        RECT 32.510 66.810 32.810 66.860 ;
        RECT 32.510 66.460 33.410 66.810 ;
        RECT 46.170 66.410 50.640 66.440 ;
        RECT 35.230 66.380 50.640 66.410 ;
        RECT 34.560 66.360 50.640 66.380 ;
        RECT 24.230 65.560 24.520 65.720 ;
        RECT 25.610 65.710 25.870 65.770 ;
        RECT 6.860 65.450 17.560 65.460 ;
        RECT 6.860 65.410 7.140 65.450 ;
        RECT 23.730 65.370 24.520 65.560 ;
        RECT 23.730 65.170 23.980 65.370 ;
        RECT 24.230 65.260 24.520 65.370 ;
        RECT 25.620 65.170 25.870 65.710 ;
        RECT 28.700 65.710 28.970 65.770 ;
        RECT 30.250 66.050 31.560 66.310 ;
        RECT 30.250 65.710 30.560 66.050 ;
        RECT 26.260 65.180 27.900 65.570 ;
        RECT 28.700 65.420 30.560 65.710 ;
        RECT 28.700 65.410 29.010 65.420 ;
        RECT 30.250 65.410 30.560 65.420 ;
        RECT 5.660 64.850 5.930 64.930 ;
        RECT 3.060 64.620 4.500 64.830 ;
        RECT 5.050 64.630 5.930 64.850 ;
        RECT 3.060 63.570 3.340 64.620 ;
        RECT 5.050 63.820 5.270 64.630 ;
        RECT 5.660 64.600 5.930 64.630 ;
        RECT 6.790 64.890 7.080 64.940 ;
        RECT 6.790 64.710 17.540 64.890 ;
        RECT 6.790 64.610 7.080 64.710 ;
        RECT 11.630 64.700 15.260 64.710 ;
        RECT 17.340 64.030 17.540 64.710 ;
        RECT 23.730 64.570 24.020 65.170 ;
        RECT 25.620 64.570 25.910 65.170 ;
        RECT 2.340 63.120 3.340 63.570 ;
        RECT 2.320 61.670 3.620 62.120 ;
        RECT 3.320 61.270 3.620 61.670 ;
        RECT 5.040 61.290 5.270 63.820 ;
        RECT 12.290 63.730 17.540 64.030 ;
        RECT 27.960 63.960 28.260 64.960 ;
        RECT 28.710 64.360 29.010 65.410 ;
        RECT 31.310 64.310 31.560 66.050 ;
        RECT 33.680 66.040 50.640 66.360 ;
        RECT 82.630 66.060 82.810 75.720 ;
        RECT 104.060 75.540 105.080 75.990 ;
        RECT 109.670 75.830 109.960 76.430 ;
        RECT 111.560 75.830 111.850 76.430 ;
        RECT 104.780 75.530 105.080 75.540 ;
        RECT 113.900 75.220 114.200 76.220 ;
        RECT 114.650 75.620 114.950 76.670 ;
        RECT 117.250 75.570 117.500 77.310 ;
        RECT 174.700 77.240 175.490 77.430 ;
        RECT 174.700 77.040 174.950 77.240 ;
        RECT 175.200 77.130 175.490 77.240 ;
        RECT 176.590 77.040 176.840 77.580 ;
        RECT 179.670 77.580 179.940 77.640 ;
        RECT 181.220 77.920 182.530 78.180 ;
        RECT 184.670 77.930 201.450 78.210 ;
        RECT 181.220 77.580 181.530 77.920 ;
        RECT 177.230 77.050 178.870 77.440 ;
        RECT 179.670 77.290 181.530 77.580 ;
        RECT 179.670 77.280 179.980 77.290 ;
        RECT 181.220 77.280 181.530 77.290 ;
        RECT 117.950 75.220 118.210 76.770 ;
        RECT 174.700 76.440 174.990 77.040 ;
        RECT 176.590 76.440 176.880 77.040 ;
        RECT 178.930 75.830 179.230 76.830 ;
        RECT 179.680 76.230 179.980 77.280 ;
        RECT 182.280 76.180 182.530 77.920 ;
        RECT 185.390 77.880 201.450 77.930 ;
        RECT 185.390 77.870 201.120 77.880 ;
        RECT 182.980 75.830 183.240 77.380 ;
        RECT 183.940 75.830 184.120 75.840 ;
        RECT 178.880 75.530 184.130 75.830 ;
        RECT 113.850 75.210 119.100 75.220 ;
        RECT 103.730 75.130 103.980 75.140 ;
        RECT 103.730 74.670 104.710 75.130 ;
        RECT 113.850 74.920 119.120 75.210 ;
        RECT 103.730 74.370 103.980 74.670 ;
        RECT 111.700 74.580 113.540 74.590 ;
        RECT 118.950 74.580 119.120 74.920 ;
        RECT 105.440 74.570 105.680 74.580 ;
        RECT 106.520 74.570 119.120 74.580 ;
        RECT 105.440 74.410 119.120 74.570 ;
        RECT 105.440 74.400 116.950 74.410 ;
        RECT 105.430 74.390 111.750 74.400 ;
        RECT 113.300 74.390 116.950 74.400 ;
        RECT 105.430 74.380 107.300 74.390 ;
        RECT 105.430 74.370 105.680 74.380 ;
        RECT 103.730 74.200 105.680 74.370 ;
        RECT 103.730 73.900 104.000 74.200 ;
        RECT 103.740 73.640 104.000 73.900 ;
        RECT 103.720 73.250 104.020 73.640 ;
        RECT 103.710 72.850 104.020 73.250 ;
        RECT 103.700 72.090 104.010 72.850 ;
        RECT 103.600 72.070 104.010 72.090 ;
        RECT 103.570 71.120 104.020 72.070 ;
        RECT 104.430 70.830 104.890 71.770 ;
        RECT 105.630 71.180 114.900 71.190 ;
        RECT 116.780 71.180 118.700 71.190 ;
        RECT 105.630 70.990 118.700 71.180 ;
        RECT 105.630 70.980 117.990 70.990 ;
        RECT 104.470 70.510 104.770 70.830 ;
        RECT 104.470 70.180 104.760 70.510 ;
        RECT 104.480 69.380 104.740 70.180 ;
        RECT 105.630 69.970 105.840 70.980 ;
        RECT 114.890 70.970 116.790 70.980 ;
        RECT 118.520 70.240 118.700 70.990 ;
        RECT 104.480 68.780 104.730 69.380 ;
        RECT 105.630 68.960 105.830 69.970 ;
        RECT 113.440 69.940 118.700 70.240 ;
        RECT 103.690 68.330 104.730 68.780 ;
        RECT 103.670 66.880 104.630 67.330 ;
        RECT 104.380 66.830 104.630 66.880 ;
        RECT 105.640 66.830 105.830 68.960 ;
        RECT 104.380 66.630 105.830 66.830 ;
        RECT 109.360 68.300 109.620 69.500 ;
        RECT 109.360 67.790 109.610 68.300 ;
        RECT 111.250 68.290 111.510 69.500 ;
        RECT 113.640 68.390 113.890 69.940 ;
        RECT 111.250 68.130 111.640 68.290 ;
        RECT 111.240 68.000 111.640 68.130 ;
        RECT 114.340 68.000 114.600 69.610 ;
        RECT 116.890 68.540 117.190 69.590 ;
        RECT 117.640 68.990 117.940 69.940 ;
        RECT 118.140 69.040 118.440 69.090 ;
        RECT 118.140 68.690 119.040 69.040 ;
        RECT 120.750 68.910 120.970 68.920 ;
        RECT 120.750 68.720 134.430 68.910 ;
        RECT 120.750 68.590 120.970 68.720 ;
        RECT 109.860 67.790 110.150 67.950 ;
        RECT 111.240 67.940 111.500 68.000 ;
        RECT 109.360 67.600 110.150 67.790 ;
        RECT 109.360 67.400 109.610 67.600 ;
        RECT 109.860 67.490 110.150 67.600 ;
        RECT 111.250 67.400 111.500 67.940 ;
        RECT 114.330 67.940 114.600 68.000 ;
        RECT 115.880 68.280 117.190 68.540 ;
        RECT 119.290 68.290 120.970 68.590 ;
        RECT 119.290 68.280 120.950 68.290 ;
        RECT 115.880 67.940 116.190 68.280 ;
        RECT 111.890 67.410 113.530 67.800 ;
        RECT 114.330 67.650 116.190 67.940 ;
        RECT 114.330 67.640 114.640 67.650 ;
        RECT 115.880 67.640 116.190 67.650 ;
        RECT 109.360 66.800 109.650 67.400 ;
        RECT 111.250 66.800 111.540 67.400 ;
        RECT 104.380 66.540 104.630 66.630 ;
        RECT 103.650 66.090 104.630 66.540 ;
        RECT 113.590 66.190 113.890 67.190 ;
        RECT 114.340 66.590 114.640 67.640 ;
        RECT 116.940 66.540 117.190 68.280 ;
        RECT 134.180 67.820 134.430 68.720 ;
        RECT 117.640 66.190 117.900 67.740 ;
        RECT 129.120 67.520 134.430 67.820 ;
        RECT 113.540 66.170 118.790 66.190 ;
        RECT 34.560 66.030 50.640 66.040 ;
        RECT 34.560 66.000 46.540 66.030 ;
        RECT 34.560 65.990 35.450 66.000 ;
        RECT 32.010 63.960 32.270 65.510 ;
        RECT 33.100 63.960 33.300 63.970 ;
        RECT 4.110 61.270 5.270 61.290 ;
        RECT 3.320 61.090 5.270 61.270 ;
        RECT 8.210 62.090 8.470 63.290 ;
        RECT 8.210 61.580 8.460 62.090 ;
        RECT 10.100 62.080 10.360 63.290 ;
        RECT 12.490 62.180 12.740 63.730 ;
        RECT 10.100 61.920 10.490 62.080 ;
        RECT 10.090 61.790 10.490 61.920 ;
        RECT 13.190 61.790 13.450 63.400 ;
        RECT 15.740 62.330 16.040 63.380 ;
        RECT 16.490 62.780 16.790 63.730 ;
        RECT 17.340 63.720 17.540 63.730 ;
        RECT 27.910 63.660 33.300 63.960 ;
        RECT 16.990 62.830 17.290 62.880 ;
        RECT 16.990 62.480 17.890 62.830 ;
        RECT 33.100 62.420 33.300 63.660 ;
        RECT 50.260 62.460 50.620 66.030 ;
        RECT 25.540 62.400 26.730 62.410 ;
        RECT 27.720 62.400 28.910 62.410 ;
        RECT 29.940 62.400 31.130 62.410 ;
        RECT 32.120 62.400 33.310 62.420 ;
        RECT 23.330 62.390 33.310 62.400 ;
        RECT 19.940 62.370 21.130 62.380 ;
        RECT 22.220 62.370 33.310 62.390 ;
        RECT 8.710 61.580 9.000 61.740 ;
        RECT 10.090 61.730 10.350 61.790 ;
        RECT 8.210 61.390 9.000 61.580 ;
        RECT 8.210 61.190 8.460 61.390 ;
        RECT 8.710 61.280 9.000 61.390 ;
        RECT 10.100 61.190 10.350 61.730 ;
        RECT 13.180 61.730 13.450 61.790 ;
        RECT 14.730 62.070 16.040 62.330 ;
        RECT 18.100 62.140 33.310 62.370 ;
        RECT 45.390 62.160 50.640 62.460 ;
        RECT 18.100 62.130 32.260 62.140 ;
        RECT 18.100 62.120 25.630 62.130 ;
        RECT 26.640 62.120 27.830 62.130 ;
        RECT 28.790 62.120 29.980 62.130 ;
        RECT 31.070 62.120 32.260 62.130 ;
        RECT 18.100 62.110 23.410 62.120 ;
        RECT 18.100 62.100 22.270 62.110 ;
        RECT 18.100 62.090 19.990 62.100 ;
        RECT 21.080 62.090 22.270 62.100 ;
        RECT 18.100 62.080 18.820 62.090 ;
        RECT 14.730 61.730 15.040 62.070 ;
        RECT 10.740 61.200 12.380 61.590 ;
        RECT 13.180 61.440 15.040 61.730 ;
        RECT 13.180 61.430 13.490 61.440 ;
        RECT 14.730 61.430 15.040 61.440 ;
        RECT 3.320 61.080 3.970 61.090 ;
        RECT 3.320 60.750 3.620 61.080 ;
        RECT 2.600 60.300 3.620 60.750 ;
        RECT 8.210 60.590 8.500 61.190 ;
        RECT 10.100 60.590 10.390 61.190 ;
        RECT 3.320 60.290 3.620 60.300 ;
        RECT 12.440 59.980 12.740 60.980 ;
        RECT 13.190 60.380 13.490 61.430 ;
        RECT 15.790 60.330 16.040 62.070 ;
        RECT 16.490 59.980 16.750 61.530 ;
        RECT 41.310 60.520 41.570 61.720 ;
        RECT 41.310 60.010 41.560 60.520 ;
        RECT 43.200 60.510 43.460 61.720 ;
        RECT 45.590 60.610 45.840 62.160 ;
        RECT 43.200 60.350 43.590 60.510 ;
        RECT 43.190 60.220 43.590 60.350 ;
        RECT 46.290 60.220 46.550 61.830 ;
        RECT 48.840 60.760 49.140 61.810 ;
        RECT 49.590 61.210 49.890 62.160 ;
        RECT 50.090 61.260 50.390 61.310 ;
        RECT 50.090 60.910 50.990 61.260 ;
        RECT 41.810 60.010 42.100 60.170 ;
        RECT 43.190 60.160 43.450 60.220 ;
        RECT 12.390 59.970 17.640 59.980 ;
        RECT 2.270 59.890 2.520 59.900 ;
        RECT 2.270 59.430 3.250 59.890 ;
        RECT 12.390 59.680 17.660 59.970 ;
        RECT 2.270 59.130 2.520 59.430 ;
        RECT 10.240 59.340 12.080 59.350 ;
        RECT 17.490 59.340 17.660 59.680 ;
        RECT 3.980 59.330 4.220 59.340 ;
        RECT 5.060 59.330 17.660 59.340 ;
        RECT 3.980 59.170 17.660 59.330 ;
        RECT 41.310 59.820 42.100 60.010 ;
        RECT 41.310 59.620 41.560 59.820 ;
        RECT 41.810 59.710 42.100 59.820 ;
        RECT 43.200 59.620 43.450 60.160 ;
        RECT 46.280 60.160 46.550 60.220 ;
        RECT 47.830 60.500 49.140 60.760 ;
        RECT 51.200 60.800 52.870 60.830 ;
        RECT 67.950 60.800 68.200 60.810 ;
        RECT 51.200 60.530 68.200 60.800 ;
        RECT 51.200 60.520 64.700 60.530 ;
        RECT 52.480 60.500 64.700 60.520 ;
        RECT 47.830 60.160 48.140 60.500 ;
        RECT 43.840 59.630 45.480 60.020 ;
        RECT 46.280 59.870 48.140 60.160 ;
        RECT 46.280 59.860 46.590 59.870 ;
        RECT 47.830 59.860 48.140 59.870 ;
        RECT 3.980 59.160 15.490 59.170 ;
        RECT 3.970 59.150 10.290 59.160 ;
        RECT 11.840 59.150 15.490 59.160 ;
        RECT 3.970 59.140 5.840 59.150 ;
        RECT 3.970 59.130 4.220 59.140 ;
        RECT 2.270 58.960 4.220 59.130 ;
        RECT 41.310 59.020 41.600 59.620 ;
        RECT 43.200 59.020 43.490 59.620 ;
        RECT 2.270 58.740 2.520 58.960 ;
        RECT 2.270 58.570 3.310 58.740 ;
        RECT 3.120 57.710 3.310 58.570 ;
        RECT 45.540 58.410 45.840 59.410 ;
        RECT 46.290 58.810 46.590 59.860 ;
        RECT 48.890 58.760 49.140 60.500 ;
        RECT 49.590 58.410 49.850 59.960 ;
        RECT 50.470 58.410 50.810 58.480 ;
        RECT 45.490 58.110 50.810 58.410 ;
        RECT 2.330 57.270 3.310 57.710 ;
        RECT 2.330 57.260 3.280 57.270 ;
        RECT 4.150 56.950 13.420 56.960 ;
        RECT 15.300 56.950 17.220 56.960 ;
        RECT 2.000 56.850 2.190 56.860 ;
        RECT 2.000 56.390 2.980 56.850 ;
        RECT 4.150 56.760 17.220 56.950 ;
        RECT 4.150 56.750 16.510 56.760 ;
        RECT 2.000 55.600 2.190 56.390 ;
        RECT 4.150 55.740 4.360 56.750 ;
        RECT 13.410 56.740 15.310 56.750 ;
        RECT 17.040 56.010 17.220 56.760 ;
        RECT 3.000 55.600 3.270 55.610 ;
        RECT 2.000 55.390 3.270 55.600 ;
        RECT 3.000 55.180 3.270 55.390 ;
        RECT 3.000 54.550 3.250 55.180 ;
        RECT 4.150 54.730 4.350 55.740 ;
        RECT 11.960 55.710 17.220 56.010 ;
        RECT 2.210 54.100 3.250 54.550 ;
        RECT 2.190 52.650 3.150 53.100 ;
        RECT 2.900 52.600 3.150 52.650 ;
        RECT 4.160 52.600 4.350 54.730 ;
        RECT 2.900 52.400 4.350 52.600 ;
        RECT 7.880 54.070 8.140 55.270 ;
        RECT 7.880 53.560 8.130 54.070 ;
        RECT 9.770 54.060 10.030 55.270 ;
        RECT 12.160 54.160 12.410 55.710 ;
        RECT 9.770 53.900 10.160 54.060 ;
        RECT 9.760 53.770 10.160 53.900 ;
        RECT 12.860 53.770 13.120 55.380 ;
        RECT 15.410 54.310 15.710 55.360 ;
        RECT 16.160 54.760 16.460 55.710 ;
        RECT 16.660 54.810 16.960 54.860 ;
        RECT 16.660 54.460 17.560 54.810 ;
        RECT 19.270 54.680 19.490 54.690 ;
        RECT 19.270 54.490 32.950 54.680 ;
        RECT 19.270 54.360 19.490 54.490 ;
        RECT 8.380 53.560 8.670 53.720 ;
        RECT 9.760 53.710 10.020 53.770 ;
        RECT 7.880 53.370 8.670 53.560 ;
        RECT 7.880 53.170 8.130 53.370 ;
        RECT 8.380 53.260 8.670 53.370 ;
        RECT 9.770 53.170 10.020 53.710 ;
        RECT 12.850 53.710 13.120 53.770 ;
        RECT 14.400 54.050 15.710 54.310 ;
        RECT 17.810 54.060 19.490 54.360 ;
        RECT 17.810 54.050 19.470 54.060 ;
        RECT 14.400 53.710 14.710 54.050 ;
        RECT 10.410 53.180 12.050 53.570 ;
        RECT 12.850 53.420 14.710 53.710 ;
        RECT 12.850 53.410 13.160 53.420 ;
        RECT 14.400 53.410 14.710 53.420 ;
        RECT 7.880 52.570 8.170 53.170 ;
        RECT 9.770 52.570 10.060 53.170 ;
        RECT 2.900 52.310 3.150 52.400 ;
        RECT 2.170 51.860 3.150 52.310 ;
        RECT 12.110 51.960 12.410 52.960 ;
        RECT 12.860 52.360 13.160 53.410 ;
        RECT 15.460 52.310 15.710 54.050 ;
        RECT 32.700 53.590 32.950 54.490 ;
        RECT 16.160 51.960 16.420 53.510 ;
        RECT 27.640 53.290 32.950 53.590 ;
        RECT 12.060 51.940 17.310 51.960 ;
        RECT 12.060 51.660 17.430 51.940 ;
        RECT 5.510 51.260 5.790 51.330 ;
        RECT 6.690 51.290 6.970 51.320 ;
        RECT 17.140 51.290 17.430 51.660 ;
        RECT 6.690 51.280 17.430 51.290 ;
        RECT 4.100 51.060 5.790 51.260 ;
        RECT 2.890 50.860 3.170 50.870 ;
        RECT 2.150 50.410 3.170 50.860 ;
        RECT 4.100 50.410 4.330 51.060 ;
        RECT 5.510 51.000 5.790 51.060 ;
        RECT 6.670 51.050 17.430 51.280 ;
        RECT 6.690 51.040 17.430 51.050 ;
        RECT 23.560 51.650 23.820 52.850 ;
        RECT 23.560 51.140 23.810 51.650 ;
        RECT 25.450 51.640 25.710 52.850 ;
        RECT 27.840 51.740 28.090 53.290 ;
        RECT 25.450 51.480 25.840 51.640 ;
        RECT 25.440 51.350 25.840 51.480 ;
        RECT 28.540 51.350 28.800 52.960 ;
        RECT 31.090 51.890 31.390 52.940 ;
        RECT 31.840 52.340 32.140 53.290 ;
        RECT 32.340 52.390 32.640 52.440 ;
        RECT 32.340 52.040 33.240 52.390 ;
        RECT 50.470 51.990 50.810 58.110 ;
        RECT 49.900 51.970 50.860 51.990 ;
        RECT 34.380 51.950 38.660 51.960 ;
        RECT 46.060 51.950 50.860 51.970 ;
        RECT 34.380 51.940 50.860 51.950 ;
        RECT 24.060 51.140 24.350 51.300 ;
        RECT 25.440 51.290 25.700 51.350 ;
        RECT 6.690 51.030 17.390 51.040 ;
        RECT 6.690 50.990 6.970 51.030 ;
        RECT 23.560 50.950 24.350 51.140 ;
        RECT 23.560 50.750 23.810 50.950 ;
        RECT 24.060 50.840 24.350 50.950 ;
        RECT 25.450 50.750 25.700 51.290 ;
        RECT 28.530 51.290 28.800 51.350 ;
        RECT 30.080 51.630 31.390 51.890 ;
        RECT 30.080 51.290 30.390 51.630 ;
        RECT 26.090 50.760 27.730 51.150 ;
        RECT 28.530 51.000 30.390 51.290 ;
        RECT 28.530 50.990 28.840 51.000 ;
        RECT 30.080 50.990 30.390 51.000 ;
        RECT 5.490 50.430 5.760 50.510 ;
        RECT 2.890 50.200 4.330 50.410 ;
        RECT 4.880 50.210 5.760 50.430 ;
        RECT 2.890 49.150 3.170 50.200 ;
        RECT 4.880 49.400 5.100 50.210 ;
        RECT 5.490 50.180 5.760 50.210 ;
        RECT 6.620 50.470 6.910 50.520 ;
        RECT 6.620 50.290 17.370 50.470 ;
        RECT 6.620 50.190 6.910 50.290 ;
        RECT 11.460 50.280 15.090 50.290 ;
        RECT 17.170 49.610 17.370 50.290 ;
        RECT 23.560 50.150 23.850 50.750 ;
        RECT 25.450 50.150 25.740 50.750 ;
        RECT 2.170 48.700 3.170 49.150 ;
        RECT 2.150 47.250 3.450 47.700 ;
        RECT 3.150 46.850 3.450 47.250 ;
        RECT 4.870 46.870 5.100 49.400 ;
        RECT 12.120 49.310 17.370 49.610 ;
        RECT 27.790 49.540 28.090 50.540 ;
        RECT 28.540 49.940 28.840 50.990 ;
        RECT 31.140 49.890 31.390 51.630 ;
        RECT 33.510 51.630 50.860 51.940 ;
        RECT 33.510 51.620 46.520 51.630 ;
        RECT 38.370 51.610 46.520 51.620 ;
        RECT 49.900 51.590 50.860 51.630 ;
        RECT 50.470 51.580 50.810 51.590 ;
        RECT 31.840 49.540 32.100 51.090 ;
        RECT 32.930 49.540 33.130 49.550 ;
        RECT 3.940 46.850 5.100 46.870 ;
        RECT 3.150 46.670 5.100 46.850 ;
        RECT 8.040 47.670 8.300 48.870 ;
        RECT 8.040 47.160 8.290 47.670 ;
        RECT 9.930 47.660 10.190 48.870 ;
        RECT 12.320 47.760 12.570 49.310 ;
        RECT 9.930 47.500 10.320 47.660 ;
        RECT 9.920 47.370 10.320 47.500 ;
        RECT 13.020 47.370 13.280 48.980 ;
        RECT 15.570 47.910 15.870 48.960 ;
        RECT 16.320 48.360 16.620 49.310 ;
        RECT 17.170 49.300 17.370 49.310 ;
        RECT 27.740 49.240 33.130 49.540 ;
        RECT 16.820 48.410 17.120 48.460 ;
        RECT 16.820 48.060 17.720 48.410 ;
        RECT 32.930 48.000 33.130 49.240 ;
        RECT 25.370 47.980 26.560 47.990 ;
        RECT 27.550 47.980 28.740 47.990 ;
        RECT 29.770 47.980 30.960 47.990 ;
        RECT 31.950 47.980 33.140 48.000 ;
        RECT 23.160 47.970 33.140 47.980 ;
        RECT 19.770 47.950 20.960 47.960 ;
        RECT 22.050 47.950 33.140 47.970 ;
        RECT 8.540 47.160 8.830 47.320 ;
        RECT 9.920 47.310 10.180 47.370 ;
        RECT 8.040 46.970 8.830 47.160 ;
        RECT 8.040 46.770 8.290 46.970 ;
        RECT 8.540 46.860 8.830 46.970 ;
        RECT 9.930 46.770 10.180 47.310 ;
        RECT 13.010 47.310 13.280 47.370 ;
        RECT 14.560 47.650 15.870 47.910 ;
        RECT 17.930 47.720 33.140 47.950 ;
        RECT 17.930 47.710 32.090 47.720 ;
        RECT 17.930 47.700 25.460 47.710 ;
        RECT 26.470 47.700 27.660 47.710 ;
        RECT 28.620 47.700 29.810 47.710 ;
        RECT 30.900 47.700 32.090 47.710 ;
        RECT 17.930 47.690 23.240 47.700 ;
        RECT 17.930 47.680 22.100 47.690 ;
        RECT 17.930 47.670 19.820 47.680 ;
        RECT 20.910 47.670 22.100 47.680 ;
        RECT 17.930 47.660 18.650 47.670 ;
        RECT 14.560 47.310 14.870 47.650 ;
        RECT 10.570 46.780 12.210 47.170 ;
        RECT 13.010 47.020 14.870 47.310 ;
        RECT 13.010 47.010 13.320 47.020 ;
        RECT 14.560 47.010 14.870 47.020 ;
        RECT 3.150 46.660 3.800 46.670 ;
        RECT 3.150 46.330 3.450 46.660 ;
        RECT 2.430 45.880 3.450 46.330 ;
        RECT 8.040 46.170 8.330 46.770 ;
        RECT 9.930 46.170 10.220 46.770 ;
        RECT 3.150 45.870 3.450 45.880 ;
        RECT 12.270 45.560 12.570 46.560 ;
        RECT 13.020 45.960 13.320 47.010 ;
        RECT 15.620 45.910 15.870 47.650 ;
        RECT 67.950 47.390 68.210 60.530 ;
        RECT 67.940 47.270 68.210 47.390 ;
        RECT 82.540 56.540 82.810 66.060 ;
        RECT 113.540 65.890 118.910 66.170 ;
        RECT 106.990 65.490 107.270 65.560 ;
        RECT 108.170 65.520 108.450 65.550 ;
        RECT 118.620 65.520 118.910 65.890 ;
        RECT 108.170 65.510 118.910 65.520 ;
        RECT 105.580 65.290 107.270 65.490 ;
        RECT 104.370 65.090 104.650 65.100 ;
        RECT 103.630 64.640 104.650 65.090 ;
        RECT 105.580 64.640 105.810 65.290 ;
        RECT 106.990 65.230 107.270 65.290 ;
        RECT 108.150 65.280 118.910 65.510 ;
        RECT 108.170 65.270 118.910 65.280 ;
        RECT 125.040 65.880 125.300 67.080 ;
        RECT 125.040 65.370 125.290 65.880 ;
        RECT 126.930 65.870 127.190 67.080 ;
        RECT 129.320 65.970 129.570 67.520 ;
        RECT 126.930 65.710 127.320 65.870 ;
        RECT 126.920 65.580 127.320 65.710 ;
        RECT 130.020 65.580 130.280 67.190 ;
        RECT 132.570 66.120 132.870 67.170 ;
        RECT 133.320 66.570 133.620 67.520 ;
        RECT 133.820 66.620 134.120 66.670 ;
        RECT 133.820 66.270 134.720 66.620 ;
        RECT 147.480 66.220 151.950 66.250 ;
        RECT 136.540 66.190 151.950 66.220 ;
        RECT 135.870 66.170 151.950 66.190 ;
        RECT 125.540 65.370 125.830 65.530 ;
        RECT 126.920 65.520 127.180 65.580 ;
        RECT 108.170 65.260 118.870 65.270 ;
        RECT 108.170 65.220 108.450 65.260 ;
        RECT 125.040 65.180 125.830 65.370 ;
        RECT 125.040 64.980 125.290 65.180 ;
        RECT 125.540 65.070 125.830 65.180 ;
        RECT 126.930 64.980 127.180 65.520 ;
        RECT 130.010 65.520 130.280 65.580 ;
        RECT 131.560 65.860 132.870 66.120 ;
        RECT 131.560 65.520 131.870 65.860 ;
        RECT 127.570 64.990 129.210 65.380 ;
        RECT 130.010 65.230 131.870 65.520 ;
        RECT 130.010 65.220 130.320 65.230 ;
        RECT 131.560 65.220 131.870 65.230 ;
        RECT 106.970 64.660 107.240 64.740 ;
        RECT 104.370 64.430 105.810 64.640 ;
        RECT 106.360 64.440 107.240 64.660 ;
        RECT 104.370 63.380 104.650 64.430 ;
        RECT 106.360 63.630 106.580 64.440 ;
        RECT 106.970 64.410 107.240 64.440 ;
        RECT 108.100 64.700 108.390 64.750 ;
        RECT 108.100 64.520 118.850 64.700 ;
        RECT 108.100 64.420 108.390 64.520 ;
        RECT 112.940 64.510 116.570 64.520 ;
        RECT 118.650 63.840 118.850 64.520 ;
        RECT 125.040 64.380 125.330 64.980 ;
        RECT 126.930 64.380 127.220 64.980 ;
        RECT 103.650 62.930 104.650 63.380 ;
        RECT 103.630 61.480 104.930 61.930 ;
        RECT 104.630 61.080 104.930 61.480 ;
        RECT 106.350 61.100 106.580 63.630 ;
        RECT 113.600 63.540 118.850 63.840 ;
        RECT 129.270 63.770 129.570 64.770 ;
        RECT 130.020 64.170 130.320 65.220 ;
        RECT 132.620 64.120 132.870 65.860 ;
        RECT 134.990 65.850 151.950 66.170 ;
        RECT 183.940 65.870 184.120 75.530 ;
        RECT 135.870 65.840 151.950 65.850 ;
        RECT 135.870 65.810 147.850 65.840 ;
        RECT 135.870 65.800 136.760 65.810 ;
        RECT 133.320 63.770 133.580 65.320 ;
        RECT 134.410 63.770 134.610 63.780 ;
        RECT 105.420 61.080 106.580 61.100 ;
        RECT 104.630 60.900 106.580 61.080 ;
        RECT 109.520 61.900 109.780 63.100 ;
        RECT 109.520 61.390 109.770 61.900 ;
        RECT 111.410 61.890 111.670 63.100 ;
        RECT 113.800 61.990 114.050 63.540 ;
        RECT 111.410 61.730 111.800 61.890 ;
        RECT 111.400 61.600 111.800 61.730 ;
        RECT 114.500 61.600 114.760 63.210 ;
        RECT 117.050 62.140 117.350 63.190 ;
        RECT 117.800 62.590 118.100 63.540 ;
        RECT 118.650 63.530 118.850 63.540 ;
        RECT 129.220 63.470 134.610 63.770 ;
        RECT 118.300 62.640 118.600 62.690 ;
        RECT 118.300 62.290 119.200 62.640 ;
        RECT 134.410 62.230 134.610 63.470 ;
        RECT 151.570 62.270 151.930 65.840 ;
        RECT 126.850 62.210 128.040 62.220 ;
        RECT 129.030 62.210 130.220 62.220 ;
        RECT 131.250 62.210 132.440 62.220 ;
        RECT 133.430 62.210 134.620 62.230 ;
        RECT 124.640 62.200 134.620 62.210 ;
        RECT 121.250 62.180 122.440 62.190 ;
        RECT 123.530 62.180 134.620 62.200 ;
        RECT 110.020 61.390 110.310 61.550 ;
        RECT 111.400 61.540 111.660 61.600 ;
        RECT 109.520 61.200 110.310 61.390 ;
        RECT 109.520 61.000 109.770 61.200 ;
        RECT 110.020 61.090 110.310 61.200 ;
        RECT 111.410 61.000 111.660 61.540 ;
        RECT 114.490 61.540 114.760 61.600 ;
        RECT 116.040 61.880 117.350 62.140 ;
        RECT 119.410 61.950 134.620 62.180 ;
        RECT 146.700 61.970 151.950 62.270 ;
        RECT 119.410 61.940 133.570 61.950 ;
        RECT 119.410 61.930 126.940 61.940 ;
        RECT 127.950 61.930 129.140 61.940 ;
        RECT 130.100 61.930 131.290 61.940 ;
        RECT 132.380 61.930 133.570 61.940 ;
        RECT 119.410 61.920 124.720 61.930 ;
        RECT 119.410 61.910 123.580 61.920 ;
        RECT 119.410 61.900 121.300 61.910 ;
        RECT 122.390 61.900 123.580 61.910 ;
        RECT 119.410 61.890 120.130 61.900 ;
        RECT 116.040 61.540 116.350 61.880 ;
        RECT 112.050 61.010 113.690 61.400 ;
        RECT 114.490 61.250 116.350 61.540 ;
        RECT 114.490 61.240 114.800 61.250 ;
        RECT 116.040 61.240 116.350 61.250 ;
        RECT 104.630 60.890 105.280 60.900 ;
        RECT 104.630 60.560 104.930 60.890 ;
        RECT 103.910 60.110 104.930 60.560 ;
        RECT 109.520 60.400 109.810 61.000 ;
        RECT 111.410 60.400 111.700 61.000 ;
        RECT 104.630 60.100 104.930 60.110 ;
        RECT 113.750 59.790 114.050 60.790 ;
        RECT 114.500 60.190 114.800 61.240 ;
        RECT 117.100 60.140 117.350 61.880 ;
        RECT 117.800 59.790 118.060 61.340 ;
        RECT 142.620 60.330 142.880 61.530 ;
        RECT 142.620 59.820 142.870 60.330 ;
        RECT 144.510 60.320 144.770 61.530 ;
        RECT 146.900 60.420 147.150 61.970 ;
        RECT 144.510 60.160 144.900 60.320 ;
        RECT 144.500 60.030 144.900 60.160 ;
        RECT 147.600 60.030 147.860 61.640 ;
        RECT 150.150 60.570 150.450 61.620 ;
        RECT 150.900 61.020 151.200 61.970 ;
        RECT 151.400 61.070 151.700 61.120 ;
        RECT 151.400 60.720 152.300 61.070 ;
        RECT 143.120 59.820 143.410 59.980 ;
        RECT 144.500 59.970 144.760 60.030 ;
        RECT 113.700 59.780 118.950 59.790 ;
        RECT 103.580 59.700 103.830 59.710 ;
        RECT 103.580 59.240 104.560 59.700 ;
        RECT 113.700 59.490 118.970 59.780 ;
        RECT 103.580 58.940 103.830 59.240 ;
        RECT 111.550 59.150 113.390 59.160 ;
        RECT 118.800 59.150 118.970 59.490 ;
        RECT 105.290 59.140 105.530 59.150 ;
        RECT 106.370 59.140 118.970 59.150 ;
        RECT 105.290 58.980 118.970 59.140 ;
        RECT 142.620 59.630 143.410 59.820 ;
        RECT 142.620 59.430 142.870 59.630 ;
        RECT 143.120 59.520 143.410 59.630 ;
        RECT 144.510 59.430 144.760 59.970 ;
        RECT 147.590 59.970 147.860 60.030 ;
        RECT 149.140 60.310 150.450 60.570 ;
        RECT 152.510 60.610 154.180 60.640 ;
        RECT 169.260 60.610 169.510 60.620 ;
        RECT 152.510 60.340 169.510 60.610 ;
        RECT 152.510 60.330 166.010 60.340 ;
        RECT 153.790 60.310 166.010 60.330 ;
        RECT 149.140 59.970 149.450 60.310 ;
        RECT 145.150 59.440 146.790 59.830 ;
        RECT 147.590 59.680 149.450 59.970 ;
        RECT 147.590 59.670 147.900 59.680 ;
        RECT 149.140 59.670 149.450 59.680 ;
        RECT 105.290 58.970 116.800 58.980 ;
        RECT 105.280 58.960 111.600 58.970 ;
        RECT 113.150 58.960 116.800 58.970 ;
        RECT 105.280 58.950 107.150 58.960 ;
        RECT 105.280 58.940 105.530 58.950 ;
        RECT 103.580 58.770 105.530 58.940 ;
        RECT 142.620 58.830 142.910 59.430 ;
        RECT 144.510 58.830 144.800 59.430 ;
        RECT 103.580 58.550 103.830 58.770 ;
        RECT 103.580 58.380 104.620 58.550 ;
        RECT 104.430 57.520 104.620 58.380 ;
        RECT 146.850 58.220 147.150 59.220 ;
        RECT 147.600 58.620 147.900 59.670 ;
        RECT 150.200 58.570 150.450 60.310 ;
        RECT 150.900 58.220 151.160 59.770 ;
        RECT 151.780 58.220 152.120 58.290 ;
        RECT 146.800 57.920 152.120 58.220 ;
        RECT 103.640 57.080 104.620 57.520 ;
        RECT 103.640 57.070 104.590 57.080 ;
        RECT 105.460 56.760 114.730 56.770 ;
        RECT 116.610 56.760 118.530 56.770 ;
        RECT 103.310 56.660 103.500 56.670 ;
        RECT 16.320 45.560 16.580 47.110 ;
        RECT 67.940 46.440 68.200 47.270 ;
        RECT 82.540 46.590 82.720 56.540 ;
        RECT 103.310 56.200 104.290 56.660 ;
        RECT 105.460 56.570 118.530 56.760 ;
        RECT 105.460 56.560 117.820 56.570 ;
        RECT 103.310 55.410 103.500 56.200 ;
        RECT 105.460 55.550 105.670 56.560 ;
        RECT 114.720 56.550 116.620 56.560 ;
        RECT 118.350 55.820 118.530 56.570 ;
        RECT 104.310 55.410 104.580 55.420 ;
        RECT 103.310 55.200 104.580 55.410 ;
        RECT 104.310 54.990 104.580 55.200 ;
        RECT 104.310 54.360 104.560 54.990 ;
        RECT 105.460 54.540 105.660 55.550 ;
        RECT 113.270 55.520 118.530 55.820 ;
        RECT 103.520 53.910 104.560 54.360 ;
        RECT 103.500 52.460 104.460 52.910 ;
        RECT 104.210 52.410 104.460 52.460 ;
        RECT 105.470 52.410 105.660 54.540 ;
        RECT 104.210 52.210 105.660 52.410 ;
        RECT 109.190 53.880 109.450 55.080 ;
        RECT 109.190 53.370 109.440 53.880 ;
        RECT 111.080 53.870 111.340 55.080 ;
        RECT 113.470 53.970 113.720 55.520 ;
        RECT 111.080 53.710 111.470 53.870 ;
        RECT 111.070 53.580 111.470 53.710 ;
        RECT 114.170 53.580 114.430 55.190 ;
        RECT 116.720 54.120 117.020 55.170 ;
        RECT 117.470 54.570 117.770 55.520 ;
        RECT 117.970 54.620 118.270 54.670 ;
        RECT 117.970 54.270 118.870 54.620 ;
        RECT 120.580 54.490 120.800 54.500 ;
        RECT 120.580 54.300 134.260 54.490 ;
        RECT 120.580 54.170 120.800 54.300 ;
        RECT 109.690 53.370 109.980 53.530 ;
        RECT 111.070 53.520 111.330 53.580 ;
        RECT 109.190 53.180 109.980 53.370 ;
        RECT 109.190 52.980 109.440 53.180 ;
        RECT 109.690 53.070 109.980 53.180 ;
        RECT 111.080 52.980 111.330 53.520 ;
        RECT 114.160 53.520 114.430 53.580 ;
        RECT 115.710 53.860 117.020 54.120 ;
        RECT 119.120 53.870 120.800 54.170 ;
        RECT 119.120 53.860 120.780 53.870 ;
        RECT 115.710 53.520 116.020 53.860 ;
        RECT 111.720 52.990 113.360 53.380 ;
        RECT 114.160 53.230 116.020 53.520 ;
        RECT 114.160 53.220 114.470 53.230 ;
        RECT 115.710 53.220 116.020 53.230 ;
        RECT 109.190 52.380 109.480 52.980 ;
        RECT 111.080 52.380 111.370 52.980 ;
        RECT 104.210 52.120 104.460 52.210 ;
        RECT 103.480 51.670 104.460 52.120 ;
        RECT 113.420 51.770 113.720 52.770 ;
        RECT 114.170 52.170 114.470 53.220 ;
        RECT 116.770 52.120 117.020 53.860 ;
        RECT 134.010 53.400 134.260 54.300 ;
        RECT 117.470 51.770 117.730 53.320 ;
        RECT 128.950 53.100 134.260 53.400 ;
        RECT 113.370 51.750 118.620 51.770 ;
        RECT 113.370 51.470 118.740 51.750 ;
        RECT 106.820 51.070 107.100 51.140 ;
        RECT 108.000 51.100 108.280 51.130 ;
        RECT 118.450 51.100 118.740 51.470 ;
        RECT 108.000 51.090 118.740 51.100 ;
        RECT 105.410 50.870 107.100 51.070 ;
        RECT 104.200 50.670 104.480 50.680 ;
        RECT 103.460 50.220 104.480 50.670 ;
        RECT 105.410 50.220 105.640 50.870 ;
        RECT 106.820 50.810 107.100 50.870 ;
        RECT 107.980 50.860 118.740 51.090 ;
        RECT 108.000 50.850 118.740 50.860 ;
        RECT 124.870 51.460 125.130 52.660 ;
        RECT 124.870 50.950 125.120 51.460 ;
        RECT 126.760 51.450 127.020 52.660 ;
        RECT 129.150 51.550 129.400 53.100 ;
        RECT 126.760 51.290 127.150 51.450 ;
        RECT 126.750 51.160 127.150 51.290 ;
        RECT 129.850 51.160 130.110 52.770 ;
        RECT 132.400 51.700 132.700 52.750 ;
        RECT 133.150 52.150 133.450 53.100 ;
        RECT 133.650 52.200 133.950 52.250 ;
        RECT 133.650 51.850 134.550 52.200 ;
        RECT 151.780 51.800 152.120 57.920 ;
        RECT 151.210 51.780 152.170 51.800 ;
        RECT 135.690 51.760 139.970 51.770 ;
        RECT 147.370 51.760 152.170 51.780 ;
        RECT 135.690 51.750 152.170 51.760 ;
        RECT 125.370 50.950 125.660 51.110 ;
        RECT 126.750 51.100 127.010 51.160 ;
        RECT 108.000 50.840 118.700 50.850 ;
        RECT 108.000 50.800 108.280 50.840 ;
        RECT 124.870 50.760 125.660 50.950 ;
        RECT 124.870 50.560 125.120 50.760 ;
        RECT 125.370 50.650 125.660 50.760 ;
        RECT 126.760 50.560 127.010 51.100 ;
        RECT 129.840 51.100 130.110 51.160 ;
        RECT 131.390 51.440 132.700 51.700 ;
        RECT 131.390 51.100 131.700 51.440 ;
        RECT 127.400 50.570 129.040 50.960 ;
        RECT 129.840 50.810 131.700 51.100 ;
        RECT 129.840 50.800 130.150 50.810 ;
        RECT 131.390 50.800 131.700 50.810 ;
        RECT 106.800 50.240 107.070 50.320 ;
        RECT 104.200 50.010 105.640 50.220 ;
        RECT 106.190 50.020 107.070 50.240 ;
        RECT 104.200 48.960 104.480 50.010 ;
        RECT 106.190 49.210 106.410 50.020 ;
        RECT 106.800 49.990 107.070 50.020 ;
        RECT 107.930 50.280 108.220 50.330 ;
        RECT 107.930 50.100 118.680 50.280 ;
        RECT 107.930 50.000 108.220 50.100 ;
        RECT 112.770 50.090 116.400 50.100 ;
        RECT 118.480 49.420 118.680 50.100 ;
        RECT 124.870 49.960 125.160 50.560 ;
        RECT 126.760 49.960 127.050 50.560 ;
        RECT 103.480 48.510 104.480 48.960 ;
        RECT 103.460 47.060 104.760 47.510 ;
        RECT 104.460 46.660 104.760 47.060 ;
        RECT 106.180 46.680 106.410 49.210 ;
        RECT 113.430 49.120 118.680 49.420 ;
        RECT 129.100 49.350 129.400 50.350 ;
        RECT 129.850 49.750 130.150 50.800 ;
        RECT 132.450 49.700 132.700 51.440 ;
        RECT 134.820 51.440 152.170 51.750 ;
        RECT 134.820 51.430 147.830 51.440 ;
        RECT 139.680 51.420 147.830 51.430 ;
        RECT 151.210 51.400 152.170 51.440 ;
        RECT 151.780 51.390 152.120 51.400 ;
        RECT 133.150 49.350 133.410 50.900 ;
        RECT 134.240 49.350 134.440 49.360 ;
        RECT 105.250 46.660 106.410 46.680 ;
        RECT 62.920 46.140 68.200 46.440 ;
        RECT 12.220 45.550 17.470 45.560 ;
        RECT 2.100 45.470 2.350 45.480 ;
        RECT 2.100 45.010 3.080 45.470 ;
        RECT 12.220 45.260 17.490 45.550 ;
        RECT 2.100 44.710 2.350 45.010 ;
        RECT 10.070 44.920 11.910 44.930 ;
        RECT 17.320 44.920 17.490 45.260 ;
        RECT 3.810 44.910 4.050 44.920 ;
        RECT 4.890 44.910 17.490 44.920 ;
        RECT 3.810 44.750 17.490 44.910 ;
        RECT 3.810 44.740 15.320 44.750 ;
        RECT 3.800 44.730 10.120 44.740 ;
        RECT 11.670 44.730 15.320 44.740 ;
        RECT 3.800 44.720 5.670 44.730 ;
        RECT 3.800 44.710 4.050 44.720 ;
        RECT 2.100 44.540 4.050 44.710 ;
        RECT 2.100 44.240 2.370 44.540 ;
        RECT 2.110 43.980 2.370 44.240 ;
        RECT 58.840 44.500 59.100 45.700 ;
        RECT 58.840 43.990 59.090 44.500 ;
        RECT 60.730 44.490 60.990 45.700 ;
        RECT 63.120 44.590 63.370 46.140 ;
        RECT 60.730 44.330 61.120 44.490 ;
        RECT 60.720 44.200 61.120 44.330 ;
        RECT 63.820 44.200 64.080 45.810 ;
        RECT 66.370 44.740 66.670 45.790 ;
        RECT 67.120 45.190 67.420 46.140 ;
        RECT 67.620 45.240 67.920 45.290 ;
        RECT 67.620 44.890 68.520 45.240 ;
        RECT 82.530 44.780 82.730 46.590 ;
        RECT 104.460 46.480 106.410 46.660 ;
        RECT 109.350 47.480 109.610 48.680 ;
        RECT 109.350 46.970 109.600 47.480 ;
        RECT 111.240 47.470 111.500 48.680 ;
        RECT 113.630 47.570 113.880 49.120 ;
        RECT 111.240 47.310 111.630 47.470 ;
        RECT 111.230 47.180 111.630 47.310 ;
        RECT 114.330 47.180 114.590 48.790 ;
        RECT 116.880 47.720 117.180 48.770 ;
        RECT 117.630 48.170 117.930 49.120 ;
        RECT 118.480 49.110 118.680 49.120 ;
        RECT 129.050 49.050 134.440 49.350 ;
        RECT 118.130 48.220 118.430 48.270 ;
        RECT 118.130 47.870 119.030 48.220 ;
        RECT 134.240 47.810 134.440 49.050 ;
        RECT 126.680 47.790 127.870 47.800 ;
        RECT 128.860 47.790 130.050 47.800 ;
        RECT 131.080 47.790 132.270 47.800 ;
        RECT 133.260 47.790 134.450 47.810 ;
        RECT 124.470 47.780 134.450 47.790 ;
        RECT 121.080 47.760 122.270 47.770 ;
        RECT 123.360 47.760 134.450 47.780 ;
        RECT 109.850 46.970 110.140 47.130 ;
        RECT 111.230 47.120 111.490 47.180 ;
        RECT 109.350 46.780 110.140 46.970 ;
        RECT 109.350 46.580 109.600 46.780 ;
        RECT 109.850 46.670 110.140 46.780 ;
        RECT 111.240 46.580 111.490 47.120 ;
        RECT 114.320 47.120 114.590 47.180 ;
        RECT 115.870 47.460 117.180 47.720 ;
        RECT 119.240 47.530 134.450 47.760 ;
        RECT 119.240 47.520 133.400 47.530 ;
        RECT 119.240 47.510 126.770 47.520 ;
        RECT 127.780 47.510 128.970 47.520 ;
        RECT 129.930 47.510 131.120 47.520 ;
        RECT 132.210 47.510 133.400 47.520 ;
        RECT 119.240 47.500 124.550 47.510 ;
        RECT 119.240 47.490 123.410 47.500 ;
        RECT 119.240 47.480 121.130 47.490 ;
        RECT 122.220 47.480 123.410 47.490 ;
        RECT 119.240 47.470 119.960 47.480 ;
        RECT 115.870 47.120 116.180 47.460 ;
        RECT 111.880 46.590 113.520 46.980 ;
        RECT 114.320 46.830 116.180 47.120 ;
        RECT 114.320 46.820 114.630 46.830 ;
        RECT 115.870 46.820 116.180 46.830 ;
        RECT 104.460 46.470 105.110 46.480 ;
        RECT 104.460 46.140 104.760 46.470 ;
        RECT 103.740 45.690 104.760 46.140 ;
        RECT 109.350 45.980 109.640 46.580 ;
        RECT 111.240 45.980 111.530 46.580 ;
        RECT 104.460 45.680 104.760 45.690 ;
        RECT 113.580 45.370 113.880 46.370 ;
        RECT 114.330 45.770 114.630 46.820 ;
        RECT 116.930 45.720 117.180 47.460 ;
        RECT 169.260 47.200 169.520 60.340 ;
        RECT 169.250 47.080 169.520 47.200 ;
        RECT 183.850 56.350 184.120 65.870 ;
        RECT 117.630 45.370 117.890 46.920 ;
        RECT 169.250 46.250 169.510 47.080 ;
        RECT 183.850 46.400 184.030 56.350 ;
        RECT 164.230 45.950 169.510 46.250 ;
        RECT 113.530 45.360 118.780 45.370 ;
        RECT 59.340 43.990 59.630 44.150 ;
        RECT 60.720 44.140 60.980 44.200 ;
        RECT 2.090 43.590 2.390 43.980 ;
        RECT 58.840 43.800 59.630 43.990 ;
        RECT 58.840 43.600 59.090 43.800 ;
        RECT 59.340 43.690 59.630 43.800 ;
        RECT 60.730 43.600 60.980 44.140 ;
        RECT 63.810 44.140 64.080 44.200 ;
        RECT 65.360 44.480 66.670 44.740 ;
        RECT 68.790 44.490 82.730 44.780 ;
        RECT 103.410 45.280 103.660 45.290 ;
        RECT 103.410 44.820 104.390 45.280 ;
        RECT 113.530 45.070 118.800 45.360 ;
        RECT 103.410 44.520 103.660 44.820 ;
        RECT 111.380 44.730 113.220 44.740 ;
        RECT 118.630 44.730 118.800 45.070 ;
        RECT 105.120 44.720 105.360 44.730 ;
        RECT 106.200 44.720 118.800 44.730 ;
        RECT 105.120 44.560 118.800 44.720 ;
        RECT 105.120 44.550 116.630 44.560 ;
        RECT 105.110 44.540 111.430 44.550 ;
        RECT 112.980 44.540 116.630 44.550 ;
        RECT 105.110 44.530 106.980 44.540 ;
        RECT 105.110 44.520 105.360 44.530 ;
        RECT 68.790 44.480 82.690 44.490 ;
        RECT 65.360 44.140 65.670 44.480 ;
        RECT 61.370 43.610 63.010 44.000 ;
        RECT 63.810 43.850 65.670 44.140 ;
        RECT 63.810 43.840 64.120 43.850 ;
        RECT 65.360 43.840 65.670 43.850 ;
        RECT 2.090 43.360 3.580 43.590 ;
        RECT 3.330 42.430 3.580 43.360 ;
        RECT 58.840 43.000 59.130 43.600 ;
        RECT 60.730 43.000 61.020 43.600 ;
        RECT 2.530 41.970 3.580 42.430 ;
        RECT 63.070 42.390 63.370 43.390 ;
        RECT 63.820 42.790 64.120 43.840 ;
        RECT 66.420 42.740 66.670 44.480 ;
        RECT 69.380 44.470 82.690 44.480 ;
        RECT 103.410 44.350 105.360 44.520 ;
        RECT 103.410 44.050 103.680 44.350 ;
        RECT 67.120 42.390 67.380 43.940 ;
        RECT 103.420 43.790 103.680 44.050 ;
        RECT 160.150 44.310 160.410 45.510 ;
        RECT 160.150 43.800 160.400 44.310 ;
        RECT 162.040 44.300 162.300 45.510 ;
        RECT 164.430 44.400 164.680 45.950 ;
        RECT 162.040 44.140 162.430 44.300 ;
        RECT 162.030 44.010 162.430 44.140 ;
        RECT 165.130 44.010 165.390 45.620 ;
        RECT 167.680 44.550 167.980 45.600 ;
        RECT 168.430 45.000 168.730 45.950 ;
        RECT 168.930 45.050 169.230 45.100 ;
        RECT 168.930 44.700 169.830 45.050 ;
        RECT 183.840 44.590 184.040 46.400 ;
        RECT 160.650 43.800 160.940 43.960 ;
        RECT 162.030 43.950 162.290 44.010 ;
        RECT 103.400 43.400 103.700 43.790 ;
        RECT 160.150 43.610 160.940 43.800 ;
        RECT 160.150 43.410 160.400 43.610 ;
        RECT 160.650 43.500 160.940 43.610 ;
        RECT 162.040 43.410 162.290 43.950 ;
        RECT 165.120 43.950 165.390 44.010 ;
        RECT 166.670 44.290 167.980 44.550 ;
        RECT 170.100 44.300 184.040 44.590 ;
        RECT 170.100 44.290 184.000 44.300 ;
        RECT 166.670 43.950 166.980 44.290 ;
        RECT 162.680 43.420 164.320 43.810 ;
        RECT 165.120 43.660 166.980 43.950 ;
        RECT 165.120 43.650 165.430 43.660 ;
        RECT 166.670 43.650 166.980 43.660 ;
        RECT 103.400 43.170 104.890 43.400 ;
        RECT 63.020 42.090 68.290 42.390 ;
        RECT 104.640 42.240 104.890 43.170 ;
        RECT 160.150 42.810 160.440 43.410 ;
        RECT 162.040 42.810 162.330 43.410 ;
        RECT 3.330 41.960 3.580 41.970 ;
        RECT 2.200 41.560 2.450 41.570 ;
        RECT 2.200 41.110 3.180 41.560 ;
        RECT 4.290 41.300 13.560 41.310 ;
        RECT 15.440 41.300 17.360 41.310 ;
        RECT 4.290 41.110 17.360 41.300 ;
        RECT 2.200 40.500 2.450 41.110 ;
        RECT 4.290 41.100 16.650 41.110 ;
        RECT 2.200 40.250 3.410 40.500 ;
        RECT 3.140 39.500 3.400 40.250 ;
        RECT 4.290 40.090 4.500 41.100 ;
        RECT 13.550 41.090 15.450 41.100 ;
        RECT 17.180 40.360 17.360 41.110 ;
        RECT 3.140 38.900 3.390 39.500 ;
        RECT 4.290 39.080 4.490 40.090 ;
        RECT 12.100 40.060 17.360 40.360 ;
        RECT 2.350 38.450 3.390 38.900 ;
        RECT 2.330 37.000 3.290 37.450 ;
        RECT 3.040 36.950 3.290 37.000 ;
        RECT 4.300 36.950 4.490 39.080 ;
        RECT 3.040 36.750 4.490 36.950 ;
        RECT 8.020 38.420 8.280 39.620 ;
        RECT 8.020 37.910 8.270 38.420 ;
        RECT 9.910 38.410 10.170 39.620 ;
        RECT 12.300 38.510 12.550 40.060 ;
        RECT 9.910 38.250 10.300 38.410 ;
        RECT 9.900 38.120 10.300 38.250 ;
        RECT 13.000 38.120 13.260 39.730 ;
        RECT 15.550 38.660 15.850 39.710 ;
        RECT 16.300 39.110 16.600 40.060 ;
        RECT 16.800 39.160 17.100 39.210 ;
        RECT 16.800 38.810 17.700 39.160 ;
        RECT 19.410 39.030 19.630 39.040 ;
        RECT 19.410 38.840 33.090 39.030 ;
        RECT 19.410 38.710 19.630 38.840 ;
        RECT 8.520 37.910 8.810 38.070 ;
        RECT 9.900 38.060 10.160 38.120 ;
        RECT 8.020 37.720 8.810 37.910 ;
        RECT 8.020 37.520 8.270 37.720 ;
        RECT 8.520 37.610 8.810 37.720 ;
        RECT 9.910 37.520 10.160 38.060 ;
        RECT 12.990 38.060 13.260 38.120 ;
        RECT 14.540 38.400 15.850 38.660 ;
        RECT 17.950 38.410 19.630 38.710 ;
        RECT 17.950 38.400 19.610 38.410 ;
        RECT 14.540 38.060 14.850 38.400 ;
        RECT 10.550 37.530 12.190 37.920 ;
        RECT 12.990 37.770 14.850 38.060 ;
        RECT 12.990 37.760 13.300 37.770 ;
        RECT 14.540 37.760 14.850 37.770 ;
        RECT 8.020 36.920 8.310 37.520 ;
        RECT 9.910 36.920 10.200 37.520 ;
        RECT 3.040 36.660 3.290 36.750 ;
        RECT 2.310 36.210 3.290 36.660 ;
        RECT 12.250 36.310 12.550 37.310 ;
        RECT 13.000 36.710 13.300 37.760 ;
        RECT 15.600 36.660 15.850 38.400 ;
        RECT 32.840 37.940 33.090 38.840 ;
        RECT 16.300 36.310 16.560 37.860 ;
        RECT 27.780 37.640 33.090 37.940 ;
        RECT 12.200 36.290 17.450 36.310 ;
        RECT 12.200 36.010 17.570 36.290 ;
        RECT 5.650 35.610 5.930 35.680 ;
        RECT 6.830 35.640 7.110 35.670 ;
        RECT 17.280 35.640 17.570 36.010 ;
        RECT 6.830 35.630 17.570 35.640 ;
        RECT 4.240 35.410 5.930 35.610 ;
        RECT 3.030 35.210 3.310 35.220 ;
        RECT 2.290 34.760 3.310 35.210 ;
        RECT 4.240 34.760 4.470 35.410 ;
        RECT 5.650 35.350 5.930 35.410 ;
        RECT 6.810 35.400 17.570 35.630 ;
        RECT 6.830 35.390 17.570 35.400 ;
        RECT 23.700 36.000 23.960 37.200 ;
        RECT 23.700 35.490 23.950 36.000 ;
        RECT 25.590 35.990 25.850 37.200 ;
        RECT 27.980 36.090 28.230 37.640 ;
        RECT 25.590 35.830 25.980 35.990 ;
        RECT 25.580 35.700 25.980 35.830 ;
        RECT 28.680 35.700 28.940 37.310 ;
        RECT 31.230 36.240 31.530 37.290 ;
        RECT 31.980 36.690 32.280 37.640 ;
        RECT 32.480 36.740 32.780 36.790 ;
        RECT 32.480 36.390 33.380 36.740 ;
        RECT 46.140 36.340 50.610 36.370 ;
        RECT 35.200 36.310 50.610 36.340 ;
        RECT 34.530 36.290 50.610 36.310 ;
        RECT 24.200 35.490 24.490 35.650 ;
        RECT 25.580 35.640 25.840 35.700 ;
        RECT 6.830 35.380 17.530 35.390 ;
        RECT 6.830 35.340 7.110 35.380 ;
        RECT 23.700 35.300 24.490 35.490 ;
        RECT 23.700 35.100 23.950 35.300 ;
        RECT 24.200 35.190 24.490 35.300 ;
        RECT 25.590 35.100 25.840 35.640 ;
        RECT 28.670 35.640 28.940 35.700 ;
        RECT 30.220 35.980 31.530 36.240 ;
        RECT 30.220 35.640 30.530 35.980 ;
        RECT 26.230 35.110 27.870 35.500 ;
        RECT 28.670 35.350 30.530 35.640 ;
        RECT 28.670 35.340 28.980 35.350 ;
        RECT 30.220 35.340 30.530 35.350 ;
        RECT 5.630 34.780 5.900 34.860 ;
        RECT 3.030 34.550 4.470 34.760 ;
        RECT 5.020 34.560 5.900 34.780 ;
        RECT 3.030 33.500 3.310 34.550 ;
        RECT 5.020 33.750 5.240 34.560 ;
        RECT 5.630 34.530 5.900 34.560 ;
        RECT 6.760 34.820 7.050 34.870 ;
        RECT 6.760 34.640 17.510 34.820 ;
        RECT 6.760 34.540 7.050 34.640 ;
        RECT 11.600 34.630 15.230 34.640 ;
        RECT 17.310 33.960 17.510 34.640 ;
        RECT 23.700 34.500 23.990 35.100 ;
        RECT 25.590 34.500 25.880 35.100 ;
        RECT 2.310 33.050 3.310 33.500 ;
        RECT 2.290 31.600 3.590 32.050 ;
        RECT 3.290 31.200 3.590 31.600 ;
        RECT 5.010 31.220 5.240 33.750 ;
        RECT 12.260 33.660 17.510 33.960 ;
        RECT 27.930 33.890 28.230 34.890 ;
        RECT 28.680 34.290 28.980 35.340 ;
        RECT 31.280 34.240 31.530 35.980 ;
        RECT 33.650 35.970 50.610 36.290 ;
        RECT 34.530 35.960 50.610 35.970 ;
        RECT 34.530 35.930 46.510 35.960 ;
        RECT 34.530 35.920 35.420 35.930 ;
        RECT 31.980 33.890 32.240 35.440 ;
        RECT 33.070 33.890 33.270 33.900 ;
        RECT 4.080 31.200 5.240 31.220 ;
        RECT 3.290 31.020 5.240 31.200 ;
        RECT 8.180 32.020 8.440 33.220 ;
        RECT 8.180 31.510 8.430 32.020 ;
        RECT 10.070 32.010 10.330 33.220 ;
        RECT 12.460 32.110 12.710 33.660 ;
        RECT 10.070 31.850 10.460 32.010 ;
        RECT 10.060 31.720 10.460 31.850 ;
        RECT 13.160 31.720 13.420 33.330 ;
        RECT 15.710 32.260 16.010 33.310 ;
        RECT 16.460 32.710 16.760 33.660 ;
        RECT 17.310 33.650 17.510 33.660 ;
        RECT 27.880 33.590 33.270 33.890 ;
        RECT 16.960 32.760 17.260 32.810 ;
        RECT 16.960 32.410 17.860 32.760 ;
        RECT 33.070 32.350 33.270 33.590 ;
        RECT 50.230 32.390 50.590 35.960 ;
        RECT 25.510 32.330 26.700 32.340 ;
        RECT 27.690 32.330 28.880 32.340 ;
        RECT 29.910 32.330 31.100 32.340 ;
        RECT 32.090 32.330 33.280 32.350 ;
        RECT 23.300 32.320 33.280 32.330 ;
        RECT 19.910 32.300 21.100 32.310 ;
        RECT 22.190 32.300 33.280 32.320 ;
        RECT 8.680 31.510 8.970 31.670 ;
        RECT 10.060 31.660 10.320 31.720 ;
        RECT 8.180 31.320 8.970 31.510 ;
        RECT 8.180 31.120 8.430 31.320 ;
        RECT 8.680 31.210 8.970 31.320 ;
        RECT 10.070 31.120 10.320 31.660 ;
        RECT 13.150 31.660 13.420 31.720 ;
        RECT 14.700 32.000 16.010 32.260 ;
        RECT 18.070 32.070 33.280 32.300 ;
        RECT 45.360 32.090 50.610 32.390 ;
        RECT 18.070 32.060 32.230 32.070 ;
        RECT 18.070 32.050 25.600 32.060 ;
        RECT 26.610 32.050 27.800 32.060 ;
        RECT 28.760 32.050 29.950 32.060 ;
        RECT 31.040 32.050 32.230 32.060 ;
        RECT 18.070 32.040 23.380 32.050 ;
        RECT 18.070 32.030 22.240 32.040 ;
        RECT 18.070 32.020 19.960 32.030 ;
        RECT 21.050 32.020 22.240 32.030 ;
        RECT 18.070 32.010 18.790 32.020 ;
        RECT 14.700 31.660 15.010 32.000 ;
        RECT 10.710 31.130 12.350 31.520 ;
        RECT 13.150 31.370 15.010 31.660 ;
        RECT 13.150 31.360 13.460 31.370 ;
        RECT 14.700 31.360 15.010 31.370 ;
        RECT 3.290 31.010 3.940 31.020 ;
        RECT 3.290 30.680 3.590 31.010 ;
        RECT 2.570 30.230 3.590 30.680 ;
        RECT 8.180 30.520 8.470 31.120 ;
        RECT 10.070 30.520 10.360 31.120 ;
        RECT 3.290 30.220 3.590 30.230 ;
        RECT 12.410 29.910 12.710 30.910 ;
        RECT 13.160 30.310 13.460 31.360 ;
        RECT 15.760 30.260 16.010 32.000 ;
        RECT 16.460 29.910 16.720 31.460 ;
        RECT 41.280 30.450 41.540 31.650 ;
        RECT 41.280 29.940 41.530 30.450 ;
        RECT 43.170 30.440 43.430 31.650 ;
        RECT 45.560 30.540 45.810 32.090 ;
        RECT 43.170 30.280 43.560 30.440 ;
        RECT 43.160 30.150 43.560 30.280 ;
        RECT 46.260 30.150 46.520 31.760 ;
        RECT 48.810 30.690 49.110 31.740 ;
        RECT 49.560 31.140 49.860 32.090 ;
        RECT 50.060 31.190 50.360 31.240 ;
        RECT 50.060 30.840 50.960 31.190 ;
        RECT 41.780 29.940 42.070 30.100 ;
        RECT 43.160 30.090 43.420 30.150 ;
        RECT 12.360 29.900 17.610 29.910 ;
        RECT 2.240 29.820 2.490 29.830 ;
        RECT 2.240 29.360 3.220 29.820 ;
        RECT 12.360 29.610 17.630 29.900 ;
        RECT 2.240 29.060 2.490 29.360 ;
        RECT 10.210 29.270 12.050 29.280 ;
        RECT 17.460 29.270 17.630 29.610 ;
        RECT 3.950 29.260 4.190 29.270 ;
        RECT 5.030 29.260 17.630 29.270 ;
        RECT 3.950 29.100 17.630 29.260 ;
        RECT 41.280 29.750 42.070 29.940 ;
        RECT 41.280 29.550 41.530 29.750 ;
        RECT 41.780 29.640 42.070 29.750 ;
        RECT 43.170 29.550 43.420 30.090 ;
        RECT 46.250 30.090 46.520 30.150 ;
        RECT 47.800 30.430 49.110 30.690 ;
        RECT 51.170 30.740 52.840 30.760 ;
        RECT 67.980 30.740 68.290 42.090 ;
        RECT 103.840 41.780 104.890 42.240 ;
        RECT 164.380 42.200 164.680 43.200 ;
        RECT 165.130 42.600 165.430 43.650 ;
        RECT 167.730 42.550 167.980 44.290 ;
        RECT 170.690 44.280 184.000 44.290 ;
        RECT 168.430 42.200 168.690 43.750 ;
        RECT 164.330 41.900 169.600 42.200 ;
        RECT 104.640 41.770 104.890 41.780 ;
        RECT 103.510 41.370 103.760 41.380 ;
        RECT 103.510 40.920 104.490 41.370 ;
        RECT 105.600 41.110 114.870 41.120 ;
        RECT 116.750 41.110 118.670 41.120 ;
        RECT 105.600 40.920 118.670 41.110 ;
        RECT 103.510 40.310 103.760 40.920 ;
        RECT 105.600 40.910 117.960 40.920 ;
        RECT 103.510 40.060 104.720 40.310 ;
        RECT 104.450 39.310 104.710 40.060 ;
        RECT 105.600 39.900 105.810 40.910 ;
        RECT 114.860 40.900 116.760 40.910 ;
        RECT 118.490 40.170 118.670 40.920 ;
        RECT 104.450 38.710 104.700 39.310 ;
        RECT 105.600 38.890 105.800 39.900 ;
        RECT 113.410 39.870 118.670 40.170 ;
        RECT 103.660 38.260 104.700 38.710 ;
        RECT 103.640 36.810 104.600 37.260 ;
        RECT 104.350 36.760 104.600 36.810 ;
        RECT 105.610 36.760 105.800 38.890 ;
        RECT 104.350 36.560 105.800 36.760 ;
        RECT 109.330 38.230 109.590 39.430 ;
        RECT 109.330 37.720 109.580 38.230 ;
        RECT 111.220 38.220 111.480 39.430 ;
        RECT 113.610 38.320 113.860 39.870 ;
        RECT 111.220 38.060 111.610 38.220 ;
        RECT 111.210 37.930 111.610 38.060 ;
        RECT 114.310 37.930 114.570 39.540 ;
        RECT 116.860 38.470 117.160 39.520 ;
        RECT 117.610 38.920 117.910 39.870 ;
        RECT 118.110 38.970 118.410 39.020 ;
        RECT 118.110 38.620 119.010 38.970 ;
        RECT 120.720 38.840 120.940 38.850 ;
        RECT 120.720 38.650 134.400 38.840 ;
        RECT 120.720 38.520 120.940 38.650 ;
        RECT 109.830 37.720 110.120 37.880 ;
        RECT 111.210 37.870 111.470 37.930 ;
        RECT 109.330 37.530 110.120 37.720 ;
        RECT 109.330 37.330 109.580 37.530 ;
        RECT 109.830 37.420 110.120 37.530 ;
        RECT 111.220 37.330 111.470 37.870 ;
        RECT 114.300 37.870 114.570 37.930 ;
        RECT 115.850 38.210 117.160 38.470 ;
        RECT 119.260 38.220 120.940 38.520 ;
        RECT 119.260 38.210 120.920 38.220 ;
        RECT 115.850 37.870 116.160 38.210 ;
        RECT 111.860 37.340 113.500 37.730 ;
        RECT 114.300 37.580 116.160 37.870 ;
        RECT 114.300 37.570 114.610 37.580 ;
        RECT 115.850 37.570 116.160 37.580 ;
        RECT 109.330 36.730 109.620 37.330 ;
        RECT 111.220 36.730 111.510 37.330 ;
        RECT 104.350 36.470 104.600 36.560 ;
        RECT 103.620 36.020 104.600 36.470 ;
        RECT 113.560 36.120 113.860 37.120 ;
        RECT 114.310 36.520 114.610 37.570 ;
        RECT 116.910 36.470 117.160 38.210 ;
        RECT 134.150 37.750 134.400 38.650 ;
        RECT 117.610 36.120 117.870 37.670 ;
        RECT 129.090 37.450 134.400 37.750 ;
        RECT 113.510 36.100 118.760 36.120 ;
        RECT 113.510 35.820 118.880 36.100 ;
        RECT 106.960 35.420 107.240 35.490 ;
        RECT 108.140 35.450 108.420 35.480 ;
        RECT 118.590 35.450 118.880 35.820 ;
        RECT 108.140 35.440 118.880 35.450 ;
        RECT 105.550 35.220 107.240 35.420 ;
        RECT 104.340 35.020 104.620 35.030 ;
        RECT 103.600 34.570 104.620 35.020 ;
        RECT 105.550 34.570 105.780 35.220 ;
        RECT 106.960 35.160 107.240 35.220 ;
        RECT 108.120 35.210 118.880 35.440 ;
        RECT 108.140 35.200 118.880 35.210 ;
        RECT 125.010 35.810 125.270 37.010 ;
        RECT 125.010 35.300 125.260 35.810 ;
        RECT 126.900 35.800 127.160 37.010 ;
        RECT 129.290 35.900 129.540 37.450 ;
        RECT 126.900 35.640 127.290 35.800 ;
        RECT 126.890 35.510 127.290 35.640 ;
        RECT 129.990 35.510 130.250 37.120 ;
        RECT 132.540 36.050 132.840 37.100 ;
        RECT 133.290 36.500 133.590 37.450 ;
        RECT 133.790 36.550 134.090 36.600 ;
        RECT 133.790 36.200 134.690 36.550 ;
        RECT 147.450 36.150 151.920 36.180 ;
        RECT 136.510 36.120 151.920 36.150 ;
        RECT 135.840 36.100 151.920 36.120 ;
        RECT 125.510 35.300 125.800 35.460 ;
        RECT 126.890 35.450 127.150 35.510 ;
        RECT 108.140 35.190 118.840 35.200 ;
        RECT 108.140 35.150 108.420 35.190 ;
        RECT 125.010 35.110 125.800 35.300 ;
        RECT 125.010 34.910 125.260 35.110 ;
        RECT 125.510 35.000 125.800 35.110 ;
        RECT 126.900 34.910 127.150 35.450 ;
        RECT 129.980 35.450 130.250 35.510 ;
        RECT 131.530 35.790 132.840 36.050 ;
        RECT 131.530 35.450 131.840 35.790 ;
        RECT 127.540 34.920 129.180 35.310 ;
        RECT 129.980 35.160 131.840 35.450 ;
        RECT 129.980 35.150 130.290 35.160 ;
        RECT 131.530 35.150 131.840 35.160 ;
        RECT 106.940 34.590 107.210 34.670 ;
        RECT 104.340 34.360 105.780 34.570 ;
        RECT 106.330 34.370 107.210 34.590 ;
        RECT 104.340 33.310 104.620 34.360 ;
        RECT 106.330 33.560 106.550 34.370 ;
        RECT 106.940 34.340 107.210 34.370 ;
        RECT 108.070 34.630 108.360 34.680 ;
        RECT 108.070 34.450 118.820 34.630 ;
        RECT 108.070 34.350 108.360 34.450 ;
        RECT 112.910 34.440 116.540 34.450 ;
        RECT 118.620 33.770 118.820 34.450 ;
        RECT 125.010 34.310 125.300 34.910 ;
        RECT 126.900 34.310 127.190 34.910 ;
        RECT 103.620 32.860 104.620 33.310 ;
        RECT 103.600 31.410 104.900 31.860 ;
        RECT 104.600 31.010 104.900 31.410 ;
        RECT 106.320 31.030 106.550 33.560 ;
        RECT 113.570 33.470 118.820 33.770 ;
        RECT 129.240 33.700 129.540 34.700 ;
        RECT 129.990 34.100 130.290 35.150 ;
        RECT 132.590 34.050 132.840 35.790 ;
        RECT 134.960 35.780 151.920 36.100 ;
        RECT 135.840 35.770 151.920 35.780 ;
        RECT 135.840 35.740 147.820 35.770 ;
        RECT 135.840 35.730 136.730 35.740 ;
        RECT 133.290 33.700 133.550 35.250 ;
        RECT 134.380 33.700 134.580 33.710 ;
        RECT 105.390 31.010 106.550 31.030 ;
        RECT 104.600 30.830 106.550 31.010 ;
        RECT 109.490 31.830 109.750 33.030 ;
        RECT 109.490 31.320 109.740 31.830 ;
        RECT 111.380 31.820 111.640 33.030 ;
        RECT 113.770 31.920 114.020 33.470 ;
        RECT 111.380 31.660 111.770 31.820 ;
        RECT 111.370 31.530 111.770 31.660 ;
        RECT 114.470 31.530 114.730 33.140 ;
        RECT 117.020 32.070 117.320 33.120 ;
        RECT 117.770 32.520 118.070 33.470 ;
        RECT 118.620 33.460 118.820 33.470 ;
        RECT 129.190 33.400 134.580 33.700 ;
        RECT 118.270 32.570 118.570 32.620 ;
        RECT 118.270 32.220 119.170 32.570 ;
        RECT 134.380 32.160 134.580 33.400 ;
        RECT 151.540 32.200 151.900 35.770 ;
        RECT 126.820 32.140 128.010 32.150 ;
        RECT 129.000 32.140 130.190 32.150 ;
        RECT 131.220 32.140 132.410 32.150 ;
        RECT 133.400 32.140 134.590 32.160 ;
        RECT 124.610 32.130 134.590 32.140 ;
        RECT 121.220 32.110 122.410 32.120 ;
        RECT 123.500 32.110 134.590 32.130 ;
        RECT 109.990 31.320 110.280 31.480 ;
        RECT 111.370 31.470 111.630 31.530 ;
        RECT 109.490 31.130 110.280 31.320 ;
        RECT 109.490 30.930 109.740 31.130 ;
        RECT 109.990 31.020 110.280 31.130 ;
        RECT 111.380 30.930 111.630 31.470 ;
        RECT 114.460 31.470 114.730 31.530 ;
        RECT 116.010 31.810 117.320 32.070 ;
        RECT 119.380 31.880 134.590 32.110 ;
        RECT 146.670 31.900 151.920 32.200 ;
        RECT 119.380 31.870 133.540 31.880 ;
        RECT 119.380 31.860 126.910 31.870 ;
        RECT 127.920 31.860 129.110 31.870 ;
        RECT 130.070 31.860 131.260 31.870 ;
        RECT 132.350 31.860 133.540 31.870 ;
        RECT 119.380 31.850 124.690 31.860 ;
        RECT 119.380 31.840 123.550 31.850 ;
        RECT 119.380 31.830 121.270 31.840 ;
        RECT 122.360 31.830 123.550 31.840 ;
        RECT 119.380 31.820 120.100 31.830 ;
        RECT 116.010 31.470 116.320 31.810 ;
        RECT 112.020 30.940 113.660 31.330 ;
        RECT 114.460 31.180 116.320 31.470 ;
        RECT 114.460 31.170 114.770 31.180 ;
        RECT 116.010 31.170 116.320 31.180 ;
        RECT 104.600 30.820 105.250 30.830 ;
        RECT 51.170 30.450 68.330 30.740 ;
        RECT 104.600 30.490 104.900 30.820 ;
        RECT 51.860 30.440 68.330 30.450 ;
        RECT 47.800 30.090 48.110 30.430 ;
        RECT 43.810 29.560 45.450 29.950 ;
        RECT 46.250 29.800 48.110 30.090 ;
        RECT 46.250 29.790 46.560 29.800 ;
        RECT 47.800 29.790 48.110 29.800 ;
        RECT 3.950 29.090 15.460 29.100 ;
        RECT 3.940 29.080 10.260 29.090 ;
        RECT 11.810 29.080 15.460 29.090 ;
        RECT 3.940 29.070 5.810 29.080 ;
        RECT 3.940 29.060 4.190 29.070 ;
        RECT 2.240 28.890 4.190 29.060 ;
        RECT 41.280 28.950 41.570 29.550 ;
        RECT 43.170 28.950 43.460 29.550 ;
        RECT 2.240 28.670 2.490 28.890 ;
        RECT 2.240 28.500 3.280 28.670 ;
        RECT 3.090 27.640 3.280 28.500 ;
        RECT 45.510 28.340 45.810 29.340 ;
        RECT 46.260 28.740 46.560 29.790 ;
        RECT 48.860 28.690 49.110 30.430 ;
        RECT 103.880 30.040 104.900 30.490 ;
        RECT 109.490 30.330 109.780 30.930 ;
        RECT 111.380 30.330 111.670 30.930 ;
        RECT 104.600 30.030 104.900 30.040 ;
        RECT 49.560 28.340 49.820 29.890 ;
        RECT 113.720 29.720 114.020 30.720 ;
        RECT 114.470 30.120 114.770 31.170 ;
        RECT 117.070 30.070 117.320 31.810 ;
        RECT 117.770 29.720 118.030 31.270 ;
        RECT 142.590 30.260 142.850 31.460 ;
        RECT 142.590 29.750 142.840 30.260 ;
        RECT 144.480 30.250 144.740 31.460 ;
        RECT 146.870 30.350 147.120 31.900 ;
        RECT 144.480 30.090 144.870 30.250 ;
        RECT 144.470 29.960 144.870 30.090 ;
        RECT 147.570 29.960 147.830 31.570 ;
        RECT 150.120 30.500 150.420 31.550 ;
        RECT 150.870 30.950 151.170 31.900 ;
        RECT 151.370 31.000 151.670 31.050 ;
        RECT 151.370 30.650 152.270 31.000 ;
        RECT 143.090 29.750 143.380 29.910 ;
        RECT 144.470 29.900 144.730 29.960 ;
        RECT 113.670 29.710 118.920 29.720 ;
        RECT 103.550 29.630 103.800 29.640 ;
        RECT 103.550 29.170 104.530 29.630 ;
        RECT 113.670 29.420 118.940 29.710 ;
        RECT 103.550 28.870 103.800 29.170 ;
        RECT 111.520 29.080 113.360 29.090 ;
        RECT 118.770 29.080 118.940 29.420 ;
        RECT 105.260 29.070 105.500 29.080 ;
        RECT 106.340 29.070 118.940 29.080 ;
        RECT 105.260 28.910 118.940 29.070 ;
        RECT 142.590 29.560 143.380 29.750 ;
        RECT 142.590 29.360 142.840 29.560 ;
        RECT 143.090 29.450 143.380 29.560 ;
        RECT 144.480 29.360 144.730 29.900 ;
        RECT 147.560 29.900 147.830 29.960 ;
        RECT 149.110 30.240 150.420 30.500 ;
        RECT 152.480 30.550 154.150 30.570 ;
        RECT 169.290 30.550 169.600 41.900 ;
        RECT 152.480 30.260 169.640 30.550 ;
        RECT 153.170 30.250 169.640 30.260 ;
        RECT 149.110 29.900 149.420 30.240 ;
        RECT 145.120 29.370 146.760 29.760 ;
        RECT 147.560 29.610 149.420 29.900 ;
        RECT 147.560 29.600 147.870 29.610 ;
        RECT 149.110 29.600 149.420 29.610 ;
        RECT 105.260 28.900 116.770 28.910 ;
        RECT 105.250 28.890 111.570 28.900 ;
        RECT 113.120 28.890 116.770 28.900 ;
        RECT 105.250 28.880 107.120 28.890 ;
        RECT 105.250 28.870 105.500 28.880 ;
        RECT 103.550 28.700 105.500 28.870 ;
        RECT 142.590 28.760 142.880 29.360 ;
        RECT 144.480 28.760 144.770 29.360 ;
        RECT 103.550 28.480 103.800 28.700 ;
        RECT 50.440 28.340 50.780 28.410 ;
        RECT 45.460 28.040 50.780 28.340 ;
        RECT 103.550 28.310 104.590 28.480 ;
        RECT 2.300 27.200 3.280 27.640 ;
        RECT 2.300 27.190 3.250 27.200 ;
        RECT 4.120 26.880 13.390 26.890 ;
        RECT 15.270 26.880 17.190 26.890 ;
        RECT 1.970 26.780 2.160 26.790 ;
        RECT 1.970 26.320 2.950 26.780 ;
        RECT 4.120 26.690 17.190 26.880 ;
        RECT 4.120 26.680 16.480 26.690 ;
        RECT 1.970 25.530 2.160 26.320 ;
        RECT 4.120 25.670 4.330 26.680 ;
        RECT 13.380 26.670 15.280 26.680 ;
        RECT 17.010 25.940 17.190 26.690 ;
        RECT 2.970 25.530 3.240 25.540 ;
        RECT 1.970 25.320 3.240 25.530 ;
        RECT 2.970 25.110 3.240 25.320 ;
        RECT 2.970 24.480 3.220 25.110 ;
        RECT 4.120 24.660 4.320 25.670 ;
        RECT 11.930 25.640 17.190 25.940 ;
        RECT 2.180 24.030 3.220 24.480 ;
        RECT 2.160 22.580 3.120 23.030 ;
        RECT 2.870 22.530 3.120 22.580 ;
        RECT 4.130 22.530 4.320 24.660 ;
        RECT 2.870 22.330 4.320 22.530 ;
        RECT 7.850 24.000 8.110 25.200 ;
        RECT 7.850 23.490 8.100 24.000 ;
        RECT 9.740 23.990 10.000 25.200 ;
        RECT 12.130 24.090 12.380 25.640 ;
        RECT 9.740 23.830 10.130 23.990 ;
        RECT 9.730 23.700 10.130 23.830 ;
        RECT 12.830 23.700 13.090 25.310 ;
        RECT 15.380 24.240 15.680 25.290 ;
        RECT 16.130 24.690 16.430 25.640 ;
        RECT 16.630 24.740 16.930 24.790 ;
        RECT 16.630 24.390 17.530 24.740 ;
        RECT 19.240 24.610 19.460 24.620 ;
        RECT 19.240 24.420 32.920 24.610 ;
        RECT 19.240 24.290 19.460 24.420 ;
        RECT 8.350 23.490 8.640 23.650 ;
        RECT 9.730 23.640 9.990 23.700 ;
        RECT 7.850 23.300 8.640 23.490 ;
        RECT 7.850 23.100 8.100 23.300 ;
        RECT 8.350 23.190 8.640 23.300 ;
        RECT 9.740 23.100 9.990 23.640 ;
        RECT 12.820 23.640 13.090 23.700 ;
        RECT 14.370 23.980 15.680 24.240 ;
        RECT 17.780 23.990 19.460 24.290 ;
        RECT 17.780 23.980 19.440 23.990 ;
        RECT 14.370 23.640 14.680 23.980 ;
        RECT 10.380 23.110 12.020 23.500 ;
        RECT 12.820 23.350 14.680 23.640 ;
        RECT 12.820 23.340 13.130 23.350 ;
        RECT 14.370 23.340 14.680 23.350 ;
        RECT 7.850 22.500 8.140 23.100 ;
        RECT 9.740 22.500 10.030 23.100 ;
        RECT 2.870 22.240 3.120 22.330 ;
        RECT 2.140 21.790 3.120 22.240 ;
        RECT 12.080 21.890 12.380 22.890 ;
        RECT 12.830 22.290 13.130 23.340 ;
        RECT 15.430 22.240 15.680 23.980 ;
        RECT 32.670 23.520 32.920 24.420 ;
        RECT 16.130 21.890 16.390 23.440 ;
        RECT 27.610 23.220 32.920 23.520 ;
        RECT 12.030 21.870 17.280 21.890 ;
        RECT 12.030 21.590 17.400 21.870 ;
        RECT 5.480 21.190 5.760 21.260 ;
        RECT 6.660 21.220 6.940 21.250 ;
        RECT 17.110 21.220 17.400 21.590 ;
        RECT 6.660 21.210 17.400 21.220 ;
        RECT 4.070 20.990 5.760 21.190 ;
        RECT 2.860 20.790 3.140 20.800 ;
        RECT 2.120 20.340 3.140 20.790 ;
        RECT 4.070 20.340 4.300 20.990 ;
        RECT 5.480 20.930 5.760 20.990 ;
        RECT 6.640 20.980 17.400 21.210 ;
        RECT 6.660 20.970 17.400 20.980 ;
        RECT 23.530 21.580 23.790 22.780 ;
        RECT 23.530 21.070 23.780 21.580 ;
        RECT 25.420 21.570 25.680 22.780 ;
        RECT 27.810 21.670 28.060 23.220 ;
        RECT 25.420 21.410 25.810 21.570 ;
        RECT 25.410 21.280 25.810 21.410 ;
        RECT 28.510 21.280 28.770 22.890 ;
        RECT 31.060 21.820 31.360 22.870 ;
        RECT 31.810 22.270 32.110 23.220 ;
        RECT 32.310 22.320 32.610 22.370 ;
        RECT 32.310 21.970 33.210 22.320 ;
        RECT 50.440 21.920 50.780 28.040 ;
        RECT 104.400 27.450 104.590 28.310 ;
        RECT 146.820 28.150 147.120 29.150 ;
        RECT 147.570 28.550 147.870 29.600 ;
        RECT 150.170 28.500 150.420 30.240 ;
        RECT 150.870 28.150 151.130 29.700 ;
        RECT 151.750 28.150 152.090 28.220 ;
        RECT 146.770 27.850 152.090 28.150 ;
        RECT 103.610 27.010 104.590 27.450 ;
        RECT 103.610 27.000 104.560 27.010 ;
        RECT 105.430 26.690 114.700 26.700 ;
        RECT 116.580 26.690 118.500 26.700 ;
        RECT 103.280 26.590 103.470 26.600 ;
        RECT 103.280 26.130 104.260 26.590 ;
        RECT 105.430 26.500 118.500 26.690 ;
        RECT 105.430 26.490 117.790 26.500 ;
        RECT 103.280 25.340 103.470 26.130 ;
        RECT 105.430 25.480 105.640 26.490 ;
        RECT 114.690 26.480 116.590 26.490 ;
        RECT 118.320 25.750 118.500 26.500 ;
        RECT 104.280 25.340 104.550 25.350 ;
        RECT 103.280 25.130 104.550 25.340 ;
        RECT 104.280 24.920 104.550 25.130 ;
        RECT 104.280 24.290 104.530 24.920 ;
        RECT 105.430 24.470 105.630 25.480 ;
        RECT 113.240 25.450 118.500 25.750 ;
        RECT 103.490 23.840 104.530 24.290 ;
        RECT 103.470 22.390 104.430 22.840 ;
        RECT 104.180 22.340 104.430 22.390 ;
        RECT 105.440 22.340 105.630 24.470 ;
        RECT 104.180 22.140 105.630 22.340 ;
        RECT 109.160 23.810 109.420 25.010 ;
        RECT 109.160 23.300 109.410 23.810 ;
        RECT 111.050 23.800 111.310 25.010 ;
        RECT 113.440 23.900 113.690 25.450 ;
        RECT 111.050 23.640 111.440 23.800 ;
        RECT 111.040 23.510 111.440 23.640 ;
        RECT 114.140 23.510 114.400 25.120 ;
        RECT 116.690 24.050 116.990 25.100 ;
        RECT 117.440 24.500 117.740 25.450 ;
        RECT 117.940 24.550 118.240 24.600 ;
        RECT 117.940 24.200 118.840 24.550 ;
        RECT 120.550 24.420 120.770 24.430 ;
        RECT 120.550 24.230 134.230 24.420 ;
        RECT 120.550 24.100 120.770 24.230 ;
        RECT 109.660 23.300 109.950 23.460 ;
        RECT 111.040 23.450 111.300 23.510 ;
        RECT 109.160 23.110 109.950 23.300 ;
        RECT 109.160 22.910 109.410 23.110 ;
        RECT 109.660 23.000 109.950 23.110 ;
        RECT 111.050 22.910 111.300 23.450 ;
        RECT 114.130 23.450 114.400 23.510 ;
        RECT 115.680 23.790 116.990 24.050 ;
        RECT 119.090 23.800 120.770 24.100 ;
        RECT 119.090 23.790 120.750 23.800 ;
        RECT 115.680 23.450 115.990 23.790 ;
        RECT 111.690 22.920 113.330 23.310 ;
        RECT 114.130 23.160 115.990 23.450 ;
        RECT 114.130 23.150 114.440 23.160 ;
        RECT 115.680 23.150 115.990 23.160 ;
        RECT 109.160 22.310 109.450 22.910 ;
        RECT 111.050 22.310 111.340 22.910 ;
        RECT 104.180 22.050 104.430 22.140 ;
        RECT 49.870 21.900 50.830 21.920 ;
        RECT 34.350 21.880 38.630 21.890 ;
        RECT 46.030 21.880 50.830 21.900 ;
        RECT 34.350 21.870 50.830 21.880 ;
        RECT 24.030 21.070 24.320 21.230 ;
        RECT 25.410 21.220 25.670 21.280 ;
        RECT 6.660 20.960 17.360 20.970 ;
        RECT 6.660 20.920 6.940 20.960 ;
        RECT 23.530 20.880 24.320 21.070 ;
        RECT 23.530 20.680 23.780 20.880 ;
        RECT 24.030 20.770 24.320 20.880 ;
        RECT 25.420 20.680 25.670 21.220 ;
        RECT 28.500 21.220 28.770 21.280 ;
        RECT 30.050 21.560 31.360 21.820 ;
        RECT 30.050 21.220 30.360 21.560 ;
        RECT 26.060 20.690 27.700 21.080 ;
        RECT 28.500 20.930 30.360 21.220 ;
        RECT 28.500 20.920 28.810 20.930 ;
        RECT 30.050 20.920 30.360 20.930 ;
        RECT 5.460 20.360 5.730 20.440 ;
        RECT 2.860 20.130 4.300 20.340 ;
        RECT 4.850 20.140 5.730 20.360 ;
        RECT 2.860 19.080 3.140 20.130 ;
        RECT 4.850 19.330 5.070 20.140 ;
        RECT 5.460 20.110 5.730 20.140 ;
        RECT 6.590 20.400 6.880 20.450 ;
        RECT 6.590 20.220 17.340 20.400 ;
        RECT 6.590 20.120 6.880 20.220 ;
        RECT 11.430 20.210 15.060 20.220 ;
        RECT 17.140 19.540 17.340 20.220 ;
        RECT 23.530 20.080 23.820 20.680 ;
        RECT 25.420 20.080 25.710 20.680 ;
        RECT 2.140 18.630 3.140 19.080 ;
        RECT 2.120 17.180 3.420 17.630 ;
        RECT 3.120 16.780 3.420 17.180 ;
        RECT 4.840 16.800 5.070 19.330 ;
        RECT 12.090 19.240 17.340 19.540 ;
        RECT 27.760 19.470 28.060 20.470 ;
        RECT 28.510 19.870 28.810 20.920 ;
        RECT 31.110 19.820 31.360 21.560 ;
        RECT 33.480 21.560 50.830 21.870 ;
        RECT 103.450 21.600 104.430 22.050 ;
        RECT 113.390 21.700 113.690 22.700 ;
        RECT 114.140 22.100 114.440 23.150 ;
        RECT 116.740 22.050 116.990 23.790 ;
        RECT 133.980 23.330 134.230 24.230 ;
        RECT 117.440 21.700 117.700 23.250 ;
        RECT 128.920 23.030 134.230 23.330 ;
        RECT 113.340 21.680 118.590 21.700 ;
        RECT 33.480 21.550 46.490 21.560 ;
        RECT 38.340 21.540 46.490 21.550 ;
        RECT 49.870 21.520 50.830 21.560 ;
        RECT 50.440 21.510 50.780 21.520 ;
        RECT 113.340 21.400 118.710 21.680 ;
        RECT 31.810 19.470 32.070 21.020 ;
        RECT 106.790 21.000 107.070 21.070 ;
        RECT 107.970 21.030 108.250 21.060 ;
        RECT 118.420 21.030 118.710 21.400 ;
        RECT 107.970 21.020 118.710 21.030 ;
        RECT 105.380 20.800 107.070 21.000 ;
        RECT 104.170 20.600 104.450 20.610 ;
        RECT 103.430 20.150 104.450 20.600 ;
        RECT 105.380 20.150 105.610 20.800 ;
        RECT 106.790 20.740 107.070 20.800 ;
        RECT 107.950 20.790 118.710 21.020 ;
        RECT 107.970 20.780 118.710 20.790 ;
        RECT 124.840 21.390 125.100 22.590 ;
        RECT 124.840 20.880 125.090 21.390 ;
        RECT 126.730 21.380 126.990 22.590 ;
        RECT 129.120 21.480 129.370 23.030 ;
        RECT 126.730 21.220 127.120 21.380 ;
        RECT 126.720 21.090 127.120 21.220 ;
        RECT 129.820 21.090 130.080 22.700 ;
        RECT 132.370 21.630 132.670 22.680 ;
        RECT 133.120 22.080 133.420 23.030 ;
        RECT 133.620 22.130 133.920 22.180 ;
        RECT 133.620 21.780 134.520 22.130 ;
        RECT 151.750 21.730 152.090 27.850 ;
        RECT 151.180 21.710 152.140 21.730 ;
        RECT 135.660 21.690 139.940 21.700 ;
        RECT 147.340 21.690 152.140 21.710 ;
        RECT 135.660 21.680 152.140 21.690 ;
        RECT 125.340 20.880 125.630 21.040 ;
        RECT 126.720 21.030 126.980 21.090 ;
        RECT 107.970 20.770 118.670 20.780 ;
        RECT 107.970 20.730 108.250 20.770 ;
        RECT 124.840 20.690 125.630 20.880 ;
        RECT 124.840 20.490 125.090 20.690 ;
        RECT 125.340 20.580 125.630 20.690 ;
        RECT 126.730 20.490 126.980 21.030 ;
        RECT 129.810 21.030 130.080 21.090 ;
        RECT 131.360 21.370 132.670 21.630 ;
        RECT 131.360 21.030 131.670 21.370 ;
        RECT 127.370 20.500 129.010 20.890 ;
        RECT 129.810 20.740 131.670 21.030 ;
        RECT 129.810 20.730 130.120 20.740 ;
        RECT 131.360 20.730 131.670 20.740 ;
        RECT 106.770 20.170 107.040 20.250 ;
        RECT 104.170 19.940 105.610 20.150 ;
        RECT 106.160 19.950 107.040 20.170 ;
        RECT 32.900 19.470 33.100 19.480 ;
        RECT 3.910 16.780 5.070 16.800 ;
        RECT 3.120 16.600 5.070 16.780 ;
        RECT 8.010 17.600 8.270 18.800 ;
        RECT 8.010 17.090 8.260 17.600 ;
        RECT 9.900 17.590 10.160 18.800 ;
        RECT 12.290 17.690 12.540 19.240 ;
        RECT 9.900 17.430 10.290 17.590 ;
        RECT 9.890 17.300 10.290 17.430 ;
        RECT 12.990 17.300 13.250 18.910 ;
        RECT 15.540 17.840 15.840 18.890 ;
        RECT 16.290 18.290 16.590 19.240 ;
        RECT 17.140 19.230 17.340 19.240 ;
        RECT 27.710 19.170 33.100 19.470 ;
        RECT 16.790 18.340 17.090 18.390 ;
        RECT 16.790 17.990 17.690 18.340 ;
        RECT 32.900 17.930 33.100 19.170 ;
        RECT 104.170 18.890 104.450 19.940 ;
        RECT 106.160 19.140 106.380 19.950 ;
        RECT 106.770 19.920 107.040 19.950 ;
        RECT 107.900 20.210 108.190 20.260 ;
        RECT 107.900 20.030 118.650 20.210 ;
        RECT 107.900 19.930 108.190 20.030 ;
        RECT 112.740 20.020 116.370 20.030 ;
        RECT 118.450 19.350 118.650 20.030 ;
        RECT 124.840 19.890 125.130 20.490 ;
        RECT 126.730 19.890 127.020 20.490 ;
        RECT 103.450 18.440 104.450 18.890 ;
        RECT 25.340 17.910 26.530 17.920 ;
        RECT 27.520 17.910 28.710 17.920 ;
        RECT 29.740 17.910 30.930 17.920 ;
        RECT 31.920 17.910 33.110 17.930 ;
        RECT 23.130 17.900 33.110 17.910 ;
        RECT 19.740 17.880 20.930 17.890 ;
        RECT 22.020 17.880 33.110 17.900 ;
        RECT 8.510 17.090 8.800 17.250 ;
        RECT 9.890 17.240 10.150 17.300 ;
        RECT 8.010 16.900 8.800 17.090 ;
        RECT 8.010 16.700 8.260 16.900 ;
        RECT 8.510 16.790 8.800 16.900 ;
        RECT 9.900 16.700 10.150 17.240 ;
        RECT 12.980 17.240 13.250 17.300 ;
        RECT 14.530 17.580 15.840 17.840 ;
        RECT 17.900 17.650 33.110 17.880 ;
        RECT 17.900 17.640 32.060 17.650 ;
        RECT 17.900 17.630 25.430 17.640 ;
        RECT 26.440 17.630 27.630 17.640 ;
        RECT 28.590 17.630 29.780 17.640 ;
        RECT 30.870 17.630 32.060 17.640 ;
        RECT 17.900 17.620 23.210 17.630 ;
        RECT 17.900 17.610 22.070 17.620 ;
        RECT 17.900 17.600 19.790 17.610 ;
        RECT 20.880 17.600 22.070 17.610 ;
        RECT 17.900 17.590 18.620 17.600 ;
        RECT 14.530 17.240 14.840 17.580 ;
        RECT 10.540 16.710 12.180 17.100 ;
        RECT 12.980 16.950 14.840 17.240 ;
        RECT 12.980 16.940 13.290 16.950 ;
        RECT 14.530 16.940 14.840 16.950 ;
        RECT 3.120 16.590 3.770 16.600 ;
        RECT 3.120 16.260 3.420 16.590 ;
        RECT 2.400 15.810 3.420 16.260 ;
        RECT 8.010 16.100 8.300 16.700 ;
        RECT 9.900 16.100 10.190 16.700 ;
        RECT 3.120 15.800 3.420 15.810 ;
        RECT 12.240 15.490 12.540 16.490 ;
        RECT 12.990 15.890 13.290 16.940 ;
        RECT 15.590 15.840 15.840 17.580 ;
        RECT 16.290 15.490 16.550 17.040 ;
        RECT 103.430 16.990 104.730 17.440 ;
        RECT 104.430 16.590 104.730 16.990 ;
        RECT 106.150 16.610 106.380 19.140 ;
        RECT 113.400 19.050 118.650 19.350 ;
        RECT 129.070 19.280 129.370 20.280 ;
        RECT 129.820 19.680 130.120 20.730 ;
        RECT 132.420 19.630 132.670 21.370 ;
        RECT 134.790 21.370 152.140 21.680 ;
        RECT 134.790 21.360 147.800 21.370 ;
        RECT 139.650 21.350 147.800 21.360 ;
        RECT 151.180 21.330 152.140 21.370 ;
        RECT 151.750 21.320 152.090 21.330 ;
        RECT 133.120 19.280 133.380 20.830 ;
        RECT 134.210 19.280 134.410 19.290 ;
        RECT 105.220 16.590 106.380 16.610 ;
        RECT 104.430 16.410 106.380 16.590 ;
        RECT 109.320 17.410 109.580 18.610 ;
        RECT 109.320 16.900 109.570 17.410 ;
        RECT 111.210 17.400 111.470 18.610 ;
        RECT 113.600 17.500 113.850 19.050 ;
        RECT 111.210 17.240 111.600 17.400 ;
        RECT 111.200 17.110 111.600 17.240 ;
        RECT 114.300 17.110 114.560 18.720 ;
        RECT 116.850 17.650 117.150 18.700 ;
        RECT 117.600 18.100 117.900 19.050 ;
        RECT 118.450 19.040 118.650 19.050 ;
        RECT 129.020 18.980 134.410 19.280 ;
        RECT 118.100 18.150 118.400 18.200 ;
        RECT 118.100 17.800 119.000 18.150 ;
        RECT 134.210 17.740 134.410 18.980 ;
        RECT 126.650 17.720 127.840 17.730 ;
        RECT 128.830 17.720 130.020 17.730 ;
        RECT 131.050 17.720 132.240 17.730 ;
        RECT 133.230 17.720 134.420 17.740 ;
        RECT 124.440 17.710 134.420 17.720 ;
        RECT 121.050 17.690 122.240 17.700 ;
        RECT 123.330 17.690 134.420 17.710 ;
        RECT 109.820 16.900 110.110 17.060 ;
        RECT 111.200 17.050 111.460 17.110 ;
        RECT 109.320 16.710 110.110 16.900 ;
        RECT 109.320 16.510 109.570 16.710 ;
        RECT 109.820 16.600 110.110 16.710 ;
        RECT 111.210 16.510 111.460 17.050 ;
        RECT 114.290 17.050 114.560 17.110 ;
        RECT 115.840 17.390 117.150 17.650 ;
        RECT 119.210 17.460 134.420 17.690 ;
        RECT 119.210 17.450 133.370 17.460 ;
        RECT 119.210 17.440 126.740 17.450 ;
        RECT 127.750 17.440 128.940 17.450 ;
        RECT 129.900 17.440 131.090 17.450 ;
        RECT 132.180 17.440 133.370 17.450 ;
        RECT 119.210 17.430 124.520 17.440 ;
        RECT 119.210 17.420 123.380 17.430 ;
        RECT 119.210 17.410 121.100 17.420 ;
        RECT 122.190 17.410 123.380 17.420 ;
        RECT 119.210 17.400 119.930 17.410 ;
        RECT 115.840 17.050 116.150 17.390 ;
        RECT 111.850 16.520 113.490 16.910 ;
        RECT 114.290 16.760 116.150 17.050 ;
        RECT 114.290 16.750 114.600 16.760 ;
        RECT 115.840 16.750 116.150 16.760 ;
        RECT 104.430 16.400 105.080 16.410 ;
        RECT 104.430 16.070 104.730 16.400 ;
        RECT 103.710 15.620 104.730 16.070 ;
        RECT 109.320 15.910 109.610 16.510 ;
        RECT 111.210 15.910 111.500 16.510 ;
        RECT 114.300 15.700 114.600 16.750 ;
        RECT 116.900 15.650 117.150 17.390 ;
        RECT 104.430 15.610 104.730 15.620 ;
        RECT 12.190 15.480 17.440 15.490 ;
        RECT 2.070 15.400 2.320 15.410 ;
        RECT 2.070 14.940 3.050 15.400 ;
        RECT 12.190 15.190 17.460 15.480 ;
        RECT 2.070 14.640 2.320 14.940 ;
        RECT 10.040 14.850 11.880 14.860 ;
        RECT 17.290 14.850 17.460 15.190 ;
        RECT 3.780 14.840 4.020 14.850 ;
        RECT 4.860 14.840 17.460 14.850 ;
        RECT 3.780 14.680 17.460 14.840 ;
        RECT 3.780 14.670 15.290 14.680 ;
        RECT 3.770 14.660 10.090 14.670 ;
        RECT 11.640 14.660 15.290 14.670 ;
        RECT 3.770 14.650 5.640 14.660 ;
        RECT 3.770 14.640 4.020 14.650 ;
        RECT 2.070 14.470 4.020 14.640 ;
        RECT 2.070 14.170 2.340 14.470 ;
        RECT 2.080 13.910 2.340 14.170 ;
        RECT 2.060 13.520 2.360 13.910 ;
        RECT 2.050 13.120 2.360 13.520 ;
        RECT 2.050 12.860 2.340 13.120 ;
        RECT 2.030 12.690 2.340 12.860 ;
        RECT 2.030 12.450 2.320 12.690 ;
        RECT 1.470 12.270 2.330 12.450 ;
        RECT 1.470 11.730 1.780 12.270 ;
        RECT 1.470 11.710 1.830 11.730 ;
        RECT 0.030 10.480 0.300 11.460 ;
        RECT 1.470 10.760 1.920 11.710 ;
        RECT 2.330 10.530 2.790 11.410 ;
        RECT 236.560 11.400 236.820 252.420 ;
        RECT 337.370 251.920 337.670 252.170 ;
        RECT 241.700 251.470 250.970 251.480 ;
        RECT 252.850 251.470 254.770 251.480 ;
        RECT 241.700 251.280 254.770 251.470 ;
        RECT 241.700 251.270 254.060 251.280 ;
        RECT 241.700 250.260 241.910 251.270 ;
        RECT 250.960 251.260 252.860 251.270 ;
        RECT 254.590 250.530 254.770 251.280 ;
        RECT 241.700 249.250 241.900 250.260 ;
        RECT 249.510 250.230 254.770 250.530 ;
        RECT 239.740 247.170 240.700 247.620 ;
        RECT 240.450 247.120 240.700 247.170 ;
        RECT 241.710 247.120 241.900 249.250 ;
        RECT 240.450 246.920 241.900 247.120 ;
        RECT 245.430 248.590 245.690 249.790 ;
        RECT 245.430 248.080 245.680 248.590 ;
        RECT 247.320 248.580 247.580 249.790 ;
        RECT 249.710 248.680 249.960 250.230 ;
        RECT 247.320 248.420 247.710 248.580 ;
        RECT 247.310 248.290 247.710 248.420 ;
        RECT 250.410 248.290 250.670 249.900 ;
        RECT 252.960 248.830 253.260 249.880 ;
        RECT 253.710 249.280 254.010 250.230 ;
        RECT 254.210 249.330 254.510 249.380 ;
        RECT 254.210 248.980 255.110 249.330 ;
        RECT 256.820 249.200 257.040 249.210 ;
        RECT 256.820 249.010 270.500 249.200 ;
        RECT 256.820 248.880 257.040 249.010 ;
        RECT 245.930 248.080 246.220 248.240 ;
        RECT 247.310 248.230 247.570 248.290 ;
        RECT 245.430 247.890 246.220 248.080 ;
        RECT 245.430 247.690 245.680 247.890 ;
        RECT 245.930 247.780 246.220 247.890 ;
        RECT 247.320 247.690 247.570 248.230 ;
        RECT 250.400 248.230 250.670 248.290 ;
        RECT 251.950 248.570 253.260 248.830 ;
        RECT 255.360 248.580 257.040 248.880 ;
        RECT 255.360 248.570 257.020 248.580 ;
        RECT 251.950 248.230 252.260 248.570 ;
        RECT 247.960 247.700 249.600 248.090 ;
        RECT 250.400 247.940 252.260 248.230 ;
        RECT 250.400 247.930 250.710 247.940 ;
        RECT 251.950 247.930 252.260 247.940 ;
        RECT 245.430 247.090 245.720 247.690 ;
        RECT 247.320 247.090 247.610 247.690 ;
        RECT 240.450 246.830 240.700 246.920 ;
        RECT 239.720 246.380 240.700 246.830 ;
        RECT 249.660 246.480 249.960 247.480 ;
        RECT 250.410 246.880 250.710 247.930 ;
        RECT 253.010 246.830 253.260 248.570 ;
        RECT 270.250 248.110 270.500 249.010 ;
        RECT 253.710 246.480 253.970 248.030 ;
        RECT 265.190 247.810 270.500 248.110 ;
        RECT 249.610 246.460 254.860 246.480 ;
        RECT 249.610 246.180 254.980 246.460 ;
        RECT 243.060 245.780 243.340 245.850 ;
        RECT 244.240 245.810 244.520 245.840 ;
        RECT 254.690 245.810 254.980 246.180 ;
        RECT 244.240 245.800 254.980 245.810 ;
        RECT 241.650 245.580 243.340 245.780 ;
        RECT 240.440 245.380 240.720 245.390 ;
        RECT 239.700 244.930 240.720 245.380 ;
        RECT 241.650 244.930 241.880 245.580 ;
        RECT 243.060 245.520 243.340 245.580 ;
        RECT 244.220 245.570 254.980 245.800 ;
        RECT 244.240 245.560 254.980 245.570 ;
        RECT 261.110 246.170 261.370 247.370 ;
        RECT 261.110 245.660 261.360 246.170 ;
        RECT 263.000 246.160 263.260 247.370 ;
        RECT 265.390 246.260 265.640 247.810 ;
        RECT 263.000 246.000 263.390 246.160 ;
        RECT 262.990 245.870 263.390 246.000 ;
        RECT 266.090 245.870 266.350 247.480 ;
        RECT 268.640 246.410 268.940 247.460 ;
        RECT 269.390 246.860 269.690 247.810 ;
        RECT 269.890 246.910 270.190 246.960 ;
        RECT 269.890 246.560 270.790 246.910 ;
        RECT 283.550 246.510 288.020 246.540 ;
        RECT 272.610 246.480 288.020 246.510 ;
        RECT 271.940 246.460 288.020 246.480 ;
        RECT 261.610 245.660 261.900 245.820 ;
        RECT 262.990 245.810 263.250 245.870 ;
        RECT 244.240 245.550 254.940 245.560 ;
        RECT 244.240 245.510 244.520 245.550 ;
        RECT 261.110 245.470 261.900 245.660 ;
        RECT 261.110 245.270 261.360 245.470 ;
        RECT 261.610 245.360 261.900 245.470 ;
        RECT 263.000 245.270 263.250 245.810 ;
        RECT 266.080 245.810 266.350 245.870 ;
        RECT 267.630 246.150 268.940 246.410 ;
        RECT 267.630 245.810 267.940 246.150 ;
        RECT 263.640 245.280 265.280 245.670 ;
        RECT 266.080 245.520 267.940 245.810 ;
        RECT 266.080 245.510 266.390 245.520 ;
        RECT 267.630 245.510 267.940 245.520 ;
        RECT 243.040 244.950 243.310 245.030 ;
        RECT 240.440 244.720 241.880 244.930 ;
        RECT 242.430 244.730 243.310 244.950 ;
        RECT 240.440 243.670 240.720 244.720 ;
        RECT 242.430 243.920 242.650 244.730 ;
        RECT 243.040 244.700 243.310 244.730 ;
        RECT 244.170 244.990 244.460 245.040 ;
        RECT 244.170 244.810 254.920 244.990 ;
        RECT 244.170 244.710 244.460 244.810 ;
        RECT 249.010 244.800 252.640 244.810 ;
        RECT 254.720 244.130 254.920 244.810 ;
        RECT 261.110 244.670 261.400 245.270 ;
        RECT 263.000 244.670 263.290 245.270 ;
        RECT 239.720 243.220 240.720 243.670 ;
        RECT 239.700 241.770 241.000 242.220 ;
        RECT 240.700 241.370 241.000 241.770 ;
        RECT 242.420 241.390 242.650 243.920 ;
        RECT 249.670 243.830 254.920 244.130 ;
        RECT 265.340 244.060 265.640 245.060 ;
        RECT 266.090 244.460 266.390 245.510 ;
        RECT 268.690 244.410 268.940 246.150 ;
        RECT 271.060 246.140 288.020 246.460 ;
        RECT 271.940 246.130 288.020 246.140 ;
        RECT 271.940 246.100 283.920 246.130 ;
        RECT 271.940 246.090 272.830 246.100 ;
        RECT 269.390 244.060 269.650 245.610 ;
        RECT 270.480 244.060 270.680 244.070 ;
        RECT 241.490 241.370 242.650 241.390 ;
        RECT 240.700 241.190 242.650 241.370 ;
        RECT 245.590 242.190 245.850 243.390 ;
        RECT 245.590 241.680 245.840 242.190 ;
        RECT 247.480 242.180 247.740 243.390 ;
        RECT 249.870 242.280 250.120 243.830 ;
        RECT 247.480 242.020 247.870 242.180 ;
        RECT 247.470 241.890 247.870 242.020 ;
        RECT 250.570 241.890 250.830 243.500 ;
        RECT 253.120 242.430 253.420 243.480 ;
        RECT 253.870 242.880 254.170 243.830 ;
        RECT 254.720 243.820 254.920 243.830 ;
        RECT 265.290 243.760 270.680 244.060 ;
        RECT 254.370 242.930 254.670 242.980 ;
        RECT 254.370 242.580 255.270 242.930 ;
        RECT 270.480 242.520 270.680 243.760 ;
        RECT 287.640 242.560 288.000 246.130 ;
        RECT 262.920 242.500 264.110 242.510 ;
        RECT 265.100 242.500 266.290 242.510 ;
        RECT 267.320 242.500 268.510 242.510 ;
        RECT 269.500 242.500 270.690 242.520 ;
        RECT 260.710 242.490 270.690 242.500 ;
        RECT 257.320 242.470 258.510 242.480 ;
        RECT 259.600 242.470 270.690 242.490 ;
        RECT 246.090 241.680 246.380 241.840 ;
        RECT 247.470 241.830 247.730 241.890 ;
        RECT 245.590 241.490 246.380 241.680 ;
        RECT 245.590 241.290 245.840 241.490 ;
        RECT 246.090 241.380 246.380 241.490 ;
        RECT 247.480 241.290 247.730 241.830 ;
        RECT 250.560 241.830 250.830 241.890 ;
        RECT 252.110 242.170 253.420 242.430 ;
        RECT 255.480 242.240 270.690 242.470 ;
        RECT 282.770 242.260 288.020 242.560 ;
        RECT 255.480 242.230 269.640 242.240 ;
        RECT 255.480 242.220 263.010 242.230 ;
        RECT 264.020 242.220 265.210 242.230 ;
        RECT 266.170 242.220 267.360 242.230 ;
        RECT 268.450 242.220 269.640 242.230 ;
        RECT 255.480 242.210 260.790 242.220 ;
        RECT 255.480 242.200 259.650 242.210 ;
        RECT 255.480 242.190 257.370 242.200 ;
        RECT 258.460 242.190 259.650 242.200 ;
        RECT 255.480 242.180 256.200 242.190 ;
        RECT 252.110 241.830 252.420 242.170 ;
        RECT 248.120 241.300 249.760 241.690 ;
        RECT 250.560 241.540 252.420 241.830 ;
        RECT 250.560 241.530 250.870 241.540 ;
        RECT 252.110 241.530 252.420 241.540 ;
        RECT 240.700 241.180 241.350 241.190 ;
        RECT 240.700 240.850 241.000 241.180 ;
        RECT 239.980 240.400 241.000 240.850 ;
        RECT 245.590 240.690 245.880 241.290 ;
        RECT 247.480 240.690 247.770 241.290 ;
        RECT 240.700 240.390 241.000 240.400 ;
        RECT 249.820 240.080 250.120 241.080 ;
        RECT 250.570 240.480 250.870 241.530 ;
        RECT 253.170 240.430 253.420 242.170 ;
        RECT 253.870 240.080 254.130 241.630 ;
        RECT 278.690 240.620 278.950 241.820 ;
        RECT 278.690 240.110 278.940 240.620 ;
        RECT 280.580 240.610 280.840 241.820 ;
        RECT 282.970 240.710 283.220 242.260 ;
        RECT 280.580 240.450 280.970 240.610 ;
        RECT 280.570 240.320 280.970 240.450 ;
        RECT 283.670 240.320 283.930 241.930 ;
        RECT 286.220 240.860 286.520 241.910 ;
        RECT 286.970 241.310 287.270 242.260 ;
        RECT 287.470 241.360 287.770 241.410 ;
        RECT 287.470 241.010 288.370 241.360 ;
        RECT 279.190 240.110 279.480 240.270 ;
        RECT 280.570 240.260 280.830 240.320 ;
        RECT 249.770 240.070 255.020 240.080 ;
        RECT 239.650 239.990 239.900 240.000 ;
        RECT 239.650 239.530 240.630 239.990 ;
        RECT 249.770 239.780 255.040 240.070 ;
        RECT 239.650 239.230 239.900 239.530 ;
        RECT 247.620 239.440 249.460 239.450 ;
        RECT 254.870 239.440 255.040 239.780 ;
        RECT 241.360 239.430 241.600 239.440 ;
        RECT 242.440 239.430 255.040 239.440 ;
        RECT 241.360 239.270 255.040 239.430 ;
        RECT 278.690 239.920 279.480 240.110 ;
        RECT 278.690 239.720 278.940 239.920 ;
        RECT 279.190 239.810 279.480 239.920 ;
        RECT 280.580 239.720 280.830 240.260 ;
        RECT 283.660 240.260 283.930 240.320 ;
        RECT 285.210 240.600 286.520 240.860 ;
        RECT 288.580 240.900 290.250 240.930 ;
        RECT 305.330 240.900 305.580 240.910 ;
        RECT 288.580 240.630 305.580 240.900 ;
        RECT 288.580 240.620 302.080 240.630 ;
        RECT 289.860 240.600 302.080 240.620 ;
        RECT 285.210 240.260 285.520 240.600 ;
        RECT 281.220 239.730 282.860 240.120 ;
        RECT 283.660 239.970 285.520 240.260 ;
        RECT 283.660 239.960 283.970 239.970 ;
        RECT 285.210 239.960 285.520 239.970 ;
        RECT 241.360 239.260 252.870 239.270 ;
        RECT 241.350 239.250 247.670 239.260 ;
        RECT 249.220 239.250 252.870 239.260 ;
        RECT 241.350 239.240 243.220 239.250 ;
        RECT 241.350 239.230 241.600 239.240 ;
        RECT 239.650 239.060 241.600 239.230 ;
        RECT 278.690 239.120 278.980 239.720 ;
        RECT 280.580 239.120 280.870 239.720 ;
        RECT 239.650 238.840 239.900 239.060 ;
        RECT 239.650 238.670 240.690 238.840 ;
        RECT 240.500 237.810 240.690 238.670 ;
        RECT 282.920 238.510 283.220 239.510 ;
        RECT 283.670 238.910 283.970 239.960 ;
        RECT 286.270 238.860 286.520 240.600 ;
        RECT 286.970 238.510 287.230 240.060 ;
        RECT 287.850 238.510 288.190 238.580 ;
        RECT 282.870 238.210 288.190 238.510 ;
        RECT 239.710 237.370 240.690 237.810 ;
        RECT 239.710 237.360 240.660 237.370 ;
        RECT 241.530 237.050 250.800 237.060 ;
        RECT 252.680 237.050 254.600 237.060 ;
        RECT 239.380 236.950 239.570 236.960 ;
        RECT 239.380 236.490 240.360 236.950 ;
        RECT 241.530 236.860 254.600 237.050 ;
        RECT 241.530 236.850 253.890 236.860 ;
        RECT 239.380 235.700 239.570 236.490 ;
        RECT 241.530 235.840 241.740 236.850 ;
        RECT 250.790 236.840 252.690 236.850 ;
        RECT 254.420 236.110 254.600 236.860 ;
        RECT 240.380 235.700 240.650 235.710 ;
        RECT 239.380 235.490 240.650 235.700 ;
        RECT 240.380 235.280 240.650 235.490 ;
        RECT 240.380 234.650 240.630 235.280 ;
        RECT 241.530 234.830 241.730 235.840 ;
        RECT 249.340 235.810 254.600 236.110 ;
        RECT 239.590 234.200 240.630 234.650 ;
        RECT 239.570 232.750 240.530 233.200 ;
        RECT 240.280 232.700 240.530 232.750 ;
        RECT 241.540 232.700 241.730 234.830 ;
        RECT 240.280 232.500 241.730 232.700 ;
        RECT 245.260 234.170 245.520 235.370 ;
        RECT 245.260 233.660 245.510 234.170 ;
        RECT 247.150 234.160 247.410 235.370 ;
        RECT 249.540 234.260 249.790 235.810 ;
        RECT 247.150 234.000 247.540 234.160 ;
        RECT 247.140 233.870 247.540 234.000 ;
        RECT 250.240 233.870 250.500 235.480 ;
        RECT 252.790 234.410 253.090 235.460 ;
        RECT 253.540 234.860 253.840 235.810 ;
        RECT 254.040 234.910 254.340 234.960 ;
        RECT 254.040 234.560 254.940 234.910 ;
        RECT 256.650 234.780 256.870 234.790 ;
        RECT 256.650 234.590 270.330 234.780 ;
        RECT 256.650 234.460 256.870 234.590 ;
        RECT 245.760 233.660 246.050 233.820 ;
        RECT 247.140 233.810 247.400 233.870 ;
        RECT 245.260 233.470 246.050 233.660 ;
        RECT 245.260 233.270 245.510 233.470 ;
        RECT 245.760 233.360 246.050 233.470 ;
        RECT 247.150 233.270 247.400 233.810 ;
        RECT 250.230 233.810 250.500 233.870 ;
        RECT 251.780 234.150 253.090 234.410 ;
        RECT 255.190 234.160 256.870 234.460 ;
        RECT 255.190 234.150 256.850 234.160 ;
        RECT 251.780 233.810 252.090 234.150 ;
        RECT 247.790 233.280 249.430 233.670 ;
        RECT 250.230 233.520 252.090 233.810 ;
        RECT 250.230 233.510 250.540 233.520 ;
        RECT 251.780 233.510 252.090 233.520 ;
        RECT 245.260 232.670 245.550 233.270 ;
        RECT 247.150 232.670 247.440 233.270 ;
        RECT 240.280 232.410 240.530 232.500 ;
        RECT 239.550 231.960 240.530 232.410 ;
        RECT 249.490 232.060 249.790 233.060 ;
        RECT 250.240 232.460 250.540 233.510 ;
        RECT 252.840 232.410 253.090 234.150 ;
        RECT 270.080 233.690 270.330 234.590 ;
        RECT 253.540 232.060 253.800 233.610 ;
        RECT 265.020 233.390 270.330 233.690 ;
        RECT 249.440 232.040 254.690 232.060 ;
        RECT 249.440 231.760 254.810 232.040 ;
        RECT 242.890 231.360 243.170 231.430 ;
        RECT 244.070 231.390 244.350 231.420 ;
        RECT 254.520 231.390 254.810 231.760 ;
        RECT 244.070 231.380 254.810 231.390 ;
        RECT 241.480 231.160 243.170 231.360 ;
        RECT 240.270 230.960 240.550 230.970 ;
        RECT 239.530 230.510 240.550 230.960 ;
        RECT 241.480 230.510 241.710 231.160 ;
        RECT 242.890 231.100 243.170 231.160 ;
        RECT 244.050 231.150 254.810 231.380 ;
        RECT 244.070 231.140 254.810 231.150 ;
        RECT 260.940 231.750 261.200 232.950 ;
        RECT 260.940 231.240 261.190 231.750 ;
        RECT 262.830 231.740 263.090 232.950 ;
        RECT 265.220 231.840 265.470 233.390 ;
        RECT 262.830 231.580 263.220 231.740 ;
        RECT 262.820 231.450 263.220 231.580 ;
        RECT 265.920 231.450 266.180 233.060 ;
        RECT 268.470 231.990 268.770 233.040 ;
        RECT 269.220 232.440 269.520 233.390 ;
        RECT 269.720 232.490 270.020 232.540 ;
        RECT 269.720 232.140 270.620 232.490 ;
        RECT 287.850 232.090 288.190 238.210 ;
        RECT 287.280 232.070 288.240 232.090 ;
        RECT 271.760 232.050 276.040 232.060 ;
        RECT 283.440 232.050 288.240 232.070 ;
        RECT 271.760 232.040 288.240 232.050 ;
        RECT 261.440 231.240 261.730 231.400 ;
        RECT 262.820 231.390 263.080 231.450 ;
        RECT 244.070 231.130 254.770 231.140 ;
        RECT 244.070 231.090 244.350 231.130 ;
        RECT 260.940 231.050 261.730 231.240 ;
        RECT 260.940 230.850 261.190 231.050 ;
        RECT 261.440 230.940 261.730 231.050 ;
        RECT 262.830 230.850 263.080 231.390 ;
        RECT 265.910 231.390 266.180 231.450 ;
        RECT 267.460 231.730 268.770 231.990 ;
        RECT 267.460 231.390 267.770 231.730 ;
        RECT 263.470 230.860 265.110 231.250 ;
        RECT 265.910 231.100 267.770 231.390 ;
        RECT 265.910 231.090 266.220 231.100 ;
        RECT 267.460 231.090 267.770 231.100 ;
        RECT 242.870 230.530 243.140 230.610 ;
        RECT 240.270 230.300 241.710 230.510 ;
        RECT 242.260 230.310 243.140 230.530 ;
        RECT 240.270 229.250 240.550 230.300 ;
        RECT 242.260 229.500 242.480 230.310 ;
        RECT 242.870 230.280 243.140 230.310 ;
        RECT 244.000 230.570 244.290 230.620 ;
        RECT 244.000 230.390 254.750 230.570 ;
        RECT 244.000 230.290 244.290 230.390 ;
        RECT 248.840 230.380 252.470 230.390 ;
        RECT 254.550 229.710 254.750 230.390 ;
        RECT 260.940 230.250 261.230 230.850 ;
        RECT 262.830 230.250 263.120 230.850 ;
        RECT 239.550 228.800 240.550 229.250 ;
        RECT 239.530 227.350 240.830 227.800 ;
        RECT 240.530 226.950 240.830 227.350 ;
        RECT 242.250 226.970 242.480 229.500 ;
        RECT 249.500 229.410 254.750 229.710 ;
        RECT 265.170 229.640 265.470 230.640 ;
        RECT 265.920 230.040 266.220 231.090 ;
        RECT 268.520 229.990 268.770 231.730 ;
        RECT 270.890 231.730 288.240 232.040 ;
        RECT 270.890 231.720 283.900 231.730 ;
        RECT 275.750 231.710 283.900 231.720 ;
        RECT 287.280 231.690 288.240 231.730 ;
        RECT 287.850 231.680 288.190 231.690 ;
        RECT 269.220 229.640 269.480 231.190 ;
        RECT 270.310 229.640 270.510 229.650 ;
        RECT 241.320 226.950 242.480 226.970 ;
        RECT 240.530 226.770 242.480 226.950 ;
        RECT 245.420 227.770 245.680 228.970 ;
        RECT 245.420 227.260 245.670 227.770 ;
        RECT 247.310 227.760 247.570 228.970 ;
        RECT 249.700 227.860 249.950 229.410 ;
        RECT 247.310 227.600 247.700 227.760 ;
        RECT 247.300 227.470 247.700 227.600 ;
        RECT 250.400 227.470 250.660 229.080 ;
        RECT 252.950 228.010 253.250 229.060 ;
        RECT 253.700 228.460 254.000 229.410 ;
        RECT 254.550 229.400 254.750 229.410 ;
        RECT 265.120 229.340 270.510 229.640 ;
        RECT 254.200 228.510 254.500 228.560 ;
        RECT 254.200 228.160 255.100 228.510 ;
        RECT 270.310 228.100 270.510 229.340 ;
        RECT 262.750 228.080 263.940 228.090 ;
        RECT 264.930 228.080 266.120 228.090 ;
        RECT 267.150 228.080 268.340 228.090 ;
        RECT 269.330 228.080 270.520 228.100 ;
        RECT 260.540 228.070 270.520 228.080 ;
        RECT 257.150 228.050 258.340 228.060 ;
        RECT 259.430 228.050 270.520 228.070 ;
        RECT 245.920 227.260 246.210 227.420 ;
        RECT 247.300 227.410 247.560 227.470 ;
        RECT 245.420 227.070 246.210 227.260 ;
        RECT 245.420 226.870 245.670 227.070 ;
        RECT 245.920 226.960 246.210 227.070 ;
        RECT 247.310 226.870 247.560 227.410 ;
        RECT 250.390 227.410 250.660 227.470 ;
        RECT 251.940 227.750 253.250 228.010 ;
        RECT 255.310 227.820 270.520 228.050 ;
        RECT 255.310 227.810 269.470 227.820 ;
        RECT 255.310 227.800 262.840 227.810 ;
        RECT 263.850 227.800 265.040 227.810 ;
        RECT 266.000 227.800 267.190 227.810 ;
        RECT 268.280 227.800 269.470 227.810 ;
        RECT 255.310 227.790 260.620 227.800 ;
        RECT 255.310 227.780 259.480 227.790 ;
        RECT 255.310 227.770 257.200 227.780 ;
        RECT 258.290 227.770 259.480 227.780 ;
        RECT 255.310 227.760 256.030 227.770 ;
        RECT 251.940 227.410 252.250 227.750 ;
        RECT 247.950 226.880 249.590 227.270 ;
        RECT 250.390 227.120 252.250 227.410 ;
        RECT 250.390 227.110 250.700 227.120 ;
        RECT 251.940 227.110 252.250 227.120 ;
        RECT 240.530 226.760 241.180 226.770 ;
        RECT 240.530 226.430 240.830 226.760 ;
        RECT 239.810 225.980 240.830 226.430 ;
        RECT 245.420 226.270 245.710 226.870 ;
        RECT 247.310 226.270 247.600 226.870 ;
        RECT 240.530 225.970 240.830 225.980 ;
        RECT 249.650 225.660 249.950 226.660 ;
        RECT 250.400 226.060 250.700 227.110 ;
        RECT 253.000 226.010 253.250 227.750 ;
        RECT 305.330 227.490 305.590 240.630 ;
        RECT 305.320 227.370 305.590 227.490 ;
        RECT 253.700 225.660 253.960 227.210 ;
        RECT 305.320 226.540 305.580 227.370 ;
        RECT 300.300 226.240 305.580 226.540 ;
        RECT 249.600 225.650 254.850 225.660 ;
        RECT 239.480 225.570 239.730 225.580 ;
        RECT 239.480 225.110 240.460 225.570 ;
        RECT 249.600 225.360 254.870 225.650 ;
        RECT 239.480 224.810 239.730 225.110 ;
        RECT 247.450 225.020 249.290 225.030 ;
        RECT 254.700 225.020 254.870 225.360 ;
        RECT 241.190 225.010 241.430 225.020 ;
        RECT 242.270 225.010 254.870 225.020 ;
        RECT 241.190 224.850 254.870 225.010 ;
        RECT 241.190 224.840 252.700 224.850 ;
        RECT 241.180 224.830 247.500 224.840 ;
        RECT 249.050 224.830 252.700 224.840 ;
        RECT 241.180 224.820 243.050 224.830 ;
        RECT 241.180 224.810 241.430 224.820 ;
        RECT 239.480 224.640 241.430 224.810 ;
        RECT 239.480 224.340 239.750 224.640 ;
        RECT 239.490 224.080 239.750 224.340 ;
        RECT 296.220 224.600 296.480 225.800 ;
        RECT 296.220 224.090 296.470 224.600 ;
        RECT 298.110 224.590 298.370 225.800 ;
        RECT 300.500 224.690 300.750 226.240 ;
        RECT 298.110 224.430 298.500 224.590 ;
        RECT 298.100 224.300 298.500 224.430 ;
        RECT 301.200 224.300 301.460 225.910 ;
        RECT 303.750 224.840 304.050 225.890 ;
        RECT 304.500 225.290 304.800 226.240 ;
        RECT 305.000 225.340 305.300 225.390 ;
        RECT 305.000 224.990 305.900 225.340 ;
        RECT 296.720 224.090 297.010 224.250 ;
        RECT 298.100 224.240 298.360 224.300 ;
        RECT 239.470 223.690 239.770 224.080 ;
        RECT 296.220 223.900 297.010 224.090 ;
        RECT 296.220 223.700 296.470 223.900 ;
        RECT 296.720 223.790 297.010 223.900 ;
        RECT 298.110 223.700 298.360 224.240 ;
        RECT 301.190 224.240 301.460 224.300 ;
        RECT 302.740 224.580 304.050 224.840 ;
        RECT 306.170 224.780 306.950 224.880 ;
        RECT 306.170 224.610 319.750 224.780 ;
        RECT 306.170 224.600 319.740 224.610 ;
        RECT 306.170 224.580 306.950 224.600 ;
        RECT 302.740 224.240 303.050 224.580 ;
        RECT 298.750 223.710 300.390 224.100 ;
        RECT 301.190 223.950 303.050 224.240 ;
        RECT 301.190 223.940 301.500 223.950 ;
        RECT 302.740 223.940 303.050 223.950 ;
        RECT 239.470 223.460 240.960 223.690 ;
        RECT 240.710 222.530 240.960 223.460 ;
        RECT 296.220 223.100 296.510 223.700 ;
        RECT 298.110 223.100 298.400 223.700 ;
        RECT 239.910 222.070 240.960 222.530 ;
        RECT 300.450 222.490 300.750 223.490 ;
        RECT 301.200 222.890 301.500 223.940 ;
        RECT 303.800 222.840 304.050 224.580 ;
        RECT 304.500 222.490 304.760 224.040 ;
        RECT 300.400 222.190 305.670 222.490 ;
        RECT 240.710 222.060 240.960 222.070 ;
        RECT 239.580 221.660 239.830 221.670 ;
        RECT 239.580 221.210 240.560 221.660 ;
        RECT 241.670 221.400 250.940 221.410 ;
        RECT 252.820 221.400 254.740 221.410 ;
        RECT 241.670 221.210 254.740 221.400 ;
        RECT 239.580 220.600 239.830 221.210 ;
        RECT 241.670 221.200 254.030 221.210 ;
        RECT 239.580 220.350 240.790 220.600 ;
        RECT 240.520 219.600 240.780 220.350 ;
        RECT 241.670 220.190 241.880 221.200 ;
        RECT 250.930 221.190 252.830 221.200 ;
        RECT 254.560 220.460 254.740 221.210 ;
        RECT 240.520 219.000 240.770 219.600 ;
        RECT 241.670 219.180 241.870 220.190 ;
        RECT 249.480 220.160 254.740 220.460 ;
        RECT 239.730 218.550 240.770 219.000 ;
        RECT 239.710 217.100 240.670 217.550 ;
        RECT 240.420 217.050 240.670 217.100 ;
        RECT 241.680 217.050 241.870 219.180 ;
        RECT 240.420 216.850 241.870 217.050 ;
        RECT 245.400 218.520 245.660 219.720 ;
        RECT 245.400 218.010 245.650 218.520 ;
        RECT 247.290 218.510 247.550 219.720 ;
        RECT 249.680 218.610 249.930 220.160 ;
        RECT 247.290 218.350 247.680 218.510 ;
        RECT 247.280 218.220 247.680 218.350 ;
        RECT 250.380 218.220 250.640 219.830 ;
        RECT 252.930 218.760 253.230 219.810 ;
        RECT 253.680 219.210 253.980 220.160 ;
        RECT 254.180 219.260 254.480 219.310 ;
        RECT 254.180 218.910 255.080 219.260 ;
        RECT 256.790 219.130 257.010 219.140 ;
        RECT 256.790 218.940 270.470 219.130 ;
        RECT 256.790 218.810 257.010 218.940 ;
        RECT 245.900 218.010 246.190 218.170 ;
        RECT 247.280 218.160 247.540 218.220 ;
        RECT 245.400 217.820 246.190 218.010 ;
        RECT 245.400 217.620 245.650 217.820 ;
        RECT 245.900 217.710 246.190 217.820 ;
        RECT 247.290 217.620 247.540 218.160 ;
        RECT 250.370 218.160 250.640 218.220 ;
        RECT 251.920 218.500 253.230 218.760 ;
        RECT 255.330 218.510 257.010 218.810 ;
        RECT 255.330 218.500 256.990 218.510 ;
        RECT 251.920 218.160 252.230 218.500 ;
        RECT 247.930 217.630 249.570 218.020 ;
        RECT 250.370 217.870 252.230 218.160 ;
        RECT 250.370 217.860 250.680 217.870 ;
        RECT 251.920 217.860 252.230 217.870 ;
        RECT 245.400 217.020 245.690 217.620 ;
        RECT 247.290 217.020 247.580 217.620 ;
        RECT 240.420 216.760 240.670 216.850 ;
        RECT 239.690 216.310 240.670 216.760 ;
        RECT 249.630 216.410 249.930 217.410 ;
        RECT 250.380 216.810 250.680 217.860 ;
        RECT 252.980 216.760 253.230 218.500 ;
        RECT 270.220 218.040 270.470 218.940 ;
        RECT 253.680 216.410 253.940 217.960 ;
        RECT 265.160 217.740 270.470 218.040 ;
        RECT 249.580 216.390 254.830 216.410 ;
        RECT 249.580 216.110 254.950 216.390 ;
        RECT 243.030 215.710 243.310 215.780 ;
        RECT 244.210 215.740 244.490 215.770 ;
        RECT 254.660 215.740 254.950 216.110 ;
        RECT 244.210 215.730 254.950 215.740 ;
        RECT 241.620 215.510 243.310 215.710 ;
        RECT 240.410 215.310 240.690 215.320 ;
        RECT 239.670 214.860 240.690 215.310 ;
        RECT 241.620 214.860 241.850 215.510 ;
        RECT 243.030 215.450 243.310 215.510 ;
        RECT 244.190 215.500 254.950 215.730 ;
        RECT 244.210 215.490 254.950 215.500 ;
        RECT 261.080 216.100 261.340 217.300 ;
        RECT 261.080 215.590 261.330 216.100 ;
        RECT 262.970 216.090 263.230 217.300 ;
        RECT 265.360 216.190 265.610 217.740 ;
        RECT 262.970 215.930 263.360 216.090 ;
        RECT 262.960 215.800 263.360 215.930 ;
        RECT 266.060 215.800 266.320 217.410 ;
        RECT 268.610 216.340 268.910 217.390 ;
        RECT 269.360 216.790 269.660 217.740 ;
        RECT 269.860 216.840 270.160 216.890 ;
        RECT 269.860 216.490 270.760 216.840 ;
        RECT 283.520 216.440 287.990 216.470 ;
        RECT 272.580 216.410 287.990 216.440 ;
        RECT 271.910 216.390 287.990 216.410 ;
        RECT 261.580 215.590 261.870 215.750 ;
        RECT 262.960 215.740 263.220 215.800 ;
        RECT 244.210 215.480 254.910 215.490 ;
        RECT 244.210 215.440 244.490 215.480 ;
        RECT 261.080 215.400 261.870 215.590 ;
        RECT 261.080 215.200 261.330 215.400 ;
        RECT 261.580 215.290 261.870 215.400 ;
        RECT 262.970 215.200 263.220 215.740 ;
        RECT 266.050 215.740 266.320 215.800 ;
        RECT 267.600 216.080 268.910 216.340 ;
        RECT 267.600 215.740 267.910 216.080 ;
        RECT 263.610 215.210 265.250 215.600 ;
        RECT 266.050 215.450 267.910 215.740 ;
        RECT 266.050 215.440 266.360 215.450 ;
        RECT 267.600 215.440 267.910 215.450 ;
        RECT 243.010 214.880 243.280 214.960 ;
        RECT 240.410 214.650 241.850 214.860 ;
        RECT 242.400 214.660 243.280 214.880 ;
        RECT 240.410 213.600 240.690 214.650 ;
        RECT 242.400 213.850 242.620 214.660 ;
        RECT 243.010 214.630 243.280 214.660 ;
        RECT 244.140 214.920 244.430 214.970 ;
        RECT 244.140 214.740 254.890 214.920 ;
        RECT 244.140 214.640 244.430 214.740 ;
        RECT 248.980 214.730 252.610 214.740 ;
        RECT 254.690 214.060 254.890 214.740 ;
        RECT 261.080 214.600 261.370 215.200 ;
        RECT 262.970 214.600 263.260 215.200 ;
        RECT 239.690 213.150 240.690 213.600 ;
        RECT 239.670 211.700 240.970 212.150 ;
        RECT 240.670 211.300 240.970 211.700 ;
        RECT 242.390 211.320 242.620 213.850 ;
        RECT 249.640 213.760 254.890 214.060 ;
        RECT 265.310 213.990 265.610 214.990 ;
        RECT 266.060 214.390 266.360 215.440 ;
        RECT 268.660 214.340 268.910 216.080 ;
        RECT 271.030 216.070 287.990 216.390 ;
        RECT 271.910 216.060 287.990 216.070 ;
        RECT 271.910 216.030 283.890 216.060 ;
        RECT 271.910 216.020 272.800 216.030 ;
        RECT 269.360 213.990 269.620 215.540 ;
        RECT 270.450 213.990 270.650 214.000 ;
        RECT 241.460 211.300 242.620 211.320 ;
        RECT 240.670 211.120 242.620 211.300 ;
        RECT 245.560 212.120 245.820 213.320 ;
        RECT 245.560 211.610 245.810 212.120 ;
        RECT 247.450 212.110 247.710 213.320 ;
        RECT 249.840 212.210 250.090 213.760 ;
        RECT 247.450 211.950 247.840 212.110 ;
        RECT 247.440 211.820 247.840 211.950 ;
        RECT 250.540 211.820 250.800 213.430 ;
        RECT 253.090 212.360 253.390 213.410 ;
        RECT 253.840 212.810 254.140 213.760 ;
        RECT 254.690 213.750 254.890 213.760 ;
        RECT 265.260 213.690 270.650 213.990 ;
        RECT 254.340 212.860 254.640 212.910 ;
        RECT 254.340 212.510 255.240 212.860 ;
        RECT 270.450 212.450 270.650 213.690 ;
        RECT 287.610 212.490 287.970 216.060 ;
        RECT 262.890 212.430 264.080 212.440 ;
        RECT 265.070 212.430 266.260 212.440 ;
        RECT 267.290 212.430 268.480 212.440 ;
        RECT 269.470 212.430 270.660 212.450 ;
        RECT 260.680 212.420 270.660 212.430 ;
        RECT 257.290 212.400 258.480 212.410 ;
        RECT 259.570 212.400 270.660 212.420 ;
        RECT 246.060 211.610 246.350 211.770 ;
        RECT 247.440 211.760 247.700 211.820 ;
        RECT 245.560 211.420 246.350 211.610 ;
        RECT 245.560 211.220 245.810 211.420 ;
        RECT 246.060 211.310 246.350 211.420 ;
        RECT 247.450 211.220 247.700 211.760 ;
        RECT 250.530 211.760 250.800 211.820 ;
        RECT 252.080 212.100 253.390 212.360 ;
        RECT 255.450 212.170 270.660 212.400 ;
        RECT 282.740 212.190 287.990 212.490 ;
        RECT 255.450 212.160 269.610 212.170 ;
        RECT 255.450 212.150 262.980 212.160 ;
        RECT 263.990 212.150 265.180 212.160 ;
        RECT 266.140 212.150 267.330 212.160 ;
        RECT 268.420 212.150 269.610 212.160 ;
        RECT 255.450 212.140 260.760 212.150 ;
        RECT 255.450 212.130 259.620 212.140 ;
        RECT 255.450 212.120 257.340 212.130 ;
        RECT 258.430 212.120 259.620 212.130 ;
        RECT 255.450 212.110 256.170 212.120 ;
        RECT 252.080 211.760 252.390 212.100 ;
        RECT 248.090 211.230 249.730 211.620 ;
        RECT 250.530 211.470 252.390 211.760 ;
        RECT 250.530 211.460 250.840 211.470 ;
        RECT 252.080 211.460 252.390 211.470 ;
        RECT 240.670 211.110 241.320 211.120 ;
        RECT 240.670 210.780 240.970 211.110 ;
        RECT 239.950 210.330 240.970 210.780 ;
        RECT 245.560 210.620 245.850 211.220 ;
        RECT 247.450 210.620 247.740 211.220 ;
        RECT 240.670 210.320 240.970 210.330 ;
        RECT 249.790 210.010 250.090 211.010 ;
        RECT 250.540 210.410 250.840 211.460 ;
        RECT 253.140 210.360 253.390 212.100 ;
        RECT 253.840 210.010 254.100 211.560 ;
        RECT 278.660 210.550 278.920 211.750 ;
        RECT 278.660 210.040 278.910 210.550 ;
        RECT 280.550 210.540 280.810 211.750 ;
        RECT 282.940 210.640 283.190 212.190 ;
        RECT 280.550 210.380 280.940 210.540 ;
        RECT 280.540 210.250 280.940 210.380 ;
        RECT 283.640 210.250 283.900 211.860 ;
        RECT 286.190 210.790 286.490 211.840 ;
        RECT 286.940 211.240 287.240 212.190 ;
        RECT 287.440 211.290 287.740 211.340 ;
        RECT 287.440 210.940 288.340 211.290 ;
        RECT 279.160 210.040 279.450 210.200 ;
        RECT 280.540 210.190 280.800 210.250 ;
        RECT 249.740 210.000 254.990 210.010 ;
        RECT 239.620 209.920 239.870 209.930 ;
        RECT 239.620 209.460 240.600 209.920 ;
        RECT 249.740 209.710 255.010 210.000 ;
        RECT 239.620 209.160 239.870 209.460 ;
        RECT 247.590 209.370 249.430 209.380 ;
        RECT 254.840 209.370 255.010 209.710 ;
        RECT 241.330 209.360 241.570 209.370 ;
        RECT 242.410 209.360 255.010 209.370 ;
        RECT 241.330 209.200 255.010 209.360 ;
        RECT 278.660 209.850 279.450 210.040 ;
        RECT 278.660 209.650 278.910 209.850 ;
        RECT 279.160 209.740 279.450 209.850 ;
        RECT 280.550 209.650 280.800 210.190 ;
        RECT 283.630 210.190 283.900 210.250 ;
        RECT 285.180 210.530 286.490 210.790 ;
        RECT 288.550 210.840 290.220 210.860 ;
        RECT 305.360 210.840 305.670 222.190 ;
        RECT 288.550 210.550 305.710 210.840 ;
        RECT 289.240 210.540 305.710 210.550 ;
        RECT 285.180 210.190 285.490 210.530 ;
        RECT 281.190 209.660 282.830 210.050 ;
        RECT 283.630 209.900 285.490 210.190 ;
        RECT 283.630 209.890 283.940 209.900 ;
        RECT 285.180 209.890 285.490 209.900 ;
        RECT 241.330 209.190 252.840 209.200 ;
        RECT 241.320 209.180 247.640 209.190 ;
        RECT 249.190 209.180 252.840 209.190 ;
        RECT 241.320 209.170 243.190 209.180 ;
        RECT 241.320 209.160 241.570 209.170 ;
        RECT 239.620 208.990 241.570 209.160 ;
        RECT 278.660 209.050 278.950 209.650 ;
        RECT 280.550 209.050 280.840 209.650 ;
        RECT 239.620 208.770 239.870 208.990 ;
        RECT 239.620 208.600 240.660 208.770 ;
        RECT 240.470 207.740 240.660 208.600 ;
        RECT 282.890 208.440 283.190 209.440 ;
        RECT 283.640 208.840 283.940 209.890 ;
        RECT 286.240 208.790 286.490 210.530 ;
        RECT 286.940 208.440 287.200 209.990 ;
        RECT 287.820 208.440 288.160 208.510 ;
        RECT 282.840 208.140 288.160 208.440 ;
        RECT 239.680 207.300 240.660 207.740 ;
        RECT 239.680 207.290 240.630 207.300 ;
        RECT 241.500 206.980 250.770 206.990 ;
        RECT 252.650 206.980 254.570 206.990 ;
        RECT 239.350 206.880 239.540 206.890 ;
        RECT 239.350 206.420 240.330 206.880 ;
        RECT 241.500 206.790 254.570 206.980 ;
        RECT 241.500 206.780 253.860 206.790 ;
        RECT 239.350 205.630 239.540 206.420 ;
        RECT 241.500 205.770 241.710 206.780 ;
        RECT 250.760 206.770 252.660 206.780 ;
        RECT 254.390 206.040 254.570 206.790 ;
        RECT 240.350 205.630 240.620 205.640 ;
        RECT 239.350 205.420 240.620 205.630 ;
        RECT 240.350 205.210 240.620 205.420 ;
        RECT 240.350 204.580 240.600 205.210 ;
        RECT 241.500 204.760 241.700 205.770 ;
        RECT 249.310 205.740 254.570 206.040 ;
        RECT 239.560 204.130 240.600 204.580 ;
        RECT 239.540 202.680 240.500 203.130 ;
        RECT 240.250 202.630 240.500 202.680 ;
        RECT 241.510 202.630 241.700 204.760 ;
        RECT 240.250 202.430 241.700 202.630 ;
        RECT 245.230 204.100 245.490 205.300 ;
        RECT 245.230 203.590 245.480 204.100 ;
        RECT 247.120 204.090 247.380 205.300 ;
        RECT 249.510 204.190 249.760 205.740 ;
        RECT 247.120 203.930 247.510 204.090 ;
        RECT 247.110 203.800 247.510 203.930 ;
        RECT 250.210 203.800 250.470 205.410 ;
        RECT 252.760 204.340 253.060 205.390 ;
        RECT 253.510 204.790 253.810 205.740 ;
        RECT 254.010 204.840 254.310 204.890 ;
        RECT 254.010 204.490 254.910 204.840 ;
        RECT 256.620 204.710 256.840 204.720 ;
        RECT 256.620 204.520 270.300 204.710 ;
        RECT 256.620 204.390 256.840 204.520 ;
        RECT 245.730 203.590 246.020 203.750 ;
        RECT 247.110 203.740 247.370 203.800 ;
        RECT 245.230 203.400 246.020 203.590 ;
        RECT 245.230 203.200 245.480 203.400 ;
        RECT 245.730 203.290 246.020 203.400 ;
        RECT 247.120 203.200 247.370 203.740 ;
        RECT 250.200 203.740 250.470 203.800 ;
        RECT 251.750 204.080 253.060 204.340 ;
        RECT 255.160 204.090 256.840 204.390 ;
        RECT 255.160 204.080 256.820 204.090 ;
        RECT 251.750 203.740 252.060 204.080 ;
        RECT 247.760 203.210 249.400 203.600 ;
        RECT 250.200 203.450 252.060 203.740 ;
        RECT 250.200 203.440 250.510 203.450 ;
        RECT 251.750 203.440 252.060 203.450 ;
        RECT 245.230 202.600 245.520 203.200 ;
        RECT 247.120 202.600 247.410 203.200 ;
        RECT 240.250 202.340 240.500 202.430 ;
        RECT 239.520 201.890 240.500 202.340 ;
        RECT 249.460 201.990 249.760 202.990 ;
        RECT 250.210 202.390 250.510 203.440 ;
        RECT 252.810 202.340 253.060 204.080 ;
        RECT 270.050 203.620 270.300 204.520 ;
        RECT 253.510 201.990 253.770 203.540 ;
        RECT 264.990 203.320 270.300 203.620 ;
        RECT 249.410 201.970 254.660 201.990 ;
        RECT 249.410 201.690 254.780 201.970 ;
        RECT 242.860 201.290 243.140 201.360 ;
        RECT 244.040 201.320 244.320 201.350 ;
        RECT 254.490 201.320 254.780 201.690 ;
        RECT 244.040 201.310 254.780 201.320 ;
        RECT 241.450 201.090 243.140 201.290 ;
        RECT 240.240 200.890 240.520 200.900 ;
        RECT 239.500 200.440 240.520 200.890 ;
        RECT 241.450 200.440 241.680 201.090 ;
        RECT 242.860 201.030 243.140 201.090 ;
        RECT 244.020 201.080 254.780 201.310 ;
        RECT 244.040 201.070 254.780 201.080 ;
        RECT 260.910 201.680 261.170 202.880 ;
        RECT 260.910 201.170 261.160 201.680 ;
        RECT 262.800 201.670 263.060 202.880 ;
        RECT 265.190 201.770 265.440 203.320 ;
        RECT 262.800 201.510 263.190 201.670 ;
        RECT 262.790 201.380 263.190 201.510 ;
        RECT 265.890 201.380 266.150 202.990 ;
        RECT 268.440 201.920 268.740 202.970 ;
        RECT 269.190 202.370 269.490 203.320 ;
        RECT 269.690 202.420 269.990 202.470 ;
        RECT 269.690 202.070 270.590 202.420 ;
        RECT 287.820 202.020 288.160 208.140 ;
        RECT 319.560 205.340 319.740 224.600 ;
        RECT 319.540 204.290 319.750 205.340 ;
        RECT 319.540 204.210 319.760 204.290 ;
        RECT 319.550 202.140 319.760 204.210 ;
        RECT 319.540 202.100 319.760 202.140 ;
        RECT 287.250 202.000 288.210 202.020 ;
        RECT 271.730 201.980 276.010 201.990 ;
        RECT 283.410 201.980 288.210 202.000 ;
        RECT 271.730 201.970 288.210 201.980 ;
        RECT 261.410 201.170 261.700 201.330 ;
        RECT 262.790 201.320 263.050 201.380 ;
        RECT 244.040 201.060 254.740 201.070 ;
        RECT 244.040 201.020 244.320 201.060 ;
        RECT 260.910 200.980 261.700 201.170 ;
        RECT 260.910 200.780 261.160 200.980 ;
        RECT 261.410 200.870 261.700 200.980 ;
        RECT 262.800 200.780 263.050 201.320 ;
        RECT 265.880 201.320 266.150 201.380 ;
        RECT 267.430 201.660 268.740 201.920 ;
        RECT 267.430 201.320 267.740 201.660 ;
        RECT 263.440 200.790 265.080 201.180 ;
        RECT 265.880 201.030 267.740 201.320 ;
        RECT 265.880 201.020 266.190 201.030 ;
        RECT 267.430 201.020 267.740 201.030 ;
        RECT 242.840 200.460 243.110 200.540 ;
        RECT 240.240 200.230 241.680 200.440 ;
        RECT 242.230 200.240 243.110 200.460 ;
        RECT 240.240 199.180 240.520 200.230 ;
        RECT 242.230 199.430 242.450 200.240 ;
        RECT 242.840 200.210 243.110 200.240 ;
        RECT 243.970 200.500 244.260 200.550 ;
        RECT 243.970 200.320 254.720 200.500 ;
        RECT 243.970 200.220 244.260 200.320 ;
        RECT 248.810 200.310 252.440 200.320 ;
        RECT 254.520 199.640 254.720 200.320 ;
        RECT 260.910 200.180 261.200 200.780 ;
        RECT 262.800 200.180 263.090 200.780 ;
        RECT 239.520 198.730 240.520 199.180 ;
        RECT 239.500 197.280 240.800 197.730 ;
        RECT 240.500 196.880 240.800 197.280 ;
        RECT 242.220 196.900 242.450 199.430 ;
        RECT 249.470 199.340 254.720 199.640 ;
        RECT 265.140 199.570 265.440 200.570 ;
        RECT 265.890 199.970 266.190 201.020 ;
        RECT 268.490 199.920 268.740 201.660 ;
        RECT 270.860 201.660 288.210 201.970 ;
        RECT 270.860 201.650 283.870 201.660 ;
        RECT 275.720 201.640 283.870 201.650 ;
        RECT 287.250 201.620 288.210 201.660 ;
        RECT 287.820 201.610 288.160 201.620 ;
        RECT 269.190 199.570 269.450 201.120 ;
        RECT 319.540 200.250 319.750 202.100 ;
        RECT 314.500 199.950 319.750 200.250 ;
        RECT 270.280 199.570 270.480 199.580 ;
        RECT 241.290 196.880 242.450 196.900 ;
        RECT 240.500 196.700 242.450 196.880 ;
        RECT 245.390 197.700 245.650 198.900 ;
        RECT 245.390 197.190 245.640 197.700 ;
        RECT 247.280 197.690 247.540 198.900 ;
        RECT 249.670 197.790 249.920 199.340 ;
        RECT 247.280 197.530 247.670 197.690 ;
        RECT 247.270 197.400 247.670 197.530 ;
        RECT 250.370 197.400 250.630 199.010 ;
        RECT 252.920 197.940 253.220 198.990 ;
        RECT 253.670 198.390 253.970 199.340 ;
        RECT 254.520 199.330 254.720 199.340 ;
        RECT 265.090 199.270 270.480 199.570 ;
        RECT 254.170 198.440 254.470 198.490 ;
        RECT 254.170 198.090 255.070 198.440 ;
        RECT 270.280 198.030 270.480 199.270 ;
        RECT 310.420 198.310 310.680 199.510 ;
        RECT 262.720 198.010 263.910 198.020 ;
        RECT 264.900 198.010 266.090 198.020 ;
        RECT 267.120 198.010 268.310 198.020 ;
        RECT 269.300 198.010 270.490 198.030 ;
        RECT 260.510 198.000 270.490 198.010 ;
        RECT 257.120 197.980 258.310 197.990 ;
        RECT 259.400 197.980 270.490 198.000 ;
        RECT 245.890 197.190 246.180 197.350 ;
        RECT 247.270 197.340 247.530 197.400 ;
        RECT 245.390 197.000 246.180 197.190 ;
        RECT 245.390 196.800 245.640 197.000 ;
        RECT 245.890 196.890 246.180 197.000 ;
        RECT 247.280 196.800 247.530 197.340 ;
        RECT 250.360 197.340 250.630 197.400 ;
        RECT 251.910 197.680 253.220 197.940 ;
        RECT 255.280 197.750 270.490 197.980 ;
        RECT 310.420 197.800 310.670 198.310 ;
        RECT 312.310 198.300 312.570 199.510 ;
        RECT 314.700 198.400 314.950 199.950 ;
        RECT 312.310 198.140 312.700 198.300 ;
        RECT 312.300 198.010 312.700 198.140 ;
        RECT 315.400 198.010 315.660 199.620 ;
        RECT 317.950 198.550 318.250 199.600 ;
        RECT 318.700 199.000 319.000 199.950 ;
        RECT 319.540 199.940 319.750 199.950 ;
        RECT 319.200 199.050 319.500 199.100 ;
        RECT 319.200 198.700 320.100 199.050 ;
        RECT 321.060 198.580 336.050 198.650 ;
        RECT 310.920 197.800 311.210 197.960 ;
        RECT 312.300 197.950 312.560 198.010 ;
        RECT 255.280 197.740 269.440 197.750 ;
        RECT 255.280 197.730 262.810 197.740 ;
        RECT 263.820 197.730 265.010 197.740 ;
        RECT 265.970 197.730 267.160 197.740 ;
        RECT 268.250 197.730 269.440 197.740 ;
        RECT 255.280 197.720 260.590 197.730 ;
        RECT 255.280 197.710 259.450 197.720 ;
        RECT 255.280 197.700 257.170 197.710 ;
        RECT 258.260 197.700 259.450 197.710 ;
        RECT 255.280 197.690 256.000 197.700 ;
        RECT 251.910 197.340 252.220 197.680 ;
        RECT 247.920 196.810 249.560 197.200 ;
        RECT 250.360 197.050 252.220 197.340 ;
        RECT 250.360 197.040 250.670 197.050 ;
        RECT 251.910 197.040 252.220 197.050 ;
        RECT 240.500 196.690 241.150 196.700 ;
        RECT 240.500 196.360 240.800 196.690 ;
        RECT 239.780 195.910 240.800 196.360 ;
        RECT 245.390 196.200 245.680 196.800 ;
        RECT 247.280 196.200 247.570 196.800 ;
        RECT 240.500 195.900 240.800 195.910 ;
        RECT 249.620 195.590 249.920 196.590 ;
        RECT 250.370 195.990 250.670 197.040 ;
        RECT 252.970 195.940 253.220 197.680 ;
        RECT 310.420 197.610 311.210 197.800 ;
        RECT 310.420 197.410 310.670 197.610 ;
        RECT 310.920 197.500 311.210 197.610 ;
        RECT 312.310 197.410 312.560 197.950 ;
        RECT 315.390 197.950 315.660 198.010 ;
        RECT 316.940 198.290 318.250 198.550 ;
        RECT 320.390 198.330 336.050 198.580 ;
        RECT 320.390 198.300 321.210 198.330 ;
        RECT 316.940 197.950 317.250 198.290 ;
        RECT 312.950 197.420 314.590 197.810 ;
        RECT 315.390 197.660 317.250 197.950 ;
        RECT 315.390 197.650 315.700 197.660 ;
        RECT 316.940 197.650 317.250 197.660 ;
        RECT 253.670 195.590 253.930 197.140 ;
        RECT 310.420 196.810 310.710 197.410 ;
        RECT 312.310 196.810 312.600 197.410 ;
        RECT 314.650 196.200 314.950 197.200 ;
        RECT 315.400 196.600 315.700 197.650 ;
        RECT 318.000 196.550 318.250 198.290 ;
        RECT 335.800 198.120 336.050 198.330 ;
        RECT 318.700 196.200 318.960 197.750 ;
        RECT 335.800 196.280 336.070 198.120 ;
        RECT 319.660 196.200 319.840 196.210 ;
        RECT 314.600 195.900 319.850 196.200 ;
        RECT 249.570 195.580 254.820 195.590 ;
        RECT 239.450 195.500 239.700 195.510 ;
        RECT 239.450 195.040 240.430 195.500 ;
        RECT 249.570 195.290 254.840 195.580 ;
        RECT 239.450 194.740 239.700 195.040 ;
        RECT 247.420 194.950 249.260 194.960 ;
        RECT 254.670 194.950 254.840 195.290 ;
        RECT 241.160 194.940 241.400 194.950 ;
        RECT 242.240 194.940 254.840 194.950 ;
        RECT 241.160 194.780 254.840 194.940 ;
        RECT 241.160 194.770 252.670 194.780 ;
        RECT 241.150 194.760 247.470 194.770 ;
        RECT 249.020 194.760 252.670 194.770 ;
        RECT 241.150 194.750 243.020 194.760 ;
        RECT 241.150 194.740 241.400 194.750 ;
        RECT 239.450 194.570 241.400 194.740 ;
        RECT 239.450 194.270 239.720 194.570 ;
        RECT 239.460 194.010 239.720 194.270 ;
        RECT 239.440 193.620 239.740 194.010 ;
        RECT 239.430 193.220 239.740 193.620 ;
        RECT 239.420 192.460 239.730 193.220 ;
        RECT 239.320 192.440 239.730 192.460 ;
        RECT 239.290 191.490 239.740 192.440 ;
        RECT 240.150 191.200 240.610 192.140 ;
        RECT 241.350 191.550 250.620 191.560 ;
        RECT 252.500 191.550 254.420 191.560 ;
        RECT 241.350 191.360 254.420 191.550 ;
        RECT 241.350 191.350 253.710 191.360 ;
        RECT 240.190 190.880 240.490 191.200 ;
        RECT 240.190 190.550 240.480 190.880 ;
        RECT 240.200 189.750 240.460 190.550 ;
        RECT 241.350 190.340 241.560 191.350 ;
        RECT 250.610 191.340 252.510 191.350 ;
        RECT 254.240 190.610 254.420 191.360 ;
        RECT 240.200 189.150 240.450 189.750 ;
        RECT 241.350 189.330 241.550 190.340 ;
        RECT 249.160 190.310 254.420 190.610 ;
        RECT 239.410 188.700 240.450 189.150 ;
        RECT 239.390 187.250 240.350 187.700 ;
        RECT 240.100 187.200 240.350 187.250 ;
        RECT 241.360 187.200 241.550 189.330 ;
        RECT 240.100 187.000 241.550 187.200 ;
        RECT 245.080 188.670 245.340 189.870 ;
        RECT 245.080 188.160 245.330 188.670 ;
        RECT 246.970 188.660 247.230 189.870 ;
        RECT 249.360 188.760 249.610 190.310 ;
        RECT 246.970 188.500 247.360 188.660 ;
        RECT 246.960 188.370 247.360 188.500 ;
        RECT 250.060 188.370 250.320 189.980 ;
        RECT 252.610 188.910 252.910 189.960 ;
        RECT 253.360 189.360 253.660 190.310 ;
        RECT 253.860 189.410 254.160 189.460 ;
        RECT 253.860 189.060 254.760 189.410 ;
        RECT 256.470 189.280 256.690 189.290 ;
        RECT 256.470 189.090 270.150 189.280 ;
        RECT 256.470 188.960 256.690 189.090 ;
        RECT 245.580 188.160 245.870 188.320 ;
        RECT 246.960 188.310 247.220 188.370 ;
        RECT 245.080 187.970 245.870 188.160 ;
        RECT 245.080 187.770 245.330 187.970 ;
        RECT 245.580 187.860 245.870 187.970 ;
        RECT 246.970 187.770 247.220 188.310 ;
        RECT 250.050 188.310 250.320 188.370 ;
        RECT 251.600 188.650 252.910 188.910 ;
        RECT 255.010 188.660 256.690 188.960 ;
        RECT 255.010 188.650 256.670 188.660 ;
        RECT 251.600 188.310 251.910 188.650 ;
        RECT 247.610 187.780 249.250 188.170 ;
        RECT 250.050 188.020 251.910 188.310 ;
        RECT 250.050 188.010 250.360 188.020 ;
        RECT 251.600 188.010 251.910 188.020 ;
        RECT 245.080 187.170 245.370 187.770 ;
        RECT 246.970 187.170 247.260 187.770 ;
        RECT 240.100 186.910 240.350 187.000 ;
        RECT 239.370 186.460 240.350 186.910 ;
        RECT 249.310 186.560 249.610 187.560 ;
        RECT 250.060 186.960 250.360 188.010 ;
        RECT 252.660 186.910 252.910 188.650 ;
        RECT 269.900 188.190 270.150 189.090 ;
        RECT 253.360 186.560 253.620 188.110 ;
        RECT 264.840 187.890 270.150 188.190 ;
        RECT 249.260 186.540 254.510 186.560 ;
        RECT 249.260 186.260 254.630 186.540 ;
        RECT 242.710 185.860 242.990 185.930 ;
        RECT 243.890 185.890 244.170 185.920 ;
        RECT 254.340 185.890 254.630 186.260 ;
        RECT 243.890 185.880 254.630 185.890 ;
        RECT 241.300 185.660 242.990 185.860 ;
        RECT 240.090 185.460 240.370 185.470 ;
        RECT 239.350 185.010 240.370 185.460 ;
        RECT 241.300 185.010 241.530 185.660 ;
        RECT 242.710 185.600 242.990 185.660 ;
        RECT 243.870 185.650 254.630 185.880 ;
        RECT 243.890 185.640 254.630 185.650 ;
        RECT 260.760 186.250 261.020 187.450 ;
        RECT 260.760 185.740 261.010 186.250 ;
        RECT 262.650 186.240 262.910 187.450 ;
        RECT 265.040 186.340 265.290 187.890 ;
        RECT 262.650 186.080 263.040 186.240 ;
        RECT 262.640 185.950 263.040 186.080 ;
        RECT 265.740 185.950 266.000 187.560 ;
        RECT 268.290 186.490 268.590 187.540 ;
        RECT 269.040 186.940 269.340 187.890 ;
        RECT 269.540 186.990 269.840 187.040 ;
        RECT 269.540 186.640 270.440 186.990 ;
        RECT 283.200 186.590 287.670 186.620 ;
        RECT 272.260 186.560 287.670 186.590 ;
        RECT 271.590 186.540 287.670 186.560 ;
        RECT 261.260 185.740 261.550 185.900 ;
        RECT 262.640 185.890 262.900 185.950 ;
        RECT 243.890 185.630 254.590 185.640 ;
        RECT 243.890 185.590 244.170 185.630 ;
        RECT 260.760 185.550 261.550 185.740 ;
        RECT 260.760 185.350 261.010 185.550 ;
        RECT 261.260 185.440 261.550 185.550 ;
        RECT 262.650 185.350 262.900 185.890 ;
        RECT 265.730 185.890 266.000 185.950 ;
        RECT 267.280 186.230 268.590 186.490 ;
        RECT 267.280 185.890 267.590 186.230 ;
        RECT 263.290 185.360 264.930 185.750 ;
        RECT 265.730 185.600 267.590 185.890 ;
        RECT 265.730 185.590 266.040 185.600 ;
        RECT 267.280 185.590 267.590 185.600 ;
        RECT 242.690 185.030 242.960 185.110 ;
        RECT 240.090 184.800 241.530 185.010 ;
        RECT 242.080 184.810 242.960 185.030 ;
        RECT 240.090 183.750 240.370 184.800 ;
        RECT 242.080 184.000 242.300 184.810 ;
        RECT 242.690 184.780 242.960 184.810 ;
        RECT 243.820 185.070 244.110 185.120 ;
        RECT 243.820 184.890 254.570 185.070 ;
        RECT 243.820 184.790 244.110 184.890 ;
        RECT 248.660 184.880 252.290 184.890 ;
        RECT 254.370 184.210 254.570 184.890 ;
        RECT 260.760 184.750 261.050 185.350 ;
        RECT 262.650 184.750 262.940 185.350 ;
        RECT 239.370 183.300 240.370 183.750 ;
        RECT 239.350 181.850 240.650 182.300 ;
        RECT 240.350 181.450 240.650 181.850 ;
        RECT 242.070 181.470 242.300 184.000 ;
        RECT 249.320 183.910 254.570 184.210 ;
        RECT 264.990 184.140 265.290 185.140 ;
        RECT 265.740 184.540 266.040 185.590 ;
        RECT 268.340 184.490 268.590 186.230 ;
        RECT 270.710 186.220 287.670 186.540 ;
        RECT 319.660 186.240 319.840 195.900 ;
        RECT 271.590 186.210 287.670 186.220 ;
        RECT 271.590 186.180 283.570 186.210 ;
        RECT 271.590 186.170 272.480 186.180 ;
        RECT 269.040 184.140 269.300 185.690 ;
        RECT 270.130 184.140 270.330 184.150 ;
        RECT 241.140 181.450 242.300 181.470 ;
        RECT 240.350 181.270 242.300 181.450 ;
        RECT 245.240 182.270 245.500 183.470 ;
        RECT 245.240 181.760 245.490 182.270 ;
        RECT 247.130 182.260 247.390 183.470 ;
        RECT 249.520 182.360 249.770 183.910 ;
        RECT 247.130 182.100 247.520 182.260 ;
        RECT 247.120 181.970 247.520 182.100 ;
        RECT 250.220 181.970 250.480 183.580 ;
        RECT 252.770 182.510 253.070 183.560 ;
        RECT 253.520 182.960 253.820 183.910 ;
        RECT 254.370 183.900 254.570 183.910 ;
        RECT 264.940 183.840 270.330 184.140 ;
        RECT 254.020 183.010 254.320 183.060 ;
        RECT 254.020 182.660 254.920 183.010 ;
        RECT 270.130 182.600 270.330 183.840 ;
        RECT 287.290 182.640 287.650 186.210 ;
        RECT 262.570 182.580 263.760 182.590 ;
        RECT 264.750 182.580 265.940 182.590 ;
        RECT 266.970 182.580 268.160 182.590 ;
        RECT 269.150 182.580 270.340 182.600 ;
        RECT 260.360 182.570 270.340 182.580 ;
        RECT 256.970 182.550 258.160 182.560 ;
        RECT 259.250 182.550 270.340 182.570 ;
        RECT 245.740 181.760 246.030 181.920 ;
        RECT 247.120 181.910 247.380 181.970 ;
        RECT 245.240 181.570 246.030 181.760 ;
        RECT 245.240 181.370 245.490 181.570 ;
        RECT 245.740 181.460 246.030 181.570 ;
        RECT 247.130 181.370 247.380 181.910 ;
        RECT 250.210 181.910 250.480 181.970 ;
        RECT 251.760 182.250 253.070 182.510 ;
        RECT 255.130 182.320 270.340 182.550 ;
        RECT 282.420 182.340 287.670 182.640 ;
        RECT 255.130 182.310 269.290 182.320 ;
        RECT 255.130 182.300 262.660 182.310 ;
        RECT 263.670 182.300 264.860 182.310 ;
        RECT 265.820 182.300 267.010 182.310 ;
        RECT 268.100 182.300 269.290 182.310 ;
        RECT 255.130 182.290 260.440 182.300 ;
        RECT 255.130 182.280 259.300 182.290 ;
        RECT 255.130 182.270 257.020 182.280 ;
        RECT 258.110 182.270 259.300 182.280 ;
        RECT 255.130 182.260 255.850 182.270 ;
        RECT 251.760 181.910 252.070 182.250 ;
        RECT 247.770 181.380 249.410 181.770 ;
        RECT 250.210 181.620 252.070 181.910 ;
        RECT 250.210 181.610 250.520 181.620 ;
        RECT 251.760 181.610 252.070 181.620 ;
        RECT 240.350 181.260 241.000 181.270 ;
        RECT 240.350 180.930 240.650 181.260 ;
        RECT 239.630 180.480 240.650 180.930 ;
        RECT 245.240 180.770 245.530 181.370 ;
        RECT 247.130 180.770 247.420 181.370 ;
        RECT 240.350 180.470 240.650 180.480 ;
        RECT 249.470 180.160 249.770 181.160 ;
        RECT 250.220 180.560 250.520 181.610 ;
        RECT 252.820 180.510 253.070 182.250 ;
        RECT 253.520 180.160 253.780 181.710 ;
        RECT 278.340 180.700 278.600 181.900 ;
        RECT 278.340 180.190 278.590 180.700 ;
        RECT 280.230 180.690 280.490 181.900 ;
        RECT 282.620 180.790 282.870 182.340 ;
        RECT 280.230 180.530 280.620 180.690 ;
        RECT 280.220 180.400 280.620 180.530 ;
        RECT 283.320 180.400 283.580 182.010 ;
        RECT 285.870 180.940 286.170 181.990 ;
        RECT 286.620 181.390 286.920 182.340 ;
        RECT 287.120 181.440 287.420 181.490 ;
        RECT 287.120 181.090 288.020 181.440 ;
        RECT 278.840 180.190 279.130 180.350 ;
        RECT 280.220 180.340 280.480 180.400 ;
        RECT 249.420 180.150 254.670 180.160 ;
        RECT 239.300 180.070 239.550 180.080 ;
        RECT 239.300 179.610 240.280 180.070 ;
        RECT 249.420 179.860 254.690 180.150 ;
        RECT 239.300 179.310 239.550 179.610 ;
        RECT 247.270 179.520 249.110 179.530 ;
        RECT 254.520 179.520 254.690 179.860 ;
        RECT 241.010 179.510 241.250 179.520 ;
        RECT 242.090 179.510 254.690 179.520 ;
        RECT 241.010 179.350 254.690 179.510 ;
        RECT 278.340 180.000 279.130 180.190 ;
        RECT 278.340 179.800 278.590 180.000 ;
        RECT 278.840 179.890 279.130 180.000 ;
        RECT 280.230 179.800 280.480 180.340 ;
        RECT 283.310 180.340 283.580 180.400 ;
        RECT 284.860 180.680 286.170 180.940 ;
        RECT 288.230 180.980 289.900 181.010 ;
        RECT 304.980 180.980 305.230 180.990 ;
        RECT 288.230 180.710 305.230 180.980 ;
        RECT 288.230 180.700 301.730 180.710 ;
        RECT 289.510 180.680 301.730 180.700 ;
        RECT 284.860 180.340 285.170 180.680 ;
        RECT 280.870 179.810 282.510 180.200 ;
        RECT 283.310 180.050 285.170 180.340 ;
        RECT 283.310 180.040 283.620 180.050 ;
        RECT 284.860 180.040 285.170 180.050 ;
        RECT 241.010 179.340 252.520 179.350 ;
        RECT 241.000 179.330 247.320 179.340 ;
        RECT 248.870 179.330 252.520 179.340 ;
        RECT 241.000 179.320 242.870 179.330 ;
        RECT 241.000 179.310 241.250 179.320 ;
        RECT 239.300 179.140 241.250 179.310 ;
        RECT 278.340 179.200 278.630 179.800 ;
        RECT 280.230 179.200 280.520 179.800 ;
        RECT 239.300 178.920 239.550 179.140 ;
        RECT 239.300 178.750 240.340 178.920 ;
        RECT 240.150 177.890 240.340 178.750 ;
        RECT 282.570 178.590 282.870 179.590 ;
        RECT 283.320 178.990 283.620 180.040 ;
        RECT 285.920 178.940 286.170 180.680 ;
        RECT 286.620 178.590 286.880 180.140 ;
        RECT 287.500 178.590 287.840 178.660 ;
        RECT 282.520 178.290 287.840 178.590 ;
        RECT 239.360 177.450 240.340 177.890 ;
        RECT 239.360 177.440 240.310 177.450 ;
        RECT 241.180 177.130 250.450 177.140 ;
        RECT 252.330 177.130 254.250 177.140 ;
        RECT 239.030 177.030 239.220 177.040 ;
        RECT 239.030 176.570 240.010 177.030 ;
        RECT 241.180 176.940 254.250 177.130 ;
        RECT 241.180 176.930 253.540 176.940 ;
        RECT 239.030 175.780 239.220 176.570 ;
        RECT 241.180 175.920 241.390 176.930 ;
        RECT 250.440 176.920 252.340 176.930 ;
        RECT 254.070 176.190 254.250 176.940 ;
        RECT 240.030 175.780 240.300 175.790 ;
        RECT 239.030 175.570 240.300 175.780 ;
        RECT 240.030 175.360 240.300 175.570 ;
        RECT 240.030 174.730 240.280 175.360 ;
        RECT 241.180 174.910 241.380 175.920 ;
        RECT 248.990 175.890 254.250 176.190 ;
        RECT 239.240 174.280 240.280 174.730 ;
        RECT 239.220 172.830 240.180 173.280 ;
        RECT 239.930 172.780 240.180 172.830 ;
        RECT 241.190 172.780 241.380 174.910 ;
        RECT 239.930 172.580 241.380 172.780 ;
        RECT 244.910 174.250 245.170 175.450 ;
        RECT 244.910 173.740 245.160 174.250 ;
        RECT 246.800 174.240 247.060 175.450 ;
        RECT 249.190 174.340 249.440 175.890 ;
        RECT 246.800 174.080 247.190 174.240 ;
        RECT 246.790 173.950 247.190 174.080 ;
        RECT 249.890 173.950 250.150 175.560 ;
        RECT 252.440 174.490 252.740 175.540 ;
        RECT 253.190 174.940 253.490 175.890 ;
        RECT 253.690 174.990 253.990 175.040 ;
        RECT 253.690 174.640 254.590 174.990 ;
        RECT 256.300 174.860 256.520 174.870 ;
        RECT 256.300 174.670 269.980 174.860 ;
        RECT 256.300 174.540 256.520 174.670 ;
        RECT 245.410 173.740 245.700 173.900 ;
        RECT 246.790 173.890 247.050 173.950 ;
        RECT 244.910 173.550 245.700 173.740 ;
        RECT 244.910 173.350 245.160 173.550 ;
        RECT 245.410 173.440 245.700 173.550 ;
        RECT 246.800 173.350 247.050 173.890 ;
        RECT 249.880 173.890 250.150 173.950 ;
        RECT 251.430 174.230 252.740 174.490 ;
        RECT 254.840 174.240 256.520 174.540 ;
        RECT 254.840 174.230 256.500 174.240 ;
        RECT 251.430 173.890 251.740 174.230 ;
        RECT 247.440 173.360 249.080 173.750 ;
        RECT 249.880 173.600 251.740 173.890 ;
        RECT 249.880 173.590 250.190 173.600 ;
        RECT 251.430 173.590 251.740 173.600 ;
        RECT 244.910 172.750 245.200 173.350 ;
        RECT 246.800 172.750 247.090 173.350 ;
        RECT 239.930 172.490 240.180 172.580 ;
        RECT 239.200 172.040 240.180 172.490 ;
        RECT 249.140 172.140 249.440 173.140 ;
        RECT 249.890 172.540 250.190 173.590 ;
        RECT 252.490 172.490 252.740 174.230 ;
        RECT 269.730 173.770 269.980 174.670 ;
        RECT 253.190 172.140 253.450 173.690 ;
        RECT 264.670 173.470 269.980 173.770 ;
        RECT 249.090 172.120 254.340 172.140 ;
        RECT 249.090 171.840 254.460 172.120 ;
        RECT 242.540 171.440 242.820 171.510 ;
        RECT 243.720 171.470 244.000 171.500 ;
        RECT 254.170 171.470 254.460 171.840 ;
        RECT 243.720 171.460 254.460 171.470 ;
        RECT 241.130 171.240 242.820 171.440 ;
        RECT 239.920 171.040 240.200 171.050 ;
        RECT 239.180 170.590 240.200 171.040 ;
        RECT 241.130 170.590 241.360 171.240 ;
        RECT 242.540 171.180 242.820 171.240 ;
        RECT 243.700 171.230 254.460 171.460 ;
        RECT 243.720 171.220 254.460 171.230 ;
        RECT 260.590 171.830 260.850 173.030 ;
        RECT 260.590 171.320 260.840 171.830 ;
        RECT 262.480 171.820 262.740 173.030 ;
        RECT 264.870 171.920 265.120 173.470 ;
        RECT 262.480 171.660 262.870 171.820 ;
        RECT 262.470 171.530 262.870 171.660 ;
        RECT 265.570 171.530 265.830 173.140 ;
        RECT 268.120 172.070 268.420 173.120 ;
        RECT 268.870 172.520 269.170 173.470 ;
        RECT 269.370 172.570 269.670 172.620 ;
        RECT 269.370 172.220 270.270 172.570 ;
        RECT 287.500 172.170 287.840 178.290 ;
        RECT 286.930 172.150 287.890 172.170 ;
        RECT 271.410 172.130 275.690 172.140 ;
        RECT 283.090 172.130 287.890 172.150 ;
        RECT 271.410 172.120 287.890 172.130 ;
        RECT 261.090 171.320 261.380 171.480 ;
        RECT 262.470 171.470 262.730 171.530 ;
        RECT 243.720 171.210 254.420 171.220 ;
        RECT 243.720 171.170 244.000 171.210 ;
        RECT 260.590 171.130 261.380 171.320 ;
        RECT 260.590 170.930 260.840 171.130 ;
        RECT 261.090 171.020 261.380 171.130 ;
        RECT 262.480 170.930 262.730 171.470 ;
        RECT 265.560 171.470 265.830 171.530 ;
        RECT 267.110 171.810 268.420 172.070 ;
        RECT 267.110 171.470 267.420 171.810 ;
        RECT 263.120 170.940 264.760 171.330 ;
        RECT 265.560 171.180 267.420 171.470 ;
        RECT 265.560 171.170 265.870 171.180 ;
        RECT 267.110 171.170 267.420 171.180 ;
        RECT 242.520 170.610 242.790 170.690 ;
        RECT 239.920 170.380 241.360 170.590 ;
        RECT 241.910 170.390 242.790 170.610 ;
        RECT 239.920 169.330 240.200 170.380 ;
        RECT 241.910 169.580 242.130 170.390 ;
        RECT 242.520 170.360 242.790 170.390 ;
        RECT 243.650 170.650 243.940 170.700 ;
        RECT 243.650 170.470 254.400 170.650 ;
        RECT 243.650 170.370 243.940 170.470 ;
        RECT 248.490 170.460 252.120 170.470 ;
        RECT 254.200 169.790 254.400 170.470 ;
        RECT 260.590 170.330 260.880 170.930 ;
        RECT 262.480 170.330 262.770 170.930 ;
        RECT 239.200 168.880 240.200 169.330 ;
        RECT 239.180 167.430 240.480 167.880 ;
        RECT 240.180 167.030 240.480 167.430 ;
        RECT 241.900 167.050 242.130 169.580 ;
        RECT 249.150 169.490 254.400 169.790 ;
        RECT 264.820 169.720 265.120 170.720 ;
        RECT 265.570 170.120 265.870 171.170 ;
        RECT 268.170 170.070 268.420 171.810 ;
        RECT 270.540 171.810 287.890 172.120 ;
        RECT 270.540 171.800 283.550 171.810 ;
        RECT 275.400 171.790 283.550 171.800 ;
        RECT 286.930 171.770 287.890 171.810 ;
        RECT 287.500 171.760 287.840 171.770 ;
        RECT 268.870 169.720 269.130 171.270 ;
        RECT 269.960 169.720 270.160 169.730 ;
        RECT 240.970 167.030 242.130 167.050 ;
        RECT 240.180 166.850 242.130 167.030 ;
        RECT 245.070 167.850 245.330 169.050 ;
        RECT 245.070 167.340 245.320 167.850 ;
        RECT 246.960 167.840 247.220 169.050 ;
        RECT 249.350 167.940 249.600 169.490 ;
        RECT 246.960 167.680 247.350 167.840 ;
        RECT 246.950 167.550 247.350 167.680 ;
        RECT 250.050 167.550 250.310 169.160 ;
        RECT 252.600 168.090 252.900 169.140 ;
        RECT 253.350 168.540 253.650 169.490 ;
        RECT 254.200 169.480 254.400 169.490 ;
        RECT 264.770 169.420 270.160 169.720 ;
        RECT 253.850 168.590 254.150 168.640 ;
        RECT 253.850 168.240 254.750 168.590 ;
        RECT 269.960 168.180 270.160 169.420 ;
        RECT 262.400 168.160 263.590 168.170 ;
        RECT 264.580 168.160 265.770 168.170 ;
        RECT 266.800 168.160 267.990 168.170 ;
        RECT 268.980 168.160 270.170 168.180 ;
        RECT 260.190 168.150 270.170 168.160 ;
        RECT 256.800 168.130 257.990 168.140 ;
        RECT 259.080 168.130 270.170 168.150 ;
        RECT 245.570 167.340 245.860 167.500 ;
        RECT 246.950 167.490 247.210 167.550 ;
        RECT 245.070 167.150 245.860 167.340 ;
        RECT 245.070 166.950 245.320 167.150 ;
        RECT 245.570 167.040 245.860 167.150 ;
        RECT 246.960 166.950 247.210 167.490 ;
        RECT 250.040 167.490 250.310 167.550 ;
        RECT 251.590 167.830 252.900 168.090 ;
        RECT 254.960 167.900 270.170 168.130 ;
        RECT 254.960 167.890 269.120 167.900 ;
        RECT 254.960 167.880 262.490 167.890 ;
        RECT 263.500 167.880 264.690 167.890 ;
        RECT 265.650 167.880 266.840 167.890 ;
        RECT 267.930 167.880 269.120 167.890 ;
        RECT 254.960 167.870 260.270 167.880 ;
        RECT 254.960 167.860 259.130 167.870 ;
        RECT 254.960 167.850 256.850 167.860 ;
        RECT 257.940 167.850 259.130 167.860 ;
        RECT 254.960 167.840 255.680 167.850 ;
        RECT 251.590 167.490 251.900 167.830 ;
        RECT 247.600 166.960 249.240 167.350 ;
        RECT 250.040 167.200 251.900 167.490 ;
        RECT 250.040 167.190 250.350 167.200 ;
        RECT 251.590 167.190 251.900 167.200 ;
        RECT 240.180 166.840 240.830 166.850 ;
        RECT 240.180 166.510 240.480 166.840 ;
        RECT 239.460 166.060 240.480 166.510 ;
        RECT 245.070 166.350 245.360 166.950 ;
        RECT 246.960 166.350 247.250 166.950 ;
        RECT 240.180 166.050 240.480 166.060 ;
        RECT 249.300 165.740 249.600 166.740 ;
        RECT 250.050 166.140 250.350 167.190 ;
        RECT 252.650 166.090 252.900 167.830 ;
        RECT 304.980 167.570 305.240 180.710 ;
        RECT 304.970 167.450 305.240 167.570 ;
        RECT 319.570 176.720 319.840 186.240 ;
        RECT 335.800 192.610 336.110 196.280 ;
        RECT 335.800 190.830 336.130 192.610 ;
        RECT 335.800 188.860 336.090 190.830 ;
        RECT 335.800 187.030 336.110 188.860 ;
        RECT 335.800 183.210 336.090 187.030 ;
        RECT 335.800 181.240 336.070 183.210 ;
        RECT 335.800 179.520 336.130 181.240 ;
        RECT 335.800 177.600 336.090 179.520 ;
        RECT 253.350 165.740 253.610 167.290 ;
        RECT 304.970 166.620 305.230 167.450 ;
        RECT 319.570 166.770 319.750 176.720 ;
        RECT 335.800 168.060 336.070 177.600 ;
        RECT 299.950 166.320 305.230 166.620 ;
        RECT 249.250 165.730 254.500 165.740 ;
        RECT 239.130 165.650 239.380 165.660 ;
        RECT 239.130 165.190 240.110 165.650 ;
        RECT 249.250 165.440 254.520 165.730 ;
        RECT 239.130 164.890 239.380 165.190 ;
        RECT 247.100 165.100 248.940 165.110 ;
        RECT 254.350 165.100 254.520 165.440 ;
        RECT 240.840 165.090 241.080 165.100 ;
        RECT 241.920 165.090 254.520 165.100 ;
        RECT 240.840 164.930 254.520 165.090 ;
        RECT 240.840 164.920 252.350 164.930 ;
        RECT 240.830 164.910 247.150 164.920 ;
        RECT 248.700 164.910 252.350 164.920 ;
        RECT 240.830 164.900 242.700 164.910 ;
        RECT 240.830 164.890 241.080 164.900 ;
        RECT 239.130 164.720 241.080 164.890 ;
        RECT 239.130 164.420 239.400 164.720 ;
        RECT 239.140 164.160 239.400 164.420 ;
        RECT 295.870 164.680 296.130 165.880 ;
        RECT 295.870 164.170 296.120 164.680 ;
        RECT 297.760 164.670 298.020 165.880 ;
        RECT 300.150 164.770 300.400 166.320 ;
        RECT 297.760 164.510 298.150 164.670 ;
        RECT 297.750 164.380 298.150 164.510 ;
        RECT 300.850 164.380 301.110 165.990 ;
        RECT 303.400 164.920 303.700 165.970 ;
        RECT 304.150 165.370 304.450 166.320 ;
        RECT 304.650 165.420 304.950 165.470 ;
        RECT 304.650 165.070 305.550 165.420 ;
        RECT 319.560 164.960 319.760 166.770 ;
        RECT 296.370 164.170 296.660 164.330 ;
        RECT 297.750 164.320 298.010 164.380 ;
        RECT 239.120 163.770 239.420 164.160 ;
        RECT 295.870 163.980 296.660 164.170 ;
        RECT 295.870 163.780 296.120 163.980 ;
        RECT 296.370 163.870 296.660 163.980 ;
        RECT 297.760 163.780 298.010 164.320 ;
        RECT 300.840 164.320 301.110 164.380 ;
        RECT 302.390 164.660 303.700 164.920 ;
        RECT 305.820 164.670 319.760 164.960 ;
        RECT 335.840 166.190 336.110 168.060 ;
        RECT 305.820 164.660 319.720 164.670 ;
        RECT 302.390 164.320 302.700 164.660 ;
        RECT 298.400 163.790 300.040 164.180 ;
        RECT 300.840 164.030 302.700 164.320 ;
        RECT 300.840 164.020 301.150 164.030 ;
        RECT 302.390 164.020 302.700 164.030 ;
        RECT 239.120 163.540 240.610 163.770 ;
        RECT 240.360 162.610 240.610 163.540 ;
        RECT 295.870 163.180 296.160 163.780 ;
        RECT 297.760 163.180 298.050 163.780 ;
        RECT 239.560 162.150 240.610 162.610 ;
        RECT 300.100 162.570 300.400 163.570 ;
        RECT 300.850 162.970 301.150 164.020 ;
        RECT 303.450 162.920 303.700 164.660 ;
        RECT 306.410 164.650 319.720 164.660 ;
        RECT 304.150 162.570 304.410 164.120 ;
        RECT 300.050 162.270 305.320 162.570 ;
        RECT 240.360 162.140 240.610 162.150 ;
        RECT 239.230 161.740 239.480 161.750 ;
        RECT 239.230 161.290 240.210 161.740 ;
        RECT 241.320 161.480 250.590 161.490 ;
        RECT 252.470 161.480 254.390 161.490 ;
        RECT 241.320 161.290 254.390 161.480 ;
        RECT 239.230 160.680 239.480 161.290 ;
        RECT 241.320 161.280 253.680 161.290 ;
        RECT 239.230 160.430 240.440 160.680 ;
        RECT 240.170 159.680 240.430 160.430 ;
        RECT 241.320 160.270 241.530 161.280 ;
        RECT 250.580 161.270 252.480 161.280 ;
        RECT 254.210 160.540 254.390 161.290 ;
        RECT 240.170 159.080 240.420 159.680 ;
        RECT 241.320 159.260 241.520 160.270 ;
        RECT 249.130 160.240 254.390 160.540 ;
        RECT 239.380 158.630 240.420 159.080 ;
        RECT 239.360 157.180 240.320 157.630 ;
        RECT 240.070 157.130 240.320 157.180 ;
        RECT 241.330 157.130 241.520 159.260 ;
        RECT 240.070 156.930 241.520 157.130 ;
        RECT 245.050 158.600 245.310 159.800 ;
        RECT 245.050 158.090 245.300 158.600 ;
        RECT 246.940 158.590 247.200 159.800 ;
        RECT 249.330 158.690 249.580 160.240 ;
        RECT 246.940 158.430 247.330 158.590 ;
        RECT 246.930 158.300 247.330 158.430 ;
        RECT 250.030 158.300 250.290 159.910 ;
        RECT 252.580 158.840 252.880 159.890 ;
        RECT 253.330 159.290 253.630 160.240 ;
        RECT 253.830 159.340 254.130 159.390 ;
        RECT 253.830 158.990 254.730 159.340 ;
        RECT 256.440 159.210 256.660 159.220 ;
        RECT 256.440 159.020 270.120 159.210 ;
        RECT 256.440 158.890 256.660 159.020 ;
        RECT 245.550 158.090 245.840 158.250 ;
        RECT 246.930 158.240 247.190 158.300 ;
        RECT 245.050 157.900 245.840 158.090 ;
        RECT 245.050 157.700 245.300 157.900 ;
        RECT 245.550 157.790 245.840 157.900 ;
        RECT 246.940 157.700 247.190 158.240 ;
        RECT 250.020 158.240 250.290 158.300 ;
        RECT 251.570 158.580 252.880 158.840 ;
        RECT 254.980 158.590 256.660 158.890 ;
        RECT 254.980 158.580 256.640 158.590 ;
        RECT 251.570 158.240 251.880 158.580 ;
        RECT 247.580 157.710 249.220 158.100 ;
        RECT 250.020 157.950 251.880 158.240 ;
        RECT 250.020 157.940 250.330 157.950 ;
        RECT 251.570 157.940 251.880 157.950 ;
        RECT 245.050 157.100 245.340 157.700 ;
        RECT 246.940 157.100 247.230 157.700 ;
        RECT 240.070 156.840 240.320 156.930 ;
        RECT 239.340 156.390 240.320 156.840 ;
        RECT 249.280 156.490 249.580 157.490 ;
        RECT 250.030 156.890 250.330 157.940 ;
        RECT 252.630 156.840 252.880 158.580 ;
        RECT 269.870 158.120 270.120 159.020 ;
        RECT 253.330 156.490 253.590 158.040 ;
        RECT 264.810 157.820 270.120 158.120 ;
        RECT 249.230 156.470 254.480 156.490 ;
        RECT 249.230 156.190 254.600 156.470 ;
        RECT 242.680 155.790 242.960 155.860 ;
        RECT 243.860 155.820 244.140 155.850 ;
        RECT 254.310 155.820 254.600 156.190 ;
        RECT 243.860 155.810 254.600 155.820 ;
        RECT 241.270 155.590 242.960 155.790 ;
        RECT 240.060 155.390 240.340 155.400 ;
        RECT 239.320 154.940 240.340 155.390 ;
        RECT 241.270 154.940 241.500 155.590 ;
        RECT 242.680 155.530 242.960 155.590 ;
        RECT 243.840 155.580 254.600 155.810 ;
        RECT 243.860 155.570 254.600 155.580 ;
        RECT 260.730 156.180 260.990 157.380 ;
        RECT 260.730 155.670 260.980 156.180 ;
        RECT 262.620 156.170 262.880 157.380 ;
        RECT 265.010 156.270 265.260 157.820 ;
        RECT 262.620 156.010 263.010 156.170 ;
        RECT 262.610 155.880 263.010 156.010 ;
        RECT 265.710 155.880 265.970 157.490 ;
        RECT 268.260 156.420 268.560 157.470 ;
        RECT 269.010 156.870 269.310 157.820 ;
        RECT 269.510 156.920 269.810 156.970 ;
        RECT 269.510 156.570 270.410 156.920 ;
        RECT 283.170 156.520 287.640 156.550 ;
        RECT 272.230 156.490 287.640 156.520 ;
        RECT 271.560 156.470 287.640 156.490 ;
        RECT 261.230 155.670 261.520 155.830 ;
        RECT 262.610 155.820 262.870 155.880 ;
        RECT 243.860 155.560 254.560 155.570 ;
        RECT 243.860 155.520 244.140 155.560 ;
        RECT 260.730 155.480 261.520 155.670 ;
        RECT 260.730 155.280 260.980 155.480 ;
        RECT 261.230 155.370 261.520 155.480 ;
        RECT 262.620 155.280 262.870 155.820 ;
        RECT 265.700 155.820 265.970 155.880 ;
        RECT 267.250 156.160 268.560 156.420 ;
        RECT 267.250 155.820 267.560 156.160 ;
        RECT 263.260 155.290 264.900 155.680 ;
        RECT 265.700 155.530 267.560 155.820 ;
        RECT 265.700 155.520 266.010 155.530 ;
        RECT 267.250 155.520 267.560 155.530 ;
        RECT 242.660 154.960 242.930 155.040 ;
        RECT 240.060 154.730 241.500 154.940 ;
        RECT 242.050 154.740 242.930 154.960 ;
        RECT 240.060 153.680 240.340 154.730 ;
        RECT 242.050 153.930 242.270 154.740 ;
        RECT 242.660 154.710 242.930 154.740 ;
        RECT 243.790 155.000 244.080 155.050 ;
        RECT 243.790 154.820 254.540 155.000 ;
        RECT 243.790 154.720 244.080 154.820 ;
        RECT 248.630 154.810 252.260 154.820 ;
        RECT 254.340 154.140 254.540 154.820 ;
        RECT 260.730 154.680 261.020 155.280 ;
        RECT 262.620 154.680 262.910 155.280 ;
        RECT 239.340 153.230 240.340 153.680 ;
        RECT 239.320 151.780 240.620 152.230 ;
        RECT 240.320 151.380 240.620 151.780 ;
        RECT 242.040 151.400 242.270 153.930 ;
        RECT 249.290 153.840 254.540 154.140 ;
        RECT 264.960 154.070 265.260 155.070 ;
        RECT 265.710 154.470 266.010 155.520 ;
        RECT 268.310 154.420 268.560 156.160 ;
        RECT 270.680 156.150 287.640 156.470 ;
        RECT 271.560 156.140 287.640 156.150 ;
        RECT 271.560 156.110 283.540 156.140 ;
        RECT 271.560 156.100 272.450 156.110 ;
        RECT 269.010 154.070 269.270 155.620 ;
        RECT 270.100 154.070 270.300 154.080 ;
        RECT 241.110 151.380 242.270 151.400 ;
        RECT 240.320 151.200 242.270 151.380 ;
        RECT 245.210 152.200 245.470 153.400 ;
        RECT 245.210 151.690 245.460 152.200 ;
        RECT 247.100 152.190 247.360 153.400 ;
        RECT 249.490 152.290 249.740 153.840 ;
        RECT 247.100 152.030 247.490 152.190 ;
        RECT 247.090 151.900 247.490 152.030 ;
        RECT 250.190 151.900 250.450 153.510 ;
        RECT 252.740 152.440 253.040 153.490 ;
        RECT 253.490 152.890 253.790 153.840 ;
        RECT 254.340 153.830 254.540 153.840 ;
        RECT 264.910 153.770 270.300 154.070 ;
        RECT 253.990 152.940 254.290 152.990 ;
        RECT 253.990 152.590 254.890 152.940 ;
        RECT 270.100 152.530 270.300 153.770 ;
        RECT 287.260 152.570 287.620 156.140 ;
        RECT 262.540 152.510 263.730 152.520 ;
        RECT 264.720 152.510 265.910 152.520 ;
        RECT 266.940 152.510 268.130 152.520 ;
        RECT 269.120 152.510 270.310 152.530 ;
        RECT 260.330 152.500 270.310 152.510 ;
        RECT 256.940 152.480 258.130 152.490 ;
        RECT 259.220 152.480 270.310 152.500 ;
        RECT 245.710 151.690 246.000 151.850 ;
        RECT 247.090 151.840 247.350 151.900 ;
        RECT 245.210 151.500 246.000 151.690 ;
        RECT 245.210 151.300 245.460 151.500 ;
        RECT 245.710 151.390 246.000 151.500 ;
        RECT 247.100 151.300 247.350 151.840 ;
        RECT 250.180 151.840 250.450 151.900 ;
        RECT 251.730 152.180 253.040 152.440 ;
        RECT 255.100 152.250 270.310 152.480 ;
        RECT 282.390 152.270 287.640 152.570 ;
        RECT 255.100 152.240 269.260 152.250 ;
        RECT 255.100 152.230 262.630 152.240 ;
        RECT 263.640 152.230 264.830 152.240 ;
        RECT 265.790 152.230 266.980 152.240 ;
        RECT 268.070 152.230 269.260 152.240 ;
        RECT 255.100 152.220 260.410 152.230 ;
        RECT 255.100 152.210 259.270 152.220 ;
        RECT 255.100 152.200 256.990 152.210 ;
        RECT 258.080 152.200 259.270 152.210 ;
        RECT 255.100 152.190 255.820 152.200 ;
        RECT 251.730 151.840 252.040 152.180 ;
        RECT 247.740 151.310 249.380 151.700 ;
        RECT 250.180 151.550 252.040 151.840 ;
        RECT 250.180 151.540 250.490 151.550 ;
        RECT 251.730 151.540 252.040 151.550 ;
        RECT 240.320 151.190 240.970 151.200 ;
        RECT 240.320 150.860 240.620 151.190 ;
        RECT 239.600 150.410 240.620 150.860 ;
        RECT 245.210 150.700 245.500 151.300 ;
        RECT 247.100 150.700 247.390 151.300 ;
        RECT 240.320 150.400 240.620 150.410 ;
        RECT 249.440 150.090 249.740 151.090 ;
        RECT 250.190 150.490 250.490 151.540 ;
        RECT 252.790 150.440 253.040 152.180 ;
        RECT 253.490 150.090 253.750 151.640 ;
        RECT 278.310 150.630 278.570 151.830 ;
        RECT 278.310 150.120 278.560 150.630 ;
        RECT 280.200 150.620 280.460 151.830 ;
        RECT 282.590 150.720 282.840 152.270 ;
        RECT 280.200 150.460 280.590 150.620 ;
        RECT 280.190 150.330 280.590 150.460 ;
        RECT 283.290 150.330 283.550 151.940 ;
        RECT 285.840 150.870 286.140 151.920 ;
        RECT 286.590 151.320 286.890 152.270 ;
        RECT 287.090 151.370 287.390 151.420 ;
        RECT 287.090 151.020 287.990 151.370 ;
        RECT 278.810 150.120 279.100 150.280 ;
        RECT 280.190 150.270 280.450 150.330 ;
        RECT 249.390 150.080 254.640 150.090 ;
        RECT 239.270 150.000 239.520 150.010 ;
        RECT 239.270 149.540 240.250 150.000 ;
        RECT 249.390 149.790 254.660 150.080 ;
        RECT 239.270 149.240 239.520 149.540 ;
        RECT 247.240 149.450 249.080 149.460 ;
        RECT 254.490 149.450 254.660 149.790 ;
        RECT 240.980 149.440 241.220 149.450 ;
        RECT 242.060 149.440 254.660 149.450 ;
        RECT 240.980 149.280 254.660 149.440 ;
        RECT 278.310 149.930 279.100 150.120 ;
        RECT 278.310 149.730 278.560 149.930 ;
        RECT 278.810 149.820 279.100 149.930 ;
        RECT 280.200 149.730 280.450 150.270 ;
        RECT 283.280 150.270 283.550 150.330 ;
        RECT 284.830 150.610 286.140 150.870 ;
        RECT 288.200 150.920 289.870 150.940 ;
        RECT 305.010 150.920 305.320 162.270 ;
        RECT 335.840 160.550 336.090 166.190 ;
        RECT 337.380 166.120 337.610 251.920 ;
        RECT 341.840 251.350 342.080 252.470 ;
        RECT 341.830 251.130 342.110 251.350 ;
        RECT 343.010 251.280 352.280 251.290 ;
        RECT 354.160 251.280 356.080 251.290 ;
        RECT 341.830 250.950 342.120 251.130 ;
        RECT 341.840 250.680 342.120 250.950 ;
        RECT 343.010 251.090 356.080 251.280 ;
        RECT 343.010 251.080 355.370 251.090 ;
        RECT 341.840 250.450 342.140 250.680 ;
        RECT 341.850 250.280 342.140 250.450 ;
        RECT 341.860 249.480 342.120 250.280 ;
        RECT 343.010 250.070 343.220 251.080 ;
        RECT 352.270 251.070 354.170 251.080 ;
        RECT 355.900 250.340 356.080 251.090 ;
        RECT 341.860 248.880 342.110 249.480 ;
        RECT 343.010 249.060 343.210 250.070 ;
        RECT 350.820 250.040 356.080 250.340 ;
        RECT 341.070 248.430 342.110 248.880 ;
        RECT 341.050 246.980 342.010 247.430 ;
        RECT 341.760 246.930 342.010 246.980 ;
        RECT 343.020 246.930 343.210 249.060 ;
        RECT 341.760 246.730 343.210 246.930 ;
        RECT 346.740 248.400 347.000 249.600 ;
        RECT 346.740 247.890 346.990 248.400 ;
        RECT 348.630 248.390 348.890 249.600 ;
        RECT 351.020 248.490 351.270 250.040 ;
        RECT 348.630 248.230 349.020 248.390 ;
        RECT 348.620 248.100 349.020 248.230 ;
        RECT 351.720 248.100 351.980 249.710 ;
        RECT 354.270 248.640 354.570 249.690 ;
        RECT 355.020 249.090 355.320 250.040 ;
        RECT 355.520 249.140 355.820 249.190 ;
        RECT 355.520 248.790 356.420 249.140 ;
        RECT 358.130 249.010 358.350 249.020 ;
        RECT 358.130 248.820 371.810 249.010 ;
        RECT 358.130 248.690 358.350 248.820 ;
        RECT 347.240 247.890 347.530 248.050 ;
        RECT 348.620 248.040 348.880 248.100 ;
        RECT 346.740 247.700 347.530 247.890 ;
        RECT 346.740 247.500 346.990 247.700 ;
        RECT 347.240 247.590 347.530 247.700 ;
        RECT 348.630 247.500 348.880 248.040 ;
        RECT 351.710 248.040 351.980 248.100 ;
        RECT 353.260 248.380 354.570 248.640 ;
        RECT 356.670 248.390 358.350 248.690 ;
        RECT 356.670 248.380 358.330 248.390 ;
        RECT 353.260 248.040 353.570 248.380 ;
        RECT 349.270 247.510 350.910 247.900 ;
        RECT 351.710 247.750 353.570 248.040 ;
        RECT 351.710 247.740 352.020 247.750 ;
        RECT 353.260 247.740 353.570 247.750 ;
        RECT 346.740 246.900 347.030 247.500 ;
        RECT 348.630 246.900 348.920 247.500 ;
        RECT 341.760 246.640 342.010 246.730 ;
        RECT 341.030 246.190 342.010 246.640 ;
        RECT 350.970 246.290 351.270 247.290 ;
        RECT 351.720 246.690 352.020 247.740 ;
        RECT 354.320 246.640 354.570 248.380 ;
        RECT 371.560 247.920 371.810 248.820 ;
        RECT 355.020 246.290 355.280 247.840 ;
        RECT 366.500 247.620 371.810 247.920 ;
        RECT 350.920 246.270 356.170 246.290 ;
        RECT 350.920 245.990 356.290 246.270 ;
        RECT 344.370 245.590 344.650 245.660 ;
        RECT 345.550 245.620 345.830 245.650 ;
        RECT 356.000 245.620 356.290 245.990 ;
        RECT 345.550 245.610 356.290 245.620 ;
        RECT 342.960 245.390 344.650 245.590 ;
        RECT 341.750 245.190 342.030 245.200 ;
        RECT 341.010 244.740 342.030 245.190 ;
        RECT 342.960 244.740 343.190 245.390 ;
        RECT 344.370 245.330 344.650 245.390 ;
        RECT 345.530 245.380 356.290 245.610 ;
        RECT 345.550 245.370 356.290 245.380 ;
        RECT 362.420 245.980 362.680 247.180 ;
        RECT 362.420 245.470 362.670 245.980 ;
        RECT 364.310 245.970 364.570 247.180 ;
        RECT 366.700 246.070 366.950 247.620 ;
        RECT 364.310 245.810 364.700 245.970 ;
        RECT 364.300 245.680 364.700 245.810 ;
        RECT 367.400 245.680 367.660 247.290 ;
        RECT 369.950 246.220 370.250 247.270 ;
        RECT 370.700 246.670 371.000 247.620 ;
        RECT 371.200 246.720 371.500 246.770 ;
        RECT 371.200 246.370 372.100 246.720 ;
        RECT 384.860 246.320 389.330 246.350 ;
        RECT 373.920 246.290 389.330 246.320 ;
        RECT 373.250 246.270 389.330 246.290 ;
        RECT 362.920 245.470 363.210 245.630 ;
        RECT 364.300 245.620 364.560 245.680 ;
        RECT 345.550 245.360 356.250 245.370 ;
        RECT 345.550 245.320 345.830 245.360 ;
        RECT 362.420 245.280 363.210 245.470 ;
        RECT 362.420 245.080 362.670 245.280 ;
        RECT 362.920 245.170 363.210 245.280 ;
        RECT 364.310 245.080 364.560 245.620 ;
        RECT 367.390 245.620 367.660 245.680 ;
        RECT 368.940 245.960 370.250 246.220 ;
        RECT 368.940 245.620 369.250 245.960 ;
        RECT 364.950 245.090 366.590 245.480 ;
        RECT 367.390 245.330 369.250 245.620 ;
        RECT 367.390 245.320 367.700 245.330 ;
        RECT 368.940 245.320 369.250 245.330 ;
        RECT 344.350 244.760 344.620 244.840 ;
        RECT 341.750 244.530 343.190 244.740 ;
        RECT 343.740 244.540 344.620 244.760 ;
        RECT 341.750 243.480 342.030 244.530 ;
        RECT 343.740 243.730 343.960 244.540 ;
        RECT 344.350 244.510 344.620 244.540 ;
        RECT 345.480 244.800 345.770 244.850 ;
        RECT 345.480 244.620 356.230 244.800 ;
        RECT 345.480 244.520 345.770 244.620 ;
        RECT 350.320 244.610 353.950 244.620 ;
        RECT 356.030 243.940 356.230 244.620 ;
        RECT 362.420 244.480 362.710 245.080 ;
        RECT 364.310 244.480 364.600 245.080 ;
        RECT 341.030 243.030 342.030 243.480 ;
        RECT 341.010 241.580 342.310 242.030 ;
        RECT 342.010 241.180 342.310 241.580 ;
        RECT 343.730 241.200 343.960 243.730 ;
        RECT 350.980 243.640 356.230 243.940 ;
        RECT 366.650 243.870 366.950 244.870 ;
        RECT 367.400 244.270 367.700 245.320 ;
        RECT 370.000 244.220 370.250 245.960 ;
        RECT 372.370 245.950 389.330 246.270 ;
        RECT 373.250 245.940 389.330 245.950 ;
        RECT 373.250 245.910 385.230 245.940 ;
        RECT 373.250 245.900 374.140 245.910 ;
        RECT 370.700 243.870 370.960 245.420 ;
        RECT 371.790 243.870 371.990 243.880 ;
        RECT 342.800 241.180 343.960 241.200 ;
        RECT 342.010 241.000 343.960 241.180 ;
        RECT 346.900 242.000 347.160 243.200 ;
        RECT 346.900 241.490 347.150 242.000 ;
        RECT 348.790 241.990 349.050 243.200 ;
        RECT 351.180 242.090 351.430 243.640 ;
        RECT 348.790 241.830 349.180 241.990 ;
        RECT 348.780 241.700 349.180 241.830 ;
        RECT 351.880 241.700 352.140 243.310 ;
        RECT 354.430 242.240 354.730 243.290 ;
        RECT 355.180 242.690 355.480 243.640 ;
        RECT 356.030 243.630 356.230 243.640 ;
        RECT 366.600 243.570 371.990 243.870 ;
        RECT 355.680 242.740 355.980 242.790 ;
        RECT 355.680 242.390 356.580 242.740 ;
        RECT 371.790 242.330 371.990 243.570 ;
        RECT 388.950 242.370 389.310 245.940 ;
        RECT 463.370 242.920 463.620 255.340 ;
        RECT 364.230 242.310 365.420 242.320 ;
        RECT 366.410 242.310 367.600 242.320 ;
        RECT 368.630 242.310 369.820 242.320 ;
        RECT 370.810 242.310 372.000 242.330 ;
        RECT 362.020 242.300 372.000 242.310 ;
        RECT 358.630 242.280 359.820 242.290 ;
        RECT 360.910 242.280 372.000 242.300 ;
        RECT 347.400 241.490 347.690 241.650 ;
        RECT 348.780 241.640 349.040 241.700 ;
        RECT 346.900 241.300 347.690 241.490 ;
        RECT 346.900 241.100 347.150 241.300 ;
        RECT 347.400 241.190 347.690 241.300 ;
        RECT 348.790 241.100 349.040 241.640 ;
        RECT 351.870 241.640 352.140 241.700 ;
        RECT 353.420 241.980 354.730 242.240 ;
        RECT 356.790 242.050 372.000 242.280 ;
        RECT 384.080 242.070 389.330 242.370 ;
        RECT 356.790 242.040 370.950 242.050 ;
        RECT 356.790 242.030 364.320 242.040 ;
        RECT 365.330 242.030 366.520 242.040 ;
        RECT 367.480 242.030 368.670 242.040 ;
        RECT 369.760 242.030 370.950 242.040 ;
        RECT 356.790 242.020 362.100 242.030 ;
        RECT 356.790 242.010 360.960 242.020 ;
        RECT 356.790 242.000 358.680 242.010 ;
        RECT 359.770 242.000 360.960 242.010 ;
        RECT 356.790 241.990 357.510 242.000 ;
        RECT 353.420 241.640 353.730 241.980 ;
        RECT 349.430 241.110 351.070 241.500 ;
        RECT 351.870 241.350 353.730 241.640 ;
        RECT 351.870 241.340 352.180 241.350 ;
        RECT 353.420 241.340 353.730 241.350 ;
        RECT 342.010 240.990 342.660 241.000 ;
        RECT 342.010 240.660 342.310 240.990 ;
        RECT 341.290 240.210 342.310 240.660 ;
        RECT 346.900 240.500 347.190 241.100 ;
        RECT 348.790 240.500 349.080 241.100 ;
        RECT 342.010 240.200 342.310 240.210 ;
        RECT 351.130 239.890 351.430 240.890 ;
        RECT 351.880 240.290 352.180 241.340 ;
        RECT 354.480 240.240 354.730 241.980 ;
        RECT 355.180 239.890 355.440 241.440 ;
        RECT 380.000 240.430 380.260 241.630 ;
        RECT 380.000 239.920 380.250 240.430 ;
        RECT 381.890 240.420 382.150 241.630 ;
        RECT 384.280 240.520 384.530 242.070 ;
        RECT 381.890 240.260 382.280 240.420 ;
        RECT 381.880 240.130 382.280 240.260 ;
        RECT 384.980 240.130 385.240 241.740 ;
        RECT 387.530 240.670 387.830 241.720 ;
        RECT 388.280 241.120 388.580 242.070 ;
        RECT 388.780 241.170 389.080 241.220 ;
        RECT 388.780 240.820 389.680 241.170 ;
        RECT 380.500 239.920 380.790 240.080 ;
        RECT 381.880 240.070 382.140 240.130 ;
        RECT 351.080 239.880 356.330 239.890 ;
        RECT 340.960 239.800 341.210 239.810 ;
        RECT 340.960 239.340 341.940 239.800 ;
        RECT 351.080 239.590 356.350 239.880 ;
        RECT 340.960 239.040 341.210 239.340 ;
        RECT 348.930 239.250 350.770 239.260 ;
        RECT 356.180 239.250 356.350 239.590 ;
        RECT 342.670 239.240 342.910 239.250 ;
        RECT 343.750 239.240 356.350 239.250 ;
        RECT 342.670 239.080 356.350 239.240 ;
        RECT 380.000 239.730 380.790 239.920 ;
        RECT 380.000 239.530 380.250 239.730 ;
        RECT 380.500 239.620 380.790 239.730 ;
        RECT 381.890 239.530 382.140 240.070 ;
        RECT 384.970 240.070 385.240 240.130 ;
        RECT 386.520 240.410 387.830 240.670 ;
        RECT 389.890 240.710 391.560 240.740 ;
        RECT 406.640 240.710 406.890 240.720 ;
        RECT 389.890 240.440 406.890 240.710 ;
        RECT 389.890 240.430 403.390 240.440 ;
        RECT 391.170 240.410 403.390 240.430 ;
        RECT 386.520 240.070 386.830 240.410 ;
        RECT 382.530 239.540 384.170 239.930 ;
        RECT 384.970 239.780 386.830 240.070 ;
        RECT 384.970 239.770 385.280 239.780 ;
        RECT 386.520 239.770 386.830 239.780 ;
        RECT 342.670 239.070 354.180 239.080 ;
        RECT 342.660 239.060 348.980 239.070 ;
        RECT 350.530 239.060 354.180 239.070 ;
        RECT 342.660 239.050 344.530 239.060 ;
        RECT 342.660 239.040 342.910 239.050 ;
        RECT 340.960 238.870 342.910 239.040 ;
        RECT 380.000 238.930 380.290 239.530 ;
        RECT 381.890 238.930 382.180 239.530 ;
        RECT 340.960 238.650 341.210 238.870 ;
        RECT 340.960 238.480 342.000 238.650 ;
        RECT 341.810 237.620 342.000 238.480 ;
        RECT 384.230 238.320 384.530 239.320 ;
        RECT 384.980 238.720 385.280 239.770 ;
        RECT 387.580 238.670 387.830 240.410 ;
        RECT 388.280 238.320 388.540 239.870 ;
        RECT 389.160 238.320 389.500 238.390 ;
        RECT 384.180 238.020 389.500 238.320 ;
        RECT 341.020 237.180 342.000 237.620 ;
        RECT 341.020 237.170 341.970 237.180 ;
        RECT 342.840 236.860 352.110 236.870 ;
        RECT 353.990 236.860 355.910 236.870 ;
        RECT 340.690 236.760 340.880 236.770 ;
        RECT 340.690 236.300 341.670 236.760 ;
        RECT 342.840 236.670 355.910 236.860 ;
        RECT 342.840 236.660 355.200 236.670 ;
        RECT 340.690 235.510 340.880 236.300 ;
        RECT 342.840 235.650 343.050 236.660 ;
        RECT 352.100 236.650 354.000 236.660 ;
        RECT 355.730 235.920 355.910 236.670 ;
        RECT 341.690 235.510 341.960 235.520 ;
        RECT 340.690 235.300 341.960 235.510 ;
        RECT 341.690 235.090 341.960 235.300 ;
        RECT 341.690 234.460 341.940 235.090 ;
        RECT 342.840 234.640 343.040 235.650 ;
        RECT 350.650 235.620 355.910 235.920 ;
        RECT 340.900 234.010 341.940 234.460 ;
        RECT 340.880 232.560 341.840 233.010 ;
        RECT 341.590 232.510 341.840 232.560 ;
        RECT 342.850 232.510 343.040 234.640 ;
        RECT 341.590 232.310 343.040 232.510 ;
        RECT 346.570 233.980 346.830 235.180 ;
        RECT 346.570 233.470 346.820 233.980 ;
        RECT 348.460 233.970 348.720 235.180 ;
        RECT 350.850 234.070 351.100 235.620 ;
        RECT 348.460 233.810 348.850 233.970 ;
        RECT 348.450 233.680 348.850 233.810 ;
        RECT 351.550 233.680 351.810 235.290 ;
        RECT 354.100 234.220 354.400 235.270 ;
        RECT 354.850 234.670 355.150 235.620 ;
        RECT 355.350 234.720 355.650 234.770 ;
        RECT 355.350 234.370 356.250 234.720 ;
        RECT 357.960 234.590 358.180 234.600 ;
        RECT 357.960 234.400 371.640 234.590 ;
        RECT 357.960 234.270 358.180 234.400 ;
        RECT 347.070 233.470 347.360 233.630 ;
        RECT 348.450 233.620 348.710 233.680 ;
        RECT 346.570 233.280 347.360 233.470 ;
        RECT 346.570 233.080 346.820 233.280 ;
        RECT 347.070 233.170 347.360 233.280 ;
        RECT 348.460 233.080 348.710 233.620 ;
        RECT 351.540 233.620 351.810 233.680 ;
        RECT 353.090 233.960 354.400 234.220 ;
        RECT 356.500 233.970 358.180 234.270 ;
        RECT 356.500 233.960 358.160 233.970 ;
        RECT 353.090 233.620 353.400 233.960 ;
        RECT 349.100 233.090 350.740 233.480 ;
        RECT 351.540 233.330 353.400 233.620 ;
        RECT 351.540 233.320 351.850 233.330 ;
        RECT 353.090 233.320 353.400 233.330 ;
        RECT 346.570 232.480 346.860 233.080 ;
        RECT 348.460 232.480 348.750 233.080 ;
        RECT 341.590 232.220 341.840 232.310 ;
        RECT 340.860 231.770 341.840 232.220 ;
        RECT 350.800 231.870 351.100 232.870 ;
        RECT 351.550 232.270 351.850 233.320 ;
        RECT 354.150 232.220 354.400 233.960 ;
        RECT 371.390 233.500 371.640 234.400 ;
        RECT 354.850 231.870 355.110 233.420 ;
        RECT 366.330 233.200 371.640 233.500 ;
        RECT 350.750 231.850 356.000 231.870 ;
        RECT 350.750 231.570 356.120 231.850 ;
        RECT 344.200 231.170 344.480 231.240 ;
        RECT 345.380 231.200 345.660 231.230 ;
        RECT 355.830 231.200 356.120 231.570 ;
        RECT 345.380 231.190 356.120 231.200 ;
        RECT 342.790 230.970 344.480 231.170 ;
        RECT 341.580 230.770 341.860 230.780 ;
        RECT 340.840 230.320 341.860 230.770 ;
        RECT 342.790 230.320 343.020 230.970 ;
        RECT 344.200 230.910 344.480 230.970 ;
        RECT 345.360 230.960 356.120 231.190 ;
        RECT 345.380 230.950 356.120 230.960 ;
        RECT 362.250 231.560 362.510 232.760 ;
        RECT 362.250 231.050 362.500 231.560 ;
        RECT 364.140 231.550 364.400 232.760 ;
        RECT 366.530 231.650 366.780 233.200 ;
        RECT 364.140 231.390 364.530 231.550 ;
        RECT 364.130 231.260 364.530 231.390 ;
        RECT 367.230 231.260 367.490 232.870 ;
        RECT 369.780 231.800 370.080 232.850 ;
        RECT 370.530 232.250 370.830 233.200 ;
        RECT 371.030 232.300 371.330 232.350 ;
        RECT 371.030 231.950 371.930 232.300 ;
        RECT 389.160 231.900 389.500 238.020 ;
        RECT 388.590 231.880 389.550 231.900 ;
        RECT 373.070 231.860 377.350 231.870 ;
        RECT 384.750 231.860 389.550 231.880 ;
        RECT 373.070 231.850 389.550 231.860 ;
        RECT 362.750 231.050 363.040 231.210 ;
        RECT 364.130 231.200 364.390 231.260 ;
        RECT 345.380 230.940 356.080 230.950 ;
        RECT 345.380 230.900 345.660 230.940 ;
        RECT 362.250 230.860 363.040 231.050 ;
        RECT 362.250 230.660 362.500 230.860 ;
        RECT 362.750 230.750 363.040 230.860 ;
        RECT 364.140 230.660 364.390 231.200 ;
        RECT 367.220 231.200 367.490 231.260 ;
        RECT 368.770 231.540 370.080 231.800 ;
        RECT 368.770 231.200 369.080 231.540 ;
        RECT 364.780 230.670 366.420 231.060 ;
        RECT 367.220 230.910 369.080 231.200 ;
        RECT 367.220 230.900 367.530 230.910 ;
        RECT 368.770 230.900 369.080 230.910 ;
        RECT 344.180 230.340 344.450 230.420 ;
        RECT 341.580 230.110 343.020 230.320 ;
        RECT 343.570 230.120 344.450 230.340 ;
        RECT 341.580 229.060 341.860 230.110 ;
        RECT 343.570 229.310 343.790 230.120 ;
        RECT 344.180 230.090 344.450 230.120 ;
        RECT 345.310 230.380 345.600 230.430 ;
        RECT 345.310 230.200 356.060 230.380 ;
        RECT 345.310 230.100 345.600 230.200 ;
        RECT 350.150 230.190 353.780 230.200 ;
        RECT 355.860 229.520 356.060 230.200 ;
        RECT 362.250 230.060 362.540 230.660 ;
        RECT 364.140 230.060 364.430 230.660 ;
        RECT 340.860 228.610 341.860 229.060 ;
        RECT 340.840 227.160 342.140 227.610 ;
        RECT 341.840 226.760 342.140 227.160 ;
        RECT 343.560 226.780 343.790 229.310 ;
        RECT 350.810 229.220 356.060 229.520 ;
        RECT 366.480 229.450 366.780 230.450 ;
        RECT 367.230 229.850 367.530 230.900 ;
        RECT 369.830 229.800 370.080 231.540 ;
        RECT 372.200 231.540 389.550 231.850 ;
        RECT 372.200 231.530 385.210 231.540 ;
        RECT 377.060 231.520 385.210 231.530 ;
        RECT 388.590 231.500 389.550 231.540 ;
        RECT 389.160 231.490 389.500 231.500 ;
        RECT 370.530 229.450 370.790 231.000 ;
        RECT 371.620 229.450 371.820 229.460 ;
        RECT 342.630 226.760 343.790 226.780 ;
        RECT 341.840 226.580 343.790 226.760 ;
        RECT 346.730 227.580 346.990 228.780 ;
        RECT 346.730 227.070 346.980 227.580 ;
        RECT 348.620 227.570 348.880 228.780 ;
        RECT 351.010 227.670 351.260 229.220 ;
        RECT 348.620 227.410 349.010 227.570 ;
        RECT 348.610 227.280 349.010 227.410 ;
        RECT 351.710 227.280 351.970 228.890 ;
        RECT 354.260 227.820 354.560 228.870 ;
        RECT 355.010 228.270 355.310 229.220 ;
        RECT 355.860 229.210 356.060 229.220 ;
        RECT 366.430 229.150 371.820 229.450 ;
        RECT 355.510 228.320 355.810 228.370 ;
        RECT 355.510 227.970 356.410 228.320 ;
        RECT 371.620 227.910 371.820 229.150 ;
        RECT 364.060 227.890 365.250 227.900 ;
        RECT 366.240 227.890 367.430 227.900 ;
        RECT 368.460 227.890 369.650 227.900 ;
        RECT 370.640 227.890 371.830 227.910 ;
        RECT 361.850 227.880 371.830 227.890 ;
        RECT 358.460 227.860 359.650 227.870 ;
        RECT 360.740 227.860 371.830 227.880 ;
        RECT 347.230 227.070 347.520 227.230 ;
        RECT 348.610 227.220 348.870 227.280 ;
        RECT 346.730 226.880 347.520 227.070 ;
        RECT 346.730 226.680 346.980 226.880 ;
        RECT 347.230 226.770 347.520 226.880 ;
        RECT 348.620 226.680 348.870 227.220 ;
        RECT 351.700 227.220 351.970 227.280 ;
        RECT 353.250 227.560 354.560 227.820 ;
        RECT 356.620 227.630 371.830 227.860 ;
        RECT 356.620 227.620 370.780 227.630 ;
        RECT 356.620 227.610 364.150 227.620 ;
        RECT 365.160 227.610 366.350 227.620 ;
        RECT 367.310 227.610 368.500 227.620 ;
        RECT 369.590 227.610 370.780 227.620 ;
        RECT 356.620 227.600 361.930 227.610 ;
        RECT 356.620 227.590 360.790 227.600 ;
        RECT 356.620 227.580 358.510 227.590 ;
        RECT 359.600 227.580 360.790 227.590 ;
        RECT 356.620 227.570 357.340 227.580 ;
        RECT 353.250 227.220 353.560 227.560 ;
        RECT 349.260 226.690 350.900 227.080 ;
        RECT 351.700 226.930 353.560 227.220 ;
        RECT 351.700 226.920 352.010 226.930 ;
        RECT 353.250 226.920 353.560 226.930 ;
        RECT 341.840 226.570 342.490 226.580 ;
        RECT 341.840 226.240 342.140 226.570 ;
        RECT 341.120 225.790 342.140 226.240 ;
        RECT 346.730 226.080 347.020 226.680 ;
        RECT 348.620 226.080 348.910 226.680 ;
        RECT 341.840 225.780 342.140 225.790 ;
        RECT 350.960 225.470 351.260 226.470 ;
        RECT 351.710 225.870 352.010 226.920 ;
        RECT 354.310 225.820 354.560 227.560 ;
        RECT 406.640 227.300 406.900 240.440 ;
        RECT 406.630 227.180 406.900 227.300 ;
        RECT 355.010 225.470 355.270 227.020 ;
        RECT 406.630 226.350 406.890 227.180 ;
        RECT 401.610 226.050 406.890 226.350 ;
        RECT 350.910 225.460 356.160 225.470 ;
        RECT 340.790 225.380 341.040 225.390 ;
        RECT 340.790 224.920 341.770 225.380 ;
        RECT 350.910 225.170 356.180 225.460 ;
        RECT 340.790 224.620 341.040 224.920 ;
        RECT 348.760 224.830 350.600 224.840 ;
        RECT 356.010 224.830 356.180 225.170 ;
        RECT 342.500 224.820 342.740 224.830 ;
        RECT 343.580 224.820 356.180 224.830 ;
        RECT 342.500 224.660 356.180 224.820 ;
        RECT 342.500 224.650 354.010 224.660 ;
        RECT 342.490 224.640 348.810 224.650 ;
        RECT 350.360 224.640 354.010 224.650 ;
        RECT 342.490 224.630 344.360 224.640 ;
        RECT 342.490 224.620 342.740 224.630 ;
        RECT 340.790 224.450 342.740 224.620 ;
        RECT 340.790 224.150 341.060 224.450 ;
        RECT 340.800 223.890 341.060 224.150 ;
        RECT 397.530 224.410 397.790 225.610 ;
        RECT 397.530 223.900 397.780 224.410 ;
        RECT 399.420 224.400 399.680 225.610 ;
        RECT 401.810 224.500 402.060 226.050 ;
        RECT 399.420 224.240 399.810 224.400 ;
        RECT 399.410 224.110 399.810 224.240 ;
        RECT 402.510 224.110 402.770 225.720 ;
        RECT 405.060 224.650 405.360 225.700 ;
        RECT 405.810 225.100 406.110 226.050 ;
        RECT 406.310 225.150 406.610 225.200 ;
        RECT 406.310 224.800 407.210 225.150 ;
        RECT 398.030 223.900 398.320 224.060 ;
        RECT 399.410 224.050 399.670 224.110 ;
        RECT 340.780 223.500 341.080 223.890 ;
        RECT 397.530 223.710 398.320 223.900 ;
        RECT 397.530 223.510 397.780 223.710 ;
        RECT 398.030 223.600 398.320 223.710 ;
        RECT 399.420 223.510 399.670 224.050 ;
        RECT 402.500 224.050 402.770 224.110 ;
        RECT 404.050 224.390 405.360 224.650 ;
        RECT 407.480 224.590 408.260 224.690 ;
        RECT 407.480 224.420 421.060 224.590 ;
        RECT 407.480 224.410 421.050 224.420 ;
        RECT 407.480 224.390 408.260 224.410 ;
        RECT 404.050 224.050 404.360 224.390 ;
        RECT 400.060 223.520 401.700 223.910 ;
        RECT 402.500 223.760 404.360 224.050 ;
        RECT 402.500 223.750 402.810 223.760 ;
        RECT 404.050 223.750 404.360 223.760 ;
        RECT 340.780 223.270 342.270 223.500 ;
        RECT 342.020 222.340 342.270 223.270 ;
        RECT 397.530 222.910 397.820 223.510 ;
        RECT 399.420 222.910 399.710 223.510 ;
        RECT 341.220 221.880 342.270 222.340 ;
        RECT 401.760 222.300 402.060 223.300 ;
        RECT 402.510 222.700 402.810 223.750 ;
        RECT 405.110 222.650 405.360 224.390 ;
        RECT 405.810 222.300 406.070 223.850 ;
        RECT 401.710 222.000 406.980 222.300 ;
        RECT 342.020 221.870 342.270 221.880 ;
        RECT 340.890 221.470 341.140 221.480 ;
        RECT 340.890 221.020 341.870 221.470 ;
        RECT 342.980 221.210 352.250 221.220 ;
        RECT 354.130 221.210 356.050 221.220 ;
        RECT 342.980 221.020 356.050 221.210 ;
        RECT 340.890 220.410 341.140 221.020 ;
        RECT 342.980 221.010 355.340 221.020 ;
        RECT 340.890 220.160 342.100 220.410 ;
        RECT 341.830 219.410 342.090 220.160 ;
        RECT 342.980 220.000 343.190 221.010 ;
        RECT 352.240 221.000 354.140 221.010 ;
        RECT 355.870 220.270 356.050 221.020 ;
        RECT 341.830 218.810 342.080 219.410 ;
        RECT 342.980 218.990 343.180 220.000 ;
        RECT 350.790 219.970 356.050 220.270 ;
        RECT 341.040 218.360 342.080 218.810 ;
        RECT 341.020 216.910 341.980 217.360 ;
        RECT 341.730 216.860 341.980 216.910 ;
        RECT 342.990 216.860 343.180 218.990 ;
        RECT 341.730 216.660 343.180 216.860 ;
        RECT 346.710 218.330 346.970 219.530 ;
        RECT 346.710 217.820 346.960 218.330 ;
        RECT 348.600 218.320 348.860 219.530 ;
        RECT 350.990 218.420 351.240 219.970 ;
        RECT 348.600 218.160 348.990 218.320 ;
        RECT 348.590 218.030 348.990 218.160 ;
        RECT 351.690 218.030 351.950 219.640 ;
        RECT 354.240 218.570 354.540 219.620 ;
        RECT 354.990 219.020 355.290 219.970 ;
        RECT 355.490 219.070 355.790 219.120 ;
        RECT 355.490 218.720 356.390 219.070 ;
        RECT 358.100 218.940 358.320 218.950 ;
        RECT 358.100 218.750 371.780 218.940 ;
        RECT 358.100 218.620 358.320 218.750 ;
        RECT 347.210 217.820 347.500 217.980 ;
        RECT 348.590 217.970 348.850 218.030 ;
        RECT 346.710 217.630 347.500 217.820 ;
        RECT 346.710 217.430 346.960 217.630 ;
        RECT 347.210 217.520 347.500 217.630 ;
        RECT 348.600 217.430 348.850 217.970 ;
        RECT 351.680 217.970 351.950 218.030 ;
        RECT 353.230 218.310 354.540 218.570 ;
        RECT 356.640 218.320 358.320 218.620 ;
        RECT 356.640 218.310 358.300 218.320 ;
        RECT 353.230 217.970 353.540 218.310 ;
        RECT 349.240 217.440 350.880 217.830 ;
        RECT 351.680 217.680 353.540 217.970 ;
        RECT 351.680 217.670 351.990 217.680 ;
        RECT 353.230 217.670 353.540 217.680 ;
        RECT 346.710 216.830 347.000 217.430 ;
        RECT 348.600 216.830 348.890 217.430 ;
        RECT 341.730 216.570 341.980 216.660 ;
        RECT 341.000 216.120 341.980 216.570 ;
        RECT 350.940 216.220 351.240 217.220 ;
        RECT 351.690 216.620 351.990 217.670 ;
        RECT 354.290 216.570 354.540 218.310 ;
        RECT 371.530 217.850 371.780 218.750 ;
        RECT 354.990 216.220 355.250 217.770 ;
        RECT 366.470 217.550 371.780 217.850 ;
        RECT 350.890 216.200 356.140 216.220 ;
        RECT 350.890 215.920 356.260 216.200 ;
        RECT 344.340 215.520 344.620 215.590 ;
        RECT 345.520 215.550 345.800 215.580 ;
        RECT 355.970 215.550 356.260 215.920 ;
        RECT 345.520 215.540 356.260 215.550 ;
        RECT 342.930 215.320 344.620 215.520 ;
        RECT 341.720 215.120 342.000 215.130 ;
        RECT 340.980 214.670 342.000 215.120 ;
        RECT 342.930 214.670 343.160 215.320 ;
        RECT 344.340 215.260 344.620 215.320 ;
        RECT 345.500 215.310 356.260 215.540 ;
        RECT 345.520 215.300 356.260 215.310 ;
        RECT 362.390 215.910 362.650 217.110 ;
        RECT 362.390 215.400 362.640 215.910 ;
        RECT 364.280 215.900 364.540 217.110 ;
        RECT 366.670 216.000 366.920 217.550 ;
        RECT 364.280 215.740 364.670 215.900 ;
        RECT 364.270 215.610 364.670 215.740 ;
        RECT 367.370 215.610 367.630 217.220 ;
        RECT 369.920 216.150 370.220 217.200 ;
        RECT 370.670 216.600 370.970 217.550 ;
        RECT 371.170 216.650 371.470 216.700 ;
        RECT 371.170 216.300 372.070 216.650 ;
        RECT 384.830 216.250 389.300 216.280 ;
        RECT 373.890 216.220 389.300 216.250 ;
        RECT 373.220 216.200 389.300 216.220 ;
        RECT 362.890 215.400 363.180 215.560 ;
        RECT 364.270 215.550 364.530 215.610 ;
        RECT 345.520 215.290 356.220 215.300 ;
        RECT 345.520 215.250 345.800 215.290 ;
        RECT 362.390 215.210 363.180 215.400 ;
        RECT 362.390 215.010 362.640 215.210 ;
        RECT 362.890 215.100 363.180 215.210 ;
        RECT 364.280 215.010 364.530 215.550 ;
        RECT 367.360 215.550 367.630 215.610 ;
        RECT 368.910 215.890 370.220 216.150 ;
        RECT 368.910 215.550 369.220 215.890 ;
        RECT 364.920 215.020 366.560 215.410 ;
        RECT 367.360 215.260 369.220 215.550 ;
        RECT 367.360 215.250 367.670 215.260 ;
        RECT 368.910 215.250 369.220 215.260 ;
        RECT 344.320 214.690 344.590 214.770 ;
        RECT 341.720 214.460 343.160 214.670 ;
        RECT 343.710 214.470 344.590 214.690 ;
        RECT 341.720 213.410 342.000 214.460 ;
        RECT 343.710 213.660 343.930 214.470 ;
        RECT 344.320 214.440 344.590 214.470 ;
        RECT 345.450 214.730 345.740 214.780 ;
        RECT 345.450 214.550 356.200 214.730 ;
        RECT 345.450 214.450 345.740 214.550 ;
        RECT 350.290 214.540 353.920 214.550 ;
        RECT 356.000 213.870 356.200 214.550 ;
        RECT 362.390 214.410 362.680 215.010 ;
        RECT 364.280 214.410 364.570 215.010 ;
        RECT 341.000 212.960 342.000 213.410 ;
        RECT 340.980 211.510 342.280 211.960 ;
        RECT 341.980 211.110 342.280 211.510 ;
        RECT 343.700 211.130 343.930 213.660 ;
        RECT 350.950 213.570 356.200 213.870 ;
        RECT 366.620 213.800 366.920 214.800 ;
        RECT 367.370 214.200 367.670 215.250 ;
        RECT 369.970 214.150 370.220 215.890 ;
        RECT 372.340 215.880 389.300 216.200 ;
        RECT 373.220 215.870 389.300 215.880 ;
        RECT 373.220 215.840 385.200 215.870 ;
        RECT 373.220 215.830 374.110 215.840 ;
        RECT 370.670 213.800 370.930 215.350 ;
        RECT 371.760 213.800 371.960 213.810 ;
        RECT 342.770 211.110 343.930 211.130 ;
        RECT 341.980 210.930 343.930 211.110 ;
        RECT 346.870 211.930 347.130 213.130 ;
        RECT 346.870 211.420 347.120 211.930 ;
        RECT 348.760 211.920 349.020 213.130 ;
        RECT 351.150 212.020 351.400 213.570 ;
        RECT 348.760 211.760 349.150 211.920 ;
        RECT 348.750 211.630 349.150 211.760 ;
        RECT 351.850 211.630 352.110 213.240 ;
        RECT 354.400 212.170 354.700 213.220 ;
        RECT 355.150 212.620 355.450 213.570 ;
        RECT 356.000 213.560 356.200 213.570 ;
        RECT 366.570 213.500 371.960 213.800 ;
        RECT 355.650 212.670 355.950 212.720 ;
        RECT 355.650 212.320 356.550 212.670 ;
        RECT 371.760 212.260 371.960 213.500 ;
        RECT 388.920 212.300 389.280 215.870 ;
        RECT 364.200 212.240 365.390 212.250 ;
        RECT 366.380 212.240 367.570 212.250 ;
        RECT 368.600 212.240 369.790 212.250 ;
        RECT 370.780 212.240 371.970 212.260 ;
        RECT 361.990 212.230 371.970 212.240 ;
        RECT 358.600 212.210 359.790 212.220 ;
        RECT 360.880 212.210 371.970 212.230 ;
        RECT 347.370 211.420 347.660 211.580 ;
        RECT 348.750 211.570 349.010 211.630 ;
        RECT 346.870 211.230 347.660 211.420 ;
        RECT 346.870 211.030 347.120 211.230 ;
        RECT 347.370 211.120 347.660 211.230 ;
        RECT 348.760 211.030 349.010 211.570 ;
        RECT 351.840 211.570 352.110 211.630 ;
        RECT 353.390 211.910 354.700 212.170 ;
        RECT 356.760 211.980 371.970 212.210 ;
        RECT 384.050 212.000 389.300 212.300 ;
        RECT 356.760 211.970 370.920 211.980 ;
        RECT 356.760 211.960 364.290 211.970 ;
        RECT 365.300 211.960 366.490 211.970 ;
        RECT 367.450 211.960 368.640 211.970 ;
        RECT 369.730 211.960 370.920 211.970 ;
        RECT 356.760 211.950 362.070 211.960 ;
        RECT 356.760 211.940 360.930 211.950 ;
        RECT 356.760 211.930 358.650 211.940 ;
        RECT 359.740 211.930 360.930 211.940 ;
        RECT 356.760 211.920 357.480 211.930 ;
        RECT 353.390 211.570 353.700 211.910 ;
        RECT 349.400 211.040 351.040 211.430 ;
        RECT 351.840 211.280 353.700 211.570 ;
        RECT 351.840 211.270 352.150 211.280 ;
        RECT 353.390 211.270 353.700 211.280 ;
        RECT 341.980 210.920 342.630 210.930 ;
        RECT 341.980 210.590 342.280 210.920 ;
        RECT 341.260 210.140 342.280 210.590 ;
        RECT 346.870 210.430 347.160 211.030 ;
        RECT 348.760 210.430 349.050 211.030 ;
        RECT 341.980 210.130 342.280 210.140 ;
        RECT 351.100 209.820 351.400 210.820 ;
        RECT 351.850 210.220 352.150 211.270 ;
        RECT 354.450 210.170 354.700 211.910 ;
        RECT 355.150 209.820 355.410 211.370 ;
        RECT 379.970 210.360 380.230 211.560 ;
        RECT 379.970 209.850 380.220 210.360 ;
        RECT 381.860 210.350 382.120 211.560 ;
        RECT 384.250 210.450 384.500 212.000 ;
        RECT 381.860 210.190 382.250 210.350 ;
        RECT 381.850 210.060 382.250 210.190 ;
        RECT 384.950 210.060 385.210 211.670 ;
        RECT 387.500 210.600 387.800 211.650 ;
        RECT 388.250 211.050 388.550 212.000 ;
        RECT 388.750 211.100 389.050 211.150 ;
        RECT 388.750 210.750 389.650 211.100 ;
        RECT 380.470 209.850 380.760 210.010 ;
        RECT 381.850 210.000 382.110 210.060 ;
        RECT 351.050 209.810 356.300 209.820 ;
        RECT 340.930 209.730 341.180 209.740 ;
        RECT 340.930 209.270 341.910 209.730 ;
        RECT 351.050 209.520 356.320 209.810 ;
        RECT 340.930 208.970 341.180 209.270 ;
        RECT 348.900 209.180 350.740 209.190 ;
        RECT 356.150 209.180 356.320 209.520 ;
        RECT 342.640 209.170 342.880 209.180 ;
        RECT 343.720 209.170 356.320 209.180 ;
        RECT 342.640 209.010 356.320 209.170 ;
        RECT 379.970 209.660 380.760 209.850 ;
        RECT 379.970 209.460 380.220 209.660 ;
        RECT 380.470 209.550 380.760 209.660 ;
        RECT 381.860 209.460 382.110 210.000 ;
        RECT 384.940 210.000 385.210 210.060 ;
        RECT 386.490 210.340 387.800 210.600 ;
        RECT 389.860 210.650 391.530 210.670 ;
        RECT 406.670 210.650 406.980 222.000 ;
        RECT 389.860 210.360 407.020 210.650 ;
        RECT 390.550 210.350 407.020 210.360 ;
        RECT 386.490 210.000 386.800 210.340 ;
        RECT 382.500 209.470 384.140 209.860 ;
        RECT 384.940 209.710 386.800 210.000 ;
        RECT 384.940 209.700 385.250 209.710 ;
        RECT 386.490 209.700 386.800 209.710 ;
        RECT 342.640 209.000 354.150 209.010 ;
        RECT 342.630 208.990 348.950 209.000 ;
        RECT 350.500 208.990 354.150 209.000 ;
        RECT 342.630 208.980 344.500 208.990 ;
        RECT 342.630 208.970 342.880 208.980 ;
        RECT 340.930 208.800 342.880 208.970 ;
        RECT 379.970 208.860 380.260 209.460 ;
        RECT 381.860 208.860 382.150 209.460 ;
        RECT 340.930 208.580 341.180 208.800 ;
        RECT 340.930 208.410 341.970 208.580 ;
        RECT 341.780 207.550 341.970 208.410 ;
        RECT 384.200 208.250 384.500 209.250 ;
        RECT 384.950 208.650 385.250 209.700 ;
        RECT 387.550 208.600 387.800 210.340 ;
        RECT 388.250 208.250 388.510 209.800 ;
        RECT 389.130 208.250 389.470 208.320 ;
        RECT 384.150 207.950 389.470 208.250 ;
        RECT 340.990 207.110 341.970 207.550 ;
        RECT 340.990 207.100 341.940 207.110 ;
        RECT 342.810 206.790 352.080 206.800 ;
        RECT 353.960 206.790 355.880 206.800 ;
        RECT 340.660 206.690 340.850 206.700 ;
        RECT 340.660 206.230 341.640 206.690 ;
        RECT 342.810 206.600 355.880 206.790 ;
        RECT 342.810 206.590 355.170 206.600 ;
        RECT 340.660 205.440 340.850 206.230 ;
        RECT 342.810 205.580 343.020 206.590 ;
        RECT 352.070 206.580 353.970 206.590 ;
        RECT 355.700 205.850 355.880 206.600 ;
        RECT 341.660 205.440 341.930 205.450 ;
        RECT 340.660 205.230 341.930 205.440 ;
        RECT 341.660 205.020 341.930 205.230 ;
        RECT 341.660 204.390 341.910 205.020 ;
        RECT 342.810 204.570 343.010 205.580 ;
        RECT 350.620 205.550 355.880 205.850 ;
        RECT 340.870 203.940 341.910 204.390 ;
        RECT 340.850 202.490 341.810 202.940 ;
        RECT 341.560 202.440 341.810 202.490 ;
        RECT 342.820 202.440 343.010 204.570 ;
        RECT 341.560 202.240 343.010 202.440 ;
        RECT 346.540 203.910 346.800 205.110 ;
        RECT 346.540 203.400 346.790 203.910 ;
        RECT 348.430 203.900 348.690 205.110 ;
        RECT 350.820 204.000 351.070 205.550 ;
        RECT 348.430 203.740 348.820 203.900 ;
        RECT 348.420 203.610 348.820 203.740 ;
        RECT 351.520 203.610 351.780 205.220 ;
        RECT 354.070 204.150 354.370 205.200 ;
        RECT 354.820 204.600 355.120 205.550 ;
        RECT 355.320 204.650 355.620 204.700 ;
        RECT 355.320 204.300 356.220 204.650 ;
        RECT 357.930 204.520 358.150 204.530 ;
        RECT 357.930 204.330 371.610 204.520 ;
        RECT 357.930 204.200 358.150 204.330 ;
        RECT 347.040 203.400 347.330 203.560 ;
        RECT 348.420 203.550 348.680 203.610 ;
        RECT 346.540 203.210 347.330 203.400 ;
        RECT 346.540 203.010 346.790 203.210 ;
        RECT 347.040 203.100 347.330 203.210 ;
        RECT 348.430 203.010 348.680 203.550 ;
        RECT 351.510 203.550 351.780 203.610 ;
        RECT 353.060 203.890 354.370 204.150 ;
        RECT 356.470 203.900 358.150 204.200 ;
        RECT 356.470 203.890 358.130 203.900 ;
        RECT 353.060 203.550 353.370 203.890 ;
        RECT 349.070 203.020 350.710 203.410 ;
        RECT 351.510 203.260 353.370 203.550 ;
        RECT 351.510 203.250 351.820 203.260 ;
        RECT 353.060 203.250 353.370 203.260 ;
        RECT 346.540 202.410 346.830 203.010 ;
        RECT 348.430 202.410 348.720 203.010 ;
        RECT 341.560 202.150 341.810 202.240 ;
        RECT 340.830 201.700 341.810 202.150 ;
        RECT 350.770 201.800 351.070 202.800 ;
        RECT 351.520 202.200 351.820 203.250 ;
        RECT 354.120 202.150 354.370 203.890 ;
        RECT 371.360 203.430 371.610 204.330 ;
        RECT 354.820 201.800 355.080 203.350 ;
        RECT 366.300 203.130 371.610 203.430 ;
        RECT 350.720 201.780 355.970 201.800 ;
        RECT 350.720 201.500 356.090 201.780 ;
        RECT 344.170 201.100 344.450 201.170 ;
        RECT 345.350 201.130 345.630 201.160 ;
        RECT 355.800 201.130 356.090 201.500 ;
        RECT 345.350 201.120 356.090 201.130 ;
        RECT 342.760 200.900 344.450 201.100 ;
        RECT 341.550 200.700 341.830 200.710 ;
        RECT 340.810 200.250 341.830 200.700 ;
        RECT 342.760 200.250 342.990 200.900 ;
        RECT 344.170 200.840 344.450 200.900 ;
        RECT 345.330 200.890 356.090 201.120 ;
        RECT 345.350 200.880 356.090 200.890 ;
        RECT 362.220 201.490 362.480 202.690 ;
        RECT 362.220 200.980 362.470 201.490 ;
        RECT 364.110 201.480 364.370 202.690 ;
        RECT 366.500 201.580 366.750 203.130 ;
        RECT 364.110 201.320 364.500 201.480 ;
        RECT 364.100 201.190 364.500 201.320 ;
        RECT 367.200 201.190 367.460 202.800 ;
        RECT 369.750 201.730 370.050 202.780 ;
        RECT 370.500 202.180 370.800 203.130 ;
        RECT 371.000 202.230 371.300 202.280 ;
        RECT 371.000 201.880 371.900 202.230 ;
        RECT 389.130 201.830 389.470 207.950 ;
        RECT 420.870 205.150 421.050 224.410 ;
        RECT 420.850 204.100 421.060 205.150 ;
        RECT 420.850 204.020 421.070 204.100 ;
        RECT 420.860 201.950 421.070 204.020 ;
        RECT 420.850 201.910 421.070 201.950 ;
        RECT 388.560 201.810 389.520 201.830 ;
        RECT 373.040 201.790 377.320 201.800 ;
        RECT 384.720 201.790 389.520 201.810 ;
        RECT 373.040 201.780 389.520 201.790 ;
        RECT 362.720 200.980 363.010 201.140 ;
        RECT 364.100 201.130 364.360 201.190 ;
        RECT 345.350 200.870 356.050 200.880 ;
        RECT 345.350 200.830 345.630 200.870 ;
        RECT 362.220 200.790 363.010 200.980 ;
        RECT 362.220 200.590 362.470 200.790 ;
        RECT 362.720 200.680 363.010 200.790 ;
        RECT 364.110 200.590 364.360 201.130 ;
        RECT 367.190 201.130 367.460 201.190 ;
        RECT 368.740 201.470 370.050 201.730 ;
        RECT 368.740 201.130 369.050 201.470 ;
        RECT 364.750 200.600 366.390 200.990 ;
        RECT 367.190 200.840 369.050 201.130 ;
        RECT 367.190 200.830 367.500 200.840 ;
        RECT 368.740 200.830 369.050 200.840 ;
        RECT 344.150 200.270 344.420 200.350 ;
        RECT 341.550 200.040 342.990 200.250 ;
        RECT 343.540 200.050 344.420 200.270 ;
        RECT 341.550 198.990 341.830 200.040 ;
        RECT 343.540 199.240 343.760 200.050 ;
        RECT 344.150 200.020 344.420 200.050 ;
        RECT 345.280 200.310 345.570 200.360 ;
        RECT 345.280 200.130 356.030 200.310 ;
        RECT 345.280 200.030 345.570 200.130 ;
        RECT 350.120 200.120 353.750 200.130 ;
        RECT 355.830 199.450 356.030 200.130 ;
        RECT 362.220 199.990 362.510 200.590 ;
        RECT 364.110 199.990 364.400 200.590 ;
        RECT 340.830 198.540 341.830 198.990 ;
        RECT 340.810 197.090 342.110 197.540 ;
        RECT 341.810 196.690 342.110 197.090 ;
        RECT 343.530 196.710 343.760 199.240 ;
        RECT 350.780 199.150 356.030 199.450 ;
        RECT 366.450 199.380 366.750 200.380 ;
        RECT 367.200 199.780 367.500 200.830 ;
        RECT 369.800 199.730 370.050 201.470 ;
        RECT 372.170 201.470 389.520 201.780 ;
        RECT 372.170 201.460 385.180 201.470 ;
        RECT 377.030 201.450 385.180 201.460 ;
        RECT 388.560 201.430 389.520 201.470 ;
        RECT 389.130 201.420 389.470 201.430 ;
        RECT 370.500 199.380 370.760 200.930 ;
        RECT 420.850 200.060 421.060 201.910 ;
        RECT 415.810 199.760 421.060 200.060 ;
        RECT 371.590 199.380 371.790 199.390 ;
        RECT 342.600 196.690 343.760 196.710 ;
        RECT 341.810 196.510 343.760 196.690 ;
        RECT 346.700 197.510 346.960 198.710 ;
        RECT 346.700 197.000 346.950 197.510 ;
        RECT 348.590 197.500 348.850 198.710 ;
        RECT 350.980 197.600 351.230 199.150 ;
        RECT 348.590 197.340 348.980 197.500 ;
        RECT 348.580 197.210 348.980 197.340 ;
        RECT 351.680 197.210 351.940 198.820 ;
        RECT 354.230 197.750 354.530 198.800 ;
        RECT 354.980 198.200 355.280 199.150 ;
        RECT 355.830 199.140 356.030 199.150 ;
        RECT 366.400 199.080 371.790 199.380 ;
        RECT 355.480 198.250 355.780 198.300 ;
        RECT 355.480 197.900 356.380 198.250 ;
        RECT 371.590 197.840 371.790 199.080 ;
        RECT 411.730 198.120 411.990 199.320 ;
        RECT 364.030 197.820 365.220 197.830 ;
        RECT 366.210 197.820 367.400 197.830 ;
        RECT 368.430 197.820 369.620 197.830 ;
        RECT 370.610 197.820 371.800 197.840 ;
        RECT 361.820 197.810 371.800 197.820 ;
        RECT 358.430 197.790 359.620 197.800 ;
        RECT 360.710 197.790 371.800 197.810 ;
        RECT 347.200 197.000 347.490 197.160 ;
        RECT 348.580 197.150 348.840 197.210 ;
        RECT 346.700 196.810 347.490 197.000 ;
        RECT 346.700 196.610 346.950 196.810 ;
        RECT 347.200 196.700 347.490 196.810 ;
        RECT 348.590 196.610 348.840 197.150 ;
        RECT 351.670 197.150 351.940 197.210 ;
        RECT 353.220 197.490 354.530 197.750 ;
        RECT 356.590 197.560 371.800 197.790 ;
        RECT 411.730 197.610 411.980 198.120 ;
        RECT 413.620 198.110 413.880 199.320 ;
        RECT 416.010 198.210 416.260 199.760 ;
        RECT 413.620 197.950 414.010 198.110 ;
        RECT 413.610 197.820 414.010 197.950 ;
        RECT 416.710 197.820 416.970 199.430 ;
        RECT 419.260 198.360 419.560 199.410 ;
        RECT 420.010 198.810 420.310 199.760 ;
        RECT 420.850 199.750 421.060 199.760 ;
        RECT 420.510 198.860 420.810 198.910 ;
        RECT 420.510 198.510 421.410 198.860 ;
        RECT 422.370 198.390 437.360 198.460 ;
        RECT 412.230 197.610 412.520 197.770 ;
        RECT 413.610 197.760 413.870 197.820 ;
        RECT 356.590 197.550 370.750 197.560 ;
        RECT 356.590 197.540 364.120 197.550 ;
        RECT 365.130 197.540 366.320 197.550 ;
        RECT 367.280 197.540 368.470 197.550 ;
        RECT 369.560 197.540 370.750 197.550 ;
        RECT 356.590 197.530 361.900 197.540 ;
        RECT 356.590 197.520 360.760 197.530 ;
        RECT 356.590 197.510 358.480 197.520 ;
        RECT 359.570 197.510 360.760 197.520 ;
        RECT 356.590 197.500 357.310 197.510 ;
        RECT 353.220 197.150 353.530 197.490 ;
        RECT 349.230 196.620 350.870 197.010 ;
        RECT 351.670 196.860 353.530 197.150 ;
        RECT 351.670 196.850 351.980 196.860 ;
        RECT 353.220 196.850 353.530 196.860 ;
        RECT 341.810 196.500 342.460 196.510 ;
        RECT 341.810 196.170 342.110 196.500 ;
        RECT 341.090 195.720 342.110 196.170 ;
        RECT 346.700 196.010 346.990 196.610 ;
        RECT 348.590 196.010 348.880 196.610 ;
        RECT 341.810 195.710 342.110 195.720 ;
        RECT 350.930 195.400 351.230 196.400 ;
        RECT 351.680 195.800 351.980 196.850 ;
        RECT 354.280 195.750 354.530 197.490 ;
        RECT 411.730 197.420 412.520 197.610 ;
        RECT 411.730 197.220 411.980 197.420 ;
        RECT 412.230 197.310 412.520 197.420 ;
        RECT 413.620 197.220 413.870 197.760 ;
        RECT 416.700 197.760 416.970 197.820 ;
        RECT 418.250 198.100 419.560 198.360 ;
        RECT 421.700 198.140 437.360 198.390 ;
        RECT 421.700 198.110 422.520 198.140 ;
        RECT 418.250 197.760 418.560 198.100 ;
        RECT 414.260 197.230 415.900 197.620 ;
        RECT 416.700 197.470 418.560 197.760 ;
        RECT 416.700 197.460 417.010 197.470 ;
        RECT 418.250 197.460 418.560 197.470 ;
        RECT 354.980 195.400 355.240 196.950 ;
        RECT 411.730 196.620 412.020 197.220 ;
        RECT 413.620 196.620 413.910 197.220 ;
        RECT 415.960 196.010 416.260 197.010 ;
        RECT 416.710 196.410 417.010 197.460 ;
        RECT 419.310 196.360 419.560 198.100 ;
        RECT 437.110 197.930 437.360 198.140 ;
        RECT 420.010 196.010 420.270 197.560 ;
        RECT 437.110 196.090 437.380 197.930 ;
        RECT 420.970 196.010 421.150 196.020 ;
        RECT 415.910 195.710 421.160 196.010 ;
        RECT 350.880 195.390 356.130 195.400 ;
        RECT 340.760 195.310 341.010 195.320 ;
        RECT 340.760 194.850 341.740 195.310 ;
        RECT 350.880 195.100 356.150 195.390 ;
        RECT 340.760 194.550 341.010 194.850 ;
        RECT 348.730 194.760 350.570 194.770 ;
        RECT 355.980 194.760 356.150 195.100 ;
        RECT 342.470 194.750 342.710 194.760 ;
        RECT 343.550 194.750 356.150 194.760 ;
        RECT 342.470 194.590 356.150 194.750 ;
        RECT 342.470 194.580 353.980 194.590 ;
        RECT 342.460 194.570 348.780 194.580 ;
        RECT 350.330 194.570 353.980 194.580 ;
        RECT 342.460 194.560 344.330 194.570 ;
        RECT 342.460 194.550 342.710 194.560 ;
        RECT 340.760 194.380 342.710 194.550 ;
        RECT 340.760 194.080 341.030 194.380 ;
        RECT 340.770 193.820 341.030 194.080 ;
        RECT 340.750 193.430 341.050 193.820 ;
        RECT 340.740 193.030 341.050 193.430 ;
        RECT 340.730 192.270 341.040 193.030 ;
        RECT 340.630 192.250 341.040 192.270 ;
        RECT 340.600 191.300 341.050 192.250 ;
        RECT 341.460 191.010 341.920 191.950 ;
        RECT 342.660 191.360 351.930 191.370 ;
        RECT 353.810 191.360 355.730 191.370 ;
        RECT 342.660 191.170 355.730 191.360 ;
        RECT 342.660 191.160 355.020 191.170 ;
        RECT 341.500 190.690 341.800 191.010 ;
        RECT 341.500 190.360 341.790 190.690 ;
        RECT 341.510 189.560 341.770 190.360 ;
        RECT 342.660 190.150 342.870 191.160 ;
        RECT 351.920 191.150 353.820 191.160 ;
        RECT 355.550 190.420 355.730 191.170 ;
        RECT 341.510 188.960 341.760 189.560 ;
        RECT 342.660 189.140 342.860 190.150 ;
        RECT 350.470 190.120 355.730 190.420 ;
        RECT 340.720 188.510 341.760 188.960 ;
        RECT 340.700 187.060 341.660 187.510 ;
        RECT 341.410 187.010 341.660 187.060 ;
        RECT 342.670 187.010 342.860 189.140 ;
        RECT 341.410 186.810 342.860 187.010 ;
        RECT 346.390 188.480 346.650 189.680 ;
        RECT 346.390 187.970 346.640 188.480 ;
        RECT 348.280 188.470 348.540 189.680 ;
        RECT 350.670 188.570 350.920 190.120 ;
        RECT 348.280 188.310 348.670 188.470 ;
        RECT 348.270 188.180 348.670 188.310 ;
        RECT 351.370 188.180 351.630 189.790 ;
        RECT 353.920 188.720 354.220 189.770 ;
        RECT 354.670 189.170 354.970 190.120 ;
        RECT 355.170 189.220 355.470 189.270 ;
        RECT 355.170 188.870 356.070 189.220 ;
        RECT 357.780 189.090 358.000 189.100 ;
        RECT 357.780 188.900 371.460 189.090 ;
        RECT 357.780 188.770 358.000 188.900 ;
        RECT 346.890 187.970 347.180 188.130 ;
        RECT 348.270 188.120 348.530 188.180 ;
        RECT 346.390 187.780 347.180 187.970 ;
        RECT 346.390 187.580 346.640 187.780 ;
        RECT 346.890 187.670 347.180 187.780 ;
        RECT 348.280 187.580 348.530 188.120 ;
        RECT 351.360 188.120 351.630 188.180 ;
        RECT 352.910 188.460 354.220 188.720 ;
        RECT 356.320 188.470 358.000 188.770 ;
        RECT 356.320 188.460 357.980 188.470 ;
        RECT 352.910 188.120 353.220 188.460 ;
        RECT 348.920 187.590 350.560 187.980 ;
        RECT 351.360 187.830 353.220 188.120 ;
        RECT 351.360 187.820 351.670 187.830 ;
        RECT 352.910 187.820 353.220 187.830 ;
        RECT 346.390 186.980 346.680 187.580 ;
        RECT 348.280 186.980 348.570 187.580 ;
        RECT 341.410 186.720 341.660 186.810 ;
        RECT 340.680 186.270 341.660 186.720 ;
        RECT 350.620 186.370 350.920 187.370 ;
        RECT 351.370 186.770 351.670 187.820 ;
        RECT 353.970 186.720 354.220 188.460 ;
        RECT 371.210 188.000 371.460 188.900 ;
        RECT 354.670 186.370 354.930 187.920 ;
        RECT 366.150 187.700 371.460 188.000 ;
        RECT 350.570 186.350 355.820 186.370 ;
        RECT 350.570 186.070 355.940 186.350 ;
        RECT 344.020 185.670 344.300 185.740 ;
        RECT 345.200 185.700 345.480 185.730 ;
        RECT 355.650 185.700 355.940 186.070 ;
        RECT 345.200 185.690 355.940 185.700 ;
        RECT 342.610 185.470 344.300 185.670 ;
        RECT 341.400 185.270 341.680 185.280 ;
        RECT 340.660 184.820 341.680 185.270 ;
        RECT 342.610 184.820 342.840 185.470 ;
        RECT 344.020 185.410 344.300 185.470 ;
        RECT 345.180 185.460 355.940 185.690 ;
        RECT 345.200 185.450 355.940 185.460 ;
        RECT 362.070 186.060 362.330 187.260 ;
        RECT 362.070 185.550 362.320 186.060 ;
        RECT 363.960 186.050 364.220 187.260 ;
        RECT 366.350 186.150 366.600 187.700 ;
        RECT 363.960 185.890 364.350 186.050 ;
        RECT 363.950 185.760 364.350 185.890 ;
        RECT 367.050 185.760 367.310 187.370 ;
        RECT 369.600 186.300 369.900 187.350 ;
        RECT 370.350 186.750 370.650 187.700 ;
        RECT 370.850 186.800 371.150 186.850 ;
        RECT 370.850 186.450 371.750 186.800 ;
        RECT 384.510 186.400 388.980 186.430 ;
        RECT 373.570 186.370 388.980 186.400 ;
        RECT 372.900 186.350 388.980 186.370 ;
        RECT 362.570 185.550 362.860 185.710 ;
        RECT 363.950 185.700 364.210 185.760 ;
        RECT 345.200 185.440 355.900 185.450 ;
        RECT 345.200 185.400 345.480 185.440 ;
        RECT 362.070 185.360 362.860 185.550 ;
        RECT 362.070 185.160 362.320 185.360 ;
        RECT 362.570 185.250 362.860 185.360 ;
        RECT 363.960 185.160 364.210 185.700 ;
        RECT 367.040 185.700 367.310 185.760 ;
        RECT 368.590 186.040 369.900 186.300 ;
        RECT 368.590 185.700 368.900 186.040 ;
        RECT 364.600 185.170 366.240 185.560 ;
        RECT 367.040 185.410 368.900 185.700 ;
        RECT 367.040 185.400 367.350 185.410 ;
        RECT 368.590 185.400 368.900 185.410 ;
        RECT 344.000 184.840 344.270 184.920 ;
        RECT 341.400 184.610 342.840 184.820 ;
        RECT 343.390 184.620 344.270 184.840 ;
        RECT 341.400 183.560 341.680 184.610 ;
        RECT 343.390 183.810 343.610 184.620 ;
        RECT 344.000 184.590 344.270 184.620 ;
        RECT 345.130 184.880 345.420 184.930 ;
        RECT 345.130 184.700 355.880 184.880 ;
        RECT 345.130 184.600 345.420 184.700 ;
        RECT 349.970 184.690 353.600 184.700 ;
        RECT 355.680 184.020 355.880 184.700 ;
        RECT 362.070 184.560 362.360 185.160 ;
        RECT 363.960 184.560 364.250 185.160 ;
        RECT 340.680 183.110 341.680 183.560 ;
        RECT 340.660 181.660 341.960 182.110 ;
        RECT 341.660 181.260 341.960 181.660 ;
        RECT 343.380 181.280 343.610 183.810 ;
        RECT 350.630 183.720 355.880 184.020 ;
        RECT 366.300 183.950 366.600 184.950 ;
        RECT 367.050 184.350 367.350 185.400 ;
        RECT 369.650 184.300 369.900 186.040 ;
        RECT 372.020 186.030 388.980 186.350 ;
        RECT 420.970 186.050 421.150 195.710 ;
        RECT 372.900 186.020 388.980 186.030 ;
        RECT 372.900 185.990 384.880 186.020 ;
        RECT 372.900 185.980 373.790 185.990 ;
        RECT 370.350 183.950 370.610 185.500 ;
        RECT 371.440 183.950 371.640 183.960 ;
        RECT 342.450 181.260 343.610 181.280 ;
        RECT 341.660 181.080 343.610 181.260 ;
        RECT 346.550 182.080 346.810 183.280 ;
        RECT 346.550 181.570 346.800 182.080 ;
        RECT 348.440 182.070 348.700 183.280 ;
        RECT 350.830 182.170 351.080 183.720 ;
        RECT 348.440 181.910 348.830 182.070 ;
        RECT 348.430 181.780 348.830 181.910 ;
        RECT 351.530 181.780 351.790 183.390 ;
        RECT 354.080 182.320 354.380 183.370 ;
        RECT 354.830 182.770 355.130 183.720 ;
        RECT 355.680 183.710 355.880 183.720 ;
        RECT 366.250 183.650 371.640 183.950 ;
        RECT 355.330 182.820 355.630 182.870 ;
        RECT 355.330 182.470 356.230 182.820 ;
        RECT 371.440 182.410 371.640 183.650 ;
        RECT 388.600 182.450 388.960 186.020 ;
        RECT 363.880 182.390 365.070 182.400 ;
        RECT 366.060 182.390 367.250 182.400 ;
        RECT 368.280 182.390 369.470 182.400 ;
        RECT 370.460 182.390 371.650 182.410 ;
        RECT 361.670 182.380 371.650 182.390 ;
        RECT 358.280 182.360 359.470 182.370 ;
        RECT 360.560 182.360 371.650 182.380 ;
        RECT 347.050 181.570 347.340 181.730 ;
        RECT 348.430 181.720 348.690 181.780 ;
        RECT 346.550 181.380 347.340 181.570 ;
        RECT 346.550 181.180 346.800 181.380 ;
        RECT 347.050 181.270 347.340 181.380 ;
        RECT 348.440 181.180 348.690 181.720 ;
        RECT 351.520 181.720 351.790 181.780 ;
        RECT 353.070 182.060 354.380 182.320 ;
        RECT 356.440 182.130 371.650 182.360 ;
        RECT 383.730 182.150 388.980 182.450 ;
        RECT 356.440 182.120 370.600 182.130 ;
        RECT 356.440 182.110 363.970 182.120 ;
        RECT 364.980 182.110 366.170 182.120 ;
        RECT 367.130 182.110 368.320 182.120 ;
        RECT 369.410 182.110 370.600 182.120 ;
        RECT 356.440 182.100 361.750 182.110 ;
        RECT 356.440 182.090 360.610 182.100 ;
        RECT 356.440 182.080 358.330 182.090 ;
        RECT 359.420 182.080 360.610 182.090 ;
        RECT 356.440 182.070 357.160 182.080 ;
        RECT 353.070 181.720 353.380 182.060 ;
        RECT 349.080 181.190 350.720 181.580 ;
        RECT 351.520 181.430 353.380 181.720 ;
        RECT 351.520 181.420 351.830 181.430 ;
        RECT 353.070 181.420 353.380 181.430 ;
        RECT 341.660 181.070 342.310 181.080 ;
        RECT 341.660 180.740 341.960 181.070 ;
        RECT 340.940 180.290 341.960 180.740 ;
        RECT 346.550 180.580 346.840 181.180 ;
        RECT 348.440 180.580 348.730 181.180 ;
        RECT 341.660 180.280 341.960 180.290 ;
        RECT 350.780 179.970 351.080 180.970 ;
        RECT 351.530 180.370 351.830 181.420 ;
        RECT 354.130 180.320 354.380 182.060 ;
        RECT 354.830 179.970 355.090 181.520 ;
        RECT 379.650 180.510 379.910 181.710 ;
        RECT 379.650 180.000 379.900 180.510 ;
        RECT 381.540 180.500 381.800 181.710 ;
        RECT 383.930 180.600 384.180 182.150 ;
        RECT 381.540 180.340 381.930 180.500 ;
        RECT 381.530 180.210 381.930 180.340 ;
        RECT 384.630 180.210 384.890 181.820 ;
        RECT 387.180 180.750 387.480 181.800 ;
        RECT 387.930 181.200 388.230 182.150 ;
        RECT 388.430 181.250 388.730 181.300 ;
        RECT 388.430 180.900 389.330 181.250 ;
        RECT 380.150 180.000 380.440 180.160 ;
        RECT 381.530 180.150 381.790 180.210 ;
        RECT 350.730 179.960 355.980 179.970 ;
        RECT 340.610 179.880 340.860 179.890 ;
        RECT 340.610 179.420 341.590 179.880 ;
        RECT 350.730 179.670 356.000 179.960 ;
        RECT 340.610 179.120 340.860 179.420 ;
        RECT 348.580 179.330 350.420 179.340 ;
        RECT 355.830 179.330 356.000 179.670 ;
        RECT 342.320 179.320 342.560 179.330 ;
        RECT 343.400 179.320 356.000 179.330 ;
        RECT 342.320 179.160 356.000 179.320 ;
        RECT 379.650 179.810 380.440 180.000 ;
        RECT 379.650 179.610 379.900 179.810 ;
        RECT 380.150 179.700 380.440 179.810 ;
        RECT 381.540 179.610 381.790 180.150 ;
        RECT 384.620 180.150 384.890 180.210 ;
        RECT 386.170 180.490 387.480 180.750 ;
        RECT 389.540 180.790 391.210 180.820 ;
        RECT 406.290 180.790 406.540 180.800 ;
        RECT 389.540 180.520 406.540 180.790 ;
        RECT 389.540 180.510 403.040 180.520 ;
        RECT 390.820 180.490 403.040 180.510 ;
        RECT 386.170 180.150 386.480 180.490 ;
        RECT 382.180 179.620 383.820 180.010 ;
        RECT 384.620 179.860 386.480 180.150 ;
        RECT 384.620 179.850 384.930 179.860 ;
        RECT 386.170 179.850 386.480 179.860 ;
        RECT 342.320 179.150 353.830 179.160 ;
        RECT 342.310 179.140 348.630 179.150 ;
        RECT 350.180 179.140 353.830 179.150 ;
        RECT 342.310 179.130 344.180 179.140 ;
        RECT 342.310 179.120 342.560 179.130 ;
        RECT 340.610 178.950 342.560 179.120 ;
        RECT 379.650 179.010 379.940 179.610 ;
        RECT 381.540 179.010 381.830 179.610 ;
        RECT 340.610 178.730 340.860 178.950 ;
        RECT 340.610 178.560 341.650 178.730 ;
        RECT 341.460 177.700 341.650 178.560 ;
        RECT 383.880 178.400 384.180 179.400 ;
        RECT 384.630 178.800 384.930 179.850 ;
        RECT 387.230 178.750 387.480 180.490 ;
        RECT 387.930 178.400 388.190 179.950 ;
        RECT 388.810 178.400 389.150 178.470 ;
        RECT 383.830 178.100 389.150 178.400 ;
        RECT 340.670 177.260 341.650 177.700 ;
        RECT 340.670 177.250 341.620 177.260 ;
        RECT 342.490 176.940 351.760 176.950 ;
        RECT 353.640 176.940 355.560 176.950 ;
        RECT 340.340 176.840 340.530 176.850 ;
        RECT 340.340 176.380 341.320 176.840 ;
        RECT 342.490 176.750 355.560 176.940 ;
        RECT 342.490 176.740 354.850 176.750 ;
        RECT 340.340 175.590 340.530 176.380 ;
        RECT 342.490 175.730 342.700 176.740 ;
        RECT 351.750 176.730 353.650 176.740 ;
        RECT 355.380 176.000 355.560 176.750 ;
        RECT 341.340 175.590 341.610 175.600 ;
        RECT 340.340 175.380 341.610 175.590 ;
        RECT 341.340 175.170 341.610 175.380 ;
        RECT 341.340 174.540 341.590 175.170 ;
        RECT 342.490 174.720 342.690 175.730 ;
        RECT 350.300 175.700 355.560 176.000 ;
        RECT 340.550 174.090 341.590 174.540 ;
        RECT 340.530 172.640 341.490 173.090 ;
        RECT 341.240 172.590 341.490 172.640 ;
        RECT 342.500 172.590 342.690 174.720 ;
        RECT 341.240 172.390 342.690 172.590 ;
        RECT 346.220 174.060 346.480 175.260 ;
        RECT 346.220 173.550 346.470 174.060 ;
        RECT 348.110 174.050 348.370 175.260 ;
        RECT 350.500 174.150 350.750 175.700 ;
        RECT 348.110 173.890 348.500 174.050 ;
        RECT 348.100 173.760 348.500 173.890 ;
        RECT 351.200 173.760 351.460 175.370 ;
        RECT 353.750 174.300 354.050 175.350 ;
        RECT 354.500 174.750 354.800 175.700 ;
        RECT 355.000 174.800 355.300 174.850 ;
        RECT 355.000 174.450 355.900 174.800 ;
        RECT 357.610 174.670 357.830 174.680 ;
        RECT 357.610 174.480 371.290 174.670 ;
        RECT 357.610 174.350 357.830 174.480 ;
        RECT 346.720 173.550 347.010 173.710 ;
        RECT 348.100 173.700 348.360 173.760 ;
        RECT 346.220 173.360 347.010 173.550 ;
        RECT 346.220 173.160 346.470 173.360 ;
        RECT 346.720 173.250 347.010 173.360 ;
        RECT 348.110 173.160 348.360 173.700 ;
        RECT 351.190 173.700 351.460 173.760 ;
        RECT 352.740 174.040 354.050 174.300 ;
        RECT 356.150 174.050 357.830 174.350 ;
        RECT 356.150 174.040 357.810 174.050 ;
        RECT 352.740 173.700 353.050 174.040 ;
        RECT 348.750 173.170 350.390 173.560 ;
        RECT 351.190 173.410 353.050 173.700 ;
        RECT 351.190 173.400 351.500 173.410 ;
        RECT 352.740 173.400 353.050 173.410 ;
        RECT 346.220 172.560 346.510 173.160 ;
        RECT 348.110 172.560 348.400 173.160 ;
        RECT 341.240 172.300 341.490 172.390 ;
        RECT 340.510 171.850 341.490 172.300 ;
        RECT 350.450 171.950 350.750 172.950 ;
        RECT 351.200 172.350 351.500 173.400 ;
        RECT 353.800 172.300 354.050 174.040 ;
        RECT 371.040 173.580 371.290 174.480 ;
        RECT 354.500 171.950 354.760 173.500 ;
        RECT 365.980 173.280 371.290 173.580 ;
        RECT 350.400 171.930 355.650 171.950 ;
        RECT 350.400 171.650 355.770 171.930 ;
        RECT 343.850 171.250 344.130 171.320 ;
        RECT 345.030 171.280 345.310 171.310 ;
        RECT 355.480 171.280 355.770 171.650 ;
        RECT 345.030 171.270 355.770 171.280 ;
        RECT 342.440 171.050 344.130 171.250 ;
        RECT 341.230 170.850 341.510 170.860 ;
        RECT 340.490 170.400 341.510 170.850 ;
        RECT 342.440 170.400 342.670 171.050 ;
        RECT 343.850 170.990 344.130 171.050 ;
        RECT 345.010 171.040 355.770 171.270 ;
        RECT 345.030 171.030 355.770 171.040 ;
        RECT 361.900 171.640 362.160 172.840 ;
        RECT 361.900 171.130 362.150 171.640 ;
        RECT 363.790 171.630 364.050 172.840 ;
        RECT 366.180 171.730 366.430 173.280 ;
        RECT 363.790 171.470 364.180 171.630 ;
        RECT 363.780 171.340 364.180 171.470 ;
        RECT 366.880 171.340 367.140 172.950 ;
        RECT 369.430 171.880 369.730 172.930 ;
        RECT 370.180 172.330 370.480 173.280 ;
        RECT 370.680 172.380 370.980 172.430 ;
        RECT 370.680 172.030 371.580 172.380 ;
        RECT 388.810 171.980 389.150 178.100 ;
        RECT 388.240 171.960 389.200 171.980 ;
        RECT 372.720 171.940 377.000 171.950 ;
        RECT 384.400 171.940 389.200 171.960 ;
        RECT 372.720 171.930 389.200 171.940 ;
        RECT 362.400 171.130 362.690 171.290 ;
        RECT 363.780 171.280 364.040 171.340 ;
        RECT 345.030 171.020 355.730 171.030 ;
        RECT 345.030 170.980 345.310 171.020 ;
        RECT 361.900 170.940 362.690 171.130 ;
        RECT 361.900 170.740 362.150 170.940 ;
        RECT 362.400 170.830 362.690 170.940 ;
        RECT 363.790 170.740 364.040 171.280 ;
        RECT 366.870 171.280 367.140 171.340 ;
        RECT 368.420 171.620 369.730 171.880 ;
        RECT 368.420 171.280 368.730 171.620 ;
        RECT 364.430 170.750 366.070 171.140 ;
        RECT 366.870 170.990 368.730 171.280 ;
        RECT 366.870 170.980 367.180 170.990 ;
        RECT 368.420 170.980 368.730 170.990 ;
        RECT 343.830 170.420 344.100 170.500 ;
        RECT 341.230 170.190 342.670 170.400 ;
        RECT 343.220 170.200 344.100 170.420 ;
        RECT 341.230 169.140 341.510 170.190 ;
        RECT 343.220 169.390 343.440 170.200 ;
        RECT 343.830 170.170 344.100 170.200 ;
        RECT 344.960 170.460 345.250 170.510 ;
        RECT 344.960 170.280 355.710 170.460 ;
        RECT 344.960 170.180 345.250 170.280 ;
        RECT 349.800 170.270 353.430 170.280 ;
        RECT 355.510 169.600 355.710 170.280 ;
        RECT 361.900 170.140 362.190 170.740 ;
        RECT 363.790 170.140 364.080 170.740 ;
        RECT 340.510 168.690 341.510 169.140 ;
        RECT 340.490 167.240 341.790 167.690 ;
        RECT 341.490 166.840 341.790 167.240 ;
        RECT 343.210 166.860 343.440 169.390 ;
        RECT 350.460 169.300 355.710 169.600 ;
        RECT 366.130 169.530 366.430 170.530 ;
        RECT 366.880 169.930 367.180 170.980 ;
        RECT 369.480 169.880 369.730 171.620 ;
        RECT 371.850 171.620 389.200 171.930 ;
        RECT 371.850 171.610 384.860 171.620 ;
        RECT 376.710 171.600 384.860 171.610 ;
        RECT 388.240 171.580 389.200 171.620 ;
        RECT 388.810 171.570 389.150 171.580 ;
        RECT 370.180 169.530 370.440 171.080 ;
        RECT 371.270 169.530 371.470 169.540 ;
        RECT 342.280 166.840 343.440 166.860 ;
        RECT 341.490 166.660 343.440 166.840 ;
        RECT 346.380 167.660 346.640 168.860 ;
        RECT 346.380 167.150 346.630 167.660 ;
        RECT 348.270 167.650 348.530 168.860 ;
        RECT 350.660 167.750 350.910 169.300 ;
        RECT 348.270 167.490 348.660 167.650 ;
        RECT 348.260 167.360 348.660 167.490 ;
        RECT 351.360 167.360 351.620 168.970 ;
        RECT 353.910 167.900 354.210 168.950 ;
        RECT 354.660 168.350 354.960 169.300 ;
        RECT 355.510 169.290 355.710 169.300 ;
        RECT 366.080 169.230 371.470 169.530 ;
        RECT 355.160 168.400 355.460 168.450 ;
        RECT 355.160 168.050 356.060 168.400 ;
        RECT 371.270 167.990 371.470 169.230 ;
        RECT 363.710 167.970 364.900 167.980 ;
        RECT 365.890 167.970 367.080 167.980 ;
        RECT 368.110 167.970 369.300 167.980 ;
        RECT 370.290 167.970 371.480 167.990 ;
        RECT 361.500 167.960 371.480 167.970 ;
        RECT 358.110 167.940 359.300 167.950 ;
        RECT 360.390 167.940 371.480 167.960 ;
        RECT 346.880 167.150 347.170 167.310 ;
        RECT 348.260 167.300 348.520 167.360 ;
        RECT 346.380 166.960 347.170 167.150 ;
        RECT 346.380 166.760 346.630 166.960 ;
        RECT 346.880 166.850 347.170 166.960 ;
        RECT 348.270 166.760 348.520 167.300 ;
        RECT 351.350 167.300 351.620 167.360 ;
        RECT 352.900 167.640 354.210 167.900 ;
        RECT 356.270 167.710 371.480 167.940 ;
        RECT 356.270 167.700 370.430 167.710 ;
        RECT 356.270 167.690 363.800 167.700 ;
        RECT 364.810 167.690 366.000 167.700 ;
        RECT 366.960 167.690 368.150 167.700 ;
        RECT 369.240 167.690 370.430 167.700 ;
        RECT 356.270 167.680 361.580 167.690 ;
        RECT 356.270 167.670 360.440 167.680 ;
        RECT 356.270 167.660 358.160 167.670 ;
        RECT 359.250 167.660 360.440 167.670 ;
        RECT 356.270 167.650 356.990 167.660 ;
        RECT 352.900 167.300 353.210 167.640 ;
        RECT 348.910 166.770 350.550 167.160 ;
        RECT 351.350 167.010 353.210 167.300 ;
        RECT 351.350 167.000 351.660 167.010 ;
        RECT 352.900 167.000 353.210 167.010 ;
        RECT 341.490 166.650 342.140 166.660 ;
        RECT 341.490 166.320 341.790 166.650 ;
        RECT 337.380 165.940 337.640 166.120 ;
        RECT 335.840 158.580 336.070 160.550 ;
        RECT 335.840 156.690 336.090 158.580 ;
        RECT 335.840 154.890 336.110 156.690 ;
        RECT 288.200 150.630 305.360 150.920 ;
        RECT 288.890 150.620 305.360 150.630 ;
        RECT 284.830 150.270 285.140 150.610 ;
        RECT 280.840 149.740 282.480 150.130 ;
        RECT 283.280 149.980 285.140 150.270 ;
        RECT 283.280 149.970 283.590 149.980 ;
        RECT 284.830 149.970 285.140 149.980 ;
        RECT 240.980 149.270 252.490 149.280 ;
        RECT 240.970 149.260 247.290 149.270 ;
        RECT 248.840 149.260 252.490 149.270 ;
        RECT 240.970 149.250 242.840 149.260 ;
        RECT 240.970 149.240 241.220 149.250 ;
        RECT 239.270 149.070 241.220 149.240 ;
        RECT 278.310 149.130 278.600 149.730 ;
        RECT 280.200 149.130 280.490 149.730 ;
        RECT 239.270 148.850 239.520 149.070 ;
        RECT 239.270 148.680 240.310 148.850 ;
        RECT 240.120 147.820 240.310 148.680 ;
        RECT 282.540 148.520 282.840 149.520 ;
        RECT 283.290 148.920 283.590 149.970 ;
        RECT 285.890 148.870 286.140 150.610 ;
        RECT 286.590 148.520 286.850 150.070 ;
        RECT 335.840 149.650 336.130 154.890 ;
        RECT 287.470 148.520 287.810 148.590 ;
        RECT 282.490 148.220 287.810 148.520 ;
        RECT 239.330 147.380 240.310 147.820 ;
        RECT 239.330 147.370 240.280 147.380 ;
        RECT 241.150 147.060 250.420 147.070 ;
        RECT 252.300 147.060 254.220 147.070 ;
        RECT 239.000 146.960 239.190 146.970 ;
        RECT 239.000 146.500 239.980 146.960 ;
        RECT 241.150 146.870 254.220 147.060 ;
        RECT 241.150 146.860 253.510 146.870 ;
        RECT 239.000 145.710 239.190 146.500 ;
        RECT 241.150 145.850 241.360 146.860 ;
        RECT 250.410 146.850 252.310 146.860 ;
        RECT 254.040 146.120 254.220 146.870 ;
        RECT 240.000 145.710 240.270 145.720 ;
        RECT 239.000 145.500 240.270 145.710 ;
        RECT 240.000 145.290 240.270 145.500 ;
        RECT 240.000 144.660 240.250 145.290 ;
        RECT 241.150 144.840 241.350 145.850 ;
        RECT 248.960 145.820 254.220 146.120 ;
        RECT 239.210 144.210 240.250 144.660 ;
        RECT 239.190 142.760 240.150 143.210 ;
        RECT 239.900 142.710 240.150 142.760 ;
        RECT 241.160 142.710 241.350 144.840 ;
        RECT 239.900 142.510 241.350 142.710 ;
        RECT 244.880 144.180 245.140 145.380 ;
        RECT 244.880 143.670 245.130 144.180 ;
        RECT 246.770 144.170 247.030 145.380 ;
        RECT 249.160 144.270 249.410 145.820 ;
        RECT 246.770 144.010 247.160 144.170 ;
        RECT 246.760 143.880 247.160 144.010 ;
        RECT 249.860 143.880 250.120 145.490 ;
        RECT 252.410 144.420 252.710 145.470 ;
        RECT 253.160 144.870 253.460 145.820 ;
        RECT 253.660 144.920 253.960 144.970 ;
        RECT 253.660 144.570 254.560 144.920 ;
        RECT 256.270 144.790 256.490 144.800 ;
        RECT 256.270 144.600 269.950 144.790 ;
        RECT 256.270 144.470 256.490 144.600 ;
        RECT 245.380 143.670 245.670 143.830 ;
        RECT 246.760 143.820 247.020 143.880 ;
        RECT 244.880 143.480 245.670 143.670 ;
        RECT 244.880 143.280 245.130 143.480 ;
        RECT 245.380 143.370 245.670 143.480 ;
        RECT 246.770 143.280 247.020 143.820 ;
        RECT 249.850 143.820 250.120 143.880 ;
        RECT 251.400 144.160 252.710 144.420 ;
        RECT 254.810 144.170 256.490 144.470 ;
        RECT 254.810 144.160 256.470 144.170 ;
        RECT 251.400 143.820 251.710 144.160 ;
        RECT 247.410 143.290 249.050 143.680 ;
        RECT 249.850 143.530 251.710 143.820 ;
        RECT 249.850 143.520 250.160 143.530 ;
        RECT 251.400 143.520 251.710 143.530 ;
        RECT 244.880 142.680 245.170 143.280 ;
        RECT 246.770 142.680 247.060 143.280 ;
        RECT 239.900 142.420 240.150 142.510 ;
        RECT 239.170 141.970 240.150 142.420 ;
        RECT 249.110 142.070 249.410 143.070 ;
        RECT 249.860 142.470 250.160 143.520 ;
        RECT 252.460 142.420 252.710 144.160 ;
        RECT 269.700 143.700 269.950 144.600 ;
        RECT 253.160 142.070 253.420 143.620 ;
        RECT 264.640 143.400 269.950 143.700 ;
        RECT 249.060 142.050 254.310 142.070 ;
        RECT 249.060 141.770 254.430 142.050 ;
        RECT 242.510 141.370 242.790 141.440 ;
        RECT 243.690 141.400 243.970 141.430 ;
        RECT 254.140 141.400 254.430 141.770 ;
        RECT 243.690 141.390 254.430 141.400 ;
        RECT 241.100 141.170 242.790 141.370 ;
        RECT 239.890 140.970 240.170 140.980 ;
        RECT 239.150 140.520 240.170 140.970 ;
        RECT 241.100 140.520 241.330 141.170 ;
        RECT 242.510 141.110 242.790 141.170 ;
        RECT 243.670 141.160 254.430 141.390 ;
        RECT 243.690 141.150 254.430 141.160 ;
        RECT 260.560 141.760 260.820 142.960 ;
        RECT 260.560 141.250 260.810 141.760 ;
        RECT 262.450 141.750 262.710 142.960 ;
        RECT 264.840 141.850 265.090 143.400 ;
        RECT 262.450 141.590 262.840 141.750 ;
        RECT 262.440 141.460 262.840 141.590 ;
        RECT 265.540 141.460 265.800 143.070 ;
        RECT 268.090 142.000 268.390 143.050 ;
        RECT 268.840 142.450 269.140 143.400 ;
        RECT 269.340 142.500 269.640 142.550 ;
        RECT 269.340 142.150 270.240 142.500 ;
        RECT 287.470 142.100 287.810 148.220 ;
        RECT 335.840 147.680 336.070 149.650 ;
        RECT 337.400 149.140 337.640 165.940 ;
        RECT 340.770 165.870 341.790 166.320 ;
        RECT 346.380 166.160 346.670 166.760 ;
        RECT 348.270 166.160 348.560 166.760 ;
        RECT 341.490 165.860 341.790 165.870 ;
        RECT 350.610 165.550 350.910 166.550 ;
        RECT 351.360 165.950 351.660 167.000 ;
        RECT 353.960 165.900 354.210 167.640 ;
        RECT 406.290 167.380 406.550 180.520 ;
        RECT 406.280 167.260 406.550 167.380 ;
        RECT 420.880 176.530 421.150 186.050 ;
        RECT 437.110 192.420 437.420 196.090 ;
        RECT 437.110 190.640 437.440 192.420 ;
        RECT 437.110 188.670 437.400 190.640 ;
        RECT 437.110 186.840 437.420 188.670 ;
        RECT 437.110 183.020 437.400 186.840 ;
        RECT 437.110 181.050 437.380 183.020 ;
        RECT 437.110 179.330 437.440 181.050 ;
        RECT 437.110 177.410 437.400 179.330 ;
        RECT 354.660 165.550 354.920 167.100 ;
        RECT 406.280 166.430 406.540 167.260 ;
        RECT 420.880 166.580 421.060 176.530 ;
        RECT 437.110 167.870 437.380 177.410 ;
        RECT 401.260 166.130 406.540 166.430 ;
        RECT 350.560 165.540 355.810 165.550 ;
        RECT 340.440 165.460 340.690 165.470 ;
        RECT 340.440 165.000 341.420 165.460 ;
        RECT 350.560 165.250 355.830 165.540 ;
        RECT 340.440 164.700 340.690 165.000 ;
        RECT 348.410 164.910 350.250 164.920 ;
        RECT 355.660 164.910 355.830 165.250 ;
        RECT 342.150 164.900 342.390 164.910 ;
        RECT 343.230 164.900 355.830 164.910 ;
        RECT 342.150 164.740 355.830 164.900 ;
        RECT 342.150 164.730 353.660 164.740 ;
        RECT 342.140 164.720 348.460 164.730 ;
        RECT 350.010 164.720 353.660 164.730 ;
        RECT 342.140 164.710 344.010 164.720 ;
        RECT 342.140 164.700 342.390 164.710 ;
        RECT 340.440 164.530 342.390 164.700 ;
        RECT 340.440 164.230 340.710 164.530 ;
        RECT 340.450 163.970 340.710 164.230 ;
        RECT 397.180 164.490 397.440 165.690 ;
        RECT 397.180 163.980 397.430 164.490 ;
        RECT 399.070 164.480 399.330 165.690 ;
        RECT 401.460 164.580 401.710 166.130 ;
        RECT 399.070 164.320 399.460 164.480 ;
        RECT 399.060 164.190 399.460 164.320 ;
        RECT 402.160 164.190 402.420 165.800 ;
        RECT 404.710 164.730 405.010 165.780 ;
        RECT 405.460 165.180 405.760 166.130 ;
        RECT 405.960 165.230 406.260 165.280 ;
        RECT 405.960 164.880 406.860 165.230 ;
        RECT 420.870 164.770 421.070 166.580 ;
        RECT 397.680 163.980 397.970 164.140 ;
        RECT 399.060 164.130 399.320 164.190 ;
        RECT 340.430 163.580 340.730 163.970 ;
        RECT 397.180 163.790 397.970 163.980 ;
        RECT 397.180 163.590 397.430 163.790 ;
        RECT 397.680 163.680 397.970 163.790 ;
        RECT 399.070 163.590 399.320 164.130 ;
        RECT 402.150 164.130 402.420 164.190 ;
        RECT 403.700 164.470 405.010 164.730 ;
        RECT 407.130 164.480 421.070 164.770 ;
        RECT 437.150 166.000 437.420 167.870 ;
        RECT 407.130 164.470 421.030 164.480 ;
        RECT 403.700 164.130 404.010 164.470 ;
        RECT 399.710 163.600 401.350 163.990 ;
        RECT 402.150 163.840 404.010 164.130 ;
        RECT 402.150 163.830 402.460 163.840 ;
        RECT 403.700 163.830 404.010 163.840 ;
        RECT 340.430 163.350 341.920 163.580 ;
        RECT 341.670 162.420 341.920 163.350 ;
        RECT 397.180 162.990 397.470 163.590 ;
        RECT 399.070 162.990 399.360 163.590 ;
        RECT 340.870 161.960 341.920 162.420 ;
        RECT 401.410 162.380 401.710 163.380 ;
        RECT 402.160 162.780 402.460 163.830 ;
        RECT 404.760 162.730 405.010 164.470 ;
        RECT 407.720 164.460 421.030 164.470 ;
        RECT 405.460 162.380 405.720 163.930 ;
        RECT 401.360 162.080 406.630 162.380 ;
        RECT 341.670 161.950 341.920 161.960 ;
        RECT 340.540 161.550 340.790 161.560 ;
        RECT 340.540 161.100 341.520 161.550 ;
        RECT 342.630 161.290 351.900 161.300 ;
        RECT 353.780 161.290 355.700 161.300 ;
        RECT 342.630 161.100 355.700 161.290 ;
        RECT 340.540 160.490 340.790 161.100 ;
        RECT 342.630 161.090 354.990 161.100 ;
        RECT 340.540 160.240 341.750 160.490 ;
        RECT 341.480 159.490 341.740 160.240 ;
        RECT 342.630 160.080 342.840 161.090 ;
        RECT 351.890 161.080 353.790 161.090 ;
        RECT 355.520 160.350 355.700 161.100 ;
        RECT 341.480 158.890 341.730 159.490 ;
        RECT 342.630 159.070 342.830 160.080 ;
        RECT 350.440 160.050 355.700 160.350 ;
        RECT 340.690 158.440 341.730 158.890 ;
        RECT 340.670 156.990 341.630 157.440 ;
        RECT 341.380 156.940 341.630 156.990 ;
        RECT 342.640 156.940 342.830 159.070 ;
        RECT 341.380 156.740 342.830 156.940 ;
        RECT 346.360 158.410 346.620 159.610 ;
        RECT 346.360 157.900 346.610 158.410 ;
        RECT 348.250 158.400 348.510 159.610 ;
        RECT 350.640 158.500 350.890 160.050 ;
        RECT 348.250 158.240 348.640 158.400 ;
        RECT 348.240 158.110 348.640 158.240 ;
        RECT 351.340 158.110 351.600 159.720 ;
        RECT 353.890 158.650 354.190 159.700 ;
        RECT 354.640 159.100 354.940 160.050 ;
        RECT 355.140 159.150 355.440 159.200 ;
        RECT 355.140 158.800 356.040 159.150 ;
        RECT 357.750 159.020 357.970 159.030 ;
        RECT 357.750 158.830 371.430 159.020 ;
        RECT 357.750 158.700 357.970 158.830 ;
        RECT 346.860 157.900 347.150 158.060 ;
        RECT 348.240 158.050 348.500 158.110 ;
        RECT 346.360 157.710 347.150 157.900 ;
        RECT 346.360 157.510 346.610 157.710 ;
        RECT 346.860 157.600 347.150 157.710 ;
        RECT 348.250 157.510 348.500 158.050 ;
        RECT 351.330 158.050 351.600 158.110 ;
        RECT 352.880 158.390 354.190 158.650 ;
        RECT 356.290 158.400 357.970 158.700 ;
        RECT 356.290 158.390 357.950 158.400 ;
        RECT 352.880 158.050 353.190 158.390 ;
        RECT 348.890 157.520 350.530 157.910 ;
        RECT 351.330 157.760 353.190 158.050 ;
        RECT 351.330 157.750 351.640 157.760 ;
        RECT 352.880 157.750 353.190 157.760 ;
        RECT 346.360 156.910 346.650 157.510 ;
        RECT 348.250 156.910 348.540 157.510 ;
        RECT 341.380 156.650 341.630 156.740 ;
        RECT 340.650 156.200 341.630 156.650 ;
        RECT 350.590 156.300 350.890 157.300 ;
        RECT 351.340 156.700 351.640 157.750 ;
        RECT 353.940 156.650 354.190 158.390 ;
        RECT 371.180 157.930 371.430 158.830 ;
        RECT 354.640 156.300 354.900 157.850 ;
        RECT 366.120 157.630 371.430 157.930 ;
        RECT 350.540 156.280 355.790 156.300 ;
        RECT 350.540 156.000 355.910 156.280 ;
        RECT 343.990 155.600 344.270 155.670 ;
        RECT 345.170 155.630 345.450 155.660 ;
        RECT 355.620 155.630 355.910 156.000 ;
        RECT 345.170 155.620 355.910 155.630 ;
        RECT 342.580 155.400 344.270 155.600 ;
        RECT 341.370 155.200 341.650 155.210 ;
        RECT 340.630 154.750 341.650 155.200 ;
        RECT 342.580 154.750 342.810 155.400 ;
        RECT 343.990 155.340 344.270 155.400 ;
        RECT 345.150 155.390 355.910 155.620 ;
        RECT 345.170 155.380 355.910 155.390 ;
        RECT 362.040 155.990 362.300 157.190 ;
        RECT 362.040 155.480 362.290 155.990 ;
        RECT 363.930 155.980 364.190 157.190 ;
        RECT 366.320 156.080 366.570 157.630 ;
        RECT 363.930 155.820 364.320 155.980 ;
        RECT 363.920 155.690 364.320 155.820 ;
        RECT 367.020 155.690 367.280 157.300 ;
        RECT 369.570 156.230 369.870 157.280 ;
        RECT 370.320 156.680 370.620 157.630 ;
        RECT 370.820 156.730 371.120 156.780 ;
        RECT 370.820 156.380 371.720 156.730 ;
        RECT 384.480 156.330 388.950 156.360 ;
        RECT 373.540 156.300 388.950 156.330 ;
        RECT 372.870 156.280 388.950 156.300 ;
        RECT 362.540 155.480 362.830 155.640 ;
        RECT 363.920 155.630 364.180 155.690 ;
        RECT 345.170 155.370 355.870 155.380 ;
        RECT 345.170 155.330 345.450 155.370 ;
        RECT 362.040 155.290 362.830 155.480 ;
        RECT 362.040 155.090 362.290 155.290 ;
        RECT 362.540 155.180 362.830 155.290 ;
        RECT 363.930 155.090 364.180 155.630 ;
        RECT 367.010 155.630 367.280 155.690 ;
        RECT 368.560 155.970 369.870 156.230 ;
        RECT 368.560 155.630 368.870 155.970 ;
        RECT 364.570 155.100 366.210 155.490 ;
        RECT 367.010 155.340 368.870 155.630 ;
        RECT 367.010 155.330 367.320 155.340 ;
        RECT 368.560 155.330 368.870 155.340 ;
        RECT 343.970 154.770 344.240 154.850 ;
        RECT 341.370 154.540 342.810 154.750 ;
        RECT 343.360 154.550 344.240 154.770 ;
        RECT 341.370 153.490 341.650 154.540 ;
        RECT 343.360 153.740 343.580 154.550 ;
        RECT 343.970 154.520 344.240 154.550 ;
        RECT 345.100 154.810 345.390 154.860 ;
        RECT 345.100 154.630 355.850 154.810 ;
        RECT 345.100 154.530 345.390 154.630 ;
        RECT 349.940 154.620 353.570 154.630 ;
        RECT 355.650 153.950 355.850 154.630 ;
        RECT 362.040 154.490 362.330 155.090 ;
        RECT 363.930 154.490 364.220 155.090 ;
        RECT 340.650 153.040 341.650 153.490 ;
        RECT 340.630 151.590 341.930 152.040 ;
        RECT 341.630 151.190 341.930 151.590 ;
        RECT 343.350 151.210 343.580 153.740 ;
        RECT 350.600 153.650 355.850 153.950 ;
        RECT 366.270 153.880 366.570 154.880 ;
        RECT 367.020 154.280 367.320 155.330 ;
        RECT 369.620 154.230 369.870 155.970 ;
        RECT 371.990 155.960 388.950 156.280 ;
        RECT 372.870 155.950 388.950 155.960 ;
        RECT 372.870 155.920 384.850 155.950 ;
        RECT 372.870 155.910 373.760 155.920 ;
        RECT 370.320 153.880 370.580 155.430 ;
        RECT 371.410 153.880 371.610 153.890 ;
        RECT 342.420 151.190 343.580 151.210 ;
        RECT 341.630 151.010 343.580 151.190 ;
        RECT 346.520 152.010 346.780 153.210 ;
        RECT 346.520 151.500 346.770 152.010 ;
        RECT 348.410 152.000 348.670 153.210 ;
        RECT 350.800 152.100 351.050 153.650 ;
        RECT 348.410 151.840 348.800 152.000 ;
        RECT 348.400 151.710 348.800 151.840 ;
        RECT 351.500 151.710 351.760 153.320 ;
        RECT 354.050 152.250 354.350 153.300 ;
        RECT 354.800 152.700 355.100 153.650 ;
        RECT 355.650 153.640 355.850 153.650 ;
        RECT 366.220 153.580 371.610 153.880 ;
        RECT 355.300 152.750 355.600 152.800 ;
        RECT 355.300 152.400 356.200 152.750 ;
        RECT 371.410 152.340 371.610 153.580 ;
        RECT 388.570 152.380 388.930 155.950 ;
        RECT 363.850 152.320 365.040 152.330 ;
        RECT 366.030 152.320 367.220 152.330 ;
        RECT 368.250 152.320 369.440 152.330 ;
        RECT 370.430 152.320 371.620 152.340 ;
        RECT 361.640 152.310 371.620 152.320 ;
        RECT 358.250 152.290 359.440 152.300 ;
        RECT 360.530 152.290 371.620 152.310 ;
        RECT 347.020 151.500 347.310 151.660 ;
        RECT 348.400 151.650 348.660 151.710 ;
        RECT 346.520 151.310 347.310 151.500 ;
        RECT 346.520 151.110 346.770 151.310 ;
        RECT 347.020 151.200 347.310 151.310 ;
        RECT 348.410 151.110 348.660 151.650 ;
        RECT 351.490 151.650 351.760 151.710 ;
        RECT 353.040 151.990 354.350 152.250 ;
        RECT 356.410 152.060 371.620 152.290 ;
        RECT 383.700 152.080 388.950 152.380 ;
        RECT 356.410 152.050 370.570 152.060 ;
        RECT 356.410 152.040 363.940 152.050 ;
        RECT 364.950 152.040 366.140 152.050 ;
        RECT 367.100 152.040 368.290 152.050 ;
        RECT 369.380 152.040 370.570 152.050 ;
        RECT 356.410 152.030 361.720 152.040 ;
        RECT 356.410 152.020 360.580 152.030 ;
        RECT 356.410 152.010 358.300 152.020 ;
        RECT 359.390 152.010 360.580 152.020 ;
        RECT 356.410 152.000 357.130 152.010 ;
        RECT 353.040 151.650 353.350 151.990 ;
        RECT 349.050 151.120 350.690 151.510 ;
        RECT 351.490 151.360 353.350 151.650 ;
        RECT 351.490 151.350 351.800 151.360 ;
        RECT 353.040 151.350 353.350 151.360 ;
        RECT 341.630 151.000 342.280 151.010 ;
        RECT 341.630 150.670 341.930 151.000 ;
        RECT 340.910 150.220 341.930 150.670 ;
        RECT 346.520 150.510 346.810 151.110 ;
        RECT 348.410 150.510 348.700 151.110 ;
        RECT 341.630 150.210 341.930 150.220 ;
        RECT 350.750 149.900 351.050 150.900 ;
        RECT 351.500 150.300 351.800 151.350 ;
        RECT 354.100 150.250 354.350 151.990 ;
        RECT 354.800 149.900 355.060 151.450 ;
        RECT 379.620 150.440 379.880 151.640 ;
        RECT 379.620 149.930 379.870 150.440 ;
        RECT 381.510 150.430 381.770 151.640 ;
        RECT 383.900 150.530 384.150 152.080 ;
        RECT 381.510 150.270 381.900 150.430 ;
        RECT 381.500 150.140 381.900 150.270 ;
        RECT 384.600 150.140 384.860 151.750 ;
        RECT 387.150 150.680 387.450 151.730 ;
        RECT 387.900 151.130 388.200 152.080 ;
        RECT 388.400 151.180 388.700 151.230 ;
        RECT 388.400 150.830 389.300 151.180 ;
        RECT 380.120 149.930 380.410 150.090 ;
        RECT 381.500 150.080 381.760 150.140 ;
        RECT 350.700 149.890 355.950 149.900 ;
        RECT 337.370 148.930 337.640 149.140 ;
        RECT 340.580 149.810 340.830 149.820 ;
        RECT 340.580 149.350 341.560 149.810 ;
        RECT 350.700 149.600 355.970 149.890 ;
        RECT 340.580 149.050 340.830 149.350 ;
        RECT 348.550 149.260 350.390 149.270 ;
        RECT 355.800 149.260 355.970 149.600 ;
        RECT 342.290 149.250 342.530 149.260 ;
        RECT 343.370 149.250 355.970 149.260 ;
        RECT 342.290 149.090 355.970 149.250 ;
        RECT 379.620 149.740 380.410 149.930 ;
        RECT 379.620 149.540 379.870 149.740 ;
        RECT 380.120 149.630 380.410 149.740 ;
        RECT 381.510 149.540 381.760 150.080 ;
        RECT 384.590 150.080 384.860 150.140 ;
        RECT 386.140 150.420 387.450 150.680 ;
        RECT 389.510 150.730 391.180 150.750 ;
        RECT 406.320 150.730 406.630 162.080 ;
        RECT 437.150 160.360 437.400 166.000 ;
        RECT 437.150 158.390 437.380 160.360 ;
        RECT 437.150 156.500 437.400 158.390 ;
        RECT 437.150 154.700 437.420 156.500 ;
        RECT 389.510 150.440 406.670 150.730 ;
        RECT 390.200 150.430 406.670 150.440 ;
        RECT 386.140 150.080 386.450 150.420 ;
        RECT 382.150 149.550 383.790 149.940 ;
        RECT 384.590 149.790 386.450 150.080 ;
        RECT 384.590 149.780 384.900 149.790 ;
        RECT 386.140 149.780 386.450 149.790 ;
        RECT 342.290 149.080 353.800 149.090 ;
        RECT 342.280 149.070 348.600 149.080 ;
        RECT 350.150 149.070 353.800 149.080 ;
        RECT 342.280 149.060 344.150 149.070 ;
        RECT 342.280 149.050 342.530 149.060 ;
        RECT 335.840 144.090 336.110 147.680 ;
        RECT 337.370 145.700 337.610 148.930 ;
        RECT 340.580 148.880 342.530 149.050 ;
        RECT 379.620 148.940 379.910 149.540 ;
        RECT 381.510 148.940 381.800 149.540 ;
        RECT 340.580 148.660 340.830 148.880 ;
        RECT 340.580 148.490 341.620 148.660 ;
        RECT 341.430 147.630 341.620 148.490 ;
        RECT 383.850 148.330 384.150 149.330 ;
        RECT 384.600 148.730 384.900 149.780 ;
        RECT 387.200 148.680 387.450 150.420 ;
        RECT 387.900 148.330 388.160 149.880 ;
        RECT 437.150 149.460 437.440 154.700 ;
        RECT 388.780 148.330 389.120 148.400 ;
        RECT 383.800 148.030 389.120 148.330 ;
        RECT 340.640 147.190 341.620 147.630 ;
        RECT 340.640 147.180 341.590 147.190 ;
        RECT 342.460 146.870 351.730 146.880 ;
        RECT 353.610 146.870 355.530 146.880 ;
        RECT 340.310 146.770 340.500 146.780 ;
        RECT 340.310 146.310 341.290 146.770 ;
        RECT 342.460 146.680 355.530 146.870 ;
        RECT 342.460 146.670 354.820 146.680 ;
        RECT 337.370 145.530 337.620 145.700 ;
        RECT 335.840 142.270 336.090 144.090 ;
        RECT 286.900 142.080 287.860 142.100 ;
        RECT 271.380 142.060 275.660 142.070 ;
        RECT 283.060 142.060 287.860 142.080 ;
        RECT 271.380 142.050 287.860 142.060 ;
        RECT 261.060 141.250 261.350 141.410 ;
        RECT 262.440 141.400 262.700 141.460 ;
        RECT 243.690 141.140 254.390 141.150 ;
        RECT 243.690 141.100 243.970 141.140 ;
        RECT 260.560 141.060 261.350 141.250 ;
        RECT 260.560 140.860 260.810 141.060 ;
        RECT 261.060 140.950 261.350 141.060 ;
        RECT 262.450 140.860 262.700 141.400 ;
        RECT 265.530 141.400 265.800 141.460 ;
        RECT 267.080 141.740 268.390 142.000 ;
        RECT 267.080 141.400 267.390 141.740 ;
        RECT 263.090 140.870 264.730 141.260 ;
        RECT 265.530 141.110 267.390 141.400 ;
        RECT 265.530 141.100 265.840 141.110 ;
        RECT 267.080 141.100 267.390 141.110 ;
        RECT 242.490 140.540 242.760 140.620 ;
        RECT 239.890 140.310 241.330 140.520 ;
        RECT 241.880 140.320 242.760 140.540 ;
        RECT 239.890 139.260 240.170 140.310 ;
        RECT 241.880 139.510 242.100 140.320 ;
        RECT 242.490 140.290 242.760 140.320 ;
        RECT 243.620 140.580 243.910 140.630 ;
        RECT 243.620 140.400 254.370 140.580 ;
        RECT 243.620 140.300 243.910 140.400 ;
        RECT 248.460 140.390 252.090 140.400 ;
        RECT 254.170 139.720 254.370 140.400 ;
        RECT 260.560 140.260 260.850 140.860 ;
        RECT 262.450 140.260 262.740 140.860 ;
        RECT 239.170 138.810 240.170 139.260 ;
        RECT 239.150 137.360 240.450 137.810 ;
        RECT 240.150 136.960 240.450 137.360 ;
        RECT 241.870 136.980 242.100 139.510 ;
        RECT 249.120 139.420 254.370 139.720 ;
        RECT 264.790 139.650 265.090 140.650 ;
        RECT 265.540 140.050 265.840 141.100 ;
        RECT 268.140 140.000 268.390 141.740 ;
        RECT 270.510 141.740 287.860 142.050 ;
        RECT 270.510 141.730 283.520 141.740 ;
        RECT 275.370 141.720 283.520 141.730 ;
        RECT 286.900 141.700 287.860 141.740 ;
        RECT 287.470 141.690 287.810 141.700 ;
        RECT 268.840 139.650 269.100 141.200 ;
        RECT 269.930 139.650 270.130 139.660 ;
        RECT 240.940 136.960 242.100 136.980 ;
        RECT 240.150 136.780 242.100 136.960 ;
        RECT 245.040 137.780 245.300 138.980 ;
        RECT 245.040 137.270 245.290 137.780 ;
        RECT 246.930 137.770 247.190 138.980 ;
        RECT 249.320 137.870 249.570 139.420 ;
        RECT 246.930 137.610 247.320 137.770 ;
        RECT 246.920 137.480 247.320 137.610 ;
        RECT 250.020 137.480 250.280 139.090 ;
        RECT 252.570 138.020 252.870 139.070 ;
        RECT 253.320 138.470 253.620 139.420 ;
        RECT 254.170 139.410 254.370 139.420 ;
        RECT 264.740 139.350 270.130 139.650 ;
        RECT 253.820 138.520 254.120 138.570 ;
        RECT 253.820 138.170 254.720 138.520 ;
        RECT 269.930 138.110 270.130 139.350 ;
        RECT 335.840 138.810 336.070 142.270 ;
        RECT 337.380 142.240 337.620 145.530 ;
        RECT 340.310 145.520 340.500 146.310 ;
        RECT 342.460 145.660 342.670 146.670 ;
        RECT 351.720 146.660 353.620 146.670 ;
        RECT 355.350 145.930 355.530 146.680 ;
        RECT 341.310 145.520 341.580 145.530 ;
        RECT 340.310 145.310 341.580 145.520 ;
        RECT 341.310 145.100 341.580 145.310 ;
        RECT 341.310 144.470 341.560 145.100 ;
        RECT 342.460 144.650 342.660 145.660 ;
        RECT 350.270 145.630 355.530 145.930 ;
        RECT 340.520 144.020 341.560 144.470 ;
        RECT 340.500 142.570 341.460 143.020 ;
        RECT 341.210 142.520 341.460 142.570 ;
        RECT 342.470 142.520 342.660 144.650 ;
        RECT 341.210 142.320 342.660 142.520 ;
        RECT 346.190 143.990 346.450 145.190 ;
        RECT 346.190 143.480 346.440 143.990 ;
        RECT 348.080 143.980 348.340 145.190 ;
        RECT 350.470 144.080 350.720 145.630 ;
        RECT 348.080 143.820 348.470 143.980 ;
        RECT 348.070 143.690 348.470 143.820 ;
        RECT 351.170 143.690 351.430 145.300 ;
        RECT 353.720 144.230 354.020 145.280 ;
        RECT 354.470 144.680 354.770 145.630 ;
        RECT 354.970 144.730 355.270 144.780 ;
        RECT 354.970 144.380 355.870 144.730 ;
        RECT 357.580 144.600 357.800 144.610 ;
        RECT 357.580 144.410 371.260 144.600 ;
        RECT 357.580 144.280 357.800 144.410 ;
        RECT 346.690 143.480 346.980 143.640 ;
        RECT 348.070 143.630 348.330 143.690 ;
        RECT 346.190 143.290 346.980 143.480 ;
        RECT 346.190 143.090 346.440 143.290 ;
        RECT 346.690 143.180 346.980 143.290 ;
        RECT 348.080 143.090 348.330 143.630 ;
        RECT 351.160 143.630 351.430 143.690 ;
        RECT 352.710 143.970 354.020 144.230 ;
        RECT 356.120 143.980 357.800 144.280 ;
        RECT 356.120 143.970 357.780 143.980 ;
        RECT 352.710 143.630 353.020 143.970 ;
        RECT 348.720 143.100 350.360 143.490 ;
        RECT 351.160 143.340 353.020 143.630 ;
        RECT 351.160 143.330 351.470 143.340 ;
        RECT 352.710 143.330 353.020 143.340 ;
        RECT 346.190 142.490 346.480 143.090 ;
        RECT 348.080 142.490 348.370 143.090 ;
        RECT 337.380 142.090 337.640 142.240 ;
        RECT 341.210 142.230 341.460 142.320 ;
        RECT 335.800 138.400 336.070 138.810 ;
        RECT 262.370 138.090 263.560 138.100 ;
        RECT 264.550 138.090 265.740 138.100 ;
        RECT 266.770 138.090 267.960 138.100 ;
        RECT 268.950 138.090 270.140 138.110 ;
        RECT 260.160 138.080 270.140 138.090 ;
        RECT 256.770 138.060 257.960 138.070 ;
        RECT 259.050 138.060 270.140 138.080 ;
        RECT 245.540 137.270 245.830 137.430 ;
        RECT 246.920 137.420 247.180 137.480 ;
        RECT 245.040 137.080 245.830 137.270 ;
        RECT 245.040 136.880 245.290 137.080 ;
        RECT 245.540 136.970 245.830 137.080 ;
        RECT 246.930 136.880 247.180 137.420 ;
        RECT 250.010 137.420 250.280 137.480 ;
        RECT 251.560 137.760 252.870 138.020 ;
        RECT 254.930 137.830 270.140 138.060 ;
        RECT 254.930 137.820 269.090 137.830 ;
        RECT 254.930 137.810 262.460 137.820 ;
        RECT 263.470 137.810 264.660 137.820 ;
        RECT 265.620 137.810 266.810 137.820 ;
        RECT 267.900 137.810 269.090 137.820 ;
        RECT 254.930 137.800 260.240 137.810 ;
        RECT 254.930 137.790 259.100 137.800 ;
        RECT 254.930 137.780 256.820 137.790 ;
        RECT 257.910 137.780 259.100 137.790 ;
        RECT 254.930 137.770 255.650 137.780 ;
        RECT 251.560 137.420 251.870 137.760 ;
        RECT 247.570 136.890 249.210 137.280 ;
        RECT 250.010 137.130 251.870 137.420 ;
        RECT 250.010 137.120 250.320 137.130 ;
        RECT 251.560 137.120 251.870 137.130 ;
        RECT 240.150 136.770 240.800 136.780 ;
        RECT 240.150 136.440 240.450 136.770 ;
        RECT 239.430 135.990 240.450 136.440 ;
        RECT 245.040 136.280 245.330 136.880 ;
        RECT 246.930 136.280 247.220 136.880 ;
        RECT 240.150 135.980 240.450 135.990 ;
        RECT 249.270 135.670 249.570 136.670 ;
        RECT 250.020 136.070 250.320 137.120 ;
        RECT 252.620 136.020 252.870 137.760 ;
        RECT 253.320 135.670 253.580 137.220 ;
        RECT 335.800 137.110 336.050 138.400 ;
        RECT 330.830 136.810 336.080 137.110 ;
        RECT 249.220 135.660 254.470 135.670 ;
        RECT 239.100 135.580 239.350 135.590 ;
        RECT 239.100 135.120 240.080 135.580 ;
        RECT 249.220 135.370 254.490 135.660 ;
        RECT 239.100 134.820 239.350 135.120 ;
        RECT 247.070 135.030 248.910 135.040 ;
        RECT 254.320 135.030 254.490 135.370 ;
        RECT 240.810 135.020 241.050 135.030 ;
        RECT 241.890 135.020 254.490 135.030 ;
        RECT 240.810 134.860 254.490 135.020 ;
        RECT 326.750 135.170 327.010 136.370 ;
        RECT 240.810 134.850 252.320 134.860 ;
        RECT 240.800 134.840 247.120 134.850 ;
        RECT 248.670 134.840 252.320 134.850 ;
        RECT 240.800 134.830 242.670 134.840 ;
        RECT 240.800 134.820 241.050 134.830 ;
        RECT 239.100 134.650 241.050 134.820 ;
        RECT 326.750 134.660 327.000 135.170 ;
        RECT 328.640 135.160 328.900 136.370 ;
        RECT 331.030 135.260 331.280 136.810 ;
        RECT 328.640 135.000 329.030 135.160 ;
        RECT 328.630 134.870 329.030 135.000 ;
        RECT 331.730 134.870 331.990 136.480 ;
        RECT 334.280 135.410 334.580 136.460 ;
        RECT 335.030 135.860 335.330 136.810 ;
        RECT 335.530 135.910 335.830 135.960 ;
        RECT 335.530 135.560 336.430 135.910 ;
        RECT 337.400 135.460 337.640 142.090 ;
        RECT 340.480 141.780 341.460 142.230 ;
        RECT 350.420 141.880 350.720 142.880 ;
        RECT 351.170 142.280 351.470 143.330 ;
        RECT 353.770 142.230 354.020 143.970 ;
        RECT 371.010 143.510 371.260 144.410 ;
        RECT 354.470 141.880 354.730 143.430 ;
        RECT 365.950 143.210 371.260 143.510 ;
        RECT 350.370 141.860 355.620 141.880 ;
        RECT 350.370 141.580 355.740 141.860 ;
        RECT 343.820 141.180 344.100 141.250 ;
        RECT 345.000 141.210 345.280 141.240 ;
        RECT 355.450 141.210 355.740 141.580 ;
        RECT 345.000 141.200 355.740 141.210 ;
        RECT 342.410 140.980 344.100 141.180 ;
        RECT 341.200 140.780 341.480 140.790 ;
        RECT 340.460 140.330 341.480 140.780 ;
        RECT 342.410 140.330 342.640 140.980 ;
        RECT 343.820 140.920 344.100 140.980 ;
        RECT 344.980 140.970 355.740 141.200 ;
        RECT 345.000 140.960 355.740 140.970 ;
        RECT 361.870 141.570 362.130 142.770 ;
        RECT 361.870 141.060 362.120 141.570 ;
        RECT 363.760 141.560 364.020 142.770 ;
        RECT 366.150 141.660 366.400 143.210 ;
        RECT 363.760 141.400 364.150 141.560 ;
        RECT 363.750 141.270 364.150 141.400 ;
        RECT 366.850 141.270 367.110 142.880 ;
        RECT 369.400 141.810 369.700 142.860 ;
        RECT 370.150 142.260 370.450 143.210 ;
        RECT 370.650 142.310 370.950 142.360 ;
        RECT 370.650 141.960 371.550 142.310 ;
        RECT 388.780 141.910 389.120 148.030 ;
        RECT 437.150 147.490 437.380 149.460 ;
        RECT 437.150 143.900 437.420 147.490 ;
        RECT 437.150 142.080 437.400 143.900 ;
        RECT 463.370 143.420 463.640 242.920 ;
        RECT 463.370 143.240 463.690 143.420 ;
        RECT 388.210 141.890 389.170 141.910 ;
        RECT 372.690 141.870 376.970 141.880 ;
        RECT 384.370 141.870 389.170 141.890 ;
        RECT 372.690 141.860 389.170 141.870 ;
        RECT 362.370 141.060 362.660 141.220 ;
        RECT 363.750 141.210 364.010 141.270 ;
        RECT 345.000 140.950 355.700 140.960 ;
        RECT 345.000 140.910 345.280 140.950 ;
        RECT 361.870 140.870 362.660 141.060 ;
        RECT 361.870 140.670 362.120 140.870 ;
        RECT 362.370 140.760 362.660 140.870 ;
        RECT 363.760 140.670 364.010 141.210 ;
        RECT 366.840 141.210 367.110 141.270 ;
        RECT 368.390 141.550 369.700 141.810 ;
        RECT 368.390 141.210 368.700 141.550 ;
        RECT 364.400 140.680 366.040 141.070 ;
        RECT 366.840 140.920 368.700 141.210 ;
        RECT 366.840 140.910 367.150 140.920 ;
        RECT 368.390 140.910 368.700 140.920 ;
        RECT 343.800 140.350 344.070 140.430 ;
        RECT 341.200 140.120 342.640 140.330 ;
        RECT 343.190 140.130 344.070 140.350 ;
        RECT 341.200 139.070 341.480 140.120 ;
        RECT 343.190 139.320 343.410 140.130 ;
        RECT 343.800 140.100 344.070 140.130 ;
        RECT 344.930 140.390 345.220 140.440 ;
        RECT 344.930 140.210 355.680 140.390 ;
        RECT 344.930 140.110 345.220 140.210 ;
        RECT 349.770 140.200 353.400 140.210 ;
        RECT 355.480 139.530 355.680 140.210 ;
        RECT 361.870 140.070 362.160 140.670 ;
        RECT 363.760 140.070 364.050 140.670 ;
        RECT 340.480 138.620 341.480 139.070 ;
        RECT 340.460 137.170 341.760 137.620 ;
        RECT 341.460 136.770 341.760 137.170 ;
        RECT 343.180 136.790 343.410 139.320 ;
        RECT 350.430 139.230 355.680 139.530 ;
        RECT 366.100 139.460 366.400 140.460 ;
        RECT 366.850 139.860 367.150 140.910 ;
        RECT 369.450 139.810 369.700 141.550 ;
        RECT 371.820 141.550 389.170 141.860 ;
        RECT 371.820 141.540 384.830 141.550 ;
        RECT 376.680 141.530 384.830 141.540 ;
        RECT 388.210 141.510 389.170 141.550 ;
        RECT 388.780 141.500 389.120 141.510 ;
        RECT 370.150 139.460 370.410 141.010 ;
        RECT 371.240 139.460 371.440 139.470 ;
        RECT 342.250 136.770 343.410 136.790 ;
        RECT 341.460 136.590 343.410 136.770 ;
        RECT 346.350 137.590 346.610 138.790 ;
        RECT 346.350 137.080 346.600 137.590 ;
        RECT 348.240 137.580 348.500 138.790 ;
        RECT 350.630 137.680 350.880 139.230 ;
        RECT 348.240 137.420 348.630 137.580 ;
        RECT 348.230 137.290 348.630 137.420 ;
        RECT 351.330 137.290 351.590 138.900 ;
        RECT 353.880 137.830 354.180 138.880 ;
        RECT 354.630 138.280 354.930 139.230 ;
        RECT 355.480 139.220 355.680 139.230 ;
        RECT 366.050 139.160 371.440 139.460 ;
        RECT 355.130 138.330 355.430 138.380 ;
        RECT 355.130 137.980 356.030 138.330 ;
        RECT 371.240 137.920 371.440 139.160 ;
        RECT 437.150 138.620 437.380 142.080 ;
        RECT 463.390 140.740 463.690 143.240 ;
        RECT 463.400 139.250 463.670 140.740 ;
        RECT 458.420 138.950 463.670 139.250 ;
        RECT 437.110 138.210 437.380 138.620 ;
        RECT 363.680 137.900 364.870 137.910 ;
        RECT 365.860 137.900 367.050 137.910 ;
        RECT 368.080 137.900 369.270 137.910 ;
        RECT 370.260 137.900 371.450 137.920 ;
        RECT 361.470 137.890 371.450 137.900 ;
        RECT 358.080 137.870 359.270 137.880 ;
        RECT 360.360 137.870 371.450 137.890 ;
        RECT 346.850 137.080 347.140 137.240 ;
        RECT 348.230 137.230 348.490 137.290 ;
        RECT 346.350 136.890 347.140 137.080 ;
        RECT 346.350 136.690 346.600 136.890 ;
        RECT 346.850 136.780 347.140 136.890 ;
        RECT 348.240 136.690 348.490 137.230 ;
        RECT 351.320 137.230 351.590 137.290 ;
        RECT 352.870 137.570 354.180 137.830 ;
        RECT 356.240 137.640 371.450 137.870 ;
        RECT 356.240 137.630 370.400 137.640 ;
        RECT 356.240 137.620 363.770 137.630 ;
        RECT 364.780 137.620 365.970 137.630 ;
        RECT 366.930 137.620 368.120 137.630 ;
        RECT 369.210 137.620 370.400 137.630 ;
        RECT 356.240 137.610 361.550 137.620 ;
        RECT 356.240 137.600 360.410 137.610 ;
        RECT 356.240 137.590 358.130 137.600 ;
        RECT 359.220 137.590 360.410 137.600 ;
        RECT 356.240 137.580 356.960 137.590 ;
        RECT 352.870 137.230 353.180 137.570 ;
        RECT 348.880 136.700 350.520 137.090 ;
        RECT 351.320 136.940 353.180 137.230 ;
        RECT 351.320 136.930 351.630 136.940 ;
        RECT 352.870 136.930 353.180 136.940 ;
        RECT 341.460 136.580 342.110 136.590 ;
        RECT 341.460 136.250 341.760 136.580 ;
        RECT 340.740 135.800 341.760 136.250 ;
        RECT 346.350 136.090 346.640 136.690 ;
        RECT 348.240 136.090 348.530 136.690 ;
        RECT 341.460 135.790 341.760 135.800 ;
        RECT 350.580 135.480 350.880 136.480 ;
        RECT 351.330 135.880 351.630 136.930 ;
        RECT 353.930 135.830 354.180 137.570 ;
        RECT 354.630 135.480 354.890 137.030 ;
        RECT 437.110 136.920 437.360 138.210 ;
        RECT 454.340 137.310 454.600 138.510 ;
        RECT 432.140 136.620 437.390 136.920 ;
        RECT 454.340 136.800 454.590 137.310 ;
        RECT 456.230 137.300 456.490 138.510 ;
        RECT 458.620 137.400 458.870 138.950 ;
        RECT 462.620 138.000 462.920 138.950 ;
        RECT 463.120 138.050 463.420 138.100 ;
        RECT 463.120 137.700 464.020 138.050 ;
        RECT 456.230 137.140 456.620 137.300 ;
        RECT 456.220 137.010 456.620 137.140 ;
        RECT 454.840 136.800 455.130 136.960 ;
        RECT 456.220 136.950 456.480 137.010 ;
        RECT 327.250 134.660 327.540 134.820 ;
        RECT 328.630 134.810 328.890 134.870 ;
        RECT 239.100 134.350 239.370 134.650 ;
        RECT 239.110 134.090 239.370 134.350 ;
        RECT 326.750 134.470 327.540 134.660 ;
        RECT 326.750 134.270 327.000 134.470 ;
        RECT 327.250 134.360 327.540 134.470 ;
        RECT 328.640 134.270 328.890 134.810 ;
        RECT 331.720 134.810 331.990 134.870 ;
        RECT 333.270 135.150 334.580 135.410 ;
        RECT 336.760 135.150 337.640 135.460 ;
        RECT 350.530 135.470 355.780 135.480 ;
        RECT 340.410 135.390 340.660 135.400 ;
        RECT 333.270 134.810 333.580 135.150 ;
        RECT 329.280 134.280 330.920 134.670 ;
        RECT 331.720 134.520 333.580 134.810 ;
        RECT 331.720 134.510 332.030 134.520 ;
        RECT 333.270 134.510 333.580 134.520 ;
        RECT 239.090 133.700 239.390 134.090 ;
        RECT 239.080 133.300 239.390 133.700 ;
        RECT 326.750 133.670 327.040 134.270 ;
        RECT 328.640 133.670 328.930 134.270 ;
        RECT 239.080 132.970 239.370 133.300 ;
        RECT 330.980 133.060 331.280 134.060 ;
        RECT 331.730 133.460 332.030 134.510 ;
        RECT 334.330 133.410 334.580 135.150 ;
        RECT 340.410 134.930 341.390 135.390 ;
        RECT 350.530 135.180 355.800 135.470 ;
        RECT 340.410 134.630 340.660 134.930 ;
        RECT 348.380 134.840 350.220 134.850 ;
        RECT 355.630 134.840 355.800 135.180 ;
        RECT 342.120 134.830 342.360 134.840 ;
        RECT 343.200 134.830 355.800 134.840 ;
        RECT 342.120 134.670 355.800 134.830 ;
        RECT 428.060 134.980 428.320 136.180 ;
        RECT 342.120 134.660 353.630 134.670 ;
        RECT 342.110 134.650 348.430 134.660 ;
        RECT 349.980 134.650 353.630 134.660 ;
        RECT 342.110 134.640 343.980 134.650 ;
        RECT 342.110 134.630 342.360 134.640 ;
        RECT 335.030 133.060 335.290 134.610 ;
        RECT 340.410 134.460 342.360 134.630 ;
        RECT 428.060 134.470 428.310 134.980 ;
        RECT 429.950 134.970 430.210 136.180 ;
        RECT 432.340 135.070 432.590 136.620 ;
        RECT 429.950 134.810 430.340 134.970 ;
        RECT 429.940 134.680 430.340 134.810 ;
        RECT 433.040 134.680 433.300 136.290 ;
        RECT 435.590 135.220 435.890 136.270 ;
        RECT 436.340 135.670 436.640 136.620 ;
        RECT 454.340 136.610 455.130 136.800 ;
        RECT 454.340 136.410 454.590 136.610 ;
        RECT 454.840 136.500 455.130 136.610 ;
        RECT 456.230 136.410 456.480 136.950 ;
        RECT 456.870 136.420 458.510 136.810 ;
        RECT 454.340 135.810 454.630 136.410 ;
        RECT 456.230 135.810 456.520 136.410 ;
        RECT 436.840 135.720 437.140 135.770 ;
        RECT 436.840 135.370 437.740 135.720 ;
        RECT 445.810 135.270 449.640 135.290 ;
        RECT 428.560 134.470 428.850 134.630 ;
        RECT 429.940 134.620 430.200 134.680 ;
        RECT 340.410 134.160 340.680 134.460 ;
        RECT 340.420 133.900 340.680 134.160 ;
        RECT 428.060 134.280 428.850 134.470 ;
        RECT 428.060 134.080 428.310 134.280 ;
        RECT 428.560 134.170 428.850 134.280 ;
        RECT 429.950 134.080 430.200 134.620 ;
        RECT 433.030 134.620 433.300 134.680 ;
        RECT 434.580 134.960 435.890 135.220 ;
        RECT 438.070 134.990 449.650 135.270 ;
        RECT 458.570 135.200 458.870 136.200 ;
        RECT 462.620 135.200 462.880 136.750 ;
        RECT 463.670 135.200 463.870 135.230 ;
        RECT 438.070 134.970 446.260 134.990 ;
        RECT 438.070 134.960 438.900 134.970 ;
        RECT 434.580 134.620 434.890 134.960 ;
        RECT 430.590 134.090 432.230 134.480 ;
        RECT 433.030 134.330 434.890 134.620 ;
        RECT 433.030 134.320 433.340 134.330 ;
        RECT 434.580 134.320 434.890 134.330 ;
        RECT 340.400 133.510 340.700 133.900 ;
        RECT 340.390 133.110 340.700 133.510 ;
        RECT 428.060 133.480 428.350 134.080 ;
        RECT 429.950 133.480 430.240 134.080 ;
        RECT 336.120 133.060 336.670 133.080 ;
        RECT 239.060 132.310 239.410 132.970 ;
        RECT 330.930 132.770 336.670 133.060 ;
        RECT 340.390 132.780 340.680 133.110 ;
        RECT 432.290 132.870 432.590 133.870 ;
        RECT 433.040 133.270 433.340 134.320 ;
        RECT 435.640 133.220 435.890 134.960 ;
        RECT 436.340 132.870 436.600 134.420 ;
        RECT 449.450 133.030 449.650 134.990 ;
        RECT 458.520 134.900 463.870 135.200 ;
        RECT 463.670 133.050 463.870 134.900 ;
        RECT 471.640 134.960 471.900 136.160 ;
        RECT 471.640 134.450 471.890 134.960 ;
        RECT 473.530 134.950 473.790 136.160 ;
        RECT 480.420 135.700 480.720 135.750 ;
        RECT 480.420 135.350 481.320 135.700 ;
        RECT 473.530 134.790 473.920 134.950 ;
        RECT 473.520 134.660 473.920 134.790 ;
        RECT 472.140 134.450 472.430 134.610 ;
        RECT 473.520 134.600 473.780 134.660 ;
        RECT 471.640 134.260 472.430 134.450 ;
        RECT 471.640 134.060 471.890 134.260 ;
        RECT 472.140 134.150 472.430 134.260 ;
        RECT 473.530 134.060 473.780 134.600 ;
        RECT 474.170 134.070 475.810 134.460 ;
        RECT 471.640 133.460 471.930 134.060 ;
        RECT 473.530 133.460 473.820 134.060 ;
        RECT 457.210 133.030 463.900 133.050 ;
        RECT 437.430 132.870 437.980 132.890 ;
        RECT 330.930 132.760 336.180 132.770 ;
        RECT 237.790 131.970 239.410 132.310 ;
        RECT 237.790 131.120 238.240 131.970 ;
        RECT 239.060 131.960 239.410 131.970 ;
        RECT 238.650 130.940 239.110 131.770 ;
        RECT 241.200 131.230 250.470 131.240 ;
        RECT 252.350 131.230 254.270 131.240 ;
        RECT 240.030 130.940 240.310 131.080 ;
        RECT 238.650 130.830 240.310 130.940 ;
        RECT 238.660 130.630 240.310 130.830 ;
        RECT 241.200 131.040 254.270 131.230 ;
        RECT 241.200 131.030 253.560 131.040 ;
        RECT 238.660 130.620 240.330 130.630 ;
        RECT 240.030 130.400 240.330 130.620 ;
        RECT 240.040 130.230 240.330 130.400 ;
        RECT 240.050 129.430 240.310 130.230 ;
        RECT 241.200 130.020 241.410 131.030 ;
        RECT 250.460 131.020 252.360 131.030 ;
        RECT 254.090 130.290 254.270 131.040 ;
        RECT 240.050 128.830 240.300 129.430 ;
        RECT 241.200 129.010 241.400 130.020 ;
        RECT 249.010 129.990 254.270 130.290 ;
        RECT 239.260 128.380 240.300 128.830 ;
        RECT 239.240 126.930 240.200 127.380 ;
        RECT 239.950 126.880 240.200 126.930 ;
        RECT 241.210 126.880 241.400 129.010 ;
        RECT 239.950 126.680 241.400 126.880 ;
        RECT 244.930 128.350 245.190 129.550 ;
        RECT 244.930 127.840 245.180 128.350 ;
        RECT 246.820 128.340 247.080 129.550 ;
        RECT 249.210 128.440 249.460 129.990 ;
        RECT 246.820 128.180 247.210 128.340 ;
        RECT 246.810 128.050 247.210 128.180 ;
        RECT 249.910 128.050 250.170 129.660 ;
        RECT 252.460 128.590 252.760 129.640 ;
        RECT 253.210 129.040 253.510 129.990 ;
        RECT 253.710 129.090 254.010 129.140 ;
        RECT 253.710 128.740 254.610 129.090 ;
        RECT 256.320 128.960 256.540 128.970 ;
        RECT 256.320 128.770 270.000 128.960 ;
        RECT 256.320 128.640 256.540 128.770 ;
        RECT 245.430 127.840 245.720 128.000 ;
        RECT 246.810 127.990 247.070 128.050 ;
        RECT 244.930 127.650 245.720 127.840 ;
        RECT 244.930 127.450 245.180 127.650 ;
        RECT 245.430 127.540 245.720 127.650 ;
        RECT 246.820 127.450 247.070 127.990 ;
        RECT 249.900 127.990 250.170 128.050 ;
        RECT 251.450 128.330 252.760 128.590 ;
        RECT 254.860 128.340 256.540 128.640 ;
        RECT 254.860 128.330 256.520 128.340 ;
        RECT 251.450 127.990 251.760 128.330 ;
        RECT 247.460 127.460 249.100 127.850 ;
        RECT 249.900 127.700 251.760 127.990 ;
        RECT 249.900 127.690 250.210 127.700 ;
        RECT 251.450 127.690 251.760 127.700 ;
        RECT 244.930 126.850 245.220 127.450 ;
        RECT 246.820 126.850 247.110 127.450 ;
        RECT 239.950 126.590 240.200 126.680 ;
        RECT 239.220 126.140 240.200 126.590 ;
        RECT 249.160 126.240 249.460 127.240 ;
        RECT 249.910 126.640 250.210 127.690 ;
        RECT 252.510 126.590 252.760 128.330 ;
        RECT 269.750 127.870 270.000 128.770 ;
        RECT 253.210 126.240 253.470 127.790 ;
        RECT 264.690 127.570 270.000 127.870 ;
        RECT 249.110 126.220 254.360 126.240 ;
        RECT 249.110 125.940 254.480 126.220 ;
        RECT 242.560 125.540 242.840 125.610 ;
        RECT 243.740 125.570 244.020 125.600 ;
        RECT 254.190 125.570 254.480 125.940 ;
        RECT 243.740 125.560 254.480 125.570 ;
        RECT 241.150 125.340 242.840 125.540 ;
        RECT 239.940 125.140 240.220 125.150 ;
        RECT 239.200 124.690 240.220 125.140 ;
        RECT 241.150 124.690 241.380 125.340 ;
        RECT 242.560 125.280 242.840 125.340 ;
        RECT 243.720 125.330 254.480 125.560 ;
        RECT 243.740 125.320 254.480 125.330 ;
        RECT 260.610 125.930 260.870 127.130 ;
        RECT 260.610 125.420 260.860 125.930 ;
        RECT 262.500 125.920 262.760 127.130 ;
        RECT 264.890 126.020 265.140 127.570 ;
        RECT 262.500 125.760 262.890 125.920 ;
        RECT 262.490 125.630 262.890 125.760 ;
        RECT 265.590 125.630 265.850 127.240 ;
        RECT 268.140 126.170 268.440 127.220 ;
        RECT 268.890 126.620 269.190 127.570 ;
        RECT 269.390 126.670 269.690 126.720 ;
        RECT 269.390 126.320 270.290 126.670 ;
        RECT 283.050 126.270 287.520 126.300 ;
        RECT 272.110 126.240 287.520 126.270 ;
        RECT 271.440 126.220 287.520 126.240 ;
        RECT 261.110 125.420 261.400 125.580 ;
        RECT 262.490 125.570 262.750 125.630 ;
        RECT 243.740 125.310 254.440 125.320 ;
        RECT 243.740 125.270 244.020 125.310 ;
        RECT 260.610 125.230 261.400 125.420 ;
        RECT 260.610 125.030 260.860 125.230 ;
        RECT 261.110 125.120 261.400 125.230 ;
        RECT 262.500 125.030 262.750 125.570 ;
        RECT 265.580 125.570 265.850 125.630 ;
        RECT 267.130 125.910 268.440 126.170 ;
        RECT 267.130 125.570 267.440 125.910 ;
        RECT 263.140 125.040 264.780 125.430 ;
        RECT 265.580 125.280 267.440 125.570 ;
        RECT 265.580 125.270 265.890 125.280 ;
        RECT 267.130 125.270 267.440 125.280 ;
        RECT 242.540 124.710 242.810 124.790 ;
        RECT 239.940 124.480 241.380 124.690 ;
        RECT 241.930 124.490 242.810 124.710 ;
        RECT 239.940 123.430 240.220 124.480 ;
        RECT 241.930 123.680 242.150 124.490 ;
        RECT 242.540 124.460 242.810 124.490 ;
        RECT 243.670 124.750 243.960 124.800 ;
        RECT 243.670 124.570 254.420 124.750 ;
        RECT 243.670 124.470 243.960 124.570 ;
        RECT 248.510 124.560 252.140 124.570 ;
        RECT 254.220 123.890 254.420 124.570 ;
        RECT 260.610 124.430 260.900 125.030 ;
        RECT 262.500 124.430 262.790 125.030 ;
        RECT 239.220 122.980 240.220 123.430 ;
        RECT 239.200 121.530 240.500 121.980 ;
        RECT 240.200 121.130 240.500 121.530 ;
        RECT 241.920 121.150 242.150 123.680 ;
        RECT 249.170 123.590 254.420 123.890 ;
        RECT 264.840 123.820 265.140 124.820 ;
        RECT 265.590 124.220 265.890 125.270 ;
        RECT 268.190 124.170 268.440 125.910 ;
        RECT 270.560 125.900 287.520 126.220 ;
        RECT 271.440 125.890 287.520 125.900 ;
        RECT 271.440 125.860 283.420 125.890 ;
        RECT 271.440 125.850 272.330 125.860 ;
        RECT 268.890 123.820 269.150 125.370 ;
        RECT 269.980 123.820 270.180 123.830 ;
        RECT 240.990 121.130 242.150 121.150 ;
        RECT 240.200 120.950 242.150 121.130 ;
        RECT 245.090 121.950 245.350 123.150 ;
        RECT 245.090 121.440 245.340 121.950 ;
        RECT 246.980 121.940 247.240 123.150 ;
        RECT 249.370 122.040 249.620 123.590 ;
        RECT 246.980 121.780 247.370 121.940 ;
        RECT 246.970 121.650 247.370 121.780 ;
        RECT 250.070 121.650 250.330 123.260 ;
        RECT 252.620 122.190 252.920 123.240 ;
        RECT 253.370 122.640 253.670 123.590 ;
        RECT 254.220 123.580 254.420 123.590 ;
        RECT 264.790 123.520 270.180 123.820 ;
        RECT 253.870 122.690 254.170 122.740 ;
        RECT 253.870 122.340 254.770 122.690 ;
        RECT 269.980 122.280 270.180 123.520 ;
        RECT 287.140 122.320 287.500 125.890 ;
        RECT 262.420 122.260 263.610 122.270 ;
        RECT 264.600 122.260 265.790 122.270 ;
        RECT 266.820 122.260 268.010 122.270 ;
        RECT 269.000 122.260 270.190 122.280 ;
        RECT 260.210 122.250 270.190 122.260 ;
        RECT 256.820 122.230 258.010 122.240 ;
        RECT 259.100 122.230 270.190 122.250 ;
        RECT 245.590 121.440 245.880 121.600 ;
        RECT 246.970 121.590 247.230 121.650 ;
        RECT 245.090 121.250 245.880 121.440 ;
        RECT 245.090 121.050 245.340 121.250 ;
        RECT 245.590 121.140 245.880 121.250 ;
        RECT 246.980 121.050 247.230 121.590 ;
        RECT 250.060 121.590 250.330 121.650 ;
        RECT 251.610 121.930 252.920 122.190 ;
        RECT 254.980 122.000 270.190 122.230 ;
        RECT 282.270 122.020 287.520 122.320 ;
        RECT 254.980 121.990 269.140 122.000 ;
        RECT 254.980 121.980 262.510 121.990 ;
        RECT 263.520 121.980 264.710 121.990 ;
        RECT 265.670 121.980 266.860 121.990 ;
        RECT 267.950 121.980 269.140 121.990 ;
        RECT 254.980 121.970 260.290 121.980 ;
        RECT 254.980 121.960 259.150 121.970 ;
        RECT 254.980 121.950 256.870 121.960 ;
        RECT 257.960 121.950 259.150 121.960 ;
        RECT 254.980 121.940 255.700 121.950 ;
        RECT 251.610 121.590 251.920 121.930 ;
        RECT 247.620 121.060 249.260 121.450 ;
        RECT 250.060 121.300 251.920 121.590 ;
        RECT 250.060 121.290 250.370 121.300 ;
        RECT 251.610 121.290 251.920 121.300 ;
        RECT 240.200 120.940 240.850 120.950 ;
        RECT 240.200 120.610 240.500 120.940 ;
        RECT 239.480 120.160 240.500 120.610 ;
        RECT 245.090 120.450 245.380 121.050 ;
        RECT 246.980 120.450 247.270 121.050 ;
        RECT 240.200 120.150 240.500 120.160 ;
        RECT 249.320 119.840 249.620 120.840 ;
        RECT 250.070 120.240 250.370 121.290 ;
        RECT 252.670 120.190 252.920 121.930 ;
        RECT 253.370 119.840 253.630 121.390 ;
        RECT 278.190 120.380 278.450 121.580 ;
        RECT 278.190 119.870 278.440 120.380 ;
        RECT 280.080 120.370 280.340 121.580 ;
        RECT 282.470 120.470 282.720 122.020 ;
        RECT 280.080 120.210 280.470 120.370 ;
        RECT 280.070 120.080 280.470 120.210 ;
        RECT 283.170 120.080 283.430 121.690 ;
        RECT 285.720 120.620 286.020 121.670 ;
        RECT 286.470 121.070 286.770 122.020 ;
        RECT 286.970 121.120 287.270 121.170 ;
        RECT 286.970 120.770 287.870 121.120 ;
        RECT 278.690 119.870 278.980 120.030 ;
        RECT 280.070 120.020 280.330 120.080 ;
        RECT 249.270 119.830 254.520 119.840 ;
        RECT 239.150 119.750 239.400 119.760 ;
        RECT 239.150 119.290 240.130 119.750 ;
        RECT 249.270 119.540 254.540 119.830 ;
        RECT 239.150 118.990 239.400 119.290 ;
        RECT 247.120 119.200 248.960 119.210 ;
        RECT 254.370 119.200 254.540 119.540 ;
        RECT 240.860 119.190 241.100 119.200 ;
        RECT 241.940 119.190 254.540 119.200 ;
        RECT 240.860 119.030 254.540 119.190 ;
        RECT 278.190 119.680 278.980 119.870 ;
        RECT 278.190 119.480 278.440 119.680 ;
        RECT 278.690 119.570 278.980 119.680 ;
        RECT 280.080 119.480 280.330 120.020 ;
        RECT 283.160 120.020 283.430 120.080 ;
        RECT 284.710 120.360 286.020 120.620 ;
        RECT 288.080 120.660 289.750 120.690 ;
        RECT 304.830 120.660 305.080 120.670 ;
        RECT 288.080 120.390 305.080 120.660 ;
        RECT 288.080 120.380 301.580 120.390 ;
        RECT 289.360 120.360 301.580 120.380 ;
        RECT 284.710 120.020 285.020 120.360 ;
        RECT 280.720 119.490 282.360 119.880 ;
        RECT 283.160 119.730 285.020 120.020 ;
        RECT 283.160 119.720 283.470 119.730 ;
        RECT 284.710 119.720 285.020 119.730 ;
        RECT 240.860 119.020 252.370 119.030 ;
        RECT 240.850 119.010 247.170 119.020 ;
        RECT 248.720 119.010 252.370 119.020 ;
        RECT 240.850 119.000 242.720 119.010 ;
        RECT 240.850 118.990 241.100 119.000 ;
        RECT 239.150 118.820 241.100 118.990 ;
        RECT 278.190 118.880 278.480 119.480 ;
        RECT 280.080 118.880 280.370 119.480 ;
        RECT 239.150 118.600 239.400 118.820 ;
        RECT 239.150 118.430 240.190 118.600 ;
        RECT 240.000 117.570 240.190 118.430 ;
        RECT 282.420 118.270 282.720 119.270 ;
        RECT 283.170 118.670 283.470 119.720 ;
        RECT 285.770 118.620 286.020 120.360 ;
        RECT 286.470 118.270 286.730 119.820 ;
        RECT 287.350 118.270 287.690 118.340 ;
        RECT 282.370 117.970 287.690 118.270 ;
        RECT 239.210 117.130 240.190 117.570 ;
        RECT 239.210 117.120 240.160 117.130 ;
        RECT 241.030 116.810 250.300 116.820 ;
        RECT 252.180 116.810 254.100 116.820 ;
        RECT 238.880 116.710 239.070 116.720 ;
        RECT 238.880 116.250 239.860 116.710 ;
        RECT 241.030 116.620 254.100 116.810 ;
        RECT 241.030 116.610 253.390 116.620 ;
        RECT 238.880 115.460 239.070 116.250 ;
        RECT 241.030 115.600 241.240 116.610 ;
        RECT 250.290 116.600 252.190 116.610 ;
        RECT 253.920 115.870 254.100 116.620 ;
        RECT 239.880 115.460 240.150 115.470 ;
        RECT 238.880 115.250 240.150 115.460 ;
        RECT 239.880 115.040 240.150 115.250 ;
        RECT 239.880 114.410 240.130 115.040 ;
        RECT 241.030 114.590 241.230 115.600 ;
        RECT 248.840 115.570 254.100 115.870 ;
        RECT 239.090 113.960 240.130 114.410 ;
        RECT 239.070 112.510 240.030 112.960 ;
        RECT 239.780 112.460 240.030 112.510 ;
        RECT 241.040 112.460 241.230 114.590 ;
        RECT 239.780 112.260 241.230 112.460 ;
        RECT 244.760 113.930 245.020 115.130 ;
        RECT 244.760 113.420 245.010 113.930 ;
        RECT 246.650 113.920 246.910 115.130 ;
        RECT 249.040 114.020 249.290 115.570 ;
        RECT 246.650 113.760 247.040 113.920 ;
        RECT 246.640 113.630 247.040 113.760 ;
        RECT 249.740 113.630 250.000 115.240 ;
        RECT 252.290 114.170 252.590 115.220 ;
        RECT 253.040 114.620 253.340 115.570 ;
        RECT 253.540 114.670 253.840 114.720 ;
        RECT 253.540 114.320 254.440 114.670 ;
        RECT 256.150 114.540 256.370 114.550 ;
        RECT 256.150 114.350 269.830 114.540 ;
        RECT 256.150 114.220 256.370 114.350 ;
        RECT 245.260 113.420 245.550 113.580 ;
        RECT 246.640 113.570 246.900 113.630 ;
        RECT 244.760 113.230 245.550 113.420 ;
        RECT 244.760 113.030 245.010 113.230 ;
        RECT 245.260 113.120 245.550 113.230 ;
        RECT 246.650 113.030 246.900 113.570 ;
        RECT 249.730 113.570 250.000 113.630 ;
        RECT 251.280 113.910 252.590 114.170 ;
        RECT 254.690 113.920 256.370 114.220 ;
        RECT 254.690 113.910 256.350 113.920 ;
        RECT 251.280 113.570 251.590 113.910 ;
        RECT 247.290 113.040 248.930 113.430 ;
        RECT 249.730 113.280 251.590 113.570 ;
        RECT 249.730 113.270 250.040 113.280 ;
        RECT 251.280 113.270 251.590 113.280 ;
        RECT 244.760 112.430 245.050 113.030 ;
        RECT 246.650 112.430 246.940 113.030 ;
        RECT 239.780 112.170 240.030 112.260 ;
        RECT 239.050 111.720 240.030 112.170 ;
        RECT 248.990 111.820 249.290 112.820 ;
        RECT 249.740 112.220 250.040 113.270 ;
        RECT 252.340 112.170 252.590 113.910 ;
        RECT 269.580 113.450 269.830 114.350 ;
        RECT 253.040 111.820 253.300 113.370 ;
        RECT 264.520 113.150 269.830 113.450 ;
        RECT 248.940 111.800 254.190 111.820 ;
        RECT 248.940 111.520 254.310 111.800 ;
        RECT 242.390 111.120 242.670 111.190 ;
        RECT 243.570 111.150 243.850 111.180 ;
        RECT 254.020 111.150 254.310 111.520 ;
        RECT 243.570 111.140 254.310 111.150 ;
        RECT 240.980 110.920 242.670 111.120 ;
        RECT 239.770 110.720 240.050 110.730 ;
        RECT 239.030 110.270 240.050 110.720 ;
        RECT 240.980 110.270 241.210 110.920 ;
        RECT 242.390 110.860 242.670 110.920 ;
        RECT 243.550 110.910 254.310 111.140 ;
        RECT 243.570 110.900 254.310 110.910 ;
        RECT 260.440 111.510 260.700 112.710 ;
        RECT 260.440 111.000 260.690 111.510 ;
        RECT 262.330 111.500 262.590 112.710 ;
        RECT 264.720 111.600 264.970 113.150 ;
        RECT 262.330 111.340 262.720 111.500 ;
        RECT 262.320 111.210 262.720 111.340 ;
        RECT 265.420 111.210 265.680 112.820 ;
        RECT 267.970 111.750 268.270 112.800 ;
        RECT 268.720 112.200 269.020 113.150 ;
        RECT 269.220 112.250 269.520 112.300 ;
        RECT 269.220 111.900 270.120 112.250 ;
        RECT 287.350 111.850 287.690 117.970 ;
        RECT 286.780 111.830 287.740 111.850 ;
        RECT 271.260 111.810 275.540 111.820 ;
        RECT 282.940 111.810 287.740 111.830 ;
        RECT 271.260 111.800 287.740 111.810 ;
        RECT 260.940 111.000 261.230 111.160 ;
        RECT 262.320 111.150 262.580 111.210 ;
        RECT 243.570 110.890 254.270 110.900 ;
        RECT 243.570 110.850 243.850 110.890 ;
        RECT 260.440 110.810 261.230 111.000 ;
        RECT 260.440 110.610 260.690 110.810 ;
        RECT 260.940 110.700 261.230 110.810 ;
        RECT 262.330 110.610 262.580 111.150 ;
        RECT 265.410 111.150 265.680 111.210 ;
        RECT 266.960 111.490 268.270 111.750 ;
        RECT 266.960 111.150 267.270 111.490 ;
        RECT 262.970 110.620 264.610 111.010 ;
        RECT 265.410 110.860 267.270 111.150 ;
        RECT 265.410 110.850 265.720 110.860 ;
        RECT 266.960 110.850 267.270 110.860 ;
        RECT 242.370 110.290 242.640 110.370 ;
        RECT 239.770 110.060 241.210 110.270 ;
        RECT 241.760 110.070 242.640 110.290 ;
        RECT 239.770 109.010 240.050 110.060 ;
        RECT 241.760 109.260 241.980 110.070 ;
        RECT 242.370 110.040 242.640 110.070 ;
        RECT 243.500 110.330 243.790 110.380 ;
        RECT 243.500 110.150 254.250 110.330 ;
        RECT 243.500 110.050 243.790 110.150 ;
        RECT 248.340 110.140 251.970 110.150 ;
        RECT 254.050 109.470 254.250 110.150 ;
        RECT 260.440 110.010 260.730 110.610 ;
        RECT 262.330 110.010 262.620 110.610 ;
        RECT 239.050 108.560 240.050 109.010 ;
        RECT 239.030 107.110 240.330 107.560 ;
        RECT 240.030 106.710 240.330 107.110 ;
        RECT 241.750 106.730 241.980 109.260 ;
        RECT 249.000 109.170 254.250 109.470 ;
        RECT 264.670 109.400 264.970 110.400 ;
        RECT 265.420 109.800 265.720 110.850 ;
        RECT 268.020 109.750 268.270 111.490 ;
        RECT 270.390 111.490 287.740 111.800 ;
        RECT 270.390 111.480 283.400 111.490 ;
        RECT 275.250 111.470 283.400 111.480 ;
        RECT 286.780 111.450 287.740 111.490 ;
        RECT 287.350 111.440 287.690 111.450 ;
        RECT 268.720 109.400 268.980 110.950 ;
        RECT 269.810 109.400 270.010 109.410 ;
        RECT 240.820 106.710 241.980 106.730 ;
        RECT 240.030 106.530 241.980 106.710 ;
        RECT 244.920 107.530 245.180 108.730 ;
        RECT 244.920 107.020 245.170 107.530 ;
        RECT 246.810 107.520 247.070 108.730 ;
        RECT 249.200 107.620 249.450 109.170 ;
        RECT 246.810 107.360 247.200 107.520 ;
        RECT 246.800 107.230 247.200 107.360 ;
        RECT 249.900 107.230 250.160 108.840 ;
        RECT 252.450 107.770 252.750 108.820 ;
        RECT 253.200 108.220 253.500 109.170 ;
        RECT 254.050 109.160 254.250 109.170 ;
        RECT 264.620 109.100 270.010 109.400 ;
        RECT 253.700 108.270 254.000 108.320 ;
        RECT 253.700 107.920 254.600 108.270 ;
        RECT 269.810 107.860 270.010 109.100 ;
        RECT 262.250 107.840 263.440 107.850 ;
        RECT 264.430 107.840 265.620 107.850 ;
        RECT 266.650 107.840 267.840 107.850 ;
        RECT 268.830 107.840 270.020 107.860 ;
        RECT 260.040 107.830 270.020 107.840 ;
        RECT 256.650 107.810 257.840 107.820 ;
        RECT 258.930 107.810 270.020 107.830 ;
        RECT 245.420 107.020 245.710 107.180 ;
        RECT 246.800 107.170 247.060 107.230 ;
        RECT 244.920 106.830 245.710 107.020 ;
        RECT 244.920 106.630 245.170 106.830 ;
        RECT 245.420 106.720 245.710 106.830 ;
        RECT 246.810 106.630 247.060 107.170 ;
        RECT 249.890 107.170 250.160 107.230 ;
        RECT 251.440 107.510 252.750 107.770 ;
        RECT 254.810 107.580 270.020 107.810 ;
        RECT 254.810 107.570 268.970 107.580 ;
        RECT 254.810 107.560 262.340 107.570 ;
        RECT 263.350 107.560 264.540 107.570 ;
        RECT 265.500 107.560 266.690 107.570 ;
        RECT 267.780 107.560 268.970 107.570 ;
        RECT 254.810 107.550 260.120 107.560 ;
        RECT 254.810 107.540 258.980 107.550 ;
        RECT 254.810 107.530 256.700 107.540 ;
        RECT 257.790 107.530 258.980 107.540 ;
        RECT 254.810 107.520 255.530 107.530 ;
        RECT 251.440 107.170 251.750 107.510 ;
        RECT 247.450 106.640 249.090 107.030 ;
        RECT 249.890 106.880 251.750 107.170 ;
        RECT 249.890 106.870 250.200 106.880 ;
        RECT 251.440 106.870 251.750 106.880 ;
        RECT 240.030 106.520 240.680 106.530 ;
        RECT 240.030 106.190 240.330 106.520 ;
        RECT 239.310 105.740 240.330 106.190 ;
        RECT 244.920 106.030 245.210 106.630 ;
        RECT 246.810 106.030 247.100 106.630 ;
        RECT 240.030 105.730 240.330 105.740 ;
        RECT 249.150 105.420 249.450 106.420 ;
        RECT 249.900 105.820 250.200 106.870 ;
        RECT 252.500 105.770 252.750 107.510 ;
        RECT 304.830 107.250 305.090 120.390 ;
        RECT 304.820 107.130 305.090 107.250 ;
        RECT 253.200 105.420 253.460 106.970 ;
        RECT 304.820 106.300 305.080 107.130 ;
        RECT 299.800 106.000 305.080 106.300 ;
        RECT 249.100 105.410 254.350 105.420 ;
        RECT 238.980 105.330 239.230 105.340 ;
        RECT 238.980 104.870 239.960 105.330 ;
        RECT 249.100 105.120 254.370 105.410 ;
        RECT 238.980 104.570 239.230 104.870 ;
        RECT 246.950 104.780 248.790 104.790 ;
        RECT 254.200 104.780 254.370 105.120 ;
        RECT 240.690 104.770 240.930 104.780 ;
        RECT 241.770 104.770 254.370 104.780 ;
        RECT 240.690 104.610 254.370 104.770 ;
        RECT 240.690 104.600 252.200 104.610 ;
        RECT 240.680 104.590 247.000 104.600 ;
        RECT 248.550 104.590 252.200 104.600 ;
        RECT 240.680 104.580 242.550 104.590 ;
        RECT 240.680 104.570 240.930 104.580 ;
        RECT 238.980 104.400 240.930 104.570 ;
        RECT 238.980 104.100 239.250 104.400 ;
        RECT 238.990 103.840 239.250 104.100 ;
        RECT 295.720 104.360 295.980 105.560 ;
        RECT 295.720 103.850 295.970 104.360 ;
        RECT 297.610 104.350 297.870 105.560 ;
        RECT 300.000 104.450 300.250 106.000 ;
        RECT 297.610 104.190 298.000 104.350 ;
        RECT 297.600 104.060 298.000 104.190 ;
        RECT 300.700 104.060 300.960 105.670 ;
        RECT 303.250 104.600 303.550 105.650 ;
        RECT 304.000 105.050 304.300 106.000 ;
        RECT 304.500 105.100 304.800 105.150 ;
        RECT 304.500 104.750 305.400 105.100 ;
        RECT 296.220 103.850 296.510 104.010 ;
        RECT 297.600 104.000 297.860 104.060 ;
        RECT 238.970 103.450 239.270 103.840 ;
        RECT 295.720 103.660 296.510 103.850 ;
        RECT 295.720 103.460 295.970 103.660 ;
        RECT 296.220 103.550 296.510 103.660 ;
        RECT 297.610 103.460 297.860 104.000 ;
        RECT 300.690 104.000 300.960 104.060 ;
        RECT 302.240 104.340 303.550 104.600 ;
        RECT 305.670 104.540 306.450 104.640 ;
        RECT 305.670 104.370 319.250 104.540 ;
        RECT 305.670 104.360 319.240 104.370 ;
        RECT 305.670 104.340 306.450 104.360 ;
        RECT 302.240 104.000 302.550 104.340 ;
        RECT 298.250 103.470 299.890 103.860 ;
        RECT 300.690 103.710 302.550 104.000 ;
        RECT 300.690 103.700 301.000 103.710 ;
        RECT 302.240 103.700 302.550 103.710 ;
        RECT 238.970 103.220 240.460 103.450 ;
        RECT 240.210 102.290 240.460 103.220 ;
        RECT 295.720 102.860 296.010 103.460 ;
        RECT 297.610 102.860 297.900 103.460 ;
        RECT 239.410 101.830 240.460 102.290 ;
        RECT 299.950 102.250 300.250 103.250 ;
        RECT 300.700 102.650 301.000 103.700 ;
        RECT 303.300 102.600 303.550 104.340 ;
        RECT 304.000 102.250 304.260 103.800 ;
        RECT 299.900 101.950 305.170 102.250 ;
        RECT 240.210 101.820 240.460 101.830 ;
        RECT 239.080 101.420 239.330 101.430 ;
        RECT 239.080 100.970 240.060 101.420 ;
        RECT 241.170 101.160 250.440 101.170 ;
        RECT 252.320 101.160 254.240 101.170 ;
        RECT 241.170 100.970 254.240 101.160 ;
        RECT 239.080 100.360 239.330 100.970 ;
        RECT 241.170 100.960 253.530 100.970 ;
        RECT 239.080 100.110 240.290 100.360 ;
        RECT 240.020 99.360 240.280 100.110 ;
        RECT 241.170 99.950 241.380 100.960 ;
        RECT 250.430 100.950 252.330 100.960 ;
        RECT 254.060 100.220 254.240 100.970 ;
        RECT 240.020 98.760 240.270 99.360 ;
        RECT 241.170 98.940 241.370 99.950 ;
        RECT 248.980 99.920 254.240 100.220 ;
        RECT 239.230 98.310 240.270 98.760 ;
        RECT 239.210 96.860 240.170 97.310 ;
        RECT 239.920 96.810 240.170 96.860 ;
        RECT 241.180 96.810 241.370 98.940 ;
        RECT 239.920 96.610 241.370 96.810 ;
        RECT 244.900 98.280 245.160 99.480 ;
        RECT 244.900 97.770 245.150 98.280 ;
        RECT 246.790 98.270 247.050 99.480 ;
        RECT 249.180 98.370 249.430 99.920 ;
        RECT 246.790 98.110 247.180 98.270 ;
        RECT 246.780 97.980 247.180 98.110 ;
        RECT 249.880 97.980 250.140 99.590 ;
        RECT 252.430 98.520 252.730 99.570 ;
        RECT 253.180 98.970 253.480 99.920 ;
        RECT 253.680 99.020 253.980 99.070 ;
        RECT 253.680 98.670 254.580 99.020 ;
        RECT 256.290 98.890 256.510 98.900 ;
        RECT 256.290 98.700 269.970 98.890 ;
        RECT 256.290 98.570 256.510 98.700 ;
        RECT 245.400 97.770 245.690 97.930 ;
        RECT 246.780 97.920 247.040 97.980 ;
        RECT 244.900 97.580 245.690 97.770 ;
        RECT 244.900 97.380 245.150 97.580 ;
        RECT 245.400 97.470 245.690 97.580 ;
        RECT 246.790 97.380 247.040 97.920 ;
        RECT 249.870 97.920 250.140 97.980 ;
        RECT 251.420 98.260 252.730 98.520 ;
        RECT 254.830 98.270 256.510 98.570 ;
        RECT 254.830 98.260 256.490 98.270 ;
        RECT 251.420 97.920 251.730 98.260 ;
        RECT 247.430 97.390 249.070 97.780 ;
        RECT 249.870 97.630 251.730 97.920 ;
        RECT 249.870 97.620 250.180 97.630 ;
        RECT 251.420 97.620 251.730 97.630 ;
        RECT 244.900 96.780 245.190 97.380 ;
        RECT 246.790 96.780 247.080 97.380 ;
        RECT 239.920 96.520 240.170 96.610 ;
        RECT 239.190 96.070 240.170 96.520 ;
        RECT 249.130 96.170 249.430 97.170 ;
        RECT 249.880 96.570 250.180 97.620 ;
        RECT 252.480 96.520 252.730 98.260 ;
        RECT 269.720 97.800 269.970 98.700 ;
        RECT 253.180 96.170 253.440 97.720 ;
        RECT 264.660 97.500 269.970 97.800 ;
        RECT 249.080 96.150 254.330 96.170 ;
        RECT 249.080 95.870 254.450 96.150 ;
        RECT 242.530 95.470 242.810 95.540 ;
        RECT 243.710 95.500 243.990 95.530 ;
        RECT 254.160 95.500 254.450 95.870 ;
        RECT 243.710 95.490 254.450 95.500 ;
        RECT 241.120 95.270 242.810 95.470 ;
        RECT 239.910 95.070 240.190 95.080 ;
        RECT 239.170 94.620 240.190 95.070 ;
        RECT 241.120 94.620 241.350 95.270 ;
        RECT 242.530 95.210 242.810 95.270 ;
        RECT 243.690 95.260 254.450 95.490 ;
        RECT 243.710 95.250 254.450 95.260 ;
        RECT 260.580 95.860 260.840 97.060 ;
        RECT 260.580 95.350 260.830 95.860 ;
        RECT 262.470 95.850 262.730 97.060 ;
        RECT 264.860 95.950 265.110 97.500 ;
        RECT 262.470 95.690 262.860 95.850 ;
        RECT 262.460 95.560 262.860 95.690 ;
        RECT 265.560 95.560 265.820 97.170 ;
        RECT 268.110 96.100 268.410 97.150 ;
        RECT 268.860 96.550 269.160 97.500 ;
        RECT 269.360 96.600 269.660 96.650 ;
        RECT 269.360 96.250 270.260 96.600 ;
        RECT 283.020 96.200 287.490 96.230 ;
        RECT 272.080 96.170 287.490 96.200 ;
        RECT 271.410 96.150 287.490 96.170 ;
        RECT 261.080 95.350 261.370 95.510 ;
        RECT 262.460 95.500 262.720 95.560 ;
        RECT 243.710 95.240 254.410 95.250 ;
        RECT 243.710 95.200 243.990 95.240 ;
        RECT 260.580 95.160 261.370 95.350 ;
        RECT 260.580 94.960 260.830 95.160 ;
        RECT 261.080 95.050 261.370 95.160 ;
        RECT 262.470 94.960 262.720 95.500 ;
        RECT 265.550 95.500 265.820 95.560 ;
        RECT 267.100 95.840 268.410 96.100 ;
        RECT 267.100 95.500 267.410 95.840 ;
        RECT 263.110 94.970 264.750 95.360 ;
        RECT 265.550 95.210 267.410 95.500 ;
        RECT 265.550 95.200 265.860 95.210 ;
        RECT 267.100 95.200 267.410 95.210 ;
        RECT 242.510 94.640 242.780 94.720 ;
        RECT 239.910 94.410 241.350 94.620 ;
        RECT 241.900 94.420 242.780 94.640 ;
        RECT 239.910 93.360 240.190 94.410 ;
        RECT 241.900 93.610 242.120 94.420 ;
        RECT 242.510 94.390 242.780 94.420 ;
        RECT 243.640 94.680 243.930 94.730 ;
        RECT 243.640 94.500 254.390 94.680 ;
        RECT 243.640 94.400 243.930 94.500 ;
        RECT 248.480 94.490 252.110 94.500 ;
        RECT 254.190 93.820 254.390 94.500 ;
        RECT 260.580 94.360 260.870 94.960 ;
        RECT 262.470 94.360 262.760 94.960 ;
        RECT 239.190 92.910 240.190 93.360 ;
        RECT 239.170 91.460 240.470 91.910 ;
        RECT 240.170 91.060 240.470 91.460 ;
        RECT 241.890 91.080 242.120 93.610 ;
        RECT 249.140 93.520 254.390 93.820 ;
        RECT 264.810 93.750 265.110 94.750 ;
        RECT 265.560 94.150 265.860 95.200 ;
        RECT 268.160 94.100 268.410 95.840 ;
        RECT 270.530 95.830 287.490 96.150 ;
        RECT 271.410 95.820 287.490 95.830 ;
        RECT 271.410 95.790 283.390 95.820 ;
        RECT 271.410 95.780 272.300 95.790 ;
        RECT 268.860 93.750 269.120 95.300 ;
        RECT 269.950 93.750 270.150 93.760 ;
        RECT 240.960 91.060 242.120 91.080 ;
        RECT 240.170 90.880 242.120 91.060 ;
        RECT 245.060 91.880 245.320 93.080 ;
        RECT 245.060 91.370 245.310 91.880 ;
        RECT 246.950 91.870 247.210 93.080 ;
        RECT 249.340 91.970 249.590 93.520 ;
        RECT 246.950 91.710 247.340 91.870 ;
        RECT 246.940 91.580 247.340 91.710 ;
        RECT 250.040 91.580 250.300 93.190 ;
        RECT 252.590 92.120 252.890 93.170 ;
        RECT 253.340 92.570 253.640 93.520 ;
        RECT 254.190 93.510 254.390 93.520 ;
        RECT 264.760 93.450 270.150 93.750 ;
        RECT 253.840 92.620 254.140 92.670 ;
        RECT 253.840 92.270 254.740 92.620 ;
        RECT 269.950 92.210 270.150 93.450 ;
        RECT 287.110 92.250 287.470 95.820 ;
        RECT 262.390 92.190 263.580 92.200 ;
        RECT 264.570 92.190 265.760 92.200 ;
        RECT 266.790 92.190 267.980 92.200 ;
        RECT 268.970 92.190 270.160 92.210 ;
        RECT 260.180 92.180 270.160 92.190 ;
        RECT 256.790 92.160 257.980 92.170 ;
        RECT 259.070 92.160 270.160 92.180 ;
        RECT 245.560 91.370 245.850 91.530 ;
        RECT 246.940 91.520 247.200 91.580 ;
        RECT 245.060 91.180 245.850 91.370 ;
        RECT 245.060 90.980 245.310 91.180 ;
        RECT 245.560 91.070 245.850 91.180 ;
        RECT 246.950 90.980 247.200 91.520 ;
        RECT 250.030 91.520 250.300 91.580 ;
        RECT 251.580 91.860 252.890 92.120 ;
        RECT 254.950 91.930 270.160 92.160 ;
        RECT 282.240 91.950 287.490 92.250 ;
        RECT 254.950 91.920 269.110 91.930 ;
        RECT 254.950 91.910 262.480 91.920 ;
        RECT 263.490 91.910 264.680 91.920 ;
        RECT 265.640 91.910 266.830 91.920 ;
        RECT 267.920 91.910 269.110 91.920 ;
        RECT 254.950 91.900 260.260 91.910 ;
        RECT 254.950 91.890 259.120 91.900 ;
        RECT 254.950 91.880 256.840 91.890 ;
        RECT 257.930 91.880 259.120 91.890 ;
        RECT 254.950 91.870 255.670 91.880 ;
        RECT 251.580 91.520 251.890 91.860 ;
        RECT 247.590 90.990 249.230 91.380 ;
        RECT 250.030 91.230 251.890 91.520 ;
        RECT 250.030 91.220 250.340 91.230 ;
        RECT 251.580 91.220 251.890 91.230 ;
        RECT 240.170 90.870 240.820 90.880 ;
        RECT 240.170 90.540 240.470 90.870 ;
        RECT 239.450 90.090 240.470 90.540 ;
        RECT 245.060 90.380 245.350 90.980 ;
        RECT 246.950 90.380 247.240 90.980 ;
        RECT 240.170 90.080 240.470 90.090 ;
        RECT 249.290 89.770 249.590 90.770 ;
        RECT 250.040 90.170 250.340 91.220 ;
        RECT 252.640 90.120 252.890 91.860 ;
        RECT 253.340 89.770 253.600 91.320 ;
        RECT 278.160 90.310 278.420 91.510 ;
        RECT 278.160 89.800 278.410 90.310 ;
        RECT 280.050 90.300 280.310 91.510 ;
        RECT 282.440 90.400 282.690 91.950 ;
        RECT 280.050 90.140 280.440 90.300 ;
        RECT 280.040 90.010 280.440 90.140 ;
        RECT 283.140 90.010 283.400 91.620 ;
        RECT 285.690 90.550 285.990 91.600 ;
        RECT 286.440 91.000 286.740 91.950 ;
        RECT 286.940 91.050 287.240 91.100 ;
        RECT 286.940 90.700 287.840 91.050 ;
        RECT 278.660 89.800 278.950 89.960 ;
        RECT 280.040 89.950 280.300 90.010 ;
        RECT 249.240 89.760 254.490 89.770 ;
        RECT 239.120 89.680 239.370 89.690 ;
        RECT 239.120 89.220 240.100 89.680 ;
        RECT 249.240 89.470 254.510 89.760 ;
        RECT 239.120 88.920 239.370 89.220 ;
        RECT 247.090 89.130 248.930 89.140 ;
        RECT 254.340 89.130 254.510 89.470 ;
        RECT 240.830 89.120 241.070 89.130 ;
        RECT 241.910 89.120 254.510 89.130 ;
        RECT 240.830 88.960 254.510 89.120 ;
        RECT 278.160 89.610 278.950 89.800 ;
        RECT 278.160 89.410 278.410 89.610 ;
        RECT 278.660 89.500 278.950 89.610 ;
        RECT 280.050 89.410 280.300 89.950 ;
        RECT 283.130 89.950 283.400 90.010 ;
        RECT 284.680 90.290 285.990 90.550 ;
        RECT 288.050 90.600 289.720 90.620 ;
        RECT 304.860 90.600 305.170 101.950 ;
        RECT 288.050 90.310 305.210 90.600 ;
        RECT 288.740 90.300 305.210 90.310 ;
        RECT 284.680 89.950 284.990 90.290 ;
        RECT 280.690 89.420 282.330 89.810 ;
        RECT 283.130 89.660 284.990 89.950 ;
        RECT 283.130 89.650 283.440 89.660 ;
        RECT 284.680 89.650 284.990 89.660 ;
        RECT 240.830 88.950 252.340 88.960 ;
        RECT 240.820 88.940 247.140 88.950 ;
        RECT 248.690 88.940 252.340 88.950 ;
        RECT 240.820 88.930 242.690 88.940 ;
        RECT 240.820 88.920 241.070 88.930 ;
        RECT 239.120 88.750 241.070 88.920 ;
        RECT 278.160 88.810 278.450 89.410 ;
        RECT 280.050 88.810 280.340 89.410 ;
        RECT 239.120 88.530 239.370 88.750 ;
        RECT 239.120 88.360 240.160 88.530 ;
        RECT 239.970 87.500 240.160 88.360 ;
        RECT 282.390 88.200 282.690 89.200 ;
        RECT 283.140 88.600 283.440 89.650 ;
        RECT 285.740 88.550 285.990 90.290 ;
        RECT 286.440 88.200 286.700 89.750 ;
        RECT 287.320 88.200 287.660 88.270 ;
        RECT 282.340 87.900 287.660 88.200 ;
        RECT 239.180 87.060 240.160 87.500 ;
        RECT 239.180 87.050 240.130 87.060 ;
        RECT 241.000 86.740 250.270 86.750 ;
        RECT 252.150 86.740 254.070 86.750 ;
        RECT 238.850 86.640 239.040 86.650 ;
        RECT 238.850 86.180 239.830 86.640 ;
        RECT 241.000 86.550 254.070 86.740 ;
        RECT 241.000 86.540 253.360 86.550 ;
        RECT 238.850 85.390 239.040 86.180 ;
        RECT 241.000 85.530 241.210 86.540 ;
        RECT 250.260 86.530 252.160 86.540 ;
        RECT 253.890 85.800 254.070 86.550 ;
        RECT 239.850 85.390 240.120 85.400 ;
        RECT 238.850 85.180 240.120 85.390 ;
        RECT 239.850 84.970 240.120 85.180 ;
        RECT 239.850 84.340 240.100 84.970 ;
        RECT 241.000 84.520 241.200 85.530 ;
        RECT 248.810 85.500 254.070 85.800 ;
        RECT 239.060 83.890 240.100 84.340 ;
        RECT 239.040 82.440 240.000 82.890 ;
        RECT 239.750 82.390 240.000 82.440 ;
        RECT 241.010 82.390 241.200 84.520 ;
        RECT 239.750 82.190 241.200 82.390 ;
        RECT 244.730 83.860 244.990 85.060 ;
        RECT 244.730 83.350 244.980 83.860 ;
        RECT 246.620 83.850 246.880 85.060 ;
        RECT 249.010 83.950 249.260 85.500 ;
        RECT 246.620 83.690 247.010 83.850 ;
        RECT 246.610 83.560 247.010 83.690 ;
        RECT 249.710 83.560 249.970 85.170 ;
        RECT 252.260 84.100 252.560 85.150 ;
        RECT 253.010 84.550 253.310 85.500 ;
        RECT 253.510 84.600 253.810 84.650 ;
        RECT 253.510 84.250 254.410 84.600 ;
        RECT 256.120 84.470 256.340 84.480 ;
        RECT 256.120 84.280 269.800 84.470 ;
        RECT 256.120 84.150 256.340 84.280 ;
        RECT 245.230 83.350 245.520 83.510 ;
        RECT 246.610 83.500 246.870 83.560 ;
        RECT 244.730 83.160 245.520 83.350 ;
        RECT 244.730 82.960 244.980 83.160 ;
        RECT 245.230 83.050 245.520 83.160 ;
        RECT 246.620 82.960 246.870 83.500 ;
        RECT 249.700 83.500 249.970 83.560 ;
        RECT 251.250 83.840 252.560 84.100 ;
        RECT 254.660 83.850 256.340 84.150 ;
        RECT 254.660 83.840 256.320 83.850 ;
        RECT 251.250 83.500 251.560 83.840 ;
        RECT 247.260 82.970 248.900 83.360 ;
        RECT 249.700 83.210 251.560 83.500 ;
        RECT 249.700 83.200 250.010 83.210 ;
        RECT 251.250 83.200 251.560 83.210 ;
        RECT 244.730 82.360 245.020 82.960 ;
        RECT 246.620 82.360 246.910 82.960 ;
        RECT 239.750 82.100 240.000 82.190 ;
        RECT 239.020 81.650 240.000 82.100 ;
        RECT 248.960 81.750 249.260 82.750 ;
        RECT 249.710 82.150 250.010 83.200 ;
        RECT 252.310 82.100 252.560 83.840 ;
        RECT 269.550 83.380 269.800 84.280 ;
        RECT 253.010 81.750 253.270 83.300 ;
        RECT 264.490 83.080 269.800 83.380 ;
        RECT 248.910 81.730 254.160 81.750 ;
        RECT 248.910 81.450 254.280 81.730 ;
        RECT 242.360 81.050 242.640 81.120 ;
        RECT 243.540 81.080 243.820 81.110 ;
        RECT 253.990 81.080 254.280 81.450 ;
        RECT 243.540 81.070 254.280 81.080 ;
        RECT 240.950 80.850 242.640 81.050 ;
        RECT 239.740 80.650 240.020 80.660 ;
        RECT 239.000 80.200 240.020 80.650 ;
        RECT 240.950 80.200 241.180 80.850 ;
        RECT 242.360 80.790 242.640 80.850 ;
        RECT 243.520 80.840 254.280 81.070 ;
        RECT 243.540 80.830 254.280 80.840 ;
        RECT 260.410 81.440 260.670 82.640 ;
        RECT 260.410 80.930 260.660 81.440 ;
        RECT 262.300 81.430 262.560 82.640 ;
        RECT 264.690 81.530 264.940 83.080 ;
        RECT 262.300 81.270 262.690 81.430 ;
        RECT 262.290 81.140 262.690 81.270 ;
        RECT 265.390 81.140 265.650 82.750 ;
        RECT 267.940 81.680 268.240 82.730 ;
        RECT 268.690 82.130 268.990 83.080 ;
        RECT 269.190 82.180 269.490 82.230 ;
        RECT 269.190 81.830 270.090 82.180 ;
        RECT 287.320 81.780 287.660 87.900 ;
        RECT 319.060 85.100 319.240 104.360 ;
        RECT 319.040 84.050 319.250 85.100 ;
        RECT 319.040 83.970 319.260 84.050 ;
        RECT 319.050 81.900 319.260 83.970 ;
        RECT 319.040 81.860 319.260 81.900 ;
        RECT 286.750 81.760 287.710 81.780 ;
        RECT 271.230 81.740 275.510 81.750 ;
        RECT 282.910 81.740 287.710 81.760 ;
        RECT 271.230 81.730 287.710 81.740 ;
        RECT 260.910 80.930 261.200 81.090 ;
        RECT 262.290 81.080 262.550 81.140 ;
        RECT 243.540 80.820 254.240 80.830 ;
        RECT 243.540 80.780 243.820 80.820 ;
        RECT 260.410 80.740 261.200 80.930 ;
        RECT 260.410 80.540 260.660 80.740 ;
        RECT 260.910 80.630 261.200 80.740 ;
        RECT 262.300 80.540 262.550 81.080 ;
        RECT 265.380 81.080 265.650 81.140 ;
        RECT 266.930 81.420 268.240 81.680 ;
        RECT 266.930 81.080 267.240 81.420 ;
        RECT 262.940 80.550 264.580 80.940 ;
        RECT 265.380 80.790 267.240 81.080 ;
        RECT 265.380 80.780 265.690 80.790 ;
        RECT 266.930 80.780 267.240 80.790 ;
        RECT 242.340 80.220 242.610 80.300 ;
        RECT 239.740 79.990 241.180 80.200 ;
        RECT 241.730 80.000 242.610 80.220 ;
        RECT 239.740 78.940 240.020 79.990 ;
        RECT 241.730 79.190 241.950 80.000 ;
        RECT 242.340 79.970 242.610 80.000 ;
        RECT 243.470 80.260 243.760 80.310 ;
        RECT 243.470 80.080 254.220 80.260 ;
        RECT 243.470 79.980 243.760 80.080 ;
        RECT 248.310 80.070 251.940 80.080 ;
        RECT 254.020 79.400 254.220 80.080 ;
        RECT 260.410 79.940 260.700 80.540 ;
        RECT 262.300 79.940 262.590 80.540 ;
        RECT 239.020 78.490 240.020 78.940 ;
        RECT 239.000 77.040 240.300 77.490 ;
        RECT 240.000 76.640 240.300 77.040 ;
        RECT 241.720 76.660 241.950 79.190 ;
        RECT 248.970 79.100 254.220 79.400 ;
        RECT 264.640 79.330 264.940 80.330 ;
        RECT 265.390 79.730 265.690 80.780 ;
        RECT 267.990 79.680 268.240 81.420 ;
        RECT 270.360 81.420 287.710 81.730 ;
        RECT 270.360 81.410 283.370 81.420 ;
        RECT 275.220 81.400 283.370 81.410 ;
        RECT 286.750 81.380 287.710 81.420 ;
        RECT 287.320 81.370 287.660 81.380 ;
        RECT 268.690 79.330 268.950 80.880 ;
        RECT 319.040 80.010 319.250 81.860 ;
        RECT 314.000 79.710 319.250 80.010 ;
        RECT 269.780 79.330 269.980 79.340 ;
        RECT 240.790 76.640 241.950 76.660 ;
        RECT 240.000 76.460 241.950 76.640 ;
        RECT 244.890 77.460 245.150 78.660 ;
        RECT 244.890 76.950 245.140 77.460 ;
        RECT 246.780 77.450 247.040 78.660 ;
        RECT 249.170 77.550 249.420 79.100 ;
        RECT 246.780 77.290 247.170 77.450 ;
        RECT 246.770 77.160 247.170 77.290 ;
        RECT 249.870 77.160 250.130 78.770 ;
        RECT 252.420 77.700 252.720 78.750 ;
        RECT 253.170 78.150 253.470 79.100 ;
        RECT 254.020 79.090 254.220 79.100 ;
        RECT 264.590 79.030 269.980 79.330 ;
        RECT 253.670 78.200 253.970 78.250 ;
        RECT 253.670 77.850 254.570 78.200 ;
        RECT 269.780 77.790 269.980 79.030 ;
        RECT 309.920 78.070 310.180 79.270 ;
        RECT 262.220 77.770 263.410 77.780 ;
        RECT 264.400 77.770 265.590 77.780 ;
        RECT 266.620 77.770 267.810 77.780 ;
        RECT 268.800 77.770 269.990 77.790 ;
        RECT 260.010 77.760 269.990 77.770 ;
        RECT 256.620 77.740 257.810 77.750 ;
        RECT 258.900 77.740 269.990 77.760 ;
        RECT 245.390 76.950 245.680 77.110 ;
        RECT 246.770 77.100 247.030 77.160 ;
        RECT 244.890 76.760 245.680 76.950 ;
        RECT 244.890 76.560 245.140 76.760 ;
        RECT 245.390 76.650 245.680 76.760 ;
        RECT 246.780 76.560 247.030 77.100 ;
        RECT 249.860 77.100 250.130 77.160 ;
        RECT 251.410 77.440 252.720 77.700 ;
        RECT 254.780 77.510 269.990 77.740 ;
        RECT 309.920 77.560 310.170 78.070 ;
        RECT 311.810 78.060 312.070 79.270 ;
        RECT 314.200 78.160 314.450 79.710 ;
        RECT 311.810 77.900 312.200 78.060 ;
        RECT 311.800 77.770 312.200 77.900 ;
        RECT 314.900 77.770 315.160 79.380 ;
        RECT 317.450 78.310 317.750 79.360 ;
        RECT 318.200 78.760 318.500 79.710 ;
        RECT 319.040 79.700 319.250 79.710 ;
        RECT 318.700 78.810 319.000 78.860 ;
        RECT 318.700 78.460 319.600 78.810 ;
        RECT 336.370 78.430 336.670 132.770 ;
        RECT 340.370 132.120 340.720 132.780 ;
        RECT 432.240 132.580 437.980 132.870 ;
        RECT 449.450 132.830 463.900 133.030 ;
        RECT 449.450 132.820 461.250 132.830 ;
        RECT 449.450 132.800 457.410 132.820 ;
        RECT 432.240 132.570 437.490 132.580 ;
        RECT 339.100 131.780 340.720 132.120 ;
        RECT 339.100 130.930 339.550 131.780 ;
        RECT 340.370 131.770 340.720 131.780 ;
        RECT 339.960 130.750 340.420 131.580 ;
        RECT 342.510 131.040 351.780 131.050 ;
        RECT 353.660 131.040 355.580 131.050 ;
        RECT 341.340 130.750 341.620 130.890 ;
        RECT 339.960 130.640 341.620 130.750 ;
        RECT 339.970 130.440 341.620 130.640 ;
        RECT 342.510 130.850 355.580 131.040 ;
        RECT 342.510 130.840 354.870 130.850 ;
        RECT 339.970 130.430 341.640 130.440 ;
        RECT 341.340 130.210 341.640 130.430 ;
        RECT 341.350 130.040 341.640 130.210 ;
        RECT 341.360 129.240 341.620 130.040 ;
        RECT 342.510 129.830 342.720 130.840 ;
        RECT 351.770 130.830 353.670 130.840 ;
        RECT 355.400 130.100 355.580 130.850 ;
        RECT 341.360 128.640 341.610 129.240 ;
        RECT 342.510 128.820 342.710 129.830 ;
        RECT 350.320 129.800 355.580 130.100 ;
        RECT 340.570 128.190 341.610 128.640 ;
        RECT 340.550 126.740 341.510 127.190 ;
        RECT 341.260 126.690 341.510 126.740 ;
        RECT 342.520 126.690 342.710 128.820 ;
        RECT 341.260 126.490 342.710 126.690 ;
        RECT 346.240 128.160 346.500 129.360 ;
        RECT 346.240 127.650 346.490 128.160 ;
        RECT 348.130 128.150 348.390 129.360 ;
        RECT 350.520 128.250 350.770 129.800 ;
        RECT 348.130 127.990 348.520 128.150 ;
        RECT 348.120 127.860 348.520 127.990 ;
        RECT 351.220 127.860 351.480 129.470 ;
        RECT 353.770 128.400 354.070 129.450 ;
        RECT 354.520 128.850 354.820 129.800 ;
        RECT 355.020 128.900 355.320 128.950 ;
        RECT 355.020 128.550 355.920 128.900 ;
        RECT 357.630 128.770 357.850 128.780 ;
        RECT 357.630 128.580 371.310 128.770 ;
        RECT 357.630 128.450 357.850 128.580 ;
        RECT 346.740 127.650 347.030 127.810 ;
        RECT 348.120 127.800 348.380 127.860 ;
        RECT 346.240 127.460 347.030 127.650 ;
        RECT 346.240 127.260 346.490 127.460 ;
        RECT 346.740 127.350 347.030 127.460 ;
        RECT 348.130 127.260 348.380 127.800 ;
        RECT 351.210 127.800 351.480 127.860 ;
        RECT 352.760 128.140 354.070 128.400 ;
        RECT 356.170 128.150 357.850 128.450 ;
        RECT 356.170 128.140 357.830 128.150 ;
        RECT 352.760 127.800 353.070 128.140 ;
        RECT 348.770 127.270 350.410 127.660 ;
        RECT 351.210 127.510 353.070 127.800 ;
        RECT 351.210 127.500 351.520 127.510 ;
        RECT 352.760 127.500 353.070 127.510 ;
        RECT 346.240 126.660 346.530 127.260 ;
        RECT 348.130 126.660 348.420 127.260 ;
        RECT 341.260 126.400 341.510 126.490 ;
        RECT 340.530 125.950 341.510 126.400 ;
        RECT 350.470 126.050 350.770 127.050 ;
        RECT 351.220 126.450 351.520 127.500 ;
        RECT 353.820 126.400 354.070 128.140 ;
        RECT 371.060 127.680 371.310 128.580 ;
        RECT 354.520 126.050 354.780 127.600 ;
        RECT 366.000 127.380 371.310 127.680 ;
        RECT 350.420 126.030 355.670 126.050 ;
        RECT 350.420 125.750 355.790 126.030 ;
        RECT 343.870 125.350 344.150 125.420 ;
        RECT 345.050 125.380 345.330 125.410 ;
        RECT 355.500 125.380 355.790 125.750 ;
        RECT 345.050 125.370 355.790 125.380 ;
        RECT 342.460 125.150 344.150 125.350 ;
        RECT 341.250 124.950 341.530 124.960 ;
        RECT 340.510 124.500 341.530 124.950 ;
        RECT 342.460 124.500 342.690 125.150 ;
        RECT 343.870 125.090 344.150 125.150 ;
        RECT 345.030 125.140 355.790 125.370 ;
        RECT 345.050 125.130 355.790 125.140 ;
        RECT 361.920 125.740 362.180 126.940 ;
        RECT 361.920 125.230 362.170 125.740 ;
        RECT 363.810 125.730 364.070 126.940 ;
        RECT 366.200 125.830 366.450 127.380 ;
        RECT 363.810 125.570 364.200 125.730 ;
        RECT 363.800 125.440 364.200 125.570 ;
        RECT 366.900 125.440 367.160 127.050 ;
        RECT 369.450 125.980 369.750 127.030 ;
        RECT 370.200 126.430 370.500 127.380 ;
        RECT 370.700 126.480 371.000 126.530 ;
        RECT 370.700 126.130 371.600 126.480 ;
        RECT 384.360 126.080 388.830 126.110 ;
        RECT 373.420 126.050 388.830 126.080 ;
        RECT 372.750 126.030 388.830 126.050 ;
        RECT 362.420 125.230 362.710 125.390 ;
        RECT 363.800 125.380 364.060 125.440 ;
        RECT 345.050 125.120 355.750 125.130 ;
        RECT 345.050 125.080 345.330 125.120 ;
        RECT 361.920 125.040 362.710 125.230 ;
        RECT 361.920 124.840 362.170 125.040 ;
        RECT 362.420 124.930 362.710 125.040 ;
        RECT 363.810 124.840 364.060 125.380 ;
        RECT 366.890 125.380 367.160 125.440 ;
        RECT 368.440 125.720 369.750 125.980 ;
        RECT 368.440 125.380 368.750 125.720 ;
        RECT 364.450 124.850 366.090 125.240 ;
        RECT 366.890 125.090 368.750 125.380 ;
        RECT 366.890 125.080 367.200 125.090 ;
        RECT 368.440 125.080 368.750 125.090 ;
        RECT 343.850 124.520 344.120 124.600 ;
        RECT 341.250 124.290 342.690 124.500 ;
        RECT 343.240 124.300 344.120 124.520 ;
        RECT 341.250 123.240 341.530 124.290 ;
        RECT 343.240 123.490 343.460 124.300 ;
        RECT 343.850 124.270 344.120 124.300 ;
        RECT 344.980 124.560 345.270 124.610 ;
        RECT 344.980 124.380 355.730 124.560 ;
        RECT 344.980 124.280 345.270 124.380 ;
        RECT 349.820 124.370 353.450 124.380 ;
        RECT 355.530 123.700 355.730 124.380 ;
        RECT 361.920 124.240 362.210 124.840 ;
        RECT 363.810 124.240 364.100 124.840 ;
        RECT 340.530 122.790 341.530 123.240 ;
        RECT 340.510 121.340 341.810 121.790 ;
        RECT 341.510 120.940 341.810 121.340 ;
        RECT 343.230 120.960 343.460 123.490 ;
        RECT 350.480 123.400 355.730 123.700 ;
        RECT 366.150 123.630 366.450 124.630 ;
        RECT 366.900 124.030 367.200 125.080 ;
        RECT 369.500 123.980 369.750 125.720 ;
        RECT 371.870 125.710 388.830 126.030 ;
        RECT 372.750 125.700 388.830 125.710 ;
        RECT 372.750 125.670 384.730 125.700 ;
        RECT 372.750 125.660 373.640 125.670 ;
        RECT 370.200 123.630 370.460 125.180 ;
        RECT 371.290 123.630 371.490 123.640 ;
        RECT 342.300 120.940 343.460 120.960 ;
        RECT 341.510 120.760 343.460 120.940 ;
        RECT 346.400 121.760 346.660 122.960 ;
        RECT 346.400 121.250 346.650 121.760 ;
        RECT 348.290 121.750 348.550 122.960 ;
        RECT 350.680 121.850 350.930 123.400 ;
        RECT 348.290 121.590 348.680 121.750 ;
        RECT 348.280 121.460 348.680 121.590 ;
        RECT 351.380 121.460 351.640 123.070 ;
        RECT 353.930 122.000 354.230 123.050 ;
        RECT 354.680 122.450 354.980 123.400 ;
        RECT 355.530 123.390 355.730 123.400 ;
        RECT 366.100 123.330 371.490 123.630 ;
        RECT 355.180 122.500 355.480 122.550 ;
        RECT 355.180 122.150 356.080 122.500 ;
        RECT 371.290 122.090 371.490 123.330 ;
        RECT 388.450 122.130 388.810 125.700 ;
        RECT 363.730 122.070 364.920 122.080 ;
        RECT 365.910 122.070 367.100 122.080 ;
        RECT 368.130 122.070 369.320 122.080 ;
        RECT 370.310 122.070 371.500 122.090 ;
        RECT 361.520 122.060 371.500 122.070 ;
        RECT 358.130 122.040 359.320 122.050 ;
        RECT 360.410 122.040 371.500 122.060 ;
        RECT 346.900 121.250 347.190 121.410 ;
        RECT 348.280 121.400 348.540 121.460 ;
        RECT 346.400 121.060 347.190 121.250 ;
        RECT 346.400 120.860 346.650 121.060 ;
        RECT 346.900 120.950 347.190 121.060 ;
        RECT 348.290 120.860 348.540 121.400 ;
        RECT 351.370 121.400 351.640 121.460 ;
        RECT 352.920 121.740 354.230 122.000 ;
        RECT 356.290 121.810 371.500 122.040 ;
        RECT 383.580 121.830 388.830 122.130 ;
        RECT 356.290 121.800 370.450 121.810 ;
        RECT 356.290 121.790 363.820 121.800 ;
        RECT 364.830 121.790 366.020 121.800 ;
        RECT 366.980 121.790 368.170 121.800 ;
        RECT 369.260 121.790 370.450 121.800 ;
        RECT 356.290 121.780 361.600 121.790 ;
        RECT 356.290 121.770 360.460 121.780 ;
        RECT 356.290 121.760 358.180 121.770 ;
        RECT 359.270 121.760 360.460 121.770 ;
        RECT 356.290 121.750 357.010 121.760 ;
        RECT 352.920 121.400 353.230 121.740 ;
        RECT 348.930 120.870 350.570 121.260 ;
        RECT 351.370 121.110 353.230 121.400 ;
        RECT 351.370 121.100 351.680 121.110 ;
        RECT 352.920 121.100 353.230 121.110 ;
        RECT 341.510 120.750 342.160 120.760 ;
        RECT 341.510 120.420 341.810 120.750 ;
        RECT 340.790 119.970 341.810 120.420 ;
        RECT 346.400 120.260 346.690 120.860 ;
        RECT 348.290 120.260 348.580 120.860 ;
        RECT 341.510 119.960 341.810 119.970 ;
        RECT 350.630 119.650 350.930 120.650 ;
        RECT 351.380 120.050 351.680 121.100 ;
        RECT 353.980 120.000 354.230 121.740 ;
        RECT 354.680 119.650 354.940 121.200 ;
        RECT 379.500 120.190 379.760 121.390 ;
        RECT 379.500 119.680 379.750 120.190 ;
        RECT 381.390 120.180 381.650 121.390 ;
        RECT 383.780 120.280 384.030 121.830 ;
        RECT 381.390 120.020 381.780 120.180 ;
        RECT 381.380 119.890 381.780 120.020 ;
        RECT 384.480 119.890 384.740 121.500 ;
        RECT 387.030 120.430 387.330 121.480 ;
        RECT 387.780 120.880 388.080 121.830 ;
        RECT 388.280 120.930 388.580 120.980 ;
        RECT 388.280 120.580 389.180 120.930 ;
        RECT 380.000 119.680 380.290 119.840 ;
        RECT 381.380 119.830 381.640 119.890 ;
        RECT 350.580 119.640 355.830 119.650 ;
        RECT 340.460 119.560 340.710 119.570 ;
        RECT 340.460 119.100 341.440 119.560 ;
        RECT 350.580 119.350 355.850 119.640 ;
        RECT 340.460 118.800 340.710 119.100 ;
        RECT 348.430 119.010 350.270 119.020 ;
        RECT 355.680 119.010 355.850 119.350 ;
        RECT 342.170 119.000 342.410 119.010 ;
        RECT 343.250 119.000 355.850 119.010 ;
        RECT 342.170 118.840 355.850 119.000 ;
        RECT 379.500 119.490 380.290 119.680 ;
        RECT 379.500 119.290 379.750 119.490 ;
        RECT 380.000 119.380 380.290 119.490 ;
        RECT 381.390 119.290 381.640 119.830 ;
        RECT 384.470 119.830 384.740 119.890 ;
        RECT 386.020 120.170 387.330 120.430 ;
        RECT 389.390 120.470 391.060 120.500 ;
        RECT 406.140 120.470 406.390 120.480 ;
        RECT 389.390 120.200 406.390 120.470 ;
        RECT 389.390 120.190 402.890 120.200 ;
        RECT 390.670 120.170 402.890 120.190 ;
        RECT 386.020 119.830 386.330 120.170 ;
        RECT 382.030 119.300 383.670 119.690 ;
        RECT 384.470 119.540 386.330 119.830 ;
        RECT 384.470 119.530 384.780 119.540 ;
        RECT 386.020 119.530 386.330 119.540 ;
        RECT 342.170 118.830 353.680 118.840 ;
        RECT 342.160 118.820 348.480 118.830 ;
        RECT 350.030 118.820 353.680 118.830 ;
        RECT 342.160 118.810 344.030 118.820 ;
        RECT 342.160 118.800 342.410 118.810 ;
        RECT 340.460 118.630 342.410 118.800 ;
        RECT 379.500 118.690 379.790 119.290 ;
        RECT 381.390 118.690 381.680 119.290 ;
        RECT 340.460 118.410 340.710 118.630 ;
        RECT 340.460 118.240 341.500 118.410 ;
        RECT 341.310 117.380 341.500 118.240 ;
        RECT 383.730 118.080 384.030 119.080 ;
        RECT 384.480 118.480 384.780 119.530 ;
        RECT 387.080 118.430 387.330 120.170 ;
        RECT 387.780 118.080 388.040 119.630 ;
        RECT 388.660 118.080 389.000 118.150 ;
        RECT 383.680 117.780 389.000 118.080 ;
        RECT 340.520 116.940 341.500 117.380 ;
        RECT 340.520 116.930 341.470 116.940 ;
        RECT 342.340 116.620 351.610 116.630 ;
        RECT 353.490 116.620 355.410 116.630 ;
        RECT 340.190 116.520 340.380 116.530 ;
        RECT 340.190 116.060 341.170 116.520 ;
        RECT 342.340 116.430 355.410 116.620 ;
        RECT 342.340 116.420 354.700 116.430 ;
        RECT 340.190 115.270 340.380 116.060 ;
        RECT 342.340 115.410 342.550 116.420 ;
        RECT 351.600 116.410 353.500 116.420 ;
        RECT 355.230 115.680 355.410 116.430 ;
        RECT 341.190 115.270 341.460 115.280 ;
        RECT 340.190 115.060 341.460 115.270 ;
        RECT 341.190 114.850 341.460 115.060 ;
        RECT 341.190 114.220 341.440 114.850 ;
        RECT 342.340 114.400 342.540 115.410 ;
        RECT 350.150 115.380 355.410 115.680 ;
        RECT 340.400 113.770 341.440 114.220 ;
        RECT 340.380 112.320 341.340 112.770 ;
        RECT 341.090 112.270 341.340 112.320 ;
        RECT 342.350 112.270 342.540 114.400 ;
        RECT 341.090 112.070 342.540 112.270 ;
        RECT 346.070 113.740 346.330 114.940 ;
        RECT 346.070 113.230 346.320 113.740 ;
        RECT 347.960 113.730 348.220 114.940 ;
        RECT 350.350 113.830 350.600 115.380 ;
        RECT 347.960 113.570 348.350 113.730 ;
        RECT 347.950 113.440 348.350 113.570 ;
        RECT 351.050 113.440 351.310 115.050 ;
        RECT 353.600 113.980 353.900 115.030 ;
        RECT 354.350 114.430 354.650 115.380 ;
        RECT 354.850 114.480 355.150 114.530 ;
        RECT 354.850 114.130 355.750 114.480 ;
        RECT 357.460 114.350 357.680 114.360 ;
        RECT 357.460 114.160 371.140 114.350 ;
        RECT 357.460 114.030 357.680 114.160 ;
        RECT 346.570 113.230 346.860 113.390 ;
        RECT 347.950 113.380 348.210 113.440 ;
        RECT 346.070 113.040 346.860 113.230 ;
        RECT 346.070 112.840 346.320 113.040 ;
        RECT 346.570 112.930 346.860 113.040 ;
        RECT 347.960 112.840 348.210 113.380 ;
        RECT 351.040 113.380 351.310 113.440 ;
        RECT 352.590 113.720 353.900 113.980 ;
        RECT 356.000 113.730 357.680 114.030 ;
        RECT 356.000 113.720 357.660 113.730 ;
        RECT 352.590 113.380 352.900 113.720 ;
        RECT 348.600 112.850 350.240 113.240 ;
        RECT 351.040 113.090 352.900 113.380 ;
        RECT 351.040 113.080 351.350 113.090 ;
        RECT 352.590 113.080 352.900 113.090 ;
        RECT 346.070 112.240 346.360 112.840 ;
        RECT 347.960 112.240 348.250 112.840 ;
        RECT 341.090 111.980 341.340 112.070 ;
        RECT 340.360 111.530 341.340 111.980 ;
        RECT 350.300 111.630 350.600 112.630 ;
        RECT 351.050 112.030 351.350 113.080 ;
        RECT 353.650 111.980 353.900 113.720 ;
        RECT 370.890 113.260 371.140 114.160 ;
        RECT 354.350 111.630 354.610 113.180 ;
        RECT 365.830 112.960 371.140 113.260 ;
        RECT 350.250 111.610 355.500 111.630 ;
        RECT 350.250 111.330 355.620 111.610 ;
        RECT 343.700 110.930 343.980 111.000 ;
        RECT 344.880 110.960 345.160 110.990 ;
        RECT 355.330 110.960 355.620 111.330 ;
        RECT 344.880 110.950 355.620 110.960 ;
        RECT 342.290 110.730 343.980 110.930 ;
        RECT 341.080 110.530 341.360 110.540 ;
        RECT 340.340 110.080 341.360 110.530 ;
        RECT 342.290 110.080 342.520 110.730 ;
        RECT 343.700 110.670 343.980 110.730 ;
        RECT 344.860 110.720 355.620 110.950 ;
        RECT 344.880 110.710 355.620 110.720 ;
        RECT 361.750 111.320 362.010 112.520 ;
        RECT 361.750 110.810 362.000 111.320 ;
        RECT 363.640 111.310 363.900 112.520 ;
        RECT 366.030 111.410 366.280 112.960 ;
        RECT 363.640 111.150 364.030 111.310 ;
        RECT 363.630 111.020 364.030 111.150 ;
        RECT 366.730 111.020 366.990 112.630 ;
        RECT 369.280 111.560 369.580 112.610 ;
        RECT 370.030 112.010 370.330 112.960 ;
        RECT 370.530 112.060 370.830 112.110 ;
        RECT 370.530 111.710 371.430 112.060 ;
        RECT 388.660 111.660 389.000 117.780 ;
        RECT 388.090 111.640 389.050 111.660 ;
        RECT 372.570 111.620 376.850 111.630 ;
        RECT 384.250 111.620 389.050 111.640 ;
        RECT 372.570 111.610 389.050 111.620 ;
        RECT 362.250 110.810 362.540 110.970 ;
        RECT 363.630 110.960 363.890 111.020 ;
        RECT 344.880 110.700 355.580 110.710 ;
        RECT 344.880 110.660 345.160 110.700 ;
        RECT 361.750 110.620 362.540 110.810 ;
        RECT 361.750 110.420 362.000 110.620 ;
        RECT 362.250 110.510 362.540 110.620 ;
        RECT 363.640 110.420 363.890 110.960 ;
        RECT 366.720 110.960 366.990 111.020 ;
        RECT 368.270 111.300 369.580 111.560 ;
        RECT 368.270 110.960 368.580 111.300 ;
        RECT 364.280 110.430 365.920 110.820 ;
        RECT 366.720 110.670 368.580 110.960 ;
        RECT 366.720 110.660 367.030 110.670 ;
        RECT 368.270 110.660 368.580 110.670 ;
        RECT 343.680 110.100 343.950 110.180 ;
        RECT 341.080 109.870 342.520 110.080 ;
        RECT 343.070 109.880 343.950 110.100 ;
        RECT 341.080 108.820 341.360 109.870 ;
        RECT 343.070 109.070 343.290 109.880 ;
        RECT 343.680 109.850 343.950 109.880 ;
        RECT 344.810 110.140 345.100 110.190 ;
        RECT 344.810 109.960 355.560 110.140 ;
        RECT 344.810 109.860 345.100 109.960 ;
        RECT 349.650 109.950 353.280 109.960 ;
        RECT 355.360 109.280 355.560 109.960 ;
        RECT 361.750 109.820 362.040 110.420 ;
        RECT 363.640 109.820 363.930 110.420 ;
        RECT 340.360 108.370 341.360 108.820 ;
        RECT 340.340 106.920 341.640 107.370 ;
        RECT 341.340 106.520 341.640 106.920 ;
        RECT 343.060 106.540 343.290 109.070 ;
        RECT 350.310 108.980 355.560 109.280 ;
        RECT 365.980 109.210 366.280 110.210 ;
        RECT 366.730 109.610 367.030 110.660 ;
        RECT 369.330 109.560 369.580 111.300 ;
        RECT 371.700 111.300 389.050 111.610 ;
        RECT 371.700 111.290 384.710 111.300 ;
        RECT 376.560 111.280 384.710 111.290 ;
        RECT 388.090 111.260 389.050 111.300 ;
        RECT 388.660 111.250 389.000 111.260 ;
        RECT 370.030 109.210 370.290 110.760 ;
        RECT 371.120 109.210 371.320 109.220 ;
        RECT 342.130 106.520 343.290 106.540 ;
        RECT 341.340 106.340 343.290 106.520 ;
        RECT 346.230 107.340 346.490 108.540 ;
        RECT 346.230 106.830 346.480 107.340 ;
        RECT 348.120 107.330 348.380 108.540 ;
        RECT 350.510 107.430 350.760 108.980 ;
        RECT 348.120 107.170 348.510 107.330 ;
        RECT 348.110 107.040 348.510 107.170 ;
        RECT 351.210 107.040 351.470 108.650 ;
        RECT 353.760 107.580 354.060 108.630 ;
        RECT 354.510 108.030 354.810 108.980 ;
        RECT 355.360 108.970 355.560 108.980 ;
        RECT 365.930 108.910 371.320 109.210 ;
        RECT 355.010 108.080 355.310 108.130 ;
        RECT 355.010 107.730 355.910 108.080 ;
        RECT 371.120 107.670 371.320 108.910 ;
        RECT 363.560 107.650 364.750 107.660 ;
        RECT 365.740 107.650 366.930 107.660 ;
        RECT 367.960 107.650 369.150 107.660 ;
        RECT 370.140 107.650 371.330 107.670 ;
        RECT 361.350 107.640 371.330 107.650 ;
        RECT 357.960 107.620 359.150 107.630 ;
        RECT 360.240 107.620 371.330 107.640 ;
        RECT 346.730 106.830 347.020 106.990 ;
        RECT 348.110 106.980 348.370 107.040 ;
        RECT 346.230 106.640 347.020 106.830 ;
        RECT 346.230 106.440 346.480 106.640 ;
        RECT 346.730 106.530 347.020 106.640 ;
        RECT 348.120 106.440 348.370 106.980 ;
        RECT 351.200 106.980 351.470 107.040 ;
        RECT 352.750 107.320 354.060 107.580 ;
        RECT 356.120 107.390 371.330 107.620 ;
        RECT 356.120 107.380 370.280 107.390 ;
        RECT 356.120 107.370 363.650 107.380 ;
        RECT 364.660 107.370 365.850 107.380 ;
        RECT 366.810 107.370 368.000 107.380 ;
        RECT 369.090 107.370 370.280 107.380 ;
        RECT 356.120 107.360 361.430 107.370 ;
        RECT 356.120 107.350 360.290 107.360 ;
        RECT 356.120 107.340 358.010 107.350 ;
        RECT 359.100 107.340 360.290 107.350 ;
        RECT 356.120 107.330 356.840 107.340 ;
        RECT 352.750 106.980 353.060 107.320 ;
        RECT 348.760 106.450 350.400 106.840 ;
        RECT 351.200 106.690 353.060 106.980 ;
        RECT 351.200 106.680 351.510 106.690 ;
        RECT 352.750 106.680 353.060 106.690 ;
        RECT 341.340 106.330 341.990 106.340 ;
        RECT 341.340 106.000 341.640 106.330 ;
        RECT 340.620 105.550 341.640 106.000 ;
        RECT 346.230 105.840 346.520 106.440 ;
        RECT 348.120 105.840 348.410 106.440 ;
        RECT 341.340 105.540 341.640 105.550 ;
        RECT 350.460 105.230 350.760 106.230 ;
        RECT 351.210 105.630 351.510 106.680 ;
        RECT 353.810 105.580 354.060 107.320 ;
        RECT 406.140 107.060 406.400 120.200 ;
        RECT 406.130 106.940 406.400 107.060 ;
        RECT 354.510 105.230 354.770 106.780 ;
        RECT 406.130 106.110 406.390 106.940 ;
        RECT 401.110 105.810 406.390 106.110 ;
        RECT 350.410 105.220 355.660 105.230 ;
        RECT 340.290 105.140 340.540 105.150 ;
        RECT 340.290 104.680 341.270 105.140 ;
        RECT 350.410 104.930 355.680 105.220 ;
        RECT 340.290 104.380 340.540 104.680 ;
        RECT 348.260 104.590 350.100 104.600 ;
        RECT 355.510 104.590 355.680 104.930 ;
        RECT 342.000 104.580 342.240 104.590 ;
        RECT 343.080 104.580 355.680 104.590 ;
        RECT 342.000 104.420 355.680 104.580 ;
        RECT 342.000 104.410 353.510 104.420 ;
        RECT 341.990 104.400 348.310 104.410 ;
        RECT 349.860 104.400 353.510 104.410 ;
        RECT 341.990 104.390 343.860 104.400 ;
        RECT 341.990 104.380 342.240 104.390 ;
        RECT 340.290 104.210 342.240 104.380 ;
        RECT 340.290 103.910 340.560 104.210 ;
        RECT 340.300 103.650 340.560 103.910 ;
        RECT 397.030 104.170 397.290 105.370 ;
        RECT 397.030 103.660 397.280 104.170 ;
        RECT 398.920 104.160 399.180 105.370 ;
        RECT 401.310 104.260 401.560 105.810 ;
        RECT 398.920 104.000 399.310 104.160 ;
        RECT 398.910 103.870 399.310 104.000 ;
        RECT 402.010 103.870 402.270 105.480 ;
        RECT 404.560 104.410 404.860 105.460 ;
        RECT 405.310 104.860 405.610 105.810 ;
        RECT 405.810 104.910 406.110 104.960 ;
        RECT 405.810 104.560 406.710 104.910 ;
        RECT 397.530 103.660 397.820 103.820 ;
        RECT 398.910 103.810 399.170 103.870 ;
        RECT 340.280 103.260 340.580 103.650 ;
        RECT 397.030 103.470 397.820 103.660 ;
        RECT 397.030 103.270 397.280 103.470 ;
        RECT 397.530 103.360 397.820 103.470 ;
        RECT 398.920 103.270 399.170 103.810 ;
        RECT 402.000 103.810 402.270 103.870 ;
        RECT 403.550 104.150 404.860 104.410 ;
        RECT 406.980 104.350 407.760 104.450 ;
        RECT 406.980 104.180 420.560 104.350 ;
        RECT 406.980 104.170 420.550 104.180 ;
        RECT 406.980 104.150 407.760 104.170 ;
        RECT 403.550 103.810 403.860 104.150 ;
        RECT 399.560 103.280 401.200 103.670 ;
        RECT 402.000 103.520 403.860 103.810 ;
        RECT 402.000 103.510 402.310 103.520 ;
        RECT 403.550 103.510 403.860 103.520 ;
        RECT 340.280 103.030 341.770 103.260 ;
        RECT 341.520 102.100 341.770 103.030 ;
        RECT 397.030 102.670 397.320 103.270 ;
        RECT 398.920 102.670 399.210 103.270 ;
        RECT 340.720 101.640 341.770 102.100 ;
        RECT 401.260 102.060 401.560 103.060 ;
        RECT 402.010 102.460 402.310 103.510 ;
        RECT 404.610 102.410 404.860 104.150 ;
        RECT 405.310 102.060 405.570 103.610 ;
        RECT 401.210 101.760 406.480 102.060 ;
        RECT 341.520 101.630 341.770 101.640 ;
        RECT 340.390 101.230 340.640 101.240 ;
        RECT 340.390 100.780 341.370 101.230 ;
        RECT 342.480 100.970 351.750 100.980 ;
        RECT 353.630 100.970 355.550 100.980 ;
        RECT 342.480 100.780 355.550 100.970 ;
        RECT 340.390 100.170 340.640 100.780 ;
        RECT 342.480 100.770 354.840 100.780 ;
        RECT 340.390 99.920 341.600 100.170 ;
        RECT 341.330 99.170 341.590 99.920 ;
        RECT 342.480 99.760 342.690 100.770 ;
        RECT 351.740 100.760 353.640 100.770 ;
        RECT 355.370 100.030 355.550 100.780 ;
        RECT 341.330 98.570 341.580 99.170 ;
        RECT 342.480 98.750 342.680 99.760 ;
        RECT 350.290 99.730 355.550 100.030 ;
        RECT 340.540 98.120 341.580 98.570 ;
        RECT 340.520 96.670 341.480 97.120 ;
        RECT 341.230 96.620 341.480 96.670 ;
        RECT 342.490 96.620 342.680 98.750 ;
        RECT 341.230 96.420 342.680 96.620 ;
        RECT 346.210 98.090 346.470 99.290 ;
        RECT 346.210 97.580 346.460 98.090 ;
        RECT 348.100 98.080 348.360 99.290 ;
        RECT 350.490 98.180 350.740 99.730 ;
        RECT 348.100 97.920 348.490 98.080 ;
        RECT 348.090 97.790 348.490 97.920 ;
        RECT 351.190 97.790 351.450 99.400 ;
        RECT 353.740 98.330 354.040 99.380 ;
        RECT 354.490 98.780 354.790 99.730 ;
        RECT 354.990 98.830 355.290 98.880 ;
        RECT 354.990 98.480 355.890 98.830 ;
        RECT 357.600 98.700 357.820 98.710 ;
        RECT 357.600 98.510 371.280 98.700 ;
        RECT 357.600 98.380 357.820 98.510 ;
        RECT 346.710 97.580 347.000 97.740 ;
        RECT 348.090 97.730 348.350 97.790 ;
        RECT 346.210 97.390 347.000 97.580 ;
        RECT 346.210 97.190 346.460 97.390 ;
        RECT 346.710 97.280 347.000 97.390 ;
        RECT 348.100 97.190 348.350 97.730 ;
        RECT 351.180 97.730 351.450 97.790 ;
        RECT 352.730 98.070 354.040 98.330 ;
        RECT 356.140 98.080 357.820 98.380 ;
        RECT 356.140 98.070 357.800 98.080 ;
        RECT 352.730 97.730 353.040 98.070 ;
        RECT 348.740 97.200 350.380 97.590 ;
        RECT 351.180 97.440 353.040 97.730 ;
        RECT 351.180 97.430 351.490 97.440 ;
        RECT 352.730 97.430 353.040 97.440 ;
        RECT 346.210 96.590 346.500 97.190 ;
        RECT 348.100 96.590 348.390 97.190 ;
        RECT 341.230 96.330 341.480 96.420 ;
        RECT 340.500 95.880 341.480 96.330 ;
        RECT 350.440 95.980 350.740 96.980 ;
        RECT 351.190 96.380 351.490 97.430 ;
        RECT 353.790 96.330 354.040 98.070 ;
        RECT 371.030 97.610 371.280 98.510 ;
        RECT 354.490 95.980 354.750 97.530 ;
        RECT 365.970 97.310 371.280 97.610 ;
        RECT 350.390 95.960 355.640 95.980 ;
        RECT 350.390 95.680 355.760 95.960 ;
        RECT 343.840 95.280 344.120 95.350 ;
        RECT 345.020 95.310 345.300 95.340 ;
        RECT 355.470 95.310 355.760 95.680 ;
        RECT 345.020 95.300 355.760 95.310 ;
        RECT 342.430 95.080 344.120 95.280 ;
        RECT 341.220 94.880 341.500 94.890 ;
        RECT 340.480 94.430 341.500 94.880 ;
        RECT 342.430 94.430 342.660 95.080 ;
        RECT 343.840 95.020 344.120 95.080 ;
        RECT 345.000 95.070 355.760 95.300 ;
        RECT 345.020 95.060 355.760 95.070 ;
        RECT 361.890 95.670 362.150 96.870 ;
        RECT 361.890 95.160 362.140 95.670 ;
        RECT 363.780 95.660 364.040 96.870 ;
        RECT 366.170 95.760 366.420 97.310 ;
        RECT 363.780 95.500 364.170 95.660 ;
        RECT 363.770 95.370 364.170 95.500 ;
        RECT 366.870 95.370 367.130 96.980 ;
        RECT 369.420 95.910 369.720 96.960 ;
        RECT 370.170 96.360 370.470 97.310 ;
        RECT 370.670 96.410 370.970 96.460 ;
        RECT 370.670 96.060 371.570 96.410 ;
        RECT 384.330 96.010 388.800 96.040 ;
        RECT 373.390 95.980 388.800 96.010 ;
        RECT 372.720 95.960 388.800 95.980 ;
        RECT 362.390 95.160 362.680 95.320 ;
        RECT 363.770 95.310 364.030 95.370 ;
        RECT 345.020 95.050 355.720 95.060 ;
        RECT 345.020 95.010 345.300 95.050 ;
        RECT 361.890 94.970 362.680 95.160 ;
        RECT 361.890 94.770 362.140 94.970 ;
        RECT 362.390 94.860 362.680 94.970 ;
        RECT 363.780 94.770 364.030 95.310 ;
        RECT 366.860 95.310 367.130 95.370 ;
        RECT 368.410 95.650 369.720 95.910 ;
        RECT 368.410 95.310 368.720 95.650 ;
        RECT 364.420 94.780 366.060 95.170 ;
        RECT 366.860 95.020 368.720 95.310 ;
        RECT 366.860 95.010 367.170 95.020 ;
        RECT 368.410 95.010 368.720 95.020 ;
        RECT 343.820 94.450 344.090 94.530 ;
        RECT 341.220 94.220 342.660 94.430 ;
        RECT 343.210 94.230 344.090 94.450 ;
        RECT 341.220 93.170 341.500 94.220 ;
        RECT 343.210 93.420 343.430 94.230 ;
        RECT 343.820 94.200 344.090 94.230 ;
        RECT 344.950 94.490 345.240 94.540 ;
        RECT 344.950 94.310 355.700 94.490 ;
        RECT 344.950 94.210 345.240 94.310 ;
        RECT 349.790 94.300 353.420 94.310 ;
        RECT 355.500 93.630 355.700 94.310 ;
        RECT 361.890 94.170 362.180 94.770 ;
        RECT 363.780 94.170 364.070 94.770 ;
        RECT 340.500 92.720 341.500 93.170 ;
        RECT 340.480 91.270 341.780 91.720 ;
        RECT 341.480 90.870 341.780 91.270 ;
        RECT 343.200 90.890 343.430 93.420 ;
        RECT 350.450 93.330 355.700 93.630 ;
        RECT 366.120 93.560 366.420 94.560 ;
        RECT 366.870 93.960 367.170 95.010 ;
        RECT 369.470 93.910 369.720 95.650 ;
        RECT 371.840 95.640 388.800 95.960 ;
        RECT 372.720 95.630 388.800 95.640 ;
        RECT 372.720 95.600 384.700 95.630 ;
        RECT 372.720 95.590 373.610 95.600 ;
        RECT 370.170 93.560 370.430 95.110 ;
        RECT 371.260 93.560 371.460 93.570 ;
        RECT 342.270 90.870 343.430 90.890 ;
        RECT 341.480 90.690 343.430 90.870 ;
        RECT 346.370 91.690 346.630 92.890 ;
        RECT 346.370 91.180 346.620 91.690 ;
        RECT 348.260 91.680 348.520 92.890 ;
        RECT 350.650 91.780 350.900 93.330 ;
        RECT 348.260 91.520 348.650 91.680 ;
        RECT 348.250 91.390 348.650 91.520 ;
        RECT 351.350 91.390 351.610 93.000 ;
        RECT 353.900 91.930 354.200 92.980 ;
        RECT 354.650 92.380 354.950 93.330 ;
        RECT 355.500 93.320 355.700 93.330 ;
        RECT 366.070 93.260 371.460 93.560 ;
        RECT 355.150 92.430 355.450 92.480 ;
        RECT 355.150 92.080 356.050 92.430 ;
        RECT 371.260 92.020 371.460 93.260 ;
        RECT 388.420 92.060 388.780 95.630 ;
        RECT 363.700 92.000 364.890 92.010 ;
        RECT 365.880 92.000 367.070 92.010 ;
        RECT 368.100 92.000 369.290 92.010 ;
        RECT 370.280 92.000 371.470 92.020 ;
        RECT 361.490 91.990 371.470 92.000 ;
        RECT 358.100 91.970 359.290 91.980 ;
        RECT 360.380 91.970 371.470 91.990 ;
        RECT 346.870 91.180 347.160 91.340 ;
        RECT 348.250 91.330 348.510 91.390 ;
        RECT 346.370 90.990 347.160 91.180 ;
        RECT 346.370 90.790 346.620 90.990 ;
        RECT 346.870 90.880 347.160 90.990 ;
        RECT 348.260 90.790 348.510 91.330 ;
        RECT 351.340 91.330 351.610 91.390 ;
        RECT 352.890 91.670 354.200 91.930 ;
        RECT 356.260 91.740 371.470 91.970 ;
        RECT 383.550 91.760 388.800 92.060 ;
        RECT 356.260 91.730 370.420 91.740 ;
        RECT 356.260 91.720 363.790 91.730 ;
        RECT 364.800 91.720 365.990 91.730 ;
        RECT 366.950 91.720 368.140 91.730 ;
        RECT 369.230 91.720 370.420 91.730 ;
        RECT 356.260 91.710 361.570 91.720 ;
        RECT 356.260 91.700 360.430 91.710 ;
        RECT 356.260 91.690 358.150 91.700 ;
        RECT 359.240 91.690 360.430 91.700 ;
        RECT 356.260 91.680 356.980 91.690 ;
        RECT 352.890 91.330 353.200 91.670 ;
        RECT 348.900 90.800 350.540 91.190 ;
        RECT 351.340 91.040 353.200 91.330 ;
        RECT 351.340 91.030 351.650 91.040 ;
        RECT 352.890 91.030 353.200 91.040 ;
        RECT 341.480 90.680 342.130 90.690 ;
        RECT 341.480 90.350 341.780 90.680 ;
        RECT 340.760 89.900 341.780 90.350 ;
        RECT 346.370 90.190 346.660 90.790 ;
        RECT 348.260 90.190 348.550 90.790 ;
        RECT 341.480 89.890 341.780 89.900 ;
        RECT 350.600 89.580 350.900 90.580 ;
        RECT 351.350 89.980 351.650 91.030 ;
        RECT 353.950 89.930 354.200 91.670 ;
        RECT 354.650 89.580 354.910 91.130 ;
        RECT 379.470 90.120 379.730 91.320 ;
        RECT 379.470 89.610 379.720 90.120 ;
        RECT 381.360 90.110 381.620 91.320 ;
        RECT 383.750 90.210 384.000 91.760 ;
        RECT 381.360 89.950 381.750 90.110 ;
        RECT 381.350 89.820 381.750 89.950 ;
        RECT 384.450 89.820 384.710 91.430 ;
        RECT 387.000 90.360 387.300 91.410 ;
        RECT 387.750 90.810 388.050 91.760 ;
        RECT 388.250 90.860 388.550 90.910 ;
        RECT 388.250 90.510 389.150 90.860 ;
        RECT 379.970 89.610 380.260 89.770 ;
        RECT 381.350 89.760 381.610 89.820 ;
        RECT 350.550 89.570 355.800 89.580 ;
        RECT 340.430 89.490 340.680 89.500 ;
        RECT 340.430 89.030 341.410 89.490 ;
        RECT 350.550 89.280 355.820 89.570 ;
        RECT 340.430 88.730 340.680 89.030 ;
        RECT 348.400 88.940 350.240 88.950 ;
        RECT 355.650 88.940 355.820 89.280 ;
        RECT 342.140 88.930 342.380 88.940 ;
        RECT 343.220 88.930 355.820 88.940 ;
        RECT 342.140 88.770 355.820 88.930 ;
        RECT 379.470 89.420 380.260 89.610 ;
        RECT 379.470 89.220 379.720 89.420 ;
        RECT 379.970 89.310 380.260 89.420 ;
        RECT 381.360 89.220 381.610 89.760 ;
        RECT 384.440 89.760 384.710 89.820 ;
        RECT 385.990 90.100 387.300 90.360 ;
        RECT 389.360 90.410 391.030 90.430 ;
        RECT 406.170 90.410 406.480 101.760 ;
        RECT 389.360 90.120 406.520 90.410 ;
        RECT 390.050 90.110 406.520 90.120 ;
        RECT 385.990 89.760 386.300 90.100 ;
        RECT 382.000 89.230 383.640 89.620 ;
        RECT 384.440 89.470 386.300 89.760 ;
        RECT 384.440 89.460 384.750 89.470 ;
        RECT 385.990 89.460 386.300 89.470 ;
        RECT 342.140 88.760 353.650 88.770 ;
        RECT 342.130 88.750 348.450 88.760 ;
        RECT 350.000 88.750 353.650 88.760 ;
        RECT 342.130 88.740 344.000 88.750 ;
        RECT 342.130 88.730 342.380 88.740 ;
        RECT 340.430 88.560 342.380 88.730 ;
        RECT 379.470 88.620 379.760 89.220 ;
        RECT 381.360 88.620 381.650 89.220 ;
        RECT 340.430 88.340 340.680 88.560 ;
        RECT 340.430 88.170 341.470 88.340 ;
        RECT 341.280 87.310 341.470 88.170 ;
        RECT 383.700 88.010 384.000 89.010 ;
        RECT 384.450 88.410 384.750 89.460 ;
        RECT 387.050 88.360 387.300 90.100 ;
        RECT 387.750 88.010 388.010 89.560 ;
        RECT 388.630 88.010 388.970 88.080 ;
        RECT 383.650 87.710 388.970 88.010 ;
        RECT 340.490 86.870 341.470 87.310 ;
        RECT 340.490 86.860 341.440 86.870 ;
        RECT 342.310 86.550 351.580 86.560 ;
        RECT 353.460 86.550 355.380 86.560 ;
        RECT 340.160 86.450 340.350 86.460 ;
        RECT 340.160 85.990 341.140 86.450 ;
        RECT 342.310 86.360 355.380 86.550 ;
        RECT 342.310 86.350 354.670 86.360 ;
        RECT 340.160 85.200 340.350 85.990 ;
        RECT 342.310 85.340 342.520 86.350 ;
        RECT 351.570 86.340 353.470 86.350 ;
        RECT 355.200 85.610 355.380 86.360 ;
        RECT 341.160 85.200 341.430 85.210 ;
        RECT 340.160 84.990 341.430 85.200 ;
        RECT 341.160 84.780 341.430 84.990 ;
        RECT 341.160 84.150 341.410 84.780 ;
        RECT 342.310 84.330 342.510 85.340 ;
        RECT 350.120 85.310 355.380 85.610 ;
        RECT 340.370 83.700 341.410 84.150 ;
        RECT 340.350 82.250 341.310 82.700 ;
        RECT 341.060 82.200 341.310 82.250 ;
        RECT 342.320 82.200 342.510 84.330 ;
        RECT 341.060 82.000 342.510 82.200 ;
        RECT 346.040 83.670 346.300 84.870 ;
        RECT 346.040 83.160 346.290 83.670 ;
        RECT 347.930 83.660 348.190 84.870 ;
        RECT 350.320 83.760 350.570 85.310 ;
        RECT 347.930 83.500 348.320 83.660 ;
        RECT 347.920 83.370 348.320 83.500 ;
        RECT 351.020 83.370 351.280 84.980 ;
        RECT 353.570 83.910 353.870 84.960 ;
        RECT 354.320 84.360 354.620 85.310 ;
        RECT 354.820 84.410 355.120 84.460 ;
        RECT 354.820 84.060 355.720 84.410 ;
        RECT 357.430 84.280 357.650 84.290 ;
        RECT 357.430 84.090 371.110 84.280 ;
        RECT 357.430 83.960 357.650 84.090 ;
        RECT 346.540 83.160 346.830 83.320 ;
        RECT 347.920 83.310 348.180 83.370 ;
        RECT 346.040 82.970 346.830 83.160 ;
        RECT 346.040 82.770 346.290 82.970 ;
        RECT 346.540 82.860 346.830 82.970 ;
        RECT 347.930 82.770 348.180 83.310 ;
        RECT 351.010 83.310 351.280 83.370 ;
        RECT 352.560 83.650 353.870 83.910 ;
        RECT 355.970 83.660 357.650 83.960 ;
        RECT 355.970 83.650 357.630 83.660 ;
        RECT 352.560 83.310 352.870 83.650 ;
        RECT 348.570 82.780 350.210 83.170 ;
        RECT 351.010 83.020 352.870 83.310 ;
        RECT 351.010 83.010 351.320 83.020 ;
        RECT 352.560 83.010 352.870 83.020 ;
        RECT 346.040 82.170 346.330 82.770 ;
        RECT 347.930 82.170 348.220 82.770 ;
        RECT 341.060 81.910 341.310 82.000 ;
        RECT 340.330 81.460 341.310 81.910 ;
        RECT 350.270 81.560 350.570 82.560 ;
        RECT 351.020 81.960 351.320 83.010 ;
        RECT 353.620 81.910 353.870 83.650 ;
        RECT 370.860 83.190 371.110 84.090 ;
        RECT 354.320 81.560 354.580 83.110 ;
        RECT 365.800 82.890 371.110 83.190 ;
        RECT 350.220 81.540 355.470 81.560 ;
        RECT 350.220 81.260 355.590 81.540 ;
        RECT 343.670 80.860 343.950 80.930 ;
        RECT 344.850 80.890 345.130 80.920 ;
        RECT 355.300 80.890 355.590 81.260 ;
        RECT 344.850 80.880 355.590 80.890 ;
        RECT 342.260 80.660 343.950 80.860 ;
        RECT 341.050 80.460 341.330 80.470 ;
        RECT 340.310 80.010 341.330 80.460 ;
        RECT 342.260 80.010 342.490 80.660 ;
        RECT 343.670 80.600 343.950 80.660 ;
        RECT 344.830 80.650 355.590 80.880 ;
        RECT 344.850 80.640 355.590 80.650 ;
        RECT 361.720 81.250 361.980 82.450 ;
        RECT 361.720 80.740 361.970 81.250 ;
        RECT 363.610 81.240 363.870 82.450 ;
        RECT 366.000 81.340 366.250 82.890 ;
        RECT 363.610 81.080 364.000 81.240 ;
        RECT 363.600 80.950 364.000 81.080 ;
        RECT 366.700 80.950 366.960 82.560 ;
        RECT 369.250 81.490 369.550 82.540 ;
        RECT 370.000 81.940 370.300 82.890 ;
        RECT 370.500 81.990 370.800 82.040 ;
        RECT 370.500 81.640 371.400 81.990 ;
        RECT 388.630 81.590 388.970 87.710 ;
        RECT 420.370 84.910 420.550 104.170 ;
        RECT 420.350 83.860 420.560 84.910 ;
        RECT 420.350 83.780 420.570 83.860 ;
        RECT 420.360 81.710 420.570 83.780 ;
        RECT 420.350 81.670 420.570 81.710 ;
        RECT 388.060 81.570 389.020 81.590 ;
        RECT 372.540 81.550 376.820 81.560 ;
        RECT 384.220 81.550 389.020 81.570 ;
        RECT 372.540 81.540 389.020 81.550 ;
        RECT 362.220 80.740 362.510 80.900 ;
        RECT 363.600 80.890 363.860 80.950 ;
        RECT 344.850 80.630 355.550 80.640 ;
        RECT 344.850 80.590 345.130 80.630 ;
        RECT 361.720 80.550 362.510 80.740 ;
        RECT 361.720 80.350 361.970 80.550 ;
        RECT 362.220 80.440 362.510 80.550 ;
        RECT 363.610 80.350 363.860 80.890 ;
        RECT 366.690 80.890 366.960 80.950 ;
        RECT 368.240 81.230 369.550 81.490 ;
        RECT 368.240 80.890 368.550 81.230 ;
        RECT 364.250 80.360 365.890 80.750 ;
        RECT 366.690 80.600 368.550 80.890 ;
        RECT 366.690 80.590 367.000 80.600 ;
        RECT 368.240 80.590 368.550 80.600 ;
        RECT 343.650 80.030 343.920 80.110 ;
        RECT 341.050 79.800 342.490 80.010 ;
        RECT 343.040 79.810 343.920 80.030 ;
        RECT 341.050 78.750 341.330 79.800 ;
        RECT 343.040 79.000 343.260 79.810 ;
        RECT 343.650 79.780 343.920 79.810 ;
        RECT 344.780 80.070 345.070 80.120 ;
        RECT 344.780 79.890 355.530 80.070 ;
        RECT 344.780 79.790 345.070 79.890 ;
        RECT 349.620 79.880 353.250 79.890 ;
        RECT 355.330 79.210 355.530 79.890 ;
        RECT 361.720 79.750 362.010 80.350 ;
        RECT 363.610 79.750 363.900 80.350 ;
        RECT 320.610 78.340 336.670 78.430 ;
        RECT 310.420 77.560 310.710 77.720 ;
        RECT 311.800 77.710 312.060 77.770 ;
        RECT 254.780 77.500 268.940 77.510 ;
        RECT 254.780 77.490 262.310 77.500 ;
        RECT 263.320 77.490 264.510 77.500 ;
        RECT 265.470 77.490 266.660 77.500 ;
        RECT 267.750 77.490 268.940 77.500 ;
        RECT 254.780 77.480 260.090 77.490 ;
        RECT 254.780 77.470 258.950 77.480 ;
        RECT 254.780 77.460 256.670 77.470 ;
        RECT 257.760 77.460 258.950 77.470 ;
        RECT 254.780 77.450 255.500 77.460 ;
        RECT 251.410 77.100 251.720 77.440 ;
        RECT 247.420 76.570 249.060 76.960 ;
        RECT 249.860 76.810 251.720 77.100 ;
        RECT 249.860 76.800 250.170 76.810 ;
        RECT 251.410 76.800 251.720 76.810 ;
        RECT 240.000 76.450 240.650 76.460 ;
        RECT 240.000 76.120 240.300 76.450 ;
        RECT 239.280 75.670 240.300 76.120 ;
        RECT 244.890 75.960 245.180 76.560 ;
        RECT 246.780 75.960 247.070 76.560 ;
        RECT 240.000 75.660 240.300 75.670 ;
        RECT 249.120 75.350 249.420 76.350 ;
        RECT 249.870 75.750 250.170 76.800 ;
        RECT 252.470 75.700 252.720 77.440 ;
        RECT 309.920 77.370 310.710 77.560 ;
        RECT 309.920 77.170 310.170 77.370 ;
        RECT 310.420 77.260 310.710 77.370 ;
        RECT 311.810 77.170 312.060 77.710 ;
        RECT 314.890 77.710 315.160 77.770 ;
        RECT 316.440 78.050 317.750 78.310 ;
        RECT 319.890 78.060 336.670 78.340 ;
        RECT 340.330 78.300 341.330 78.750 ;
        RECT 316.440 77.710 316.750 78.050 ;
        RECT 312.450 77.180 314.090 77.570 ;
        RECT 314.890 77.420 316.750 77.710 ;
        RECT 314.890 77.410 315.200 77.420 ;
        RECT 316.440 77.410 316.750 77.420 ;
        RECT 253.170 75.350 253.430 76.900 ;
        RECT 309.920 76.570 310.210 77.170 ;
        RECT 311.810 76.570 312.100 77.170 ;
        RECT 314.150 75.960 314.450 76.960 ;
        RECT 314.900 76.360 315.200 77.410 ;
        RECT 317.500 76.310 317.750 78.050 ;
        RECT 320.610 78.010 336.670 78.060 ;
        RECT 320.610 78.000 336.340 78.010 ;
        RECT 318.200 75.960 318.460 77.510 ;
        RECT 340.310 76.850 341.610 77.300 ;
        RECT 341.310 76.450 341.610 76.850 ;
        RECT 343.030 76.470 343.260 79.000 ;
        RECT 350.280 78.910 355.530 79.210 ;
        RECT 365.950 79.140 366.250 80.140 ;
        RECT 366.700 79.540 367.000 80.590 ;
        RECT 369.300 79.490 369.550 81.230 ;
        RECT 371.670 81.230 389.020 81.540 ;
        RECT 371.670 81.220 384.680 81.230 ;
        RECT 376.530 81.210 384.680 81.220 ;
        RECT 388.060 81.190 389.020 81.230 ;
        RECT 388.630 81.180 388.970 81.190 ;
        RECT 370.000 79.140 370.260 80.690 ;
        RECT 420.350 79.820 420.560 81.670 ;
        RECT 415.310 79.520 420.560 79.820 ;
        RECT 371.090 79.140 371.290 79.150 ;
        RECT 342.100 76.450 343.260 76.470 ;
        RECT 341.310 76.270 343.260 76.450 ;
        RECT 346.200 77.270 346.460 78.470 ;
        RECT 346.200 76.760 346.450 77.270 ;
        RECT 348.090 77.260 348.350 78.470 ;
        RECT 350.480 77.360 350.730 78.910 ;
        RECT 348.090 77.100 348.480 77.260 ;
        RECT 348.080 76.970 348.480 77.100 ;
        RECT 351.180 76.970 351.440 78.580 ;
        RECT 353.730 77.510 354.030 78.560 ;
        RECT 354.480 77.960 354.780 78.910 ;
        RECT 355.330 78.900 355.530 78.910 ;
        RECT 365.900 78.840 371.290 79.140 ;
        RECT 354.980 78.010 355.280 78.060 ;
        RECT 354.980 77.660 355.880 78.010 ;
        RECT 371.090 77.600 371.290 78.840 ;
        RECT 411.230 77.880 411.490 79.080 ;
        RECT 363.530 77.580 364.720 77.590 ;
        RECT 365.710 77.580 366.900 77.590 ;
        RECT 367.930 77.580 369.120 77.590 ;
        RECT 370.110 77.580 371.300 77.600 ;
        RECT 361.320 77.570 371.300 77.580 ;
        RECT 357.930 77.550 359.120 77.560 ;
        RECT 360.210 77.550 371.300 77.570 ;
        RECT 346.700 76.760 346.990 76.920 ;
        RECT 348.080 76.910 348.340 76.970 ;
        RECT 346.200 76.570 346.990 76.760 ;
        RECT 346.200 76.370 346.450 76.570 ;
        RECT 346.700 76.460 346.990 76.570 ;
        RECT 348.090 76.370 348.340 76.910 ;
        RECT 351.170 76.910 351.440 76.970 ;
        RECT 352.720 77.250 354.030 77.510 ;
        RECT 356.090 77.320 371.300 77.550 ;
        RECT 411.230 77.370 411.480 77.880 ;
        RECT 413.120 77.870 413.380 79.080 ;
        RECT 415.510 77.970 415.760 79.520 ;
        RECT 413.120 77.710 413.510 77.870 ;
        RECT 413.110 77.580 413.510 77.710 ;
        RECT 416.210 77.580 416.470 79.190 ;
        RECT 418.760 78.120 419.060 79.170 ;
        RECT 419.510 78.570 419.810 79.520 ;
        RECT 420.350 79.510 420.560 79.520 ;
        RECT 420.010 78.620 420.310 78.670 ;
        RECT 420.010 78.270 420.910 78.620 ;
        RECT 437.680 78.240 437.980 132.580 ;
        RECT 421.920 78.150 437.980 78.240 ;
        RECT 411.730 77.370 412.020 77.530 ;
        RECT 413.110 77.520 413.370 77.580 ;
        RECT 356.090 77.310 370.250 77.320 ;
        RECT 356.090 77.300 363.620 77.310 ;
        RECT 364.630 77.300 365.820 77.310 ;
        RECT 366.780 77.300 367.970 77.310 ;
        RECT 369.060 77.300 370.250 77.310 ;
        RECT 356.090 77.290 361.400 77.300 ;
        RECT 356.090 77.280 360.260 77.290 ;
        RECT 356.090 77.270 357.980 77.280 ;
        RECT 359.070 77.270 360.260 77.280 ;
        RECT 356.090 77.260 356.810 77.270 ;
        RECT 352.720 76.910 353.030 77.250 ;
        RECT 348.730 76.380 350.370 76.770 ;
        RECT 351.170 76.620 353.030 76.910 ;
        RECT 351.170 76.610 351.480 76.620 ;
        RECT 352.720 76.610 353.030 76.620 ;
        RECT 341.310 76.260 341.960 76.270 ;
        RECT 319.160 75.960 319.340 75.970 ;
        RECT 314.100 75.660 319.350 75.960 ;
        RECT 341.310 75.930 341.610 76.260 ;
        RECT 249.070 75.340 254.320 75.350 ;
        RECT 238.950 75.260 239.200 75.270 ;
        RECT 238.950 74.800 239.930 75.260 ;
        RECT 249.070 75.050 254.340 75.340 ;
        RECT 238.950 74.500 239.200 74.800 ;
        RECT 246.920 74.710 248.760 74.720 ;
        RECT 254.170 74.710 254.340 75.050 ;
        RECT 240.660 74.700 240.900 74.710 ;
        RECT 241.740 74.700 254.340 74.710 ;
        RECT 240.660 74.540 254.340 74.700 ;
        RECT 240.660 74.530 252.170 74.540 ;
        RECT 240.650 74.520 246.970 74.530 ;
        RECT 248.520 74.520 252.170 74.530 ;
        RECT 240.650 74.510 242.520 74.520 ;
        RECT 240.650 74.500 240.900 74.510 ;
        RECT 238.950 74.330 240.900 74.500 ;
        RECT 238.950 74.030 239.220 74.330 ;
        RECT 238.960 73.770 239.220 74.030 ;
        RECT 238.940 73.380 239.240 73.770 ;
        RECT 238.930 72.980 239.240 73.380 ;
        RECT 238.920 72.220 239.230 72.980 ;
        RECT 238.820 72.200 239.230 72.220 ;
        RECT 238.790 71.250 239.240 72.200 ;
        RECT 239.650 70.960 240.110 71.900 ;
        RECT 240.850 71.310 250.120 71.320 ;
        RECT 252.000 71.310 253.920 71.320 ;
        RECT 240.850 71.120 253.920 71.310 ;
        RECT 240.850 71.110 253.210 71.120 ;
        RECT 239.690 70.640 239.990 70.960 ;
        RECT 239.690 70.310 239.980 70.640 ;
        RECT 239.700 69.510 239.960 70.310 ;
        RECT 240.850 70.100 241.060 71.110 ;
        RECT 250.110 71.100 252.010 71.110 ;
        RECT 253.740 70.370 253.920 71.120 ;
        RECT 239.700 68.910 239.950 69.510 ;
        RECT 240.850 69.090 241.050 70.100 ;
        RECT 248.660 70.070 253.920 70.370 ;
        RECT 238.910 68.460 239.950 68.910 ;
        RECT 238.890 67.010 239.850 67.460 ;
        RECT 239.600 66.960 239.850 67.010 ;
        RECT 240.860 66.960 241.050 69.090 ;
        RECT 239.600 66.760 241.050 66.960 ;
        RECT 244.580 68.430 244.840 69.630 ;
        RECT 244.580 67.920 244.830 68.430 ;
        RECT 246.470 68.420 246.730 69.630 ;
        RECT 248.860 68.520 249.110 70.070 ;
        RECT 246.470 68.260 246.860 68.420 ;
        RECT 246.460 68.130 246.860 68.260 ;
        RECT 249.560 68.130 249.820 69.740 ;
        RECT 252.110 68.670 252.410 69.720 ;
        RECT 252.860 69.120 253.160 70.070 ;
        RECT 253.360 69.170 253.660 69.220 ;
        RECT 253.360 68.820 254.260 69.170 ;
        RECT 255.970 69.040 256.190 69.050 ;
        RECT 255.970 68.850 269.650 69.040 ;
        RECT 255.970 68.720 256.190 68.850 ;
        RECT 245.080 67.920 245.370 68.080 ;
        RECT 246.460 68.070 246.720 68.130 ;
        RECT 244.580 67.730 245.370 67.920 ;
        RECT 244.580 67.530 244.830 67.730 ;
        RECT 245.080 67.620 245.370 67.730 ;
        RECT 246.470 67.530 246.720 68.070 ;
        RECT 249.550 68.070 249.820 68.130 ;
        RECT 251.100 68.410 252.410 68.670 ;
        RECT 254.510 68.420 256.190 68.720 ;
        RECT 254.510 68.410 256.170 68.420 ;
        RECT 251.100 68.070 251.410 68.410 ;
        RECT 247.110 67.540 248.750 67.930 ;
        RECT 249.550 67.780 251.410 68.070 ;
        RECT 249.550 67.770 249.860 67.780 ;
        RECT 251.100 67.770 251.410 67.780 ;
        RECT 244.580 66.930 244.870 67.530 ;
        RECT 246.470 66.930 246.760 67.530 ;
        RECT 239.600 66.670 239.850 66.760 ;
        RECT 238.870 66.220 239.850 66.670 ;
        RECT 248.810 66.320 249.110 67.320 ;
        RECT 249.560 66.720 249.860 67.770 ;
        RECT 252.160 66.670 252.410 68.410 ;
        RECT 269.400 67.950 269.650 68.850 ;
        RECT 252.860 66.320 253.120 67.870 ;
        RECT 264.340 67.650 269.650 67.950 ;
        RECT 248.760 66.300 254.010 66.320 ;
        RECT 248.760 66.020 254.130 66.300 ;
        RECT 242.210 65.620 242.490 65.690 ;
        RECT 243.390 65.650 243.670 65.680 ;
        RECT 253.840 65.650 254.130 66.020 ;
        RECT 243.390 65.640 254.130 65.650 ;
        RECT 240.800 65.420 242.490 65.620 ;
        RECT 239.590 65.220 239.870 65.230 ;
        RECT 238.850 64.770 239.870 65.220 ;
        RECT 240.800 64.770 241.030 65.420 ;
        RECT 242.210 65.360 242.490 65.420 ;
        RECT 243.370 65.410 254.130 65.640 ;
        RECT 243.390 65.400 254.130 65.410 ;
        RECT 260.260 66.010 260.520 67.210 ;
        RECT 260.260 65.500 260.510 66.010 ;
        RECT 262.150 66.000 262.410 67.210 ;
        RECT 264.540 66.100 264.790 67.650 ;
        RECT 262.150 65.840 262.540 66.000 ;
        RECT 262.140 65.710 262.540 65.840 ;
        RECT 265.240 65.710 265.500 67.320 ;
        RECT 267.790 66.250 268.090 67.300 ;
        RECT 268.540 66.700 268.840 67.650 ;
        RECT 269.040 66.750 269.340 66.800 ;
        RECT 269.040 66.400 269.940 66.750 ;
        RECT 282.700 66.350 287.170 66.380 ;
        RECT 271.760 66.320 287.170 66.350 ;
        RECT 271.090 66.300 287.170 66.320 ;
        RECT 260.760 65.500 261.050 65.660 ;
        RECT 262.140 65.650 262.400 65.710 ;
        RECT 243.390 65.390 254.090 65.400 ;
        RECT 243.390 65.350 243.670 65.390 ;
        RECT 260.260 65.310 261.050 65.500 ;
        RECT 260.260 65.110 260.510 65.310 ;
        RECT 260.760 65.200 261.050 65.310 ;
        RECT 262.150 65.110 262.400 65.650 ;
        RECT 265.230 65.650 265.500 65.710 ;
        RECT 266.780 65.990 268.090 66.250 ;
        RECT 266.780 65.650 267.090 65.990 ;
        RECT 262.790 65.120 264.430 65.510 ;
        RECT 265.230 65.360 267.090 65.650 ;
        RECT 265.230 65.350 265.540 65.360 ;
        RECT 266.780 65.350 267.090 65.360 ;
        RECT 242.190 64.790 242.460 64.870 ;
        RECT 239.590 64.560 241.030 64.770 ;
        RECT 241.580 64.570 242.460 64.790 ;
        RECT 239.590 63.510 239.870 64.560 ;
        RECT 241.580 63.760 241.800 64.570 ;
        RECT 242.190 64.540 242.460 64.570 ;
        RECT 243.320 64.830 243.610 64.880 ;
        RECT 243.320 64.650 254.070 64.830 ;
        RECT 243.320 64.550 243.610 64.650 ;
        RECT 248.160 64.640 251.790 64.650 ;
        RECT 253.870 63.970 254.070 64.650 ;
        RECT 260.260 64.510 260.550 65.110 ;
        RECT 262.150 64.510 262.440 65.110 ;
        RECT 238.870 63.060 239.870 63.510 ;
        RECT 238.850 61.610 240.150 62.060 ;
        RECT 239.850 61.210 240.150 61.610 ;
        RECT 241.570 61.230 241.800 63.760 ;
        RECT 248.820 63.670 254.070 63.970 ;
        RECT 264.490 63.900 264.790 64.900 ;
        RECT 265.240 64.300 265.540 65.350 ;
        RECT 267.840 64.250 268.090 65.990 ;
        RECT 270.210 65.980 287.170 66.300 ;
        RECT 319.160 66.000 319.340 75.660 ;
        RECT 340.590 75.480 341.610 75.930 ;
        RECT 346.200 75.770 346.490 76.370 ;
        RECT 348.090 75.770 348.380 76.370 ;
        RECT 341.310 75.470 341.610 75.480 ;
        RECT 350.430 75.160 350.730 76.160 ;
        RECT 351.180 75.560 351.480 76.610 ;
        RECT 353.780 75.510 354.030 77.250 ;
        RECT 411.230 77.180 412.020 77.370 ;
        RECT 411.230 76.980 411.480 77.180 ;
        RECT 411.730 77.070 412.020 77.180 ;
        RECT 413.120 76.980 413.370 77.520 ;
        RECT 416.200 77.520 416.470 77.580 ;
        RECT 417.750 77.860 419.060 78.120 ;
        RECT 421.200 77.870 437.980 78.150 ;
        RECT 417.750 77.520 418.060 77.860 ;
        RECT 413.760 76.990 415.400 77.380 ;
        RECT 416.200 77.230 418.060 77.520 ;
        RECT 416.200 77.220 416.510 77.230 ;
        RECT 417.750 77.220 418.060 77.230 ;
        RECT 354.480 75.160 354.740 76.710 ;
        RECT 411.230 76.380 411.520 76.980 ;
        RECT 413.120 76.380 413.410 76.980 ;
        RECT 415.460 75.770 415.760 76.770 ;
        RECT 416.210 76.170 416.510 77.220 ;
        RECT 418.810 76.120 419.060 77.860 ;
        RECT 421.920 77.820 437.980 77.870 ;
        RECT 421.920 77.810 437.650 77.820 ;
        RECT 419.510 75.770 419.770 77.320 ;
        RECT 420.470 75.770 420.650 75.780 ;
        RECT 415.410 75.470 420.660 75.770 ;
        RECT 350.380 75.150 355.630 75.160 ;
        RECT 340.260 75.070 340.510 75.080 ;
        RECT 340.260 74.610 341.240 75.070 ;
        RECT 350.380 74.860 355.650 75.150 ;
        RECT 340.260 74.310 340.510 74.610 ;
        RECT 348.230 74.520 350.070 74.530 ;
        RECT 355.480 74.520 355.650 74.860 ;
        RECT 341.970 74.510 342.210 74.520 ;
        RECT 343.050 74.510 355.650 74.520 ;
        RECT 341.970 74.350 355.650 74.510 ;
        RECT 341.970 74.340 353.480 74.350 ;
        RECT 341.960 74.330 348.280 74.340 ;
        RECT 349.830 74.330 353.480 74.340 ;
        RECT 341.960 74.320 343.830 74.330 ;
        RECT 341.960 74.310 342.210 74.320 ;
        RECT 340.260 74.140 342.210 74.310 ;
        RECT 340.260 73.840 340.530 74.140 ;
        RECT 340.270 73.580 340.530 73.840 ;
        RECT 340.250 73.190 340.550 73.580 ;
        RECT 340.240 72.790 340.550 73.190 ;
        RECT 340.230 72.030 340.540 72.790 ;
        RECT 340.130 72.010 340.540 72.030 ;
        RECT 340.100 71.060 340.550 72.010 ;
        RECT 340.960 70.770 341.420 71.710 ;
        RECT 342.160 71.120 351.430 71.130 ;
        RECT 353.310 71.120 355.230 71.130 ;
        RECT 342.160 70.930 355.230 71.120 ;
        RECT 342.160 70.920 354.520 70.930 ;
        RECT 341.000 70.450 341.300 70.770 ;
        RECT 341.000 70.120 341.290 70.450 ;
        RECT 341.010 69.320 341.270 70.120 ;
        RECT 342.160 69.910 342.370 70.920 ;
        RECT 351.420 70.910 353.320 70.920 ;
        RECT 355.050 70.180 355.230 70.930 ;
        RECT 341.010 68.720 341.260 69.320 ;
        RECT 342.160 68.900 342.360 69.910 ;
        RECT 349.970 69.880 355.230 70.180 ;
        RECT 340.220 68.270 341.260 68.720 ;
        RECT 340.200 66.820 341.160 67.270 ;
        RECT 340.910 66.770 341.160 66.820 ;
        RECT 342.170 66.770 342.360 68.900 ;
        RECT 340.910 66.570 342.360 66.770 ;
        RECT 345.890 68.240 346.150 69.440 ;
        RECT 345.890 67.730 346.140 68.240 ;
        RECT 347.780 68.230 348.040 69.440 ;
        RECT 350.170 68.330 350.420 69.880 ;
        RECT 347.780 68.070 348.170 68.230 ;
        RECT 347.770 67.940 348.170 68.070 ;
        RECT 350.870 67.940 351.130 69.550 ;
        RECT 353.420 68.480 353.720 69.530 ;
        RECT 354.170 68.930 354.470 69.880 ;
        RECT 354.670 68.980 354.970 69.030 ;
        RECT 354.670 68.630 355.570 68.980 ;
        RECT 357.280 68.850 357.500 68.860 ;
        RECT 357.280 68.660 370.960 68.850 ;
        RECT 357.280 68.530 357.500 68.660 ;
        RECT 346.390 67.730 346.680 67.890 ;
        RECT 347.770 67.880 348.030 67.940 ;
        RECT 345.890 67.540 346.680 67.730 ;
        RECT 345.890 67.340 346.140 67.540 ;
        RECT 346.390 67.430 346.680 67.540 ;
        RECT 347.780 67.340 348.030 67.880 ;
        RECT 350.860 67.880 351.130 67.940 ;
        RECT 352.410 68.220 353.720 68.480 ;
        RECT 355.820 68.230 357.500 68.530 ;
        RECT 355.820 68.220 357.480 68.230 ;
        RECT 352.410 67.880 352.720 68.220 ;
        RECT 348.420 67.350 350.060 67.740 ;
        RECT 350.860 67.590 352.720 67.880 ;
        RECT 350.860 67.580 351.170 67.590 ;
        RECT 352.410 67.580 352.720 67.590 ;
        RECT 345.890 66.740 346.180 67.340 ;
        RECT 347.780 66.740 348.070 67.340 ;
        RECT 340.910 66.480 341.160 66.570 ;
        RECT 340.180 66.030 341.160 66.480 ;
        RECT 350.120 66.130 350.420 67.130 ;
        RECT 350.870 66.530 351.170 67.580 ;
        RECT 353.470 66.480 353.720 68.220 ;
        RECT 370.710 67.760 370.960 68.660 ;
        RECT 354.170 66.130 354.430 67.680 ;
        RECT 365.650 67.460 370.960 67.760 ;
        RECT 350.070 66.110 355.320 66.130 ;
        RECT 271.090 65.970 287.170 65.980 ;
        RECT 271.090 65.940 283.070 65.970 ;
        RECT 271.090 65.930 271.980 65.940 ;
        RECT 268.540 63.900 268.800 65.450 ;
        RECT 269.630 63.900 269.830 63.910 ;
        RECT 240.640 61.210 241.800 61.230 ;
        RECT 239.850 61.030 241.800 61.210 ;
        RECT 244.740 62.030 245.000 63.230 ;
        RECT 244.740 61.520 244.990 62.030 ;
        RECT 246.630 62.020 246.890 63.230 ;
        RECT 249.020 62.120 249.270 63.670 ;
        RECT 246.630 61.860 247.020 62.020 ;
        RECT 246.620 61.730 247.020 61.860 ;
        RECT 249.720 61.730 249.980 63.340 ;
        RECT 252.270 62.270 252.570 63.320 ;
        RECT 253.020 62.720 253.320 63.670 ;
        RECT 253.870 63.660 254.070 63.670 ;
        RECT 264.440 63.600 269.830 63.900 ;
        RECT 253.520 62.770 253.820 62.820 ;
        RECT 253.520 62.420 254.420 62.770 ;
        RECT 269.630 62.360 269.830 63.600 ;
        RECT 286.790 62.400 287.150 65.970 ;
        RECT 262.070 62.340 263.260 62.350 ;
        RECT 264.250 62.340 265.440 62.350 ;
        RECT 266.470 62.340 267.660 62.350 ;
        RECT 268.650 62.340 269.840 62.360 ;
        RECT 259.860 62.330 269.840 62.340 ;
        RECT 256.470 62.310 257.660 62.320 ;
        RECT 258.750 62.310 269.840 62.330 ;
        RECT 245.240 61.520 245.530 61.680 ;
        RECT 246.620 61.670 246.880 61.730 ;
        RECT 244.740 61.330 245.530 61.520 ;
        RECT 244.740 61.130 244.990 61.330 ;
        RECT 245.240 61.220 245.530 61.330 ;
        RECT 246.630 61.130 246.880 61.670 ;
        RECT 249.710 61.670 249.980 61.730 ;
        RECT 251.260 62.010 252.570 62.270 ;
        RECT 254.630 62.080 269.840 62.310 ;
        RECT 281.920 62.100 287.170 62.400 ;
        RECT 254.630 62.070 268.790 62.080 ;
        RECT 254.630 62.060 262.160 62.070 ;
        RECT 263.170 62.060 264.360 62.070 ;
        RECT 265.320 62.060 266.510 62.070 ;
        RECT 267.600 62.060 268.790 62.070 ;
        RECT 254.630 62.050 259.940 62.060 ;
        RECT 254.630 62.040 258.800 62.050 ;
        RECT 254.630 62.030 256.520 62.040 ;
        RECT 257.610 62.030 258.800 62.040 ;
        RECT 254.630 62.020 255.350 62.030 ;
        RECT 251.260 61.670 251.570 62.010 ;
        RECT 247.270 61.140 248.910 61.530 ;
        RECT 249.710 61.380 251.570 61.670 ;
        RECT 249.710 61.370 250.020 61.380 ;
        RECT 251.260 61.370 251.570 61.380 ;
        RECT 239.850 61.020 240.500 61.030 ;
        RECT 239.850 60.690 240.150 61.020 ;
        RECT 239.130 60.240 240.150 60.690 ;
        RECT 244.740 60.530 245.030 61.130 ;
        RECT 246.630 60.530 246.920 61.130 ;
        RECT 239.850 60.230 240.150 60.240 ;
        RECT 248.970 59.920 249.270 60.920 ;
        RECT 249.720 60.320 250.020 61.370 ;
        RECT 252.320 60.270 252.570 62.010 ;
        RECT 253.020 59.920 253.280 61.470 ;
        RECT 277.840 60.460 278.100 61.660 ;
        RECT 277.840 59.950 278.090 60.460 ;
        RECT 279.730 60.450 279.990 61.660 ;
        RECT 282.120 60.550 282.370 62.100 ;
        RECT 279.730 60.290 280.120 60.450 ;
        RECT 279.720 60.160 280.120 60.290 ;
        RECT 282.820 60.160 283.080 61.770 ;
        RECT 285.370 60.700 285.670 61.750 ;
        RECT 286.120 61.150 286.420 62.100 ;
        RECT 286.620 61.200 286.920 61.250 ;
        RECT 286.620 60.850 287.520 61.200 ;
        RECT 278.340 59.950 278.630 60.110 ;
        RECT 279.720 60.100 279.980 60.160 ;
        RECT 248.920 59.910 254.170 59.920 ;
        RECT 238.800 59.830 239.050 59.840 ;
        RECT 238.800 59.370 239.780 59.830 ;
        RECT 248.920 59.620 254.190 59.910 ;
        RECT 238.800 59.070 239.050 59.370 ;
        RECT 246.770 59.280 248.610 59.290 ;
        RECT 254.020 59.280 254.190 59.620 ;
        RECT 240.510 59.270 240.750 59.280 ;
        RECT 241.590 59.270 254.190 59.280 ;
        RECT 240.510 59.110 254.190 59.270 ;
        RECT 277.840 59.760 278.630 59.950 ;
        RECT 277.840 59.560 278.090 59.760 ;
        RECT 278.340 59.650 278.630 59.760 ;
        RECT 279.730 59.560 279.980 60.100 ;
        RECT 282.810 60.100 283.080 60.160 ;
        RECT 284.360 60.440 285.670 60.700 ;
        RECT 287.730 60.740 289.400 60.770 ;
        RECT 304.480 60.740 304.730 60.750 ;
        RECT 287.730 60.470 304.730 60.740 ;
        RECT 287.730 60.460 301.230 60.470 ;
        RECT 289.010 60.440 301.230 60.460 ;
        RECT 284.360 60.100 284.670 60.440 ;
        RECT 280.370 59.570 282.010 59.960 ;
        RECT 282.810 59.810 284.670 60.100 ;
        RECT 282.810 59.800 283.120 59.810 ;
        RECT 284.360 59.800 284.670 59.810 ;
        RECT 240.510 59.100 252.020 59.110 ;
        RECT 240.500 59.090 246.820 59.100 ;
        RECT 248.370 59.090 252.020 59.100 ;
        RECT 240.500 59.080 242.370 59.090 ;
        RECT 240.500 59.070 240.750 59.080 ;
        RECT 238.800 58.900 240.750 59.070 ;
        RECT 277.840 58.960 278.130 59.560 ;
        RECT 279.730 58.960 280.020 59.560 ;
        RECT 238.800 58.680 239.050 58.900 ;
        RECT 238.800 58.510 239.840 58.680 ;
        RECT 239.650 57.650 239.840 58.510 ;
        RECT 282.070 58.350 282.370 59.350 ;
        RECT 282.820 58.750 283.120 59.800 ;
        RECT 285.420 58.700 285.670 60.440 ;
        RECT 286.120 58.350 286.380 59.900 ;
        RECT 287.000 58.350 287.340 58.420 ;
        RECT 282.020 58.050 287.340 58.350 ;
        RECT 238.860 57.210 239.840 57.650 ;
        RECT 238.860 57.200 239.810 57.210 ;
        RECT 240.680 56.890 249.950 56.900 ;
        RECT 251.830 56.890 253.750 56.900 ;
        RECT 238.530 56.790 238.720 56.800 ;
        RECT 238.530 56.330 239.510 56.790 ;
        RECT 240.680 56.700 253.750 56.890 ;
        RECT 240.680 56.690 253.040 56.700 ;
        RECT 238.530 55.540 238.720 56.330 ;
        RECT 240.680 55.680 240.890 56.690 ;
        RECT 249.940 56.680 251.840 56.690 ;
        RECT 253.570 55.950 253.750 56.700 ;
        RECT 239.530 55.540 239.800 55.550 ;
        RECT 238.530 55.330 239.800 55.540 ;
        RECT 239.530 55.120 239.800 55.330 ;
        RECT 239.530 54.490 239.780 55.120 ;
        RECT 240.680 54.670 240.880 55.680 ;
        RECT 248.490 55.650 253.750 55.950 ;
        RECT 238.740 54.040 239.780 54.490 ;
        RECT 238.720 52.590 239.680 53.040 ;
        RECT 239.430 52.540 239.680 52.590 ;
        RECT 240.690 52.540 240.880 54.670 ;
        RECT 239.430 52.340 240.880 52.540 ;
        RECT 244.410 54.010 244.670 55.210 ;
        RECT 244.410 53.500 244.660 54.010 ;
        RECT 246.300 54.000 246.560 55.210 ;
        RECT 248.690 54.100 248.940 55.650 ;
        RECT 246.300 53.840 246.690 54.000 ;
        RECT 246.290 53.710 246.690 53.840 ;
        RECT 249.390 53.710 249.650 55.320 ;
        RECT 251.940 54.250 252.240 55.300 ;
        RECT 252.690 54.700 252.990 55.650 ;
        RECT 253.190 54.750 253.490 54.800 ;
        RECT 253.190 54.400 254.090 54.750 ;
        RECT 255.800 54.620 256.020 54.630 ;
        RECT 255.800 54.430 269.480 54.620 ;
        RECT 255.800 54.300 256.020 54.430 ;
        RECT 244.910 53.500 245.200 53.660 ;
        RECT 246.290 53.650 246.550 53.710 ;
        RECT 244.410 53.310 245.200 53.500 ;
        RECT 244.410 53.110 244.660 53.310 ;
        RECT 244.910 53.200 245.200 53.310 ;
        RECT 246.300 53.110 246.550 53.650 ;
        RECT 249.380 53.650 249.650 53.710 ;
        RECT 250.930 53.990 252.240 54.250 ;
        RECT 254.340 54.000 256.020 54.300 ;
        RECT 254.340 53.990 256.000 54.000 ;
        RECT 250.930 53.650 251.240 53.990 ;
        RECT 246.940 53.120 248.580 53.510 ;
        RECT 249.380 53.360 251.240 53.650 ;
        RECT 249.380 53.350 249.690 53.360 ;
        RECT 250.930 53.350 251.240 53.360 ;
        RECT 244.410 52.510 244.700 53.110 ;
        RECT 246.300 52.510 246.590 53.110 ;
        RECT 239.430 52.250 239.680 52.340 ;
        RECT 238.700 51.800 239.680 52.250 ;
        RECT 248.640 51.900 248.940 52.900 ;
        RECT 249.390 52.300 249.690 53.350 ;
        RECT 251.990 52.250 252.240 53.990 ;
        RECT 269.230 53.530 269.480 54.430 ;
        RECT 252.690 51.900 252.950 53.450 ;
        RECT 264.170 53.230 269.480 53.530 ;
        RECT 248.590 51.880 253.840 51.900 ;
        RECT 248.590 51.600 253.960 51.880 ;
        RECT 242.040 51.200 242.320 51.270 ;
        RECT 243.220 51.230 243.500 51.260 ;
        RECT 253.670 51.230 253.960 51.600 ;
        RECT 243.220 51.220 253.960 51.230 ;
        RECT 240.630 51.000 242.320 51.200 ;
        RECT 239.420 50.800 239.700 50.810 ;
        RECT 238.680 50.350 239.700 50.800 ;
        RECT 240.630 50.350 240.860 51.000 ;
        RECT 242.040 50.940 242.320 51.000 ;
        RECT 243.200 50.990 253.960 51.220 ;
        RECT 243.220 50.980 253.960 50.990 ;
        RECT 260.090 51.590 260.350 52.790 ;
        RECT 260.090 51.080 260.340 51.590 ;
        RECT 261.980 51.580 262.240 52.790 ;
        RECT 264.370 51.680 264.620 53.230 ;
        RECT 261.980 51.420 262.370 51.580 ;
        RECT 261.970 51.290 262.370 51.420 ;
        RECT 265.070 51.290 265.330 52.900 ;
        RECT 267.620 51.830 267.920 52.880 ;
        RECT 268.370 52.280 268.670 53.230 ;
        RECT 268.870 52.330 269.170 52.380 ;
        RECT 268.870 51.980 269.770 52.330 ;
        RECT 287.000 51.930 287.340 58.050 ;
        RECT 286.430 51.910 287.390 51.930 ;
        RECT 270.910 51.890 275.190 51.900 ;
        RECT 282.590 51.890 287.390 51.910 ;
        RECT 270.910 51.880 287.390 51.890 ;
        RECT 260.590 51.080 260.880 51.240 ;
        RECT 261.970 51.230 262.230 51.290 ;
        RECT 243.220 50.970 253.920 50.980 ;
        RECT 243.220 50.930 243.500 50.970 ;
        RECT 260.090 50.890 260.880 51.080 ;
        RECT 260.090 50.690 260.340 50.890 ;
        RECT 260.590 50.780 260.880 50.890 ;
        RECT 261.980 50.690 262.230 51.230 ;
        RECT 265.060 51.230 265.330 51.290 ;
        RECT 266.610 51.570 267.920 51.830 ;
        RECT 266.610 51.230 266.920 51.570 ;
        RECT 262.620 50.700 264.260 51.090 ;
        RECT 265.060 50.940 266.920 51.230 ;
        RECT 265.060 50.930 265.370 50.940 ;
        RECT 266.610 50.930 266.920 50.940 ;
        RECT 242.020 50.370 242.290 50.450 ;
        RECT 239.420 50.140 240.860 50.350 ;
        RECT 241.410 50.150 242.290 50.370 ;
        RECT 239.420 49.090 239.700 50.140 ;
        RECT 241.410 49.340 241.630 50.150 ;
        RECT 242.020 50.120 242.290 50.150 ;
        RECT 243.150 50.410 243.440 50.460 ;
        RECT 243.150 50.230 253.900 50.410 ;
        RECT 243.150 50.130 243.440 50.230 ;
        RECT 247.990 50.220 251.620 50.230 ;
        RECT 253.700 49.550 253.900 50.230 ;
        RECT 260.090 50.090 260.380 50.690 ;
        RECT 261.980 50.090 262.270 50.690 ;
        RECT 238.700 48.640 239.700 49.090 ;
        RECT 238.680 47.190 239.980 47.640 ;
        RECT 239.680 46.790 239.980 47.190 ;
        RECT 241.400 46.810 241.630 49.340 ;
        RECT 248.650 49.250 253.900 49.550 ;
        RECT 264.320 49.480 264.620 50.480 ;
        RECT 265.070 49.880 265.370 50.930 ;
        RECT 267.670 49.830 267.920 51.570 ;
        RECT 270.040 51.570 287.390 51.880 ;
        RECT 270.040 51.560 283.050 51.570 ;
        RECT 274.900 51.550 283.050 51.560 ;
        RECT 286.430 51.530 287.390 51.570 ;
        RECT 287.000 51.520 287.340 51.530 ;
        RECT 268.370 49.480 268.630 51.030 ;
        RECT 269.460 49.480 269.660 49.490 ;
        RECT 240.470 46.790 241.630 46.810 ;
        RECT 239.680 46.610 241.630 46.790 ;
        RECT 244.570 47.610 244.830 48.810 ;
        RECT 244.570 47.100 244.820 47.610 ;
        RECT 246.460 47.600 246.720 48.810 ;
        RECT 248.850 47.700 249.100 49.250 ;
        RECT 246.460 47.440 246.850 47.600 ;
        RECT 246.450 47.310 246.850 47.440 ;
        RECT 249.550 47.310 249.810 48.920 ;
        RECT 252.100 47.850 252.400 48.900 ;
        RECT 252.850 48.300 253.150 49.250 ;
        RECT 253.700 49.240 253.900 49.250 ;
        RECT 264.270 49.180 269.660 49.480 ;
        RECT 253.350 48.350 253.650 48.400 ;
        RECT 253.350 48.000 254.250 48.350 ;
        RECT 269.460 47.940 269.660 49.180 ;
        RECT 261.900 47.920 263.090 47.930 ;
        RECT 264.080 47.920 265.270 47.930 ;
        RECT 266.300 47.920 267.490 47.930 ;
        RECT 268.480 47.920 269.670 47.940 ;
        RECT 259.690 47.910 269.670 47.920 ;
        RECT 256.300 47.890 257.490 47.900 ;
        RECT 258.580 47.890 269.670 47.910 ;
        RECT 245.070 47.100 245.360 47.260 ;
        RECT 246.450 47.250 246.710 47.310 ;
        RECT 244.570 46.910 245.360 47.100 ;
        RECT 244.570 46.710 244.820 46.910 ;
        RECT 245.070 46.800 245.360 46.910 ;
        RECT 246.460 46.710 246.710 47.250 ;
        RECT 249.540 47.250 249.810 47.310 ;
        RECT 251.090 47.590 252.400 47.850 ;
        RECT 254.460 47.660 269.670 47.890 ;
        RECT 254.460 47.650 268.620 47.660 ;
        RECT 254.460 47.640 261.990 47.650 ;
        RECT 263.000 47.640 264.190 47.650 ;
        RECT 265.150 47.640 266.340 47.650 ;
        RECT 267.430 47.640 268.620 47.650 ;
        RECT 254.460 47.630 259.770 47.640 ;
        RECT 254.460 47.620 258.630 47.630 ;
        RECT 254.460 47.610 256.350 47.620 ;
        RECT 257.440 47.610 258.630 47.620 ;
        RECT 254.460 47.600 255.180 47.610 ;
        RECT 251.090 47.250 251.400 47.590 ;
        RECT 247.100 46.720 248.740 47.110 ;
        RECT 249.540 46.960 251.400 47.250 ;
        RECT 249.540 46.950 249.850 46.960 ;
        RECT 251.090 46.950 251.400 46.960 ;
        RECT 239.680 46.600 240.330 46.610 ;
        RECT 239.680 46.270 239.980 46.600 ;
        RECT 238.960 45.820 239.980 46.270 ;
        RECT 244.570 46.110 244.860 46.710 ;
        RECT 246.460 46.110 246.750 46.710 ;
        RECT 239.680 45.810 239.980 45.820 ;
        RECT 248.800 45.500 249.100 46.500 ;
        RECT 249.550 45.900 249.850 46.950 ;
        RECT 252.150 45.850 252.400 47.590 ;
        RECT 304.480 47.330 304.740 60.470 ;
        RECT 304.470 47.210 304.740 47.330 ;
        RECT 319.070 56.480 319.340 66.000 ;
        RECT 350.070 65.830 355.440 66.110 ;
        RECT 343.520 65.430 343.800 65.500 ;
        RECT 344.700 65.460 344.980 65.490 ;
        RECT 355.150 65.460 355.440 65.830 ;
        RECT 344.700 65.450 355.440 65.460 ;
        RECT 342.110 65.230 343.800 65.430 ;
        RECT 340.900 65.030 341.180 65.040 ;
        RECT 340.160 64.580 341.180 65.030 ;
        RECT 342.110 64.580 342.340 65.230 ;
        RECT 343.520 65.170 343.800 65.230 ;
        RECT 344.680 65.220 355.440 65.450 ;
        RECT 344.700 65.210 355.440 65.220 ;
        RECT 361.570 65.820 361.830 67.020 ;
        RECT 361.570 65.310 361.820 65.820 ;
        RECT 363.460 65.810 363.720 67.020 ;
        RECT 365.850 65.910 366.100 67.460 ;
        RECT 363.460 65.650 363.850 65.810 ;
        RECT 363.450 65.520 363.850 65.650 ;
        RECT 366.550 65.520 366.810 67.130 ;
        RECT 369.100 66.060 369.400 67.110 ;
        RECT 369.850 66.510 370.150 67.460 ;
        RECT 370.350 66.560 370.650 66.610 ;
        RECT 370.350 66.210 371.250 66.560 ;
        RECT 384.010 66.160 388.480 66.190 ;
        RECT 373.070 66.130 388.480 66.160 ;
        RECT 372.400 66.110 388.480 66.130 ;
        RECT 362.070 65.310 362.360 65.470 ;
        RECT 363.450 65.460 363.710 65.520 ;
        RECT 344.700 65.200 355.400 65.210 ;
        RECT 344.700 65.160 344.980 65.200 ;
        RECT 361.570 65.120 362.360 65.310 ;
        RECT 361.570 64.920 361.820 65.120 ;
        RECT 362.070 65.010 362.360 65.120 ;
        RECT 363.460 64.920 363.710 65.460 ;
        RECT 366.540 65.460 366.810 65.520 ;
        RECT 368.090 65.800 369.400 66.060 ;
        RECT 368.090 65.460 368.400 65.800 ;
        RECT 364.100 64.930 365.740 65.320 ;
        RECT 366.540 65.170 368.400 65.460 ;
        RECT 366.540 65.160 366.850 65.170 ;
        RECT 368.090 65.160 368.400 65.170 ;
        RECT 343.500 64.600 343.770 64.680 ;
        RECT 340.900 64.370 342.340 64.580 ;
        RECT 342.890 64.380 343.770 64.600 ;
        RECT 340.900 63.320 341.180 64.370 ;
        RECT 342.890 63.570 343.110 64.380 ;
        RECT 343.500 64.350 343.770 64.380 ;
        RECT 344.630 64.640 344.920 64.690 ;
        RECT 344.630 64.460 355.380 64.640 ;
        RECT 344.630 64.360 344.920 64.460 ;
        RECT 349.470 64.450 353.100 64.460 ;
        RECT 355.180 63.780 355.380 64.460 ;
        RECT 361.570 64.320 361.860 64.920 ;
        RECT 363.460 64.320 363.750 64.920 ;
        RECT 340.180 62.870 341.180 63.320 ;
        RECT 340.160 61.420 341.460 61.870 ;
        RECT 341.160 61.020 341.460 61.420 ;
        RECT 342.880 61.040 343.110 63.570 ;
        RECT 350.130 63.480 355.380 63.780 ;
        RECT 365.800 63.710 366.100 64.710 ;
        RECT 366.550 64.110 366.850 65.160 ;
        RECT 369.150 64.060 369.400 65.800 ;
        RECT 371.520 65.790 388.480 66.110 ;
        RECT 420.470 65.810 420.650 75.470 ;
        RECT 372.400 65.780 388.480 65.790 ;
        RECT 372.400 65.750 384.380 65.780 ;
        RECT 372.400 65.740 373.290 65.750 ;
        RECT 369.850 63.710 370.110 65.260 ;
        RECT 370.940 63.710 371.140 63.720 ;
        RECT 341.950 61.020 343.110 61.040 ;
        RECT 341.160 60.840 343.110 61.020 ;
        RECT 346.050 61.840 346.310 63.040 ;
        RECT 346.050 61.330 346.300 61.840 ;
        RECT 347.940 61.830 348.200 63.040 ;
        RECT 350.330 61.930 350.580 63.480 ;
        RECT 347.940 61.670 348.330 61.830 ;
        RECT 347.930 61.540 348.330 61.670 ;
        RECT 351.030 61.540 351.290 63.150 ;
        RECT 353.580 62.080 353.880 63.130 ;
        RECT 354.330 62.530 354.630 63.480 ;
        RECT 355.180 63.470 355.380 63.480 ;
        RECT 365.750 63.410 371.140 63.710 ;
        RECT 354.830 62.580 355.130 62.630 ;
        RECT 354.830 62.230 355.730 62.580 ;
        RECT 370.940 62.170 371.140 63.410 ;
        RECT 388.100 62.210 388.460 65.780 ;
        RECT 363.380 62.150 364.570 62.160 ;
        RECT 365.560 62.150 366.750 62.160 ;
        RECT 367.780 62.150 368.970 62.160 ;
        RECT 369.960 62.150 371.150 62.170 ;
        RECT 361.170 62.140 371.150 62.150 ;
        RECT 357.780 62.120 358.970 62.130 ;
        RECT 360.060 62.120 371.150 62.140 ;
        RECT 346.550 61.330 346.840 61.490 ;
        RECT 347.930 61.480 348.190 61.540 ;
        RECT 346.050 61.140 346.840 61.330 ;
        RECT 346.050 60.940 346.300 61.140 ;
        RECT 346.550 61.030 346.840 61.140 ;
        RECT 347.940 60.940 348.190 61.480 ;
        RECT 351.020 61.480 351.290 61.540 ;
        RECT 352.570 61.820 353.880 62.080 ;
        RECT 355.940 61.890 371.150 62.120 ;
        RECT 383.230 61.910 388.480 62.210 ;
        RECT 355.940 61.880 370.100 61.890 ;
        RECT 355.940 61.870 363.470 61.880 ;
        RECT 364.480 61.870 365.670 61.880 ;
        RECT 366.630 61.870 367.820 61.880 ;
        RECT 368.910 61.870 370.100 61.880 ;
        RECT 355.940 61.860 361.250 61.870 ;
        RECT 355.940 61.850 360.110 61.860 ;
        RECT 355.940 61.840 357.830 61.850 ;
        RECT 358.920 61.840 360.110 61.850 ;
        RECT 355.940 61.830 356.660 61.840 ;
        RECT 352.570 61.480 352.880 61.820 ;
        RECT 348.580 60.950 350.220 61.340 ;
        RECT 351.020 61.190 352.880 61.480 ;
        RECT 351.020 61.180 351.330 61.190 ;
        RECT 352.570 61.180 352.880 61.190 ;
        RECT 341.160 60.830 341.810 60.840 ;
        RECT 341.160 60.500 341.460 60.830 ;
        RECT 340.440 60.050 341.460 60.500 ;
        RECT 346.050 60.340 346.340 60.940 ;
        RECT 347.940 60.340 348.230 60.940 ;
        RECT 341.160 60.040 341.460 60.050 ;
        RECT 350.280 59.730 350.580 60.730 ;
        RECT 351.030 60.130 351.330 61.180 ;
        RECT 353.630 60.080 353.880 61.820 ;
        RECT 354.330 59.730 354.590 61.280 ;
        RECT 379.150 60.270 379.410 61.470 ;
        RECT 379.150 59.760 379.400 60.270 ;
        RECT 381.040 60.260 381.300 61.470 ;
        RECT 383.430 60.360 383.680 61.910 ;
        RECT 381.040 60.100 381.430 60.260 ;
        RECT 381.030 59.970 381.430 60.100 ;
        RECT 384.130 59.970 384.390 61.580 ;
        RECT 386.680 60.510 386.980 61.560 ;
        RECT 387.430 60.960 387.730 61.910 ;
        RECT 387.930 61.010 388.230 61.060 ;
        RECT 387.930 60.660 388.830 61.010 ;
        RECT 379.650 59.760 379.940 59.920 ;
        RECT 381.030 59.910 381.290 59.970 ;
        RECT 350.230 59.720 355.480 59.730 ;
        RECT 340.110 59.640 340.360 59.650 ;
        RECT 340.110 59.180 341.090 59.640 ;
        RECT 350.230 59.430 355.500 59.720 ;
        RECT 340.110 58.880 340.360 59.180 ;
        RECT 348.080 59.090 349.920 59.100 ;
        RECT 355.330 59.090 355.500 59.430 ;
        RECT 341.820 59.080 342.060 59.090 ;
        RECT 342.900 59.080 355.500 59.090 ;
        RECT 341.820 58.920 355.500 59.080 ;
        RECT 379.150 59.570 379.940 59.760 ;
        RECT 379.150 59.370 379.400 59.570 ;
        RECT 379.650 59.460 379.940 59.570 ;
        RECT 381.040 59.370 381.290 59.910 ;
        RECT 384.120 59.910 384.390 59.970 ;
        RECT 385.670 60.250 386.980 60.510 ;
        RECT 389.040 60.550 390.710 60.580 ;
        RECT 405.790 60.550 406.040 60.560 ;
        RECT 389.040 60.280 406.040 60.550 ;
        RECT 389.040 60.270 402.540 60.280 ;
        RECT 390.320 60.250 402.540 60.270 ;
        RECT 385.670 59.910 385.980 60.250 ;
        RECT 381.680 59.380 383.320 59.770 ;
        RECT 384.120 59.620 385.980 59.910 ;
        RECT 384.120 59.610 384.430 59.620 ;
        RECT 385.670 59.610 385.980 59.620 ;
        RECT 341.820 58.910 353.330 58.920 ;
        RECT 341.810 58.900 348.130 58.910 ;
        RECT 349.680 58.900 353.330 58.910 ;
        RECT 341.810 58.890 343.680 58.900 ;
        RECT 341.810 58.880 342.060 58.890 ;
        RECT 340.110 58.710 342.060 58.880 ;
        RECT 379.150 58.770 379.440 59.370 ;
        RECT 381.040 58.770 381.330 59.370 ;
        RECT 340.110 58.490 340.360 58.710 ;
        RECT 340.110 58.320 341.150 58.490 ;
        RECT 340.960 57.460 341.150 58.320 ;
        RECT 383.380 58.160 383.680 59.160 ;
        RECT 384.130 58.560 384.430 59.610 ;
        RECT 386.730 58.510 386.980 60.250 ;
        RECT 387.430 58.160 387.690 59.710 ;
        RECT 388.310 58.160 388.650 58.230 ;
        RECT 383.330 57.860 388.650 58.160 ;
        RECT 340.170 57.020 341.150 57.460 ;
        RECT 340.170 57.010 341.120 57.020 ;
        RECT 341.990 56.700 351.260 56.710 ;
        RECT 353.140 56.700 355.060 56.710 ;
        RECT 339.840 56.600 340.030 56.610 ;
        RECT 252.850 45.500 253.110 47.050 ;
        RECT 304.470 46.380 304.730 47.210 ;
        RECT 319.070 46.530 319.250 56.480 ;
        RECT 339.840 56.140 340.820 56.600 ;
        RECT 341.990 56.510 355.060 56.700 ;
        RECT 341.990 56.500 354.350 56.510 ;
        RECT 339.840 55.350 340.030 56.140 ;
        RECT 341.990 55.490 342.200 56.500 ;
        RECT 351.250 56.490 353.150 56.500 ;
        RECT 354.880 55.760 355.060 56.510 ;
        RECT 340.840 55.350 341.110 55.360 ;
        RECT 339.840 55.140 341.110 55.350 ;
        RECT 340.840 54.930 341.110 55.140 ;
        RECT 340.840 54.300 341.090 54.930 ;
        RECT 341.990 54.480 342.190 55.490 ;
        RECT 349.800 55.460 355.060 55.760 ;
        RECT 340.050 53.850 341.090 54.300 ;
        RECT 340.030 52.400 340.990 52.850 ;
        RECT 340.740 52.350 340.990 52.400 ;
        RECT 342.000 52.350 342.190 54.480 ;
        RECT 340.740 52.150 342.190 52.350 ;
        RECT 345.720 53.820 345.980 55.020 ;
        RECT 345.720 53.310 345.970 53.820 ;
        RECT 347.610 53.810 347.870 55.020 ;
        RECT 350.000 53.910 350.250 55.460 ;
        RECT 347.610 53.650 348.000 53.810 ;
        RECT 347.600 53.520 348.000 53.650 ;
        RECT 350.700 53.520 350.960 55.130 ;
        RECT 353.250 54.060 353.550 55.110 ;
        RECT 354.000 54.510 354.300 55.460 ;
        RECT 354.500 54.560 354.800 54.610 ;
        RECT 354.500 54.210 355.400 54.560 ;
        RECT 357.110 54.430 357.330 54.440 ;
        RECT 357.110 54.240 370.790 54.430 ;
        RECT 357.110 54.110 357.330 54.240 ;
        RECT 346.220 53.310 346.510 53.470 ;
        RECT 347.600 53.460 347.860 53.520 ;
        RECT 345.720 53.120 346.510 53.310 ;
        RECT 345.720 52.920 345.970 53.120 ;
        RECT 346.220 53.010 346.510 53.120 ;
        RECT 347.610 52.920 347.860 53.460 ;
        RECT 350.690 53.460 350.960 53.520 ;
        RECT 352.240 53.800 353.550 54.060 ;
        RECT 355.650 53.810 357.330 54.110 ;
        RECT 355.650 53.800 357.310 53.810 ;
        RECT 352.240 53.460 352.550 53.800 ;
        RECT 348.250 52.930 349.890 53.320 ;
        RECT 350.690 53.170 352.550 53.460 ;
        RECT 350.690 53.160 351.000 53.170 ;
        RECT 352.240 53.160 352.550 53.170 ;
        RECT 345.720 52.320 346.010 52.920 ;
        RECT 347.610 52.320 347.900 52.920 ;
        RECT 340.740 52.060 340.990 52.150 ;
        RECT 340.010 51.610 340.990 52.060 ;
        RECT 349.950 51.710 350.250 52.710 ;
        RECT 350.700 52.110 351.000 53.160 ;
        RECT 353.300 52.060 353.550 53.800 ;
        RECT 370.540 53.340 370.790 54.240 ;
        RECT 354.000 51.710 354.260 53.260 ;
        RECT 365.480 53.040 370.790 53.340 ;
        RECT 349.900 51.690 355.150 51.710 ;
        RECT 349.900 51.410 355.270 51.690 ;
        RECT 343.350 51.010 343.630 51.080 ;
        RECT 344.530 51.040 344.810 51.070 ;
        RECT 354.980 51.040 355.270 51.410 ;
        RECT 344.530 51.030 355.270 51.040 ;
        RECT 341.940 50.810 343.630 51.010 ;
        RECT 340.730 50.610 341.010 50.620 ;
        RECT 339.990 50.160 341.010 50.610 ;
        RECT 341.940 50.160 342.170 50.810 ;
        RECT 343.350 50.750 343.630 50.810 ;
        RECT 344.510 50.800 355.270 51.030 ;
        RECT 344.530 50.790 355.270 50.800 ;
        RECT 361.400 51.400 361.660 52.600 ;
        RECT 361.400 50.890 361.650 51.400 ;
        RECT 363.290 51.390 363.550 52.600 ;
        RECT 365.680 51.490 365.930 53.040 ;
        RECT 363.290 51.230 363.680 51.390 ;
        RECT 363.280 51.100 363.680 51.230 ;
        RECT 366.380 51.100 366.640 52.710 ;
        RECT 368.930 51.640 369.230 52.690 ;
        RECT 369.680 52.090 369.980 53.040 ;
        RECT 370.180 52.140 370.480 52.190 ;
        RECT 370.180 51.790 371.080 52.140 ;
        RECT 388.310 51.740 388.650 57.860 ;
        RECT 387.740 51.720 388.700 51.740 ;
        RECT 372.220 51.700 376.500 51.710 ;
        RECT 383.900 51.700 388.700 51.720 ;
        RECT 372.220 51.690 388.700 51.700 ;
        RECT 361.900 50.890 362.190 51.050 ;
        RECT 363.280 51.040 363.540 51.100 ;
        RECT 344.530 50.780 355.230 50.790 ;
        RECT 344.530 50.740 344.810 50.780 ;
        RECT 361.400 50.700 362.190 50.890 ;
        RECT 361.400 50.500 361.650 50.700 ;
        RECT 361.900 50.590 362.190 50.700 ;
        RECT 363.290 50.500 363.540 51.040 ;
        RECT 366.370 51.040 366.640 51.100 ;
        RECT 367.920 51.380 369.230 51.640 ;
        RECT 367.920 51.040 368.230 51.380 ;
        RECT 363.930 50.510 365.570 50.900 ;
        RECT 366.370 50.750 368.230 51.040 ;
        RECT 366.370 50.740 366.680 50.750 ;
        RECT 367.920 50.740 368.230 50.750 ;
        RECT 343.330 50.180 343.600 50.260 ;
        RECT 340.730 49.950 342.170 50.160 ;
        RECT 342.720 49.960 343.600 50.180 ;
        RECT 340.730 48.900 341.010 49.950 ;
        RECT 342.720 49.150 342.940 49.960 ;
        RECT 343.330 49.930 343.600 49.960 ;
        RECT 344.460 50.220 344.750 50.270 ;
        RECT 344.460 50.040 355.210 50.220 ;
        RECT 344.460 49.940 344.750 50.040 ;
        RECT 349.300 50.030 352.930 50.040 ;
        RECT 355.010 49.360 355.210 50.040 ;
        RECT 361.400 49.900 361.690 50.500 ;
        RECT 363.290 49.900 363.580 50.500 ;
        RECT 340.010 48.450 341.010 48.900 ;
        RECT 339.990 47.000 341.290 47.450 ;
        RECT 340.990 46.600 341.290 47.000 ;
        RECT 342.710 46.620 342.940 49.150 ;
        RECT 349.960 49.060 355.210 49.360 ;
        RECT 365.630 49.290 365.930 50.290 ;
        RECT 366.380 49.690 366.680 50.740 ;
        RECT 368.980 49.640 369.230 51.380 ;
        RECT 371.350 51.380 388.700 51.690 ;
        RECT 371.350 51.370 384.360 51.380 ;
        RECT 376.210 51.360 384.360 51.370 ;
        RECT 387.740 51.340 388.700 51.380 ;
        RECT 388.310 51.330 388.650 51.340 ;
        RECT 369.680 49.290 369.940 50.840 ;
        RECT 370.770 49.290 370.970 49.300 ;
        RECT 341.780 46.600 342.940 46.620 ;
        RECT 299.450 46.080 304.730 46.380 ;
        RECT 248.750 45.490 254.000 45.500 ;
        RECT 238.630 45.410 238.880 45.420 ;
        RECT 238.630 44.950 239.610 45.410 ;
        RECT 248.750 45.200 254.020 45.490 ;
        RECT 238.630 44.650 238.880 44.950 ;
        RECT 246.600 44.860 248.440 44.870 ;
        RECT 253.850 44.860 254.020 45.200 ;
        RECT 240.340 44.850 240.580 44.860 ;
        RECT 241.420 44.850 254.020 44.860 ;
        RECT 240.340 44.690 254.020 44.850 ;
        RECT 240.340 44.680 251.850 44.690 ;
        RECT 240.330 44.670 246.650 44.680 ;
        RECT 248.200 44.670 251.850 44.680 ;
        RECT 240.330 44.660 242.200 44.670 ;
        RECT 240.330 44.650 240.580 44.660 ;
        RECT 238.630 44.480 240.580 44.650 ;
        RECT 238.630 44.180 238.900 44.480 ;
        RECT 238.640 43.920 238.900 44.180 ;
        RECT 295.370 44.440 295.630 45.640 ;
        RECT 295.370 43.930 295.620 44.440 ;
        RECT 297.260 44.430 297.520 45.640 ;
        RECT 299.650 44.530 299.900 46.080 ;
        RECT 297.260 44.270 297.650 44.430 ;
        RECT 297.250 44.140 297.650 44.270 ;
        RECT 300.350 44.140 300.610 45.750 ;
        RECT 302.900 44.680 303.200 45.730 ;
        RECT 303.650 45.130 303.950 46.080 ;
        RECT 304.150 45.180 304.450 45.230 ;
        RECT 304.150 44.830 305.050 45.180 ;
        RECT 319.060 44.720 319.260 46.530 ;
        RECT 340.990 46.420 342.940 46.600 ;
        RECT 345.880 47.420 346.140 48.620 ;
        RECT 345.880 46.910 346.130 47.420 ;
        RECT 347.770 47.410 348.030 48.620 ;
        RECT 350.160 47.510 350.410 49.060 ;
        RECT 347.770 47.250 348.160 47.410 ;
        RECT 347.760 47.120 348.160 47.250 ;
        RECT 350.860 47.120 351.120 48.730 ;
        RECT 353.410 47.660 353.710 48.710 ;
        RECT 354.160 48.110 354.460 49.060 ;
        RECT 355.010 49.050 355.210 49.060 ;
        RECT 365.580 48.990 370.970 49.290 ;
        RECT 354.660 48.160 354.960 48.210 ;
        RECT 354.660 47.810 355.560 48.160 ;
        RECT 370.770 47.750 370.970 48.990 ;
        RECT 363.210 47.730 364.400 47.740 ;
        RECT 365.390 47.730 366.580 47.740 ;
        RECT 367.610 47.730 368.800 47.740 ;
        RECT 369.790 47.730 370.980 47.750 ;
        RECT 361.000 47.720 370.980 47.730 ;
        RECT 357.610 47.700 358.800 47.710 ;
        RECT 359.890 47.700 370.980 47.720 ;
        RECT 346.380 46.910 346.670 47.070 ;
        RECT 347.760 47.060 348.020 47.120 ;
        RECT 345.880 46.720 346.670 46.910 ;
        RECT 345.880 46.520 346.130 46.720 ;
        RECT 346.380 46.610 346.670 46.720 ;
        RECT 347.770 46.520 348.020 47.060 ;
        RECT 350.850 47.060 351.120 47.120 ;
        RECT 352.400 47.400 353.710 47.660 ;
        RECT 355.770 47.470 370.980 47.700 ;
        RECT 355.770 47.460 369.930 47.470 ;
        RECT 355.770 47.450 363.300 47.460 ;
        RECT 364.310 47.450 365.500 47.460 ;
        RECT 366.460 47.450 367.650 47.460 ;
        RECT 368.740 47.450 369.930 47.460 ;
        RECT 355.770 47.440 361.080 47.450 ;
        RECT 355.770 47.430 359.940 47.440 ;
        RECT 355.770 47.420 357.660 47.430 ;
        RECT 358.750 47.420 359.940 47.430 ;
        RECT 355.770 47.410 356.490 47.420 ;
        RECT 352.400 47.060 352.710 47.400 ;
        RECT 348.410 46.530 350.050 46.920 ;
        RECT 350.850 46.770 352.710 47.060 ;
        RECT 350.850 46.760 351.160 46.770 ;
        RECT 352.400 46.760 352.710 46.770 ;
        RECT 340.990 46.410 341.640 46.420 ;
        RECT 340.990 46.080 341.290 46.410 ;
        RECT 340.270 45.630 341.290 46.080 ;
        RECT 345.880 45.920 346.170 46.520 ;
        RECT 347.770 45.920 348.060 46.520 ;
        RECT 340.990 45.620 341.290 45.630 ;
        RECT 350.110 45.310 350.410 46.310 ;
        RECT 350.860 45.710 351.160 46.760 ;
        RECT 353.460 45.660 353.710 47.400 ;
        RECT 405.790 47.140 406.050 60.280 ;
        RECT 405.780 47.020 406.050 47.140 ;
        RECT 420.380 56.290 420.650 65.810 ;
        RECT 354.160 45.310 354.420 46.860 ;
        RECT 405.780 46.190 406.040 47.020 ;
        RECT 420.380 46.340 420.560 56.290 ;
        RECT 400.760 45.890 406.040 46.190 ;
        RECT 350.060 45.300 355.310 45.310 ;
        RECT 295.870 43.930 296.160 44.090 ;
        RECT 297.250 44.080 297.510 44.140 ;
        RECT 238.620 43.530 238.920 43.920 ;
        RECT 295.370 43.740 296.160 43.930 ;
        RECT 295.370 43.540 295.620 43.740 ;
        RECT 295.870 43.630 296.160 43.740 ;
        RECT 297.260 43.540 297.510 44.080 ;
        RECT 300.340 44.080 300.610 44.140 ;
        RECT 301.890 44.420 303.200 44.680 ;
        RECT 305.320 44.430 319.260 44.720 ;
        RECT 339.940 45.220 340.190 45.230 ;
        RECT 339.940 44.760 340.920 45.220 ;
        RECT 350.060 45.010 355.330 45.300 ;
        RECT 339.940 44.460 340.190 44.760 ;
        RECT 347.910 44.670 349.750 44.680 ;
        RECT 355.160 44.670 355.330 45.010 ;
        RECT 341.650 44.660 341.890 44.670 ;
        RECT 342.730 44.660 355.330 44.670 ;
        RECT 341.650 44.500 355.330 44.660 ;
        RECT 341.650 44.490 353.160 44.500 ;
        RECT 341.640 44.480 347.960 44.490 ;
        RECT 349.510 44.480 353.160 44.490 ;
        RECT 341.640 44.470 343.510 44.480 ;
        RECT 341.640 44.460 341.890 44.470 ;
        RECT 305.320 44.420 319.220 44.430 ;
        RECT 301.890 44.080 302.200 44.420 ;
        RECT 297.900 43.550 299.540 43.940 ;
        RECT 300.340 43.790 302.200 44.080 ;
        RECT 300.340 43.780 300.650 43.790 ;
        RECT 301.890 43.780 302.200 43.790 ;
        RECT 238.620 43.300 240.110 43.530 ;
        RECT 239.860 42.370 240.110 43.300 ;
        RECT 295.370 42.940 295.660 43.540 ;
        RECT 297.260 42.940 297.550 43.540 ;
        RECT 239.060 41.910 240.110 42.370 ;
        RECT 299.600 42.330 299.900 43.330 ;
        RECT 300.350 42.730 300.650 43.780 ;
        RECT 302.950 42.680 303.200 44.420 ;
        RECT 305.910 44.410 319.220 44.420 ;
        RECT 339.940 44.290 341.890 44.460 ;
        RECT 339.940 43.990 340.210 44.290 ;
        RECT 303.650 42.330 303.910 43.880 ;
        RECT 339.950 43.730 340.210 43.990 ;
        RECT 396.680 44.250 396.940 45.450 ;
        RECT 396.680 43.740 396.930 44.250 ;
        RECT 398.570 44.240 398.830 45.450 ;
        RECT 400.960 44.340 401.210 45.890 ;
        RECT 398.570 44.080 398.960 44.240 ;
        RECT 398.560 43.950 398.960 44.080 ;
        RECT 401.660 43.950 401.920 45.560 ;
        RECT 404.210 44.490 404.510 45.540 ;
        RECT 404.960 44.940 405.260 45.890 ;
        RECT 405.460 44.990 405.760 45.040 ;
        RECT 405.460 44.640 406.360 44.990 ;
        RECT 420.370 44.530 420.570 46.340 ;
        RECT 397.180 43.740 397.470 43.900 ;
        RECT 398.560 43.890 398.820 43.950 ;
        RECT 339.930 43.340 340.230 43.730 ;
        RECT 396.680 43.550 397.470 43.740 ;
        RECT 396.680 43.350 396.930 43.550 ;
        RECT 397.180 43.440 397.470 43.550 ;
        RECT 398.570 43.350 398.820 43.890 ;
        RECT 401.650 43.890 401.920 43.950 ;
        RECT 403.200 44.230 404.510 44.490 ;
        RECT 406.630 44.240 420.570 44.530 ;
        RECT 406.630 44.230 420.530 44.240 ;
        RECT 403.200 43.890 403.510 44.230 ;
        RECT 399.210 43.360 400.850 43.750 ;
        RECT 401.650 43.600 403.510 43.890 ;
        RECT 401.650 43.590 401.960 43.600 ;
        RECT 403.200 43.590 403.510 43.600 ;
        RECT 339.930 43.110 341.420 43.340 ;
        RECT 299.550 42.030 304.820 42.330 ;
        RECT 341.170 42.180 341.420 43.110 ;
        RECT 396.680 42.750 396.970 43.350 ;
        RECT 398.570 42.750 398.860 43.350 ;
        RECT 239.860 41.900 240.110 41.910 ;
        RECT 238.730 41.500 238.980 41.510 ;
        RECT 238.730 41.050 239.710 41.500 ;
        RECT 240.820 41.240 250.090 41.250 ;
        RECT 251.970 41.240 253.890 41.250 ;
        RECT 240.820 41.050 253.890 41.240 ;
        RECT 238.730 40.440 238.980 41.050 ;
        RECT 240.820 41.040 253.180 41.050 ;
        RECT 238.730 40.190 239.940 40.440 ;
        RECT 239.670 39.440 239.930 40.190 ;
        RECT 240.820 40.030 241.030 41.040 ;
        RECT 250.080 41.030 251.980 41.040 ;
        RECT 253.710 40.300 253.890 41.050 ;
        RECT 239.670 38.840 239.920 39.440 ;
        RECT 240.820 39.020 241.020 40.030 ;
        RECT 248.630 40.000 253.890 40.300 ;
        RECT 238.880 38.390 239.920 38.840 ;
        RECT 238.860 36.940 239.820 37.390 ;
        RECT 239.570 36.890 239.820 36.940 ;
        RECT 240.830 36.890 241.020 39.020 ;
        RECT 239.570 36.690 241.020 36.890 ;
        RECT 244.550 38.360 244.810 39.560 ;
        RECT 244.550 37.850 244.800 38.360 ;
        RECT 246.440 38.350 246.700 39.560 ;
        RECT 248.830 38.450 249.080 40.000 ;
        RECT 246.440 38.190 246.830 38.350 ;
        RECT 246.430 38.060 246.830 38.190 ;
        RECT 249.530 38.060 249.790 39.670 ;
        RECT 252.080 38.600 252.380 39.650 ;
        RECT 252.830 39.050 253.130 40.000 ;
        RECT 253.330 39.100 253.630 39.150 ;
        RECT 253.330 38.750 254.230 39.100 ;
        RECT 255.940 38.970 256.160 38.980 ;
        RECT 255.940 38.780 269.620 38.970 ;
        RECT 255.940 38.650 256.160 38.780 ;
        RECT 245.050 37.850 245.340 38.010 ;
        RECT 246.430 38.000 246.690 38.060 ;
        RECT 244.550 37.660 245.340 37.850 ;
        RECT 244.550 37.460 244.800 37.660 ;
        RECT 245.050 37.550 245.340 37.660 ;
        RECT 246.440 37.460 246.690 38.000 ;
        RECT 249.520 38.000 249.790 38.060 ;
        RECT 251.070 38.340 252.380 38.600 ;
        RECT 254.480 38.350 256.160 38.650 ;
        RECT 254.480 38.340 256.140 38.350 ;
        RECT 251.070 38.000 251.380 38.340 ;
        RECT 247.080 37.470 248.720 37.860 ;
        RECT 249.520 37.710 251.380 38.000 ;
        RECT 249.520 37.700 249.830 37.710 ;
        RECT 251.070 37.700 251.380 37.710 ;
        RECT 244.550 36.860 244.840 37.460 ;
        RECT 246.440 36.860 246.730 37.460 ;
        RECT 239.570 36.600 239.820 36.690 ;
        RECT 238.840 36.150 239.820 36.600 ;
        RECT 248.780 36.250 249.080 37.250 ;
        RECT 249.530 36.650 249.830 37.700 ;
        RECT 252.130 36.600 252.380 38.340 ;
        RECT 269.370 37.880 269.620 38.780 ;
        RECT 252.830 36.250 253.090 37.800 ;
        RECT 264.310 37.580 269.620 37.880 ;
        RECT 248.730 36.230 253.980 36.250 ;
        RECT 248.730 35.950 254.100 36.230 ;
        RECT 242.180 35.550 242.460 35.620 ;
        RECT 243.360 35.580 243.640 35.610 ;
        RECT 253.810 35.580 254.100 35.950 ;
        RECT 243.360 35.570 254.100 35.580 ;
        RECT 240.770 35.350 242.460 35.550 ;
        RECT 239.560 35.150 239.840 35.160 ;
        RECT 238.820 34.700 239.840 35.150 ;
        RECT 240.770 34.700 241.000 35.350 ;
        RECT 242.180 35.290 242.460 35.350 ;
        RECT 243.340 35.340 254.100 35.570 ;
        RECT 243.360 35.330 254.100 35.340 ;
        RECT 260.230 35.940 260.490 37.140 ;
        RECT 260.230 35.430 260.480 35.940 ;
        RECT 262.120 35.930 262.380 37.140 ;
        RECT 264.510 36.030 264.760 37.580 ;
        RECT 262.120 35.770 262.510 35.930 ;
        RECT 262.110 35.640 262.510 35.770 ;
        RECT 265.210 35.640 265.470 37.250 ;
        RECT 267.760 36.180 268.060 37.230 ;
        RECT 268.510 36.630 268.810 37.580 ;
        RECT 269.010 36.680 269.310 36.730 ;
        RECT 269.010 36.330 269.910 36.680 ;
        RECT 282.670 36.280 287.140 36.310 ;
        RECT 271.730 36.250 287.140 36.280 ;
        RECT 271.060 36.230 287.140 36.250 ;
        RECT 260.730 35.430 261.020 35.590 ;
        RECT 262.110 35.580 262.370 35.640 ;
        RECT 243.360 35.320 254.060 35.330 ;
        RECT 243.360 35.280 243.640 35.320 ;
        RECT 260.230 35.240 261.020 35.430 ;
        RECT 260.230 35.040 260.480 35.240 ;
        RECT 260.730 35.130 261.020 35.240 ;
        RECT 262.120 35.040 262.370 35.580 ;
        RECT 265.200 35.580 265.470 35.640 ;
        RECT 266.750 35.920 268.060 36.180 ;
        RECT 266.750 35.580 267.060 35.920 ;
        RECT 262.760 35.050 264.400 35.440 ;
        RECT 265.200 35.290 267.060 35.580 ;
        RECT 265.200 35.280 265.510 35.290 ;
        RECT 266.750 35.280 267.060 35.290 ;
        RECT 242.160 34.720 242.430 34.800 ;
        RECT 239.560 34.490 241.000 34.700 ;
        RECT 241.550 34.500 242.430 34.720 ;
        RECT 239.560 33.440 239.840 34.490 ;
        RECT 241.550 33.690 241.770 34.500 ;
        RECT 242.160 34.470 242.430 34.500 ;
        RECT 243.290 34.760 243.580 34.810 ;
        RECT 243.290 34.580 254.040 34.760 ;
        RECT 243.290 34.480 243.580 34.580 ;
        RECT 248.130 34.570 251.760 34.580 ;
        RECT 253.840 33.900 254.040 34.580 ;
        RECT 260.230 34.440 260.520 35.040 ;
        RECT 262.120 34.440 262.410 35.040 ;
        RECT 238.840 32.990 239.840 33.440 ;
        RECT 238.820 31.540 240.120 31.990 ;
        RECT 239.820 31.140 240.120 31.540 ;
        RECT 241.540 31.160 241.770 33.690 ;
        RECT 248.790 33.600 254.040 33.900 ;
        RECT 264.460 33.830 264.760 34.830 ;
        RECT 265.210 34.230 265.510 35.280 ;
        RECT 267.810 34.180 268.060 35.920 ;
        RECT 270.180 35.910 287.140 36.230 ;
        RECT 271.060 35.900 287.140 35.910 ;
        RECT 271.060 35.870 283.040 35.900 ;
        RECT 271.060 35.860 271.950 35.870 ;
        RECT 268.510 33.830 268.770 35.380 ;
        RECT 269.600 33.830 269.800 33.840 ;
        RECT 240.610 31.140 241.770 31.160 ;
        RECT 239.820 30.960 241.770 31.140 ;
        RECT 244.710 31.960 244.970 33.160 ;
        RECT 244.710 31.450 244.960 31.960 ;
        RECT 246.600 31.950 246.860 33.160 ;
        RECT 248.990 32.050 249.240 33.600 ;
        RECT 246.600 31.790 246.990 31.950 ;
        RECT 246.590 31.660 246.990 31.790 ;
        RECT 249.690 31.660 249.950 33.270 ;
        RECT 252.240 32.200 252.540 33.250 ;
        RECT 252.990 32.650 253.290 33.600 ;
        RECT 253.840 33.590 254.040 33.600 ;
        RECT 264.410 33.530 269.800 33.830 ;
        RECT 253.490 32.700 253.790 32.750 ;
        RECT 253.490 32.350 254.390 32.700 ;
        RECT 269.600 32.290 269.800 33.530 ;
        RECT 286.760 32.330 287.120 35.900 ;
        RECT 262.040 32.270 263.230 32.280 ;
        RECT 264.220 32.270 265.410 32.280 ;
        RECT 266.440 32.270 267.630 32.280 ;
        RECT 268.620 32.270 269.810 32.290 ;
        RECT 259.830 32.260 269.810 32.270 ;
        RECT 256.440 32.240 257.630 32.250 ;
        RECT 258.720 32.240 269.810 32.260 ;
        RECT 245.210 31.450 245.500 31.610 ;
        RECT 246.590 31.600 246.850 31.660 ;
        RECT 244.710 31.260 245.500 31.450 ;
        RECT 244.710 31.060 244.960 31.260 ;
        RECT 245.210 31.150 245.500 31.260 ;
        RECT 246.600 31.060 246.850 31.600 ;
        RECT 249.680 31.600 249.950 31.660 ;
        RECT 251.230 31.940 252.540 32.200 ;
        RECT 254.600 32.010 269.810 32.240 ;
        RECT 281.890 32.030 287.140 32.330 ;
        RECT 254.600 32.000 268.760 32.010 ;
        RECT 254.600 31.990 262.130 32.000 ;
        RECT 263.140 31.990 264.330 32.000 ;
        RECT 265.290 31.990 266.480 32.000 ;
        RECT 267.570 31.990 268.760 32.000 ;
        RECT 254.600 31.980 259.910 31.990 ;
        RECT 254.600 31.970 258.770 31.980 ;
        RECT 254.600 31.960 256.490 31.970 ;
        RECT 257.580 31.960 258.770 31.970 ;
        RECT 254.600 31.950 255.320 31.960 ;
        RECT 251.230 31.600 251.540 31.940 ;
        RECT 247.240 31.070 248.880 31.460 ;
        RECT 249.680 31.310 251.540 31.600 ;
        RECT 249.680 31.300 249.990 31.310 ;
        RECT 251.230 31.300 251.540 31.310 ;
        RECT 239.820 30.950 240.470 30.960 ;
        RECT 239.820 30.620 240.120 30.950 ;
        RECT 239.100 30.170 240.120 30.620 ;
        RECT 244.710 30.460 245.000 31.060 ;
        RECT 246.600 30.460 246.890 31.060 ;
        RECT 239.820 30.160 240.120 30.170 ;
        RECT 248.940 29.850 249.240 30.850 ;
        RECT 249.690 30.250 249.990 31.300 ;
        RECT 252.290 30.200 252.540 31.940 ;
        RECT 252.990 29.850 253.250 31.400 ;
        RECT 277.810 30.390 278.070 31.590 ;
        RECT 277.810 29.880 278.060 30.390 ;
        RECT 279.700 30.380 279.960 31.590 ;
        RECT 282.090 30.480 282.340 32.030 ;
        RECT 279.700 30.220 280.090 30.380 ;
        RECT 279.690 30.090 280.090 30.220 ;
        RECT 282.790 30.090 283.050 31.700 ;
        RECT 285.340 30.630 285.640 31.680 ;
        RECT 286.090 31.080 286.390 32.030 ;
        RECT 286.590 31.130 286.890 31.180 ;
        RECT 286.590 30.780 287.490 31.130 ;
        RECT 278.310 29.880 278.600 30.040 ;
        RECT 279.690 30.030 279.950 30.090 ;
        RECT 248.890 29.840 254.140 29.850 ;
        RECT 238.770 29.760 239.020 29.770 ;
        RECT 238.770 29.300 239.750 29.760 ;
        RECT 248.890 29.550 254.160 29.840 ;
        RECT 238.770 29.000 239.020 29.300 ;
        RECT 246.740 29.210 248.580 29.220 ;
        RECT 253.990 29.210 254.160 29.550 ;
        RECT 240.480 29.200 240.720 29.210 ;
        RECT 241.560 29.200 254.160 29.210 ;
        RECT 240.480 29.040 254.160 29.200 ;
        RECT 277.810 29.690 278.600 29.880 ;
        RECT 277.810 29.490 278.060 29.690 ;
        RECT 278.310 29.580 278.600 29.690 ;
        RECT 279.700 29.490 279.950 30.030 ;
        RECT 282.780 30.030 283.050 30.090 ;
        RECT 284.330 30.370 285.640 30.630 ;
        RECT 287.700 30.680 289.370 30.700 ;
        RECT 304.510 30.680 304.820 42.030 ;
        RECT 340.370 41.720 341.420 42.180 ;
        RECT 400.910 42.140 401.210 43.140 ;
        RECT 401.660 42.540 401.960 43.590 ;
        RECT 404.260 42.490 404.510 44.230 ;
        RECT 407.220 44.220 420.530 44.230 ;
        RECT 404.960 42.140 405.220 43.690 ;
        RECT 400.860 41.840 406.130 42.140 ;
        RECT 341.170 41.710 341.420 41.720 ;
        RECT 340.040 41.310 340.290 41.320 ;
        RECT 340.040 40.860 341.020 41.310 ;
        RECT 342.130 41.050 351.400 41.060 ;
        RECT 353.280 41.050 355.200 41.060 ;
        RECT 342.130 40.860 355.200 41.050 ;
        RECT 340.040 40.250 340.290 40.860 ;
        RECT 342.130 40.850 354.490 40.860 ;
        RECT 340.040 40.000 341.250 40.250 ;
        RECT 340.980 39.250 341.240 40.000 ;
        RECT 342.130 39.840 342.340 40.850 ;
        RECT 351.390 40.840 353.290 40.850 ;
        RECT 355.020 40.110 355.200 40.860 ;
        RECT 340.980 38.650 341.230 39.250 ;
        RECT 342.130 38.830 342.330 39.840 ;
        RECT 349.940 39.810 355.200 40.110 ;
        RECT 340.190 38.200 341.230 38.650 ;
        RECT 340.170 36.750 341.130 37.200 ;
        RECT 340.880 36.700 341.130 36.750 ;
        RECT 342.140 36.700 342.330 38.830 ;
        RECT 340.880 36.500 342.330 36.700 ;
        RECT 345.860 38.170 346.120 39.370 ;
        RECT 345.860 37.660 346.110 38.170 ;
        RECT 347.750 38.160 348.010 39.370 ;
        RECT 350.140 38.260 350.390 39.810 ;
        RECT 347.750 38.000 348.140 38.160 ;
        RECT 347.740 37.870 348.140 38.000 ;
        RECT 350.840 37.870 351.100 39.480 ;
        RECT 353.390 38.410 353.690 39.460 ;
        RECT 354.140 38.860 354.440 39.810 ;
        RECT 354.640 38.910 354.940 38.960 ;
        RECT 354.640 38.560 355.540 38.910 ;
        RECT 357.250 38.780 357.470 38.790 ;
        RECT 357.250 38.590 370.930 38.780 ;
        RECT 357.250 38.460 357.470 38.590 ;
        RECT 346.360 37.660 346.650 37.820 ;
        RECT 347.740 37.810 348.000 37.870 ;
        RECT 345.860 37.470 346.650 37.660 ;
        RECT 345.860 37.270 346.110 37.470 ;
        RECT 346.360 37.360 346.650 37.470 ;
        RECT 347.750 37.270 348.000 37.810 ;
        RECT 350.830 37.810 351.100 37.870 ;
        RECT 352.380 38.150 353.690 38.410 ;
        RECT 355.790 38.160 357.470 38.460 ;
        RECT 355.790 38.150 357.450 38.160 ;
        RECT 352.380 37.810 352.690 38.150 ;
        RECT 348.390 37.280 350.030 37.670 ;
        RECT 350.830 37.520 352.690 37.810 ;
        RECT 350.830 37.510 351.140 37.520 ;
        RECT 352.380 37.510 352.690 37.520 ;
        RECT 345.860 36.670 346.150 37.270 ;
        RECT 347.750 36.670 348.040 37.270 ;
        RECT 340.880 36.410 341.130 36.500 ;
        RECT 340.150 35.960 341.130 36.410 ;
        RECT 350.090 36.060 350.390 37.060 ;
        RECT 350.840 36.460 351.140 37.510 ;
        RECT 353.440 36.410 353.690 38.150 ;
        RECT 370.680 37.690 370.930 38.590 ;
        RECT 354.140 36.060 354.400 37.610 ;
        RECT 365.620 37.390 370.930 37.690 ;
        RECT 350.040 36.040 355.290 36.060 ;
        RECT 350.040 35.760 355.410 36.040 ;
        RECT 343.490 35.360 343.770 35.430 ;
        RECT 344.670 35.390 344.950 35.420 ;
        RECT 355.120 35.390 355.410 35.760 ;
        RECT 344.670 35.380 355.410 35.390 ;
        RECT 342.080 35.160 343.770 35.360 ;
        RECT 340.870 34.960 341.150 34.970 ;
        RECT 340.130 34.510 341.150 34.960 ;
        RECT 342.080 34.510 342.310 35.160 ;
        RECT 343.490 35.100 343.770 35.160 ;
        RECT 344.650 35.150 355.410 35.380 ;
        RECT 344.670 35.140 355.410 35.150 ;
        RECT 361.540 35.750 361.800 36.950 ;
        RECT 361.540 35.240 361.790 35.750 ;
        RECT 363.430 35.740 363.690 36.950 ;
        RECT 365.820 35.840 366.070 37.390 ;
        RECT 363.430 35.580 363.820 35.740 ;
        RECT 363.420 35.450 363.820 35.580 ;
        RECT 366.520 35.450 366.780 37.060 ;
        RECT 369.070 35.990 369.370 37.040 ;
        RECT 369.820 36.440 370.120 37.390 ;
        RECT 370.320 36.490 370.620 36.540 ;
        RECT 370.320 36.140 371.220 36.490 ;
        RECT 383.980 36.090 388.450 36.120 ;
        RECT 373.040 36.060 388.450 36.090 ;
        RECT 372.370 36.040 388.450 36.060 ;
        RECT 362.040 35.240 362.330 35.400 ;
        RECT 363.420 35.390 363.680 35.450 ;
        RECT 344.670 35.130 355.370 35.140 ;
        RECT 344.670 35.090 344.950 35.130 ;
        RECT 361.540 35.050 362.330 35.240 ;
        RECT 361.540 34.850 361.790 35.050 ;
        RECT 362.040 34.940 362.330 35.050 ;
        RECT 363.430 34.850 363.680 35.390 ;
        RECT 366.510 35.390 366.780 35.450 ;
        RECT 368.060 35.730 369.370 35.990 ;
        RECT 368.060 35.390 368.370 35.730 ;
        RECT 364.070 34.860 365.710 35.250 ;
        RECT 366.510 35.100 368.370 35.390 ;
        RECT 366.510 35.090 366.820 35.100 ;
        RECT 368.060 35.090 368.370 35.100 ;
        RECT 343.470 34.530 343.740 34.610 ;
        RECT 340.870 34.300 342.310 34.510 ;
        RECT 342.860 34.310 343.740 34.530 ;
        RECT 340.870 33.250 341.150 34.300 ;
        RECT 342.860 33.500 343.080 34.310 ;
        RECT 343.470 34.280 343.740 34.310 ;
        RECT 344.600 34.570 344.890 34.620 ;
        RECT 344.600 34.390 355.350 34.570 ;
        RECT 344.600 34.290 344.890 34.390 ;
        RECT 349.440 34.380 353.070 34.390 ;
        RECT 355.150 33.710 355.350 34.390 ;
        RECT 361.540 34.250 361.830 34.850 ;
        RECT 363.430 34.250 363.720 34.850 ;
        RECT 340.150 32.800 341.150 33.250 ;
        RECT 340.130 31.350 341.430 31.800 ;
        RECT 341.130 30.950 341.430 31.350 ;
        RECT 342.850 30.970 343.080 33.500 ;
        RECT 350.100 33.410 355.350 33.710 ;
        RECT 365.770 33.640 366.070 34.640 ;
        RECT 366.520 34.040 366.820 35.090 ;
        RECT 369.120 33.990 369.370 35.730 ;
        RECT 371.490 35.720 388.450 36.040 ;
        RECT 372.370 35.710 388.450 35.720 ;
        RECT 372.370 35.680 384.350 35.710 ;
        RECT 372.370 35.670 373.260 35.680 ;
        RECT 369.820 33.640 370.080 35.190 ;
        RECT 370.910 33.640 371.110 33.650 ;
        RECT 341.920 30.950 343.080 30.970 ;
        RECT 341.130 30.770 343.080 30.950 ;
        RECT 346.020 31.770 346.280 32.970 ;
        RECT 346.020 31.260 346.270 31.770 ;
        RECT 347.910 31.760 348.170 32.970 ;
        RECT 350.300 31.860 350.550 33.410 ;
        RECT 347.910 31.600 348.300 31.760 ;
        RECT 347.900 31.470 348.300 31.600 ;
        RECT 351.000 31.470 351.260 33.080 ;
        RECT 353.550 32.010 353.850 33.060 ;
        RECT 354.300 32.460 354.600 33.410 ;
        RECT 355.150 33.400 355.350 33.410 ;
        RECT 365.720 33.340 371.110 33.640 ;
        RECT 354.800 32.510 355.100 32.560 ;
        RECT 354.800 32.160 355.700 32.510 ;
        RECT 370.910 32.100 371.110 33.340 ;
        RECT 388.070 32.140 388.430 35.710 ;
        RECT 363.350 32.080 364.540 32.090 ;
        RECT 365.530 32.080 366.720 32.090 ;
        RECT 367.750 32.080 368.940 32.090 ;
        RECT 369.930 32.080 371.120 32.100 ;
        RECT 361.140 32.070 371.120 32.080 ;
        RECT 357.750 32.050 358.940 32.060 ;
        RECT 360.030 32.050 371.120 32.070 ;
        RECT 346.520 31.260 346.810 31.420 ;
        RECT 347.900 31.410 348.160 31.470 ;
        RECT 346.020 31.070 346.810 31.260 ;
        RECT 346.020 30.870 346.270 31.070 ;
        RECT 346.520 30.960 346.810 31.070 ;
        RECT 347.910 30.870 348.160 31.410 ;
        RECT 350.990 31.410 351.260 31.470 ;
        RECT 352.540 31.750 353.850 32.010 ;
        RECT 355.910 31.820 371.120 32.050 ;
        RECT 383.200 31.840 388.450 32.140 ;
        RECT 355.910 31.810 370.070 31.820 ;
        RECT 355.910 31.800 363.440 31.810 ;
        RECT 364.450 31.800 365.640 31.810 ;
        RECT 366.600 31.800 367.790 31.810 ;
        RECT 368.880 31.800 370.070 31.810 ;
        RECT 355.910 31.790 361.220 31.800 ;
        RECT 355.910 31.780 360.080 31.790 ;
        RECT 355.910 31.770 357.800 31.780 ;
        RECT 358.890 31.770 360.080 31.780 ;
        RECT 355.910 31.760 356.630 31.770 ;
        RECT 352.540 31.410 352.850 31.750 ;
        RECT 348.550 30.880 350.190 31.270 ;
        RECT 350.990 31.120 352.850 31.410 ;
        RECT 350.990 31.110 351.300 31.120 ;
        RECT 352.540 31.110 352.850 31.120 ;
        RECT 341.130 30.760 341.780 30.770 ;
        RECT 287.700 30.390 304.860 30.680 ;
        RECT 341.130 30.430 341.430 30.760 ;
        RECT 288.390 30.380 304.860 30.390 ;
        RECT 284.330 30.030 284.640 30.370 ;
        RECT 280.340 29.500 281.980 29.890 ;
        RECT 282.780 29.740 284.640 30.030 ;
        RECT 282.780 29.730 283.090 29.740 ;
        RECT 284.330 29.730 284.640 29.740 ;
        RECT 240.480 29.030 251.990 29.040 ;
        RECT 240.470 29.020 246.790 29.030 ;
        RECT 248.340 29.020 251.990 29.030 ;
        RECT 240.470 29.010 242.340 29.020 ;
        RECT 240.470 29.000 240.720 29.010 ;
        RECT 238.770 28.830 240.720 29.000 ;
        RECT 277.810 28.890 278.100 29.490 ;
        RECT 279.700 28.890 279.990 29.490 ;
        RECT 238.770 28.610 239.020 28.830 ;
        RECT 238.770 28.440 239.810 28.610 ;
        RECT 239.620 27.580 239.810 28.440 ;
        RECT 282.040 28.280 282.340 29.280 ;
        RECT 282.790 28.680 283.090 29.730 ;
        RECT 285.390 28.630 285.640 30.370 ;
        RECT 340.410 29.980 341.430 30.430 ;
        RECT 346.020 30.270 346.310 30.870 ;
        RECT 347.910 30.270 348.200 30.870 ;
        RECT 341.130 29.970 341.430 29.980 ;
        RECT 286.090 28.280 286.350 29.830 ;
        RECT 350.250 29.660 350.550 30.660 ;
        RECT 351.000 30.060 351.300 31.110 ;
        RECT 353.600 30.010 353.850 31.750 ;
        RECT 354.300 29.660 354.560 31.210 ;
        RECT 379.120 30.200 379.380 31.400 ;
        RECT 379.120 29.690 379.370 30.200 ;
        RECT 381.010 30.190 381.270 31.400 ;
        RECT 383.400 30.290 383.650 31.840 ;
        RECT 381.010 30.030 381.400 30.190 ;
        RECT 381.000 29.900 381.400 30.030 ;
        RECT 384.100 29.900 384.360 31.510 ;
        RECT 386.650 30.440 386.950 31.490 ;
        RECT 387.400 30.890 387.700 31.840 ;
        RECT 387.900 30.940 388.200 30.990 ;
        RECT 387.900 30.590 388.800 30.940 ;
        RECT 379.620 29.690 379.910 29.850 ;
        RECT 381.000 29.840 381.260 29.900 ;
        RECT 350.200 29.650 355.450 29.660 ;
        RECT 340.080 29.570 340.330 29.580 ;
        RECT 340.080 29.110 341.060 29.570 ;
        RECT 350.200 29.360 355.470 29.650 ;
        RECT 340.080 28.810 340.330 29.110 ;
        RECT 348.050 29.020 349.890 29.030 ;
        RECT 355.300 29.020 355.470 29.360 ;
        RECT 341.790 29.010 342.030 29.020 ;
        RECT 342.870 29.010 355.470 29.020 ;
        RECT 341.790 28.850 355.470 29.010 ;
        RECT 379.120 29.500 379.910 29.690 ;
        RECT 379.120 29.300 379.370 29.500 ;
        RECT 379.620 29.390 379.910 29.500 ;
        RECT 381.010 29.300 381.260 29.840 ;
        RECT 384.090 29.840 384.360 29.900 ;
        RECT 385.640 30.180 386.950 30.440 ;
        RECT 389.010 30.490 390.680 30.510 ;
        RECT 405.820 30.490 406.130 41.840 ;
        RECT 389.010 30.200 406.170 30.490 ;
        RECT 389.700 30.190 406.170 30.200 ;
        RECT 385.640 29.840 385.950 30.180 ;
        RECT 381.650 29.310 383.290 29.700 ;
        RECT 384.090 29.550 385.950 29.840 ;
        RECT 384.090 29.540 384.400 29.550 ;
        RECT 385.640 29.540 385.950 29.550 ;
        RECT 341.790 28.840 353.300 28.850 ;
        RECT 341.780 28.830 348.100 28.840 ;
        RECT 349.650 28.830 353.300 28.840 ;
        RECT 341.780 28.820 343.650 28.830 ;
        RECT 341.780 28.810 342.030 28.820 ;
        RECT 340.080 28.640 342.030 28.810 ;
        RECT 379.120 28.700 379.410 29.300 ;
        RECT 381.010 28.700 381.300 29.300 ;
        RECT 340.080 28.420 340.330 28.640 ;
        RECT 286.970 28.280 287.310 28.350 ;
        RECT 281.990 27.980 287.310 28.280 ;
        RECT 340.080 28.250 341.120 28.420 ;
        RECT 238.830 27.140 239.810 27.580 ;
        RECT 238.830 27.130 239.780 27.140 ;
        RECT 240.650 26.820 249.920 26.830 ;
        RECT 251.800 26.820 253.720 26.830 ;
        RECT 238.500 26.720 238.690 26.730 ;
        RECT 238.500 26.260 239.480 26.720 ;
        RECT 240.650 26.630 253.720 26.820 ;
        RECT 240.650 26.620 253.010 26.630 ;
        RECT 238.500 25.470 238.690 26.260 ;
        RECT 240.650 25.610 240.860 26.620 ;
        RECT 249.910 26.610 251.810 26.620 ;
        RECT 253.540 25.880 253.720 26.630 ;
        RECT 239.500 25.470 239.770 25.480 ;
        RECT 238.500 25.260 239.770 25.470 ;
        RECT 239.500 25.050 239.770 25.260 ;
        RECT 239.500 24.420 239.750 25.050 ;
        RECT 240.650 24.600 240.850 25.610 ;
        RECT 248.460 25.580 253.720 25.880 ;
        RECT 238.710 23.970 239.750 24.420 ;
        RECT 238.690 22.520 239.650 22.970 ;
        RECT 239.400 22.470 239.650 22.520 ;
        RECT 240.660 22.470 240.850 24.600 ;
        RECT 239.400 22.270 240.850 22.470 ;
        RECT 244.380 23.940 244.640 25.140 ;
        RECT 244.380 23.430 244.630 23.940 ;
        RECT 246.270 23.930 246.530 25.140 ;
        RECT 248.660 24.030 248.910 25.580 ;
        RECT 246.270 23.770 246.660 23.930 ;
        RECT 246.260 23.640 246.660 23.770 ;
        RECT 249.360 23.640 249.620 25.250 ;
        RECT 251.910 24.180 252.210 25.230 ;
        RECT 252.660 24.630 252.960 25.580 ;
        RECT 253.160 24.680 253.460 24.730 ;
        RECT 253.160 24.330 254.060 24.680 ;
        RECT 255.770 24.550 255.990 24.560 ;
        RECT 255.770 24.360 269.450 24.550 ;
        RECT 255.770 24.230 255.990 24.360 ;
        RECT 244.880 23.430 245.170 23.590 ;
        RECT 246.260 23.580 246.520 23.640 ;
        RECT 244.380 23.240 245.170 23.430 ;
        RECT 244.380 23.040 244.630 23.240 ;
        RECT 244.880 23.130 245.170 23.240 ;
        RECT 246.270 23.040 246.520 23.580 ;
        RECT 249.350 23.580 249.620 23.640 ;
        RECT 250.900 23.920 252.210 24.180 ;
        RECT 254.310 23.930 255.990 24.230 ;
        RECT 254.310 23.920 255.970 23.930 ;
        RECT 250.900 23.580 251.210 23.920 ;
        RECT 246.910 23.050 248.550 23.440 ;
        RECT 249.350 23.290 251.210 23.580 ;
        RECT 249.350 23.280 249.660 23.290 ;
        RECT 250.900 23.280 251.210 23.290 ;
        RECT 244.380 22.440 244.670 23.040 ;
        RECT 246.270 22.440 246.560 23.040 ;
        RECT 239.400 22.180 239.650 22.270 ;
        RECT 238.670 21.730 239.650 22.180 ;
        RECT 248.610 21.830 248.910 22.830 ;
        RECT 249.360 22.230 249.660 23.280 ;
        RECT 251.960 22.180 252.210 23.920 ;
        RECT 269.200 23.460 269.450 24.360 ;
        RECT 252.660 21.830 252.920 23.380 ;
        RECT 264.140 23.160 269.450 23.460 ;
        RECT 248.560 21.810 253.810 21.830 ;
        RECT 248.560 21.530 253.930 21.810 ;
        RECT 242.010 21.130 242.290 21.200 ;
        RECT 243.190 21.160 243.470 21.190 ;
        RECT 253.640 21.160 253.930 21.530 ;
        RECT 243.190 21.150 253.930 21.160 ;
        RECT 240.600 20.930 242.290 21.130 ;
        RECT 239.390 20.730 239.670 20.740 ;
        RECT 238.650 20.280 239.670 20.730 ;
        RECT 240.600 20.280 240.830 20.930 ;
        RECT 242.010 20.870 242.290 20.930 ;
        RECT 243.170 20.920 253.930 21.150 ;
        RECT 243.190 20.910 253.930 20.920 ;
        RECT 260.060 21.520 260.320 22.720 ;
        RECT 260.060 21.010 260.310 21.520 ;
        RECT 261.950 21.510 262.210 22.720 ;
        RECT 264.340 21.610 264.590 23.160 ;
        RECT 261.950 21.350 262.340 21.510 ;
        RECT 261.940 21.220 262.340 21.350 ;
        RECT 265.040 21.220 265.300 22.830 ;
        RECT 267.590 21.760 267.890 22.810 ;
        RECT 268.340 22.210 268.640 23.160 ;
        RECT 268.840 22.260 269.140 22.310 ;
        RECT 268.840 21.910 269.740 22.260 ;
        RECT 286.970 21.860 287.310 27.980 ;
        RECT 340.930 27.390 341.120 28.250 ;
        RECT 383.350 28.090 383.650 29.090 ;
        RECT 384.100 28.490 384.400 29.540 ;
        RECT 386.700 28.440 386.950 30.180 ;
        RECT 387.400 28.090 387.660 29.640 ;
        RECT 388.280 28.090 388.620 28.160 ;
        RECT 383.300 27.790 388.620 28.090 ;
        RECT 340.140 26.950 341.120 27.390 ;
        RECT 340.140 26.940 341.090 26.950 ;
        RECT 341.960 26.630 351.230 26.640 ;
        RECT 353.110 26.630 355.030 26.640 ;
        RECT 339.810 26.530 340.000 26.540 ;
        RECT 339.810 26.070 340.790 26.530 ;
        RECT 341.960 26.440 355.030 26.630 ;
        RECT 341.960 26.430 354.320 26.440 ;
        RECT 339.810 25.280 340.000 26.070 ;
        RECT 341.960 25.420 342.170 26.430 ;
        RECT 351.220 26.420 353.120 26.430 ;
        RECT 354.850 25.690 355.030 26.440 ;
        RECT 340.810 25.280 341.080 25.290 ;
        RECT 339.810 25.070 341.080 25.280 ;
        RECT 340.810 24.860 341.080 25.070 ;
        RECT 340.810 24.230 341.060 24.860 ;
        RECT 341.960 24.410 342.160 25.420 ;
        RECT 349.770 25.390 355.030 25.690 ;
        RECT 340.020 23.780 341.060 24.230 ;
        RECT 340.000 22.330 340.960 22.780 ;
        RECT 340.710 22.280 340.960 22.330 ;
        RECT 341.970 22.280 342.160 24.410 ;
        RECT 340.710 22.080 342.160 22.280 ;
        RECT 345.690 23.750 345.950 24.950 ;
        RECT 345.690 23.240 345.940 23.750 ;
        RECT 347.580 23.740 347.840 24.950 ;
        RECT 349.970 23.840 350.220 25.390 ;
        RECT 347.580 23.580 347.970 23.740 ;
        RECT 347.570 23.450 347.970 23.580 ;
        RECT 350.670 23.450 350.930 25.060 ;
        RECT 353.220 23.990 353.520 25.040 ;
        RECT 353.970 24.440 354.270 25.390 ;
        RECT 354.470 24.490 354.770 24.540 ;
        RECT 354.470 24.140 355.370 24.490 ;
        RECT 357.080 24.360 357.300 24.370 ;
        RECT 357.080 24.170 370.760 24.360 ;
        RECT 357.080 24.040 357.300 24.170 ;
        RECT 346.190 23.240 346.480 23.400 ;
        RECT 347.570 23.390 347.830 23.450 ;
        RECT 345.690 23.050 346.480 23.240 ;
        RECT 345.690 22.850 345.940 23.050 ;
        RECT 346.190 22.940 346.480 23.050 ;
        RECT 347.580 22.850 347.830 23.390 ;
        RECT 350.660 23.390 350.930 23.450 ;
        RECT 352.210 23.730 353.520 23.990 ;
        RECT 355.620 23.740 357.300 24.040 ;
        RECT 355.620 23.730 357.280 23.740 ;
        RECT 352.210 23.390 352.520 23.730 ;
        RECT 348.220 22.860 349.860 23.250 ;
        RECT 350.660 23.100 352.520 23.390 ;
        RECT 350.660 23.090 350.970 23.100 ;
        RECT 352.210 23.090 352.520 23.100 ;
        RECT 345.690 22.250 345.980 22.850 ;
        RECT 347.580 22.250 347.870 22.850 ;
        RECT 340.710 21.990 340.960 22.080 ;
        RECT 286.400 21.840 287.360 21.860 ;
        RECT 270.880 21.820 275.160 21.830 ;
        RECT 282.560 21.820 287.360 21.840 ;
        RECT 270.880 21.810 287.360 21.820 ;
        RECT 260.560 21.010 260.850 21.170 ;
        RECT 261.940 21.160 262.200 21.220 ;
        RECT 243.190 20.900 253.890 20.910 ;
        RECT 243.190 20.860 243.470 20.900 ;
        RECT 260.060 20.820 260.850 21.010 ;
        RECT 260.060 20.620 260.310 20.820 ;
        RECT 260.560 20.710 260.850 20.820 ;
        RECT 261.950 20.620 262.200 21.160 ;
        RECT 265.030 21.160 265.300 21.220 ;
        RECT 266.580 21.500 267.890 21.760 ;
        RECT 266.580 21.160 266.890 21.500 ;
        RECT 262.590 20.630 264.230 21.020 ;
        RECT 265.030 20.870 266.890 21.160 ;
        RECT 265.030 20.860 265.340 20.870 ;
        RECT 266.580 20.860 266.890 20.870 ;
        RECT 241.990 20.300 242.260 20.380 ;
        RECT 239.390 20.070 240.830 20.280 ;
        RECT 241.380 20.080 242.260 20.300 ;
        RECT 239.390 19.020 239.670 20.070 ;
        RECT 241.380 19.270 241.600 20.080 ;
        RECT 241.990 20.050 242.260 20.080 ;
        RECT 243.120 20.340 243.410 20.390 ;
        RECT 243.120 20.160 253.870 20.340 ;
        RECT 243.120 20.060 243.410 20.160 ;
        RECT 247.960 20.150 251.590 20.160 ;
        RECT 253.670 19.480 253.870 20.160 ;
        RECT 260.060 20.020 260.350 20.620 ;
        RECT 261.950 20.020 262.240 20.620 ;
        RECT 238.670 18.570 239.670 19.020 ;
        RECT 238.650 17.120 239.950 17.570 ;
        RECT 239.650 16.720 239.950 17.120 ;
        RECT 241.370 16.740 241.600 19.270 ;
        RECT 248.620 19.180 253.870 19.480 ;
        RECT 264.290 19.410 264.590 20.410 ;
        RECT 265.040 19.810 265.340 20.860 ;
        RECT 267.640 19.760 267.890 21.500 ;
        RECT 270.010 21.500 287.360 21.810 ;
        RECT 339.980 21.540 340.960 21.990 ;
        RECT 349.920 21.640 350.220 22.640 ;
        RECT 350.670 22.040 350.970 23.090 ;
        RECT 353.270 21.990 353.520 23.730 ;
        RECT 370.510 23.270 370.760 24.170 ;
        RECT 353.970 21.640 354.230 23.190 ;
        RECT 365.450 22.970 370.760 23.270 ;
        RECT 349.870 21.620 355.120 21.640 ;
        RECT 270.010 21.490 283.020 21.500 ;
        RECT 274.870 21.480 283.020 21.490 ;
        RECT 286.400 21.460 287.360 21.500 ;
        RECT 286.970 21.450 287.310 21.460 ;
        RECT 349.870 21.340 355.240 21.620 ;
        RECT 268.340 19.410 268.600 20.960 ;
        RECT 343.320 20.940 343.600 21.010 ;
        RECT 344.500 20.970 344.780 21.000 ;
        RECT 354.950 20.970 355.240 21.340 ;
        RECT 344.500 20.960 355.240 20.970 ;
        RECT 341.910 20.740 343.600 20.940 ;
        RECT 340.700 20.540 340.980 20.550 ;
        RECT 339.960 20.090 340.980 20.540 ;
        RECT 341.910 20.090 342.140 20.740 ;
        RECT 343.320 20.680 343.600 20.740 ;
        RECT 344.480 20.730 355.240 20.960 ;
        RECT 344.500 20.720 355.240 20.730 ;
        RECT 361.370 21.330 361.630 22.530 ;
        RECT 361.370 20.820 361.620 21.330 ;
        RECT 363.260 21.320 363.520 22.530 ;
        RECT 365.650 21.420 365.900 22.970 ;
        RECT 363.260 21.160 363.650 21.320 ;
        RECT 363.250 21.030 363.650 21.160 ;
        RECT 366.350 21.030 366.610 22.640 ;
        RECT 368.900 21.570 369.200 22.620 ;
        RECT 369.650 22.020 369.950 22.970 ;
        RECT 370.150 22.070 370.450 22.120 ;
        RECT 370.150 21.720 371.050 22.070 ;
        RECT 388.280 21.670 388.620 27.790 ;
        RECT 387.710 21.650 388.670 21.670 ;
        RECT 372.190 21.630 376.470 21.640 ;
        RECT 383.870 21.630 388.670 21.650 ;
        RECT 372.190 21.620 388.670 21.630 ;
        RECT 361.870 20.820 362.160 20.980 ;
        RECT 363.250 20.970 363.510 21.030 ;
        RECT 344.500 20.710 355.200 20.720 ;
        RECT 344.500 20.670 344.780 20.710 ;
        RECT 361.370 20.630 362.160 20.820 ;
        RECT 361.370 20.430 361.620 20.630 ;
        RECT 361.870 20.520 362.160 20.630 ;
        RECT 363.260 20.430 363.510 20.970 ;
        RECT 366.340 20.970 366.610 21.030 ;
        RECT 367.890 21.310 369.200 21.570 ;
        RECT 367.890 20.970 368.200 21.310 ;
        RECT 363.900 20.440 365.540 20.830 ;
        RECT 366.340 20.680 368.200 20.970 ;
        RECT 366.340 20.670 366.650 20.680 ;
        RECT 367.890 20.670 368.200 20.680 ;
        RECT 343.300 20.110 343.570 20.190 ;
        RECT 340.700 19.880 342.140 20.090 ;
        RECT 342.690 19.890 343.570 20.110 ;
        RECT 269.430 19.410 269.630 19.420 ;
        RECT 240.440 16.720 241.600 16.740 ;
        RECT 239.650 16.540 241.600 16.720 ;
        RECT 244.540 17.540 244.800 18.740 ;
        RECT 244.540 17.030 244.790 17.540 ;
        RECT 246.430 17.530 246.690 18.740 ;
        RECT 248.820 17.630 249.070 19.180 ;
        RECT 246.430 17.370 246.820 17.530 ;
        RECT 246.420 17.240 246.820 17.370 ;
        RECT 249.520 17.240 249.780 18.850 ;
        RECT 252.070 17.780 252.370 18.830 ;
        RECT 252.820 18.230 253.120 19.180 ;
        RECT 253.670 19.170 253.870 19.180 ;
        RECT 264.240 19.110 269.630 19.410 ;
        RECT 253.320 18.280 253.620 18.330 ;
        RECT 253.320 17.930 254.220 18.280 ;
        RECT 269.430 17.870 269.630 19.110 ;
        RECT 340.700 18.830 340.980 19.880 ;
        RECT 342.690 19.080 342.910 19.890 ;
        RECT 343.300 19.860 343.570 19.890 ;
        RECT 344.430 20.150 344.720 20.200 ;
        RECT 344.430 19.970 355.180 20.150 ;
        RECT 344.430 19.870 344.720 19.970 ;
        RECT 349.270 19.960 352.900 19.970 ;
        RECT 354.980 19.290 355.180 19.970 ;
        RECT 361.370 19.830 361.660 20.430 ;
        RECT 363.260 19.830 363.550 20.430 ;
        RECT 339.980 18.380 340.980 18.830 ;
        RECT 261.870 17.850 263.060 17.860 ;
        RECT 264.050 17.850 265.240 17.860 ;
        RECT 266.270 17.850 267.460 17.860 ;
        RECT 268.450 17.850 269.640 17.870 ;
        RECT 259.660 17.840 269.640 17.850 ;
        RECT 256.270 17.820 257.460 17.830 ;
        RECT 258.550 17.820 269.640 17.840 ;
        RECT 245.040 17.030 245.330 17.190 ;
        RECT 246.420 17.180 246.680 17.240 ;
        RECT 244.540 16.840 245.330 17.030 ;
        RECT 244.540 16.640 244.790 16.840 ;
        RECT 245.040 16.730 245.330 16.840 ;
        RECT 246.430 16.640 246.680 17.180 ;
        RECT 249.510 17.180 249.780 17.240 ;
        RECT 251.060 17.520 252.370 17.780 ;
        RECT 254.430 17.590 269.640 17.820 ;
        RECT 254.430 17.580 268.590 17.590 ;
        RECT 254.430 17.570 261.960 17.580 ;
        RECT 262.970 17.570 264.160 17.580 ;
        RECT 265.120 17.570 266.310 17.580 ;
        RECT 267.400 17.570 268.590 17.580 ;
        RECT 254.430 17.560 259.740 17.570 ;
        RECT 254.430 17.550 258.600 17.560 ;
        RECT 254.430 17.540 256.320 17.550 ;
        RECT 257.410 17.540 258.600 17.550 ;
        RECT 254.430 17.530 255.150 17.540 ;
        RECT 251.060 17.180 251.370 17.520 ;
        RECT 247.070 16.650 248.710 17.040 ;
        RECT 249.510 16.890 251.370 17.180 ;
        RECT 249.510 16.880 249.820 16.890 ;
        RECT 251.060 16.880 251.370 16.890 ;
        RECT 239.650 16.530 240.300 16.540 ;
        RECT 239.650 16.200 239.950 16.530 ;
        RECT 238.930 15.750 239.950 16.200 ;
        RECT 244.540 16.040 244.830 16.640 ;
        RECT 246.430 16.040 246.720 16.640 ;
        RECT 239.650 15.740 239.950 15.750 ;
        RECT 248.770 15.430 249.070 16.430 ;
        RECT 249.520 15.830 249.820 16.880 ;
        RECT 252.120 15.780 252.370 17.520 ;
        RECT 252.820 15.430 253.080 16.980 ;
        RECT 339.960 16.930 341.260 17.380 ;
        RECT 340.960 16.530 341.260 16.930 ;
        RECT 342.680 16.550 342.910 19.080 ;
        RECT 349.930 18.990 355.180 19.290 ;
        RECT 365.600 19.220 365.900 20.220 ;
        RECT 366.350 19.620 366.650 20.670 ;
        RECT 368.950 19.570 369.200 21.310 ;
        RECT 371.320 21.310 388.670 21.620 ;
        RECT 371.320 21.300 384.330 21.310 ;
        RECT 376.180 21.290 384.330 21.300 ;
        RECT 387.710 21.270 388.670 21.310 ;
        RECT 388.280 21.260 388.620 21.270 ;
        RECT 369.650 19.220 369.910 20.770 ;
        RECT 370.740 19.220 370.940 19.230 ;
        RECT 341.750 16.530 342.910 16.550 ;
        RECT 340.960 16.350 342.910 16.530 ;
        RECT 345.850 17.350 346.110 18.550 ;
        RECT 345.850 16.840 346.100 17.350 ;
        RECT 347.740 17.340 348.000 18.550 ;
        RECT 350.130 17.440 350.380 18.990 ;
        RECT 347.740 17.180 348.130 17.340 ;
        RECT 347.730 17.050 348.130 17.180 ;
        RECT 350.830 17.050 351.090 18.660 ;
        RECT 353.380 17.590 353.680 18.640 ;
        RECT 354.130 18.040 354.430 18.990 ;
        RECT 354.980 18.980 355.180 18.990 ;
        RECT 365.550 18.920 370.940 19.220 ;
        RECT 354.630 18.090 354.930 18.140 ;
        RECT 354.630 17.740 355.530 18.090 ;
        RECT 370.740 17.680 370.940 18.920 ;
        RECT 363.180 17.660 364.370 17.670 ;
        RECT 365.360 17.660 366.550 17.670 ;
        RECT 367.580 17.660 368.770 17.670 ;
        RECT 369.760 17.660 370.950 17.680 ;
        RECT 360.970 17.650 370.950 17.660 ;
        RECT 357.580 17.630 358.770 17.640 ;
        RECT 359.860 17.630 370.950 17.650 ;
        RECT 346.350 16.840 346.640 17.000 ;
        RECT 347.730 16.990 347.990 17.050 ;
        RECT 345.850 16.650 346.640 16.840 ;
        RECT 345.850 16.450 346.100 16.650 ;
        RECT 346.350 16.540 346.640 16.650 ;
        RECT 347.740 16.450 347.990 16.990 ;
        RECT 350.820 16.990 351.090 17.050 ;
        RECT 352.370 17.330 353.680 17.590 ;
        RECT 355.740 17.400 370.950 17.630 ;
        RECT 355.740 17.390 369.900 17.400 ;
        RECT 355.740 17.380 363.270 17.390 ;
        RECT 364.280 17.380 365.470 17.390 ;
        RECT 366.430 17.380 367.620 17.390 ;
        RECT 368.710 17.380 369.900 17.390 ;
        RECT 355.740 17.370 361.050 17.380 ;
        RECT 355.740 17.360 359.910 17.370 ;
        RECT 355.740 17.350 357.630 17.360 ;
        RECT 358.720 17.350 359.910 17.360 ;
        RECT 355.740 17.340 356.460 17.350 ;
        RECT 352.370 16.990 352.680 17.330 ;
        RECT 348.380 16.460 350.020 16.850 ;
        RECT 350.820 16.700 352.680 16.990 ;
        RECT 350.820 16.690 351.130 16.700 ;
        RECT 352.370 16.690 352.680 16.700 ;
        RECT 340.960 16.340 341.610 16.350 ;
        RECT 340.960 16.010 341.260 16.340 ;
        RECT 340.240 15.560 341.260 16.010 ;
        RECT 345.850 15.850 346.140 16.450 ;
        RECT 347.740 15.850 348.030 16.450 ;
        RECT 350.830 15.640 351.130 16.690 ;
        RECT 353.430 15.590 353.680 17.330 ;
        RECT 340.960 15.550 341.260 15.560 ;
        RECT 248.720 15.420 253.970 15.430 ;
        RECT 238.600 15.340 238.850 15.350 ;
        RECT 238.600 14.880 239.580 15.340 ;
        RECT 248.720 15.130 253.990 15.420 ;
        RECT 238.600 14.580 238.850 14.880 ;
        RECT 246.570 14.790 248.410 14.800 ;
        RECT 253.820 14.790 253.990 15.130 ;
        RECT 240.310 14.780 240.550 14.790 ;
        RECT 241.390 14.780 253.990 14.790 ;
        RECT 240.310 14.620 253.990 14.780 ;
        RECT 240.310 14.610 251.820 14.620 ;
        RECT 240.300 14.600 246.620 14.610 ;
        RECT 248.170 14.600 251.820 14.610 ;
        RECT 240.300 14.590 242.170 14.600 ;
        RECT 240.300 14.580 240.550 14.590 ;
        RECT 238.600 14.410 240.550 14.580 ;
        RECT 238.600 14.110 238.870 14.410 ;
        RECT 238.610 13.850 238.870 14.110 ;
        RECT 238.590 13.460 238.890 13.850 ;
        RECT 238.580 13.060 238.890 13.460 ;
        RECT 238.580 12.800 238.870 13.060 ;
        RECT 238.560 12.630 238.870 12.800 ;
        RECT 238.560 12.390 238.850 12.630 ;
        RECT 238.000 12.210 238.860 12.390 ;
        RECT 238.000 11.670 238.310 12.210 ;
        RECT 238.000 11.650 238.360 11.670 ;
        RECT 0.030 10.470 2.120 10.480 ;
        RECT 2.330 10.470 2.800 10.530 ;
        RECT 0.030 10.200 2.800 10.470 ;
        RECT 0.670 10.190 2.800 10.200 ;
        RECT 2.330 10.180 2.800 10.190 ;
        RECT 236.560 10.420 236.830 11.400 ;
        RECT 238.000 10.700 238.450 11.650 ;
        RECT 238.860 10.470 239.320 11.350 ;
        RECT 236.560 10.410 238.650 10.420 ;
        RECT 238.860 10.410 239.330 10.470 ;
        RECT 236.560 10.140 239.330 10.410 ;
        RECT 237.200 10.130 239.330 10.140 ;
        RECT 238.860 10.120 239.330 10.130 ;
      LAYER mcon ;
        RECT 100.880 255.470 101.050 255.640 ;
        RECT 337.410 255.410 337.580 255.580 ;
        RECT 100.910 252.020 101.080 252.190 ;
        RECT 10.895 248.405 11.065 248.575 ;
        RECT 18.350 249.135 18.520 249.305 ;
        RECT 16.490 248.700 16.660 248.870 ;
        RECT 18.895 248.710 19.065 248.880 ;
        RECT 6.580 245.665 6.750 245.835 ;
        RECT 7.760 245.645 7.930 245.815 ;
        RECT 26.575 245.985 26.745 246.155 ;
        RECT 34.030 246.715 34.200 246.885 ;
        RECT 32.170 246.280 32.340 246.450 ;
        RECT 6.560 244.850 6.730 245.020 ;
        RECT 7.690 244.860 7.860 245.030 ;
        RECT 34.575 246.290 34.745 246.460 ;
        RECT 11.055 242.005 11.225 242.175 ;
        RECT 18.510 242.735 18.680 242.905 ;
        RECT 16.650 242.300 16.820 242.470 ;
        RECT 19.020 242.275 19.190 242.445 ;
        RECT 44.155 240.435 44.325 240.605 ;
        RECT 51.610 241.165 51.780 241.335 ;
        RECT 49.750 240.730 49.920 240.900 ;
        RECT 52.145 240.735 52.315 240.905 ;
        RECT 10.725 233.985 10.895 234.155 ;
        RECT 18.180 234.715 18.350 234.885 ;
        RECT 16.320 234.280 16.490 234.450 ;
        RECT 18.725 234.290 18.895 234.460 ;
        RECT 6.410 231.245 6.580 231.415 ;
        RECT 7.590 231.225 7.760 231.395 ;
        RECT 26.405 231.565 26.575 231.735 ;
        RECT 33.860 232.295 34.030 232.465 ;
        RECT 32.000 231.860 32.170 232.030 ;
        RECT 6.390 230.430 6.560 230.600 ;
        RECT 7.520 230.440 7.690 230.610 ;
        RECT 34.405 231.870 34.575 232.040 ;
        RECT 10.885 227.585 11.055 227.755 ;
        RECT 18.340 228.315 18.510 228.485 ;
        RECT 16.480 227.880 16.650 228.050 ;
        RECT 18.850 227.855 19.020 228.025 ;
        RECT 61.685 224.415 61.855 224.585 ;
        RECT 69.140 225.145 69.310 225.315 ;
        RECT 67.280 224.710 67.450 224.880 ;
        RECT 69.700 224.710 69.870 224.880 ;
        RECT 10.865 218.335 11.035 218.505 ;
        RECT 18.320 219.065 18.490 219.235 ;
        RECT 16.460 218.630 16.630 218.800 ;
        RECT 18.865 218.640 19.035 218.810 ;
        RECT 6.550 215.595 6.720 215.765 ;
        RECT 7.730 215.575 7.900 215.745 ;
        RECT 26.545 215.915 26.715 216.085 ;
        RECT 34.000 216.645 34.170 216.815 ;
        RECT 32.140 216.210 32.310 216.380 ;
        RECT 6.530 214.780 6.700 214.950 ;
        RECT 7.660 214.790 7.830 214.960 ;
        RECT 34.545 216.220 34.715 216.390 ;
        RECT 11.025 211.935 11.195 212.105 ;
        RECT 18.480 212.665 18.650 212.835 ;
        RECT 16.620 212.230 16.790 212.400 ;
        RECT 18.990 212.205 19.160 212.375 ;
        RECT 44.125 210.365 44.295 210.535 ;
        RECT 51.580 211.095 51.750 211.265 ;
        RECT 49.720 210.660 49.890 210.830 ;
        RECT 52.115 210.665 52.285 210.835 ;
        RECT 10.695 203.915 10.865 204.085 ;
        RECT 18.150 204.645 18.320 204.815 ;
        RECT 16.290 204.210 16.460 204.380 ;
        RECT 18.695 204.220 18.865 204.390 ;
        RECT 6.380 201.175 6.550 201.345 ;
        RECT 7.560 201.155 7.730 201.325 ;
        RECT 26.375 201.495 26.545 201.665 ;
        RECT 33.830 202.225 34.000 202.395 ;
        RECT 31.970 201.790 32.140 201.960 ;
        RECT 6.360 200.360 6.530 200.530 ;
        RECT 7.490 200.370 7.660 200.540 ;
        RECT 34.375 201.800 34.545 201.970 ;
        RECT 10.855 197.515 11.025 197.685 ;
        RECT 18.310 198.245 18.480 198.415 ;
        RECT 16.450 197.810 16.620 197.980 ;
        RECT 18.820 197.785 18.990 197.955 ;
        RECT 75.885 198.125 76.055 198.295 ;
        RECT 83.340 198.855 83.510 199.025 ;
        RECT 81.480 198.420 81.650 198.590 ;
        RECT 83.900 198.415 84.070 198.585 ;
        RECT 10.545 188.485 10.715 188.655 ;
        RECT 18.000 189.215 18.170 189.385 ;
        RECT 16.140 188.780 16.310 188.950 ;
        RECT 18.545 188.790 18.715 188.960 ;
        RECT 6.230 185.745 6.400 185.915 ;
        RECT 7.410 185.725 7.580 185.895 ;
        RECT 26.225 186.065 26.395 186.235 ;
        RECT 33.680 186.795 33.850 186.965 ;
        RECT 31.820 186.360 31.990 186.530 ;
        RECT 6.210 184.930 6.380 185.100 ;
        RECT 7.340 184.940 7.510 185.110 ;
        RECT 34.225 186.370 34.395 186.540 ;
        RECT 10.705 182.085 10.875 182.255 ;
        RECT 18.160 182.815 18.330 182.985 ;
        RECT 16.300 182.380 16.470 182.550 ;
        RECT 18.670 182.355 18.840 182.525 ;
        RECT 43.805 180.515 43.975 180.685 ;
        RECT 51.260 181.245 51.430 181.415 ;
        RECT 49.400 180.810 49.570 180.980 ;
        RECT 51.795 180.815 51.965 180.985 ;
        RECT 10.375 174.065 10.545 174.235 ;
        RECT 17.830 174.795 18.000 174.965 ;
        RECT 15.970 174.360 16.140 174.530 ;
        RECT 18.375 174.370 18.545 174.540 ;
        RECT 6.060 171.325 6.230 171.495 ;
        RECT 7.240 171.305 7.410 171.475 ;
        RECT 26.055 171.645 26.225 171.815 ;
        RECT 33.510 172.375 33.680 172.545 ;
        RECT 31.650 171.940 31.820 172.110 ;
        RECT 6.040 170.510 6.210 170.680 ;
        RECT 7.170 170.520 7.340 170.690 ;
        RECT 34.055 171.950 34.225 172.120 ;
        RECT 10.535 167.665 10.705 167.835 ;
        RECT 17.990 168.395 18.160 168.565 ;
        RECT 16.130 167.960 16.300 168.130 ;
        RECT 18.500 167.935 18.670 168.105 ;
        RECT 61.335 164.495 61.505 164.665 ;
        RECT 68.790 165.225 68.960 165.395 ;
        RECT 66.930 164.790 67.100 164.960 ;
        RECT 69.350 164.790 69.520 164.960 ;
        RECT 10.515 158.415 10.685 158.585 ;
        RECT 17.970 159.145 18.140 159.315 ;
        RECT 16.110 158.710 16.280 158.880 ;
        RECT 18.515 158.720 18.685 158.890 ;
        RECT 6.200 155.675 6.370 155.845 ;
        RECT 7.380 155.655 7.550 155.825 ;
        RECT 26.195 155.995 26.365 156.165 ;
        RECT 33.650 156.725 33.820 156.895 ;
        RECT 31.790 156.290 31.960 156.460 ;
        RECT 6.180 154.860 6.350 155.030 ;
        RECT 7.310 154.870 7.480 155.040 ;
        RECT 34.195 156.300 34.365 156.470 ;
        RECT 10.675 152.015 10.845 152.185 ;
        RECT 18.130 152.745 18.300 152.915 ;
        RECT 16.270 152.310 16.440 152.480 ;
        RECT 18.640 152.285 18.810 152.455 ;
        RECT 43.775 150.445 43.945 150.615 ;
        RECT 51.230 151.175 51.400 151.345 ;
        RECT 49.370 150.740 49.540 150.910 ;
        RECT 112.205 248.215 112.375 248.385 ;
        RECT 119.660 248.945 119.830 249.115 ;
        RECT 117.800 248.510 117.970 248.680 ;
        RECT 120.205 248.520 120.375 248.690 ;
        RECT 107.890 245.475 108.060 245.645 ;
        RECT 109.070 245.455 109.240 245.625 ;
        RECT 127.885 245.795 128.055 245.965 ;
        RECT 135.340 246.525 135.510 246.695 ;
        RECT 133.480 246.090 133.650 246.260 ;
        RECT 107.870 244.660 108.040 244.830 ;
        RECT 109.000 244.670 109.170 244.840 ;
        RECT 135.885 246.100 136.055 246.270 ;
        RECT 112.365 241.815 112.535 241.985 ;
        RECT 119.820 242.545 119.990 242.715 ;
        RECT 117.960 242.110 118.130 242.280 ;
        RECT 120.330 242.085 120.500 242.255 ;
        RECT 145.465 240.245 145.635 240.415 ;
        RECT 152.920 240.975 153.090 241.145 ;
        RECT 151.060 240.540 151.230 240.710 ;
        RECT 153.455 240.545 153.625 240.715 ;
        RECT 112.035 233.795 112.205 233.965 ;
        RECT 119.490 234.525 119.660 234.695 ;
        RECT 117.630 234.090 117.800 234.260 ;
        RECT 120.035 234.100 120.205 234.270 ;
        RECT 107.720 231.055 107.890 231.225 ;
        RECT 108.900 231.035 109.070 231.205 ;
        RECT 127.715 231.375 127.885 231.545 ;
        RECT 135.170 232.105 135.340 232.275 ;
        RECT 133.310 231.670 133.480 231.840 ;
        RECT 107.700 230.240 107.870 230.410 ;
        RECT 108.830 230.250 109.000 230.420 ;
        RECT 135.715 231.680 135.885 231.850 ;
        RECT 112.195 227.395 112.365 227.565 ;
        RECT 119.650 228.125 119.820 228.295 ;
        RECT 117.790 227.690 117.960 227.860 ;
        RECT 120.160 227.665 120.330 227.835 ;
        RECT 162.995 224.225 163.165 224.395 ;
        RECT 170.450 224.955 170.620 225.125 ;
        RECT 168.590 224.520 168.760 224.690 ;
        RECT 171.010 224.520 171.180 224.690 ;
        RECT 112.175 218.145 112.345 218.315 ;
        RECT 119.630 218.875 119.800 219.045 ;
        RECT 117.770 218.440 117.940 218.610 ;
        RECT 120.175 218.450 120.345 218.620 ;
        RECT 107.860 215.405 108.030 215.575 ;
        RECT 109.040 215.385 109.210 215.555 ;
        RECT 127.855 215.725 128.025 215.895 ;
        RECT 135.310 216.455 135.480 216.625 ;
        RECT 133.450 216.020 133.620 216.190 ;
        RECT 107.840 214.590 108.010 214.760 ;
        RECT 108.970 214.600 109.140 214.770 ;
        RECT 135.855 216.030 136.025 216.200 ;
        RECT 112.335 211.745 112.505 211.915 ;
        RECT 119.790 212.475 119.960 212.645 ;
        RECT 117.930 212.040 118.100 212.210 ;
        RECT 120.300 212.015 120.470 212.185 ;
        RECT 145.435 210.175 145.605 210.345 ;
        RECT 152.890 210.905 153.060 211.075 ;
        RECT 151.030 210.470 151.200 210.640 ;
        RECT 153.425 210.475 153.595 210.645 ;
        RECT 112.005 203.725 112.175 203.895 ;
        RECT 119.460 204.455 119.630 204.625 ;
        RECT 117.600 204.020 117.770 204.190 ;
        RECT 120.005 204.030 120.175 204.200 ;
        RECT 107.690 200.985 107.860 201.155 ;
        RECT 108.870 200.965 109.040 201.135 ;
        RECT 127.685 201.305 127.855 201.475 ;
        RECT 135.140 202.035 135.310 202.205 ;
        RECT 133.280 201.600 133.450 201.770 ;
        RECT 107.670 200.170 107.840 200.340 ;
        RECT 108.800 200.180 108.970 200.350 ;
        RECT 135.685 201.610 135.855 201.780 ;
        RECT 112.165 197.325 112.335 197.495 ;
        RECT 119.620 198.055 119.790 198.225 ;
        RECT 117.760 197.620 117.930 197.790 ;
        RECT 120.130 197.595 120.300 197.765 ;
        RECT 177.195 197.935 177.365 198.105 ;
        RECT 184.650 198.665 184.820 198.835 ;
        RECT 182.790 198.230 182.960 198.400 ;
        RECT 185.210 198.225 185.380 198.395 ;
        RECT 111.855 188.295 112.025 188.465 ;
        RECT 119.310 189.025 119.480 189.195 ;
        RECT 117.450 188.590 117.620 188.760 ;
        RECT 119.855 188.600 120.025 188.770 ;
        RECT 107.540 185.555 107.710 185.725 ;
        RECT 108.720 185.535 108.890 185.705 ;
        RECT 127.535 185.875 127.705 186.045 ;
        RECT 134.990 186.605 135.160 186.775 ;
        RECT 133.130 186.170 133.300 186.340 ;
        RECT 107.520 184.740 107.690 184.910 ;
        RECT 108.650 184.750 108.820 184.920 ;
        RECT 135.535 186.180 135.705 186.350 ;
        RECT 112.015 181.895 112.185 182.065 ;
        RECT 119.470 182.625 119.640 182.795 ;
        RECT 117.610 182.190 117.780 182.360 ;
        RECT 119.980 182.165 120.150 182.335 ;
        RECT 145.115 180.325 145.285 180.495 ;
        RECT 152.570 181.055 152.740 181.225 ;
        RECT 150.710 180.620 150.880 180.790 ;
        RECT 153.105 180.625 153.275 180.795 ;
        RECT 111.685 173.875 111.855 174.045 ;
        RECT 119.140 174.605 119.310 174.775 ;
        RECT 117.280 174.170 117.450 174.340 ;
        RECT 119.685 174.180 119.855 174.350 ;
        RECT 107.370 171.135 107.540 171.305 ;
        RECT 108.550 171.115 108.720 171.285 ;
        RECT 127.365 171.455 127.535 171.625 ;
        RECT 134.820 172.185 134.990 172.355 ;
        RECT 132.960 171.750 133.130 171.920 ;
        RECT 107.350 170.320 107.520 170.490 ;
        RECT 108.480 170.330 108.650 170.500 ;
        RECT 135.365 171.760 135.535 171.930 ;
        RECT 111.845 167.475 112.015 167.645 ;
        RECT 119.300 168.205 119.470 168.375 ;
        RECT 117.440 167.770 117.610 167.940 ;
        RECT 119.810 167.745 119.980 167.915 ;
        RECT 51.765 150.745 51.935 150.915 ;
        RECT 10.345 143.995 10.515 144.165 ;
        RECT 17.800 144.725 17.970 144.895 ;
        RECT 15.940 144.290 16.110 144.460 ;
        RECT 18.345 144.300 18.515 144.470 ;
        RECT 6.030 141.255 6.200 141.425 ;
        RECT 7.210 141.235 7.380 141.405 ;
        RECT 26.025 141.575 26.195 141.745 ;
        RECT 33.480 142.305 33.650 142.475 ;
        RECT 162.645 164.305 162.815 164.475 ;
        RECT 170.100 165.035 170.270 165.205 ;
        RECT 168.240 164.600 168.410 164.770 ;
        RECT 170.660 164.600 170.830 164.770 ;
        RECT 111.825 158.225 111.995 158.395 ;
        RECT 119.280 158.955 119.450 159.125 ;
        RECT 117.420 158.520 117.590 158.690 ;
        RECT 119.825 158.530 119.995 158.700 ;
        RECT 107.510 155.485 107.680 155.655 ;
        RECT 108.690 155.465 108.860 155.635 ;
        RECT 127.505 155.805 127.675 155.975 ;
        RECT 134.960 156.535 135.130 156.705 ;
        RECT 133.100 156.100 133.270 156.270 ;
        RECT 107.490 154.670 107.660 154.840 ;
        RECT 108.620 154.680 108.790 154.850 ;
        RECT 135.505 156.110 135.675 156.280 ;
        RECT 111.985 151.825 112.155 151.995 ;
        RECT 119.440 152.555 119.610 152.725 ;
        RECT 117.580 152.120 117.750 152.290 ;
        RECT 119.950 152.095 120.120 152.265 ;
        RECT 145.085 150.255 145.255 150.425 ;
        RECT 152.540 150.985 152.710 151.155 ;
        RECT 150.680 150.550 150.850 150.720 ;
        RECT 153.075 150.555 153.245 150.725 ;
        RECT 31.620 141.870 31.790 142.040 ;
        RECT 6.010 140.440 6.180 140.610 ;
        RECT 7.140 140.450 7.310 140.620 ;
        RECT 34.025 141.880 34.195 142.050 ;
        RECT 10.505 137.595 10.675 137.765 ;
        RECT 17.960 138.325 18.130 138.495 ;
        RECT 111.655 143.805 111.825 143.975 ;
        RECT 119.110 144.535 119.280 144.705 ;
        RECT 117.250 144.100 117.420 144.270 ;
        RECT 119.655 144.110 119.825 144.280 ;
        RECT 16.100 137.890 16.270 138.060 ;
        RECT 18.470 137.865 18.640 138.035 ;
        RECT 92.215 134.985 92.385 135.155 ;
        RECT 99.670 135.715 99.840 135.885 ;
        RECT 107.340 141.065 107.510 141.235 ;
        RECT 108.520 141.045 108.690 141.215 ;
        RECT 127.335 141.385 127.505 141.555 ;
        RECT 134.790 142.115 134.960 142.285 ;
        RECT 132.930 141.680 133.100 141.850 ;
        RECT 107.320 140.250 107.490 140.420 ;
        RECT 108.450 140.260 108.620 140.430 ;
        RECT 135.335 141.690 135.505 141.860 ;
        RECT 111.815 137.405 111.985 137.575 ;
        RECT 119.270 138.135 119.440 138.305 ;
        RECT 117.410 137.700 117.580 137.870 ;
        RECT 119.780 137.675 119.950 137.845 ;
        RECT 227.260 137.855 227.430 138.025 ;
        RECT 219.805 137.125 219.975 137.295 ;
        RECT 97.810 135.280 97.980 135.450 ;
        RECT 100.275 135.290 100.445 135.460 ;
        RECT 193.525 134.795 193.695 134.965 ;
        RECT 200.980 135.525 201.150 135.695 ;
        RECT 199.120 135.090 199.290 135.260 ;
        RECT 201.585 135.100 201.755 135.270 ;
        RECT 10.395 128.165 10.565 128.335 ;
        RECT 17.850 128.895 18.020 129.065 ;
        RECT 15.990 128.460 16.160 128.630 ;
        RECT 18.395 128.470 18.565 128.640 ;
        RECT 6.080 125.425 6.250 125.595 ;
        RECT 7.260 125.405 7.430 125.575 ;
        RECT 26.075 125.745 26.245 125.915 ;
        RECT 33.530 126.475 33.700 126.645 ;
        RECT 31.670 126.040 31.840 126.210 ;
        RECT 6.060 124.610 6.230 124.780 ;
        RECT 7.190 124.620 7.360 124.790 ;
        RECT 34.075 126.050 34.245 126.220 ;
        RECT 10.555 121.765 10.725 121.935 ;
        RECT 18.010 122.495 18.180 122.665 ;
        RECT 16.150 122.060 16.320 122.230 ;
        RECT 18.520 122.035 18.690 122.205 ;
        RECT 43.655 120.195 43.825 120.365 ;
        RECT 51.110 120.925 51.280 121.095 ;
        RECT 49.250 120.490 49.420 120.660 ;
        RECT 51.645 120.495 51.815 120.665 ;
        RECT 10.225 113.745 10.395 113.915 ;
        RECT 17.680 114.475 17.850 114.645 ;
        RECT 15.820 114.040 15.990 114.210 ;
        RECT 18.225 114.050 18.395 114.220 ;
        RECT 5.910 111.005 6.080 111.175 ;
        RECT 7.090 110.985 7.260 111.155 ;
        RECT 25.905 111.325 26.075 111.495 ;
        RECT 33.360 112.055 33.530 112.225 ;
        RECT 31.500 111.620 31.670 111.790 ;
        RECT 5.890 110.190 6.060 110.360 ;
        RECT 7.020 110.200 7.190 110.370 ;
        RECT 33.905 111.630 34.075 111.800 ;
        RECT 10.385 107.345 10.555 107.515 ;
        RECT 17.840 108.075 18.010 108.245 ;
        RECT 15.980 107.640 16.150 107.810 ;
        RECT 18.350 107.615 18.520 107.785 ;
        RECT 61.185 104.175 61.355 104.345 ;
        RECT 68.640 104.905 68.810 105.075 ;
        RECT 66.780 104.470 66.950 104.640 ;
        RECT 69.200 104.470 69.370 104.640 ;
        RECT 10.365 98.095 10.535 98.265 ;
        RECT 17.820 98.825 17.990 98.995 ;
        RECT 15.960 98.390 16.130 98.560 ;
        RECT 18.365 98.400 18.535 98.570 ;
        RECT 6.050 95.355 6.220 95.525 ;
        RECT 7.230 95.335 7.400 95.505 ;
        RECT 26.045 95.675 26.215 95.845 ;
        RECT 33.500 96.405 33.670 96.575 ;
        RECT 31.640 95.970 31.810 96.140 ;
        RECT 6.030 94.540 6.200 94.710 ;
        RECT 7.160 94.550 7.330 94.720 ;
        RECT 34.045 95.980 34.215 96.150 ;
        RECT 10.525 91.695 10.695 91.865 ;
        RECT 17.980 92.425 18.150 92.595 ;
        RECT 16.120 91.990 16.290 92.160 ;
        RECT 18.490 91.965 18.660 92.135 ;
        RECT 43.625 90.125 43.795 90.295 ;
        RECT 51.080 90.855 51.250 91.025 ;
        RECT 49.220 90.420 49.390 90.590 ;
        RECT 51.615 90.425 51.785 90.595 ;
        RECT 10.195 83.675 10.365 83.845 ;
        RECT 17.650 84.405 17.820 84.575 ;
        RECT 15.790 83.970 15.960 84.140 ;
        RECT 18.195 83.980 18.365 84.150 ;
        RECT 5.880 80.935 6.050 81.105 ;
        RECT 7.060 80.915 7.230 81.085 ;
        RECT 25.875 81.255 26.045 81.425 ;
        RECT 33.330 81.985 33.500 82.155 ;
        RECT 31.470 81.550 31.640 81.720 ;
        RECT 5.860 80.120 6.030 80.290 ;
        RECT 6.990 80.130 7.160 80.300 ;
        RECT 33.875 81.560 34.045 81.730 ;
        RECT 10.355 77.275 10.525 77.445 ;
        RECT 17.810 78.005 17.980 78.175 ;
        RECT 15.950 77.570 16.120 77.740 ;
        RECT 18.320 77.545 18.490 77.715 ;
        RECT 75.385 77.885 75.555 78.055 ;
        RECT 82.840 78.615 83.010 78.785 ;
        RECT 111.705 127.975 111.875 128.145 ;
        RECT 119.160 128.705 119.330 128.875 ;
        RECT 117.300 128.270 117.470 128.440 ;
        RECT 119.705 128.280 119.875 128.450 ;
        RECT 107.390 125.235 107.560 125.405 ;
        RECT 108.570 125.215 108.740 125.385 ;
        RECT 127.385 125.555 127.555 125.725 ;
        RECT 134.840 126.285 135.010 126.455 ;
        RECT 132.980 125.850 133.150 126.020 ;
        RECT 107.370 124.420 107.540 124.590 ;
        RECT 108.500 124.430 108.670 124.600 ;
        RECT 135.385 125.860 135.555 126.030 ;
        RECT 111.865 121.575 112.035 121.745 ;
        RECT 119.320 122.305 119.490 122.475 ;
        RECT 117.460 121.870 117.630 122.040 ;
        RECT 119.830 121.845 120.000 122.015 ;
        RECT 144.965 120.005 145.135 120.175 ;
        RECT 152.420 120.735 152.590 120.905 ;
        RECT 150.560 120.300 150.730 120.470 ;
        RECT 152.955 120.305 153.125 120.475 ;
        RECT 111.535 113.555 111.705 113.725 ;
        RECT 118.990 114.285 119.160 114.455 ;
        RECT 117.130 113.850 117.300 114.020 ;
        RECT 119.535 113.860 119.705 114.030 ;
        RECT 107.220 110.815 107.390 110.985 ;
        RECT 108.400 110.795 108.570 110.965 ;
        RECT 127.215 111.135 127.385 111.305 ;
        RECT 134.670 111.865 134.840 112.035 ;
        RECT 132.810 111.430 132.980 111.600 ;
        RECT 107.200 110.000 107.370 110.170 ;
        RECT 108.330 110.010 108.500 110.180 ;
        RECT 135.215 111.440 135.385 111.610 ;
        RECT 111.695 107.155 111.865 107.325 ;
        RECT 119.150 107.885 119.320 108.055 ;
        RECT 117.290 107.450 117.460 107.620 ;
        RECT 119.660 107.425 119.830 107.595 ;
        RECT 162.495 103.985 162.665 104.155 ;
        RECT 169.950 104.715 170.120 104.885 ;
        RECT 168.090 104.280 168.260 104.450 ;
        RECT 170.510 104.280 170.680 104.450 ;
        RECT 111.675 97.905 111.845 98.075 ;
        RECT 119.130 98.635 119.300 98.805 ;
        RECT 117.270 98.200 117.440 98.370 ;
        RECT 119.675 98.210 119.845 98.380 ;
        RECT 107.360 95.165 107.530 95.335 ;
        RECT 108.540 95.145 108.710 95.315 ;
        RECT 127.355 95.485 127.525 95.655 ;
        RECT 134.810 96.215 134.980 96.385 ;
        RECT 132.950 95.780 133.120 95.950 ;
        RECT 107.340 94.350 107.510 94.520 ;
        RECT 108.470 94.360 108.640 94.530 ;
        RECT 135.355 95.790 135.525 95.960 ;
        RECT 111.835 91.505 112.005 91.675 ;
        RECT 119.290 92.235 119.460 92.405 ;
        RECT 117.430 91.800 117.600 91.970 ;
        RECT 119.800 91.775 119.970 91.945 ;
        RECT 144.935 89.935 145.105 90.105 ;
        RECT 152.390 90.665 152.560 90.835 ;
        RECT 150.530 90.230 150.700 90.400 ;
        RECT 152.925 90.235 153.095 90.405 ;
        RECT 111.505 83.485 111.675 83.655 ;
        RECT 118.960 84.215 119.130 84.385 ;
        RECT 117.100 83.780 117.270 83.950 ;
        RECT 119.505 83.790 119.675 83.960 ;
        RECT 107.190 80.745 107.360 80.915 ;
        RECT 108.370 80.725 108.540 80.895 ;
        RECT 127.185 81.065 127.355 81.235 ;
        RECT 134.640 81.795 134.810 81.965 ;
        RECT 132.780 81.360 132.950 81.530 ;
        RECT 107.170 79.930 107.340 80.100 ;
        RECT 108.300 79.940 108.470 80.110 ;
        RECT 80.980 78.180 81.150 78.350 ;
        RECT 83.400 78.175 83.570 78.345 ;
        RECT 135.185 81.370 135.355 81.540 ;
        RECT 111.665 77.085 111.835 77.255 ;
        RECT 119.120 77.815 119.290 77.985 ;
        RECT 117.260 77.380 117.430 77.550 ;
        RECT 119.630 77.355 119.800 77.525 ;
        RECT 176.695 77.695 176.865 77.865 ;
        RECT 184.150 78.425 184.320 78.595 ;
        RECT 10.045 68.245 10.215 68.415 ;
        RECT 17.500 68.975 17.670 69.145 ;
        RECT 15.640 68.540 15.810 68.710 ;
        RECT 18.045 68.550 18.215 68.720 ;
        RECT 5.730 65.505 5.900 65.675 ;
        RECT 6.910 65.485 7.080 65.655 ;
        RECT 25.725 65.825 25.895 65.995 ;
        RECT 33.180 66.555 33.350 66.725 ;
        RECT 31.320 66.120 31.490 66.290 ;
        RECT 5.710 64.690 5.880 64.860 ;
        RECT 6.840 64.700 7.010 64.870 ;
        RECT 33.725 66.130 33.895 66.300 ;
        RECT 182.290 77.990 182.460 78.160 ;
        RECT 184.710 77.985 184.880 78.155 ;
        RECT 111.355 68.055 111.525 68.225 ;
        RECT 118.810 68.785 118.980 68.955 ;
        RECT 116.950 68.350 117.120 68.520 ;
        RECT 119.355 68.360 119.525 68.530 ;
        RECT 10.205 61.845 10.375 62.015 ;
        RECT 17.660 62.575 17.830 62.745 ;
        RECT 15.800 62.140 15.970 62.310 ;
        RECT 18.170 62.115 18.340 62.285 ;
        RECT 43.305 60.275 43.475 60.445 ;
        RECT 50.760 61.005 50.930 61.175 ;
        RECT 48.900 60.570 49.070 60.740 ;
        RECT 51.295 60.575 51.465 60.745 ;
        RECT 9.875 53.825 10.045 53.995 ;
        RECT 17.330 54.555 17.500 54.725 ;
        RECT 15.470 54.120 15.640 54.290 ;
        RECT 17.875 54.130 18.045 54.300 ;
        RECT 5.560 51.085 5.730 51.255 ;
        RECT 6.740 51.065 6.910 51.235 ;
        RECT 25.555 51.405 25.725 51.575 ;
        RECT 33.010 52.135 33.180 52.305 ;
        RECT 31.150 51.700 31.320 51.870 ;
        RECT 5.540 50.270 5.710 50.440 ;
        RECT 6.670 50.280 6.840 50.450 ;
        RECT 33.555 51.710 33.725 51.880 ;
        RECT 10.035 47.425 10.205 47.595 ;
        RECT 17.490 48.155 17.660 48.325 ;
        RECT 15.630 47.720 15.800 47.890 ;
        RECT 18.000 47.695 18.170 47.865 ;
        RECT 107.040 65.315 107.210 65.485 ;
        RECT 108.220 65.295 108.390 65.465 ;
        RECT 127.035 65.635 127.205 65.805 ;
        RECT 134.490 66.365 134.660 66.535 ;
        RECT 132.630 65.930 132.800 66.100 ;
        RECT 107.020 64.500 107.190 64.670 ;
        RECT 108.150 64.510 108.320 64.680 ;
        RECT 135.035 65.940 135.205 66.110 ;
        RECT 111.515 61.655 111.685 61.825 ;
        RECT 118.970 62.385 119.140 62.555 ;
        RECT 117.110 61.950 117.280 62.120 ;
        RECT 119.480 61.925 119.650 62.095 ;
        RECT 144.615 60.085 144.785 60.255 ;
        RECT 152.070 60.815 152.240 60.985 ;
        RECT 150.210 60.380 150.380 60.550 ;
        RECT 152.605 60.385 152.775 60.555 ;
        RECT 111.185 53.635 111.355 53.805 ;
        RECT 118.640 54.365 118.810 54.535 ;
        RECT 116.780 53.930 116.950 54.100 ;
        RECT 119.185 53.940 119.355 54.110 ;
        RECT 106.870 50.895 107.040 51.065 ;
        RECT 108.050 50.875 108.220 51.045 ;
        RECT 126.865 51.215 127.035 51.385 ;
        RECT 134.320 51.945 134.490 52.115 ;
        RECT 132.460 51.510 132.630 51.680 ;
        RECT 106.850 50.080 107.020 50.250 ;
        RECT 107.980 50.090 108.150 50.260 ;
        RECT 134.865 51.520 135.035 51.690 ;
        RECT 60.835 44.255 61.005 44.425 ;
        RECT 68.290 44.985 68.460 45.155 ;
        RECT 111.345 47.235 111.515 47.405 ;
        RECT 118.800 47.965 118.970 48.135 ;
        RECT 116.940 47.530 117.110 47.700 ;
        RECT 119.310 47.505 119.480 47.675 ;
        RECT 66.430 44.550 66.600 44.720 ;
        RECT 68.850 44.550 69.020 44.720 ;
        RECT 162.145 44.065 162.315 44.235 ;
        RECT 169.600 44.795 169.770 44.965 ;
        RECT 167.740 44.360 167.910 44.530 ;
        RECT 170.160 44.360 170.330 44.530 ;
        RECT 10.015 38.175 10.185 38.345 ;
        RECT 17.470 38.905 17.640 39.075 ;
        RECT 15.610 38.470 15.780 38.640 ;
        RECT 18.015 38.480 18.185 38.650 ;
        RECT 5.700 35.435 5.870 35.605 ;
        RECT 6.880 35.415 7.050 35.585 ;
        RECT 25.695 35.755 25.865 35.925 ;
        RECT 33.150 36.485 33.320 36.655 ;
        RECT 31.290 36.050 31.460 36.220 ;
        RECT 5.680 34.620 5.850 34.790 ;
        RECT 6.810 34.630 6.980 34.800 ;
        RECT 33.695 36.060 33.865 36.230 ;
        RECT 10.175 31.775 10.345 31.945 ;
        RECT 17.630 32.505 17.800 32.675 ;
        RECT 15.770 32.070 15.940 32.240 ;
        RECT 18.140 32.045 18.310 32.215 ;
        RECT 43.275 30.205 43.445 30.375 ;
        RECT 50.730 30.935 50.900 31.105 ;
        RECT 48.870 30.500 49.040 30.670 ;
        RECT 111.325 37.985 111.495 38.155 ;
        RECT 118.780 38.715 118.950 38.885 ;
        RECT 116.920 38.280 117.090 38.450 ;
        RECT 119.325 38.290 119.495 38.460 ;
        RECT 107.010 35.245 107.180 35.415 ;
        RECT 108.190 35.225 108.360 35.395 ;
        RECT 127.005 35.565 127.175 35.735 ;
        RECT 134.460 36.295 134.630 36.465 ;
        RECT 132.600 35.860 132.770 36.030 ;
        RECT 106.990 34.430 107.160 34.600 ;
        RECT 108.120 34.440 108.290 34.610 ;
        RECT 135.005 35.870 135.175 36.040 ;
        RECT 111.485 31.585 111.655 31.755 ;
        RECT 118.940 32.315 119.110 32.485 ;
        RECT 117.080 31.880 117.250 32.050 ;
        RECT 119.450 31.855 119.620 32.025 ;
        RECT 51.265 30.505 51.435 30.675 ;
        RECT 144.585 30.015 144.755 30.185 ;
        RECT 152.040 30.745 152.210 30.915 ;
        RECT 150.180 30.310 150.350 30.480 ;
        RECT 152.575 30.315 152.745 30.485 ;
        RECT 9.845 23.755 10.015 23.925 ;
        RECT 17.300 24.485 17.470 24.655 ;
        RECT 15.440 24.050 15.610 24.220 ;
        RECT 17.845 24.060 18.015 24.230 ;
        RECT 5.530 21.015 5.700 21.185 ;
        RECT 6.710 20.995 6.880 21.165 ;
        RECT 25.525 21.335 25.695 21.505 ;
        RECT 32.980 22.065 33.150 22.235 ;
        RECT 111.155 23.565 111.325 23.735 ;
        RECT 118.610 24.295 118.780 24.465 ;
        RECT 116.750 23.860 116.920 24.030 ;
        RECT 119.155 23.870 119.325 24.040 ;
        RECT 31.120 21.630 31.290 21.800 ;
        RECT 5.510 20.200 5.680 20.370 ;
        RECT 6.640 20.210 6.810 20.380 ;
        RECT 33.525 21.640 33.695 21.810 ;
        RECT 106.840 20.825 107.010 20.995 ;
        RECT 108.020 20.805 108.190 20.975 ;
        RECT 126.835 21.145 127.005 21.315 ;
        RECT 134.290 21.875 134.460 22.045 ;
        RECT 132.430 21.440 132.600 21.610 ;
        RECT 106.820 20.010 106.990 20.180 ;
        RECT 10.005 17.355 10.175 17.525 ;
        RECT 17.460 18.085 17.630 18.255 ;
        RECT 107.950 20.020 108.120 20.190 ;
        RECT 15.600 17.650 15.770 17.820 ;
        RECT 17.970 17.625 18.140 17.795 ;
        RECT 134.835 21.450 135.005 21.620 ;
        RECT 111.315 17.165 111.485 17.335 ;
        RECT 118.770 17.895 118.940 18.065 ;
        RECT 116.910 17.460 117.080 17.630 ;
        RECT 119.280 17.435 119.450 17.605 ;
        RECT 337.440 251.960 337.610 252.130 ;
        RECT 247.425 248.345 247.595 248.515 ;
        RECT 254.880 249.075 255.050 249.245 ;
        RECT 253.020 248.640 253.190 248.810 ;
        RECT 255.425 248.650 255.595 248.820 ;
        RECT 243.110 245.605 243.280 245.775 ;
        RECT 244.290 245.585 244.460 245.755 ;
        RECT 263.105 245.925 263.275 246.095 ;
        RECT 270.560 246.655 270.730 246.825 ;
        RECT 268.700 246.220 268.870 246.390 ;
        RECT 243.090 244.790 243.260 244.960 ;
        RECT 244.220 244.800 244.390 244.970 ;
        RECT 271.105 246.230 271.275 246.400 ;
        RECT 247.585 241.945 247.755 242.115 ;
        RECT 255.040 242.675 255.210 242.845 ;
        RECT 253.180 242.240 253.350 242.410 ;
        RECT 255.550 242.215 255.720 242.385 ;
        RECT 280.685 240.375 280.855 240.545 ;
        RECT 288.140 241.105 288.310 241.275 ;
        RECT 286.280 240.670 286.450 240.840 ;
        RECT 288.675 240.675 288.845 240.845 ;
        RECT 247.255 233.925 247.425 234.095 ;
        RECT 254.710 234.655 254.880 234.825 ;
        RECT 252.850 234.220 253.020 234.390 ;
        RECT 255.255 234.230 255.425 234.400 ;
        RECT 242.940 231.185 243.110 231.355 ;
        RECT 244.120 231.165 244.290 231.335 ;
        RECT 262.935 231.505 263.105 231.675 ;
        RECT 270.390 232.235 270.560 232.405 ;
        RECT 268.530 231.800 268.700 231.970 ;
        RECT 242.920 230.370 243.090 230.540 ;
        RECT 244.050 230.380 244.220 230.550 ;
        RECT 270.935 231.810 271.105 231.980 ;
        RECT 247.415 227.525 247.585 227.695 ;
        RECT 254.870 228.255 255.040 228.425 ;
        RECT 253.010 227.820 253.180 227.990 ;
        RECT 255.380 227.795 255.550 227.965 ;
        RECT 298.215 224.355 298.385 224.525 ;
        RECT 305.670 225.085 305.840 225.255 ;
        RECT 303.810 224.650 303.980 224.820 ;
        RECT 306.230 224.650 306.400 224.820 ;
        RECT 247.395 218.275 247.565 218.445 ;
        RECT 254.850 219.005 255.020 219.175 ;
        RECT 252.990 218.570 253.160 218.740 ;
        RECT 255.395 218.580 255.565 218.750 ;
        RECT 243.080 215.535 243.250 215.705 ;
        RECT 244.260 215.515 244.430 215.685 ;
        RECT 263.075 215.855 263.245 216.025 ;
        RECT 270.530 216.585 270.700 216.755 ;
        RECT 268.670 216.150 268.840 216.320 ;
        RECT 243.060 214.720 243.230 214.890 ;
        RECT 244.190 214.730 244.360 214.900 ;
        RECT 271.075 216.160 271.245 216.330 ;
        RECT 247.555 211.875 247.725 212.045 ;
        RECT 255.010 212.605 255.180 212.775 ;
        RECT 253.150 212.170 253.320 212.340 ;
        RECT 255.520 212.145 255.690 212.315 ;
        RECT 280.655 210.305 280.825 210.475 ;
        RECT 288.110 211.035 288.280 211.205 ;
        RECT 286.250 210.600 286.420 210.770 ;
        RECT 288.645 210.605 288.815 210.775 ;
        RECT 247.225 203.855 247.395 204.025 ;
        RECT 254.680 204.585 254.850 204.755 ;
        RECT 252.820 204.150 252.990 204.320 ;
        RECT 255.225 204.160 255.395 204.330 ;
        RECT 242.910 201.115 243.080 201.285 ;
        RECT 244.090 201.095 244.260 201.265 ;
        RECT 262.905 201.435 263.075 201.605 ;
        RECT 270.360 202.165 270.530 202.335 ;
        RECT 268.500 201.730 268.670 201.900 ;
        RECT 242.890 200.300 243.060 200.470 ;
        RECT 244.020 200.310 244.190 200.480 ;
        RECT 270.905 201.740 271.075 201.910 ;
        RECT 247.385 197.455 247.555 197.625 ;
        RECT 254.840 198.185 255.010 198.355 ;
        RECT 252.980 197.750 253.150 197.920 ;
        RECT 255.350 197.725 255.520 197.895 ;
        RECT 312.415 198.065 312.585 198.235 ;
        RECT 319.870 198.795 320.040 198.965 ;
        RECT 318.010 198.360 318.180 198.530 ;
        RECT 320.430 198.355 320.600 198.525 ;
        RECT 247.075 188.425 247.245 188.595 ;
        RECT 254.530 189.155 254.700 189.325 ;
        RECT 252.670 188.720 252.840 188.890 ;
        RECT 255.075 188.730 255.245 188.900 ;
        RECT 242.760 185.685 242.930 185.855 ;
        RECT 243.940 185.665 244.110 185.835 ;
        RECT 262.755 186.005 262.925 186.175 ;
        RECT 270.210 186.735 270.380 186.905 ;
        RECT 268.350 186.300 268.520 186.470 ;
        RECT 242.740 184.870 242.910 185.040 ;
        RECT 243.870 184.880 244.040 185.050 ;
        RECT 270.755 186.310 270.925 186.480 ;
        RECT 247.235 182.025 247.405 182.195 ;
        RECT 254.690 182.755 254.860 182.925 ;
        RECT 252.830 182.320 253.000 182.490 ;
        RECT 255.200 182.295 255.370 182.465 ;
        RECT 280.335 180.455 280.505 180.625 ;
        RECT 287.790 181.185 287.960 181.355 ;
        RECT 285.930 180.750 286.100 180.920 ;
        RECT 288.325 180.755 288.495 180.925 ;
        RECT 246.905 174.005 247.075 174.175 ;
        RECT 254.360 174.735 254.530 174.905 ;
        RECT 252.500 174.300 252.670 174.470 ;
        RECT 254.905 174.310 255.075 174.480 ;
        RECT 242.590 171.265 242.760 171.435 ;
        RECT 243.770 171.245 243.940 171.415 ;
        RECT 262.585 171.585 262.755 171.755 ;
        RECT 270.040 172.315 270.210 172.485 ;
        RECT 268.180 171.880 268.350 172.050 ;
        RECT 242.570 170.450 242.740 170.620 ;
        RECT 243.700 170.460 243.870 170.630 ;
        RECT 270.585 171.890 270.755 172.060 ;
        RECT 247.065 167.605 247.235 167.775 ;
        RECT 254.520 168.335 254.690 168.505 ;
        RECT 252.660 167.900 252.830 168.070 ;
        RECT 255.030 167.875 255.200 168.045 ;
        RECT 297.865 164.435 298.035 164.605 ;
        RECT 305.320 165.165 305.490 165.335 ;
        RECT 303.460 164.730 303.630 164.900 ;
        RECT 305.880 164.730 306.050 164.900 ;
        RECT 247.045 158.355 247.215 158.525 ;
        RECT 254.500 159.085 254.670 159.255 ;
        RECT 252.640 158.650 252.810 158.820 ;
        RECT 255.045 158.660 255.215 158.830 ;
        RECT 242.730 155.615 242.900 155.785 ;
        RECT 243.910 155.595 244.080 155.765 ;
        RECT 262.725 155.935 262.895 156.105 ;
        RECT 270.180 156.665 270.350 156.835 ;
        RECT 268.320 156.230 268.490 156.400 ;
        RECT 242.710 154.800 242.880 154.970 ;
        RECT 243.840 154.810 244.010 154.980 ;
        RECT 270.725 156.240 270.895 156.410 ;
        RECT 247.205 151.955 247.375 152.125 ;
        RECT 254.660 152.685 254.830 152.855 ;
        RECT 252.800 152.250 252.970 152.420 ;
        RECT 255.170 152.225 255.340 152.395 ;
        RECT 280.305 150.385 280.475 150.555 ;
        RECT 287.760 151.115 287.930 151.285 ;
        RECT 285.900 150.680 286.070 150.850 ;
        RECT 348.735 248.155 348.905 248.325 ;
        RECT 356.190 248.885 356.360 249.055 ;
        RECT 354.330 248.450 354.500 248.620 ;
        RECT 356.735 248.460 356.905 248.630 ;
        RECT 344.420 245.415 344.590 245.585 ;
        RECT 345.600 245.395 345.770 245.565 ;
        RECT 364.415 245.735 364.585 245.905 ;
        RECT 371.870 246.465 372.040 246.635 ;
        RECT 370.010 246.030 370.180 246.200 ;
        RECT 344.400 244.600 344.570 244.770 ;
        RECT 345.530 244.610 345.700 244.780 ;
        RECT 372.415 246.040 372.585 246.210 ;
        RECT 348.895 241.755 349.065 241.925 ;
        RECT 356.350 242.485 356.520 242.655 ;
        RECT 354.490 242.050 354.660 242.220 ;
        RECT 356.860 242.025 357.030 242.195 ;
        RECT 381.995 240.185 382.165 240.355 ;
        RECT 389.450 240.915 389.620 241.085 ;
        RECT 387.590 240.480 387.760 240.650 ;
        RECT 389.985 240.485 390.155 240.655 ;
        RECT 348.565 233.735 348.735 233.905 ;
        RECT 356.020 234.465 356.190 234.635 ;
        RECT 354.160 234.030 354.330 234.200 ;
        RECT 356.565 234.040 356.735 234.210 ;
        RECT 344.250 230.995 344.420 231.165 ;
        RECT 345.430 230.975 345.600 231.145 ;
        RECT 364.245 231.315 364.415 231.485 ;
        RECT 371.700 232.045 371.870 232.215 ;
        RECT 369.840 231.610 370.010 231.780 ;
        RECT 344.230 230.180 344.400 230.350 ;
        RECT 345.360 230.190 345.530 230.360 ;
        RECT 372.245 231.620 372.415 231.790 ;
        RECT 348.725 227.335 348.895 227.505 ;
        RECT 356.180 228.065 356.350 228.235 ;
        RECT 354.320 227.630 354.490 227.800 ;
        RECT 356.690 227.605 356.860 227.775 ;
        RECT 399.525 224.165 399.695 224.335 ;
        RECT 406.980 224.895 407.150 225.065 ;
        RECT 405.120 224.460 405.290 224.630 ;
        RECT 407.540 224.460 407.710 224.630 ;
        RECT 348.705 218.085 348.875 218.255 ;
        RECT 356.160 218.815 356.330 218.985 ;
        RECT 354.300 218.380 354.470 218.550 ;
        RECT 356.705 218.390 356.875 218.560 ;
        RECT 344.390 215.345 344.560 215.515 ;
        RECT 345.570 215.325 345.740 215.495 ;
        RECT 364.385 215.665 364.555 215.835 ;
        RECT 371.840 216.395 372.010 216.565 ;
        RECT 369.980 215.960 370.150 216.130 ;
        RECT 344.370 214.530 344.540 214.700 ;
        RECT 345.500 214.540 345.670 214.710 ;
        RECT 372.385 215.970 372.555 216.140 ;
        RECT 348.865 211.685 349.035 211.855 ;
        RECT 356.320 212.415 356.490 212.585 ;
        RECT 354.460 211.980 354.630 212.150 ;
        RECT 356.830 211.955 357.000 212.125 ;
        RECT 381.965 210.115 382.135 210.285 ;
        RECT 389.420 210.845 389.590 211.015 ;
        RECT 387.560 210.410 387.730 210.580 ;
        RECT 389.955 210.415 390.125 210.585 ;
        RECT 348.535 203.665 348.705 203.835 ;
        RECT 355.990 204.395 356.160 204.565 ;
        RECT 354.130 203.960 354.300 204.130 ;
        RECT 356.535 203.970 356.705 204.140 ;
        RECT 344.220 200.925 344.390 201.095 ;
        RECT 345.400 200.905 345.570 201.075 ;
        RECT 364.215 201.245 364.385 201.415 ;
        RECT 371.670 201.975 371.840 202.145 ;
        RECT 369.810 201.540 369.980 201.710 ;
        RECT 344.200 200.110 344.370 200.280 ;
        RECT 345.330 200.120 345.500 200.290 ;
        RECT 372.215 201.550 372.385 201.720 ;
        RECT 348.695 197.265 348.865 197.435 ;
        RECT 356.150 197.995 356.320 198.165 ;
        RECT 354.290 197.560 354.460 197.730 ;
        RECT 356.660 197.535 356.830 197.705 ;
        RECT 413.725 197.875 413.895 198.045 ;
        RECT 421.180 198.605 421.350 198.775 ;
        RECT 419.320 198.170 419.490 198.340 ;
        RECT 421.740 198.165 421.910 198.335 ;
        RECT 348.385 188.235 348.555 188.405 ;
        RECT 355.840 188.965 356.010 189.135 ;
        RECT 353.980 188.530 354.150 188.700 ;
        RECT 356.385 188.540 356.555 188.710 ;
        RECT 344.070 185.495 344.240 185.665 ;
        RECT 345.250 185.475 345.420 185.645 ;
        RECT 364.065 185.815 364.235 185.985 ;
        RECT 371.520 186.545 371.690 186.715 ;
        RECT 369.660 186.110 369.830 186.280 ;
        RECT 344.050 184.680 344.220 184.850 ;
        RECT 345.180 184.690 345.350 184.860 ;
        RECT 372.065 186.120 372.235 186.290 ;
        RECT 348.545 181.835 348.715 182.005 ;
        RECT 356.000 182.565 356.170 182.735 ;
        RECT 354.140 182.130 354.310 182.300 ;
        RECT 356.510 182.105 356.680 182.275 ;
        RECT 381.645 180.265 381.815 180.435 ;
        RECT 389.100 180.995 389.270 181.165 ;
        RECT 387.240 180.560 387.410 180.730 ;
        RECT 389.635 180.565 389.805 180.735 ;
        RECT 348.215 173.815 348.385 173.985 ;
        RECT 355.670 174.545 355.840 174.715 ;
        RECT 353.810 174.110 353.980 174.280 ;
        RECT 356.215 174.120 356.385 174.290 ;
        RECT 343.900 171.075 344.070 171.245 ;
        RECT 345.080 171.055 345.250 171.225 ;
        RECT 363.895 171.395 364.065 171.565 ;
        RECT 371.350 172.125 371.520 172.295 ;
        RECT 369.490 171.690 369.660 171.860 ;
        RECT 343.880 170.260 344.050 170.430 ;
        RECT 345.010 170.270 345.180 170.440 ;
        RECT 371.895 171.700 372.065 171.870 ;
        RECT 348.375 167.415 348.545 167.585 ;
        RECT 355.830 168.145 356.000 168.315 ;
        RECT 353.970 167.710 354.140 167.880 ;
        RECT 356.340 167.685 356.510 167.855 ;
        RECT 288.295 150.685 288.465 150.855 ;
        RECT 246.875 143.935 247.045 144.105 ;
        RECT 254.330 144.665 254.500 144.835 ;
        RECT 252.470 144.230 252.640 144.400 ;
        RECT 254.875 144.240 255.045 144.410 ;
        RECT 242.560 141.195 242.730 141.365 ;
        RECT 243.740 141.175 243.910 141.345 ;
        RECT 262.555 141.515 262.725 141.685 ;
        RECT 270.010 142.245 270.180 142.415 ;
        RECT 399.175 164.245 399.345 164.415 ;
        RECT 406.630 164.975 406.800 165.145 ;
        RECT 404.770 164.540 404.940 164.710 ;
        RECT 407.190 164.540 407.360 164.710 ;
        RECT 348.355 158.165 348.525 158.335 ;
        RECT 355.810 158.895 355.980 159.065 ;
        RECT 353.950 158.460 354.120 158.630 ;
        RECT 356.355 158.470 356.525 158.640 ;
        RECT 344.040 155.425 344.210 155.595 ;
        RECT 345.220 155.405 345.390 155.575 ;
        RECT 364.035 155.745 364.205 155.915 ;
        RECT 371.490 156.475 371.660 156.645 ;
        RECT 369.630 156.040 369.800 156.210 ;
        RECT 344.020 154.610 344.190 154.780 ;
        RECT 345.150 154.620 345.320 154.790 ;
        RECT 372.035 156.050 372.205 156.220 ;
        RECT 348.515 151.765 348.685 151.935 ;
        RECT 355.970 152.495 356.140 152.665 ;
        RECT 354.110 152.060 354.280 152.230 ;
        RECT 356.480 152.035 356.650 152.205 ;
        RECT 381.615 150.195 381.785 150.365 ;
        RECT 389.070 150.925 389.240 151.095 ;
        RECT 387.210 150.490 387.380 150.660 ;
        RECT 389.605 150.495 389.775 150.665 ;
        RECT 268.150 141.810 268.320 141.980 ;
        RECT 242.540 140.380 242.710 140.550 ;
        RECT 243.670 140.390 243.840 140.560 ;
        RECT 270.555 141.820 270.725 141.990 ;
        RECT 247.035 137.535 247.205 137.705 ;
        RECT 254.490 138.265 254.660 138.435 ;
        RECT 348.185 143.745 348.355 143.915 ;
        RECT 355.640 144.475 355.810 144.645 ;
        RECT 353.780 144.040 353.950 144.210 ;
        RECT 356.185 144.050 356.355 144.220 ;
        RECT 252.630 137.830 252.800 138.000 ;
        RECT 255.000 137.805 255.170 137.975 ;
        RECT 328.745 134.925 328.915 135.095 ;
        RECT 336.200 135.655 336.370 135.825 ;
        RECT 343.870 141.005 344.040 141.175 ;
        RECT 345.050 140.985 345.220 141.155 ;
        RECT 363.865 141.325 364.035 141.495 ;
        RECT 371.320 142.055 371.490 142.225 ;
        RECT 369.460 141.620 369.630 141.790 ;
        RECT 343.850 140.190 344.020 140.360 ;
        RECT 344.980 140.200 345.150 140.370 ;
        RECT 371.865 141.630 372.035 141.800 ;
        RECT 348.345 137.345 348.515 137.515 ;
        RECT 355.800 138.075 355.970 138.245 ;
        RECT 353.940 137.640 354.110 137.810 ;
        RECT 356.310 137.615 356.480 137.785 ;
        RECT 463.790 137.795 463.960 137.965 ;
        RECT 456.335 137.065 456.505 137.235 ;
        RECT 334.340 135.220 334.510 135.390 ;
        RECT 336.805 135.230 336.975 135.400 ;
        RECT 430.055 134.735 430.225 134.905 ;
        RECT 437.510 135.465 437.680 135.635 ;
        RECT 435.650 135.030 435.820 135.200 ;
        RECT 438.115 135.040 438.285 135.210 ;
        RECT 481.090 135.445 481.260 135.615 ;
        RECT 473.635 134.715 473.805 134.885 ;
        RECT 246.925 128.105 247.095 128.275 ;
        RECT 254.380 128.835 254.550 129.005 ;
        RECT 252.520 128.400 252.690 128.570 ;
        RECT 254.925 128.410 255.095 128.580 ;
        RECT 242.610 125.365 242.780 125.535 ;
        RECT 243.790 125.345 243.960 125.515 ;
        RECT 262.605 125.685 262.775 125.855 ;
        RECT 270.060 126.415 270.230 126.585 ;
        RECT 268.200 125.980 268.370 126.150 ;
        RECT 242.590 124.550 242.760 124.720 ;
        RECT 243.720 124.560 243.890 124.730 ;
        RECT 270.605 125.990 270.775 126.160 ;
        RECT 247.085 121.705 247.255 121.875 ;
        RECT 254.540 122.435 254.710 122.605 ;
        RECT 252.680 122.000 252.850 122.170 ;
        RECT 255.050 121.975 255.220 122.145 ;
        RECT 280.185 120.135 280.355 120.305 ;
        RECT 287.640 120.865 287.810 121.035 ;
        RECT 285.780 120.430 285.950 120.600 ;
        RECT 288.175 120.435 288.345 120.605 ;
        RECT 246.755 113.685 246.925 113.855 ;
        RECT 254.210 114.415 254.380 114.585 ;
        RECT 252.350 113.980 252.520 114.150 ;
        RECT 254.755 113.990 254.925 114.160 ;
        RECT 242.440 110.945 242.610 111.115 ;
        RECT 243.620 110.925 243.790 111.095 ;
        RECT 262.435 111.265 262.605 111.435 ;
        RECT 269.890 111.995 270.060 112.165 ;
        RECT 268.030 111.560 268.200 111.730 ;
        RECT 242.420 110.130 242.590 110.300 ;
        RECT 243.550 110.140 243.720 110.310 ;
        RECT 270.435 111.570 270.605 111.740 ;
        RECT 246.915 107.285 247.085 107.455 ;
        RECT 254.370 108.015 254.540 108.185 ;
        RECT 252.510 107.580 252.680 107.750 ;
        RECT 254.880 107.555 255.050 107.725 ;
        RECT 297.715 104.115 297.885 104.285 ;
        RECT 305.170 104.845 305.340 105.015 ;
        RECT 303.310 104.410 303.480 104.580 ;
        RECT 305.730 104.410 305.900 104.580 ;
        RECT 246.895 98.035 247.065 98.205 ;
        RECT 254.350 98.765 254.520 98.935 ;
        RECT 252.490 98.330 252.660 98.500 ;
        RECT 254.895 98.340 255.065 98.510 ;
        RECT 242.580 95.295 242.750 95.465 ;
        RECT 243.760 95.275 243.930 95.445 ;
        RECT 262.575 95.615 262.745 95.785 ;
        RECT 270.030 96.345 270.200 96.515 ;
        RECT 268.170 95.910 268.340 96.080 ;
        RECT 242.560 94.480 242.730 94.650 ;
        RECT 243.690 94.490 243.860 94.660 ;
        RECT 270.575 95.920 270.745 96.090 ;
        RECT 247.055 91.635 247.225 91.805 ;
        RECT 254.510 92.365 254.680 92.535 ;
        RECT 252.650 91.930 252.820 92.100 ;
        RECT 255.020 91.905 255.190 92.075 ;
        RECT 280.155 90.065 280.325 90.235 ;
        RECT 287.610 90.795 287.780 90.965 ;
        RECT 285.750 90.360 285.920 90.530 ;
        RECT 288.145 90.365 288.315 90.535 ;
        RECT 246.725 83.615 246.895 83.785 ;
        RECT 254.180 84.345 254.350 84.515 ;
        RECT 252.320 83.910 252.490 84.080 ;
        RECT 254.725 83.920 254.895 84.090 ;
        RECT 242.410 80.875 242.580 81.045 ;
        RECT 243.590 80.855 243.760 81.025 ;
        RECT 262.405 81.195 262.575 81.365 ;
        RECT 269.860 81.925 270.030 82.095 ;
        RECT 268.000 81.490 268.170 81.660 ;
        RECT 242.390 80.060 242.560 80.230 ;
        RECT 243.520 80.070 243.690 80.240 ;
        RECT 270.405 81.500 270.575 81.670 ;
        RECT 246.885 77.215 247.055 77.385 ;
        RECT 254.340 77.945 254.510 78.115 ;
        RECT 252.480 77.510 252.650 77.680 ;
        RECT 254.850 77.485 255.020 77.655 ;
        RECT 311.915 77.825 312.085 77.995 ;
        RECT 319.370 78.555 319.540 78.725 ;
        RECT 348.235 127.915 348.405 128.085 ;
        RECT 355.690 128.645 355.860 128.815 ;
        RECT 353.830 128.210 354.000 128.380 ;
        RECT 356.235 128.220 356.405 128.390 ;
        RECT 343.920 125.175 344.090 125.345 ;
        RECT 345.100 125.155 345.270 125.325 ;
        RECT 363.915 125.495 364.085 125.665 ;
        RECT 371.370 126.225 371.540 126.395 ;
        RECT 369.510 125.790 369.680 125.960 ;
        RECT 343.900 124.360 344.070 124.530 ;
        RECT 345.030 124.370 345.200 124.540 ;
        RECT 371.915 125.800 372.085 125.970 ;
        RECT 348.395 121.515 348.565 121.685 ;
        RECT 355.850 122.245 356.020 122.415 ;
        RECT 353.990 121.810 354.160 121.980 ;
        RECT 356.360 121.785 356.530 121.955 ;
        RECT 381.495 119.945 381.665 120.115 ;
        RECT 388.950 120.675 389.120 120.845 ;
        RECT 387.090 120.240 387.260 120.410 ;
        RECT 389.485 120.245 389.655 120.415 ;
        RECT 348.065 113.495 348.235 113.665 ;
        RECT 355.520 114.225 355.690 114.395 ;
        RECT 353.660 113.790 353.830 113.960 ;
        RECT 356.065 113.800 356.235 113.970 ;
        RECT 343.750 110.755 343.920 110.925 ;
        RECT 344.930 110.735 345.100 110.905 ;
        RECT 363.745 111.075 363.915 111.245 ;
        RECT 371.200 111.805 371.370 111.975 ;
        RECT 369.340 111.370 369.510 111.540 ;
        RECT 343.730 109.940 343.900 110.110 ;
        RECT 344.860 109.950 345.030 110.120 ;
        RECT 371.745 111.380 371.915 111.550 ;
        RECT 348.225 107.095 348.395 107.265 ;
        RECT 355.680 107.825 355.850 107.995 ;
        RECT 353.820 107.390 353.990 107.560 ;
        RECT 356.190 107.365 356.360 107.535 ;
        RECT 399.025 103.925 399.195 104.095 ;
        RECT 406.480 104.655 406.650 104.825 ;
        RECT 404.620 104.220 404.790 104.390 ;
        RECT 407.040 104.220 407.210 104.390 ;
        RECT 348.205 97.845 348.375 98.015 ;
        RECT 355.660 98.575 355.830 98.745 ;
        RECT 353.800 98.140 353.970 98.310 ;
        RECT 356.205 98.150 356.375 98.320 ;
        RECT 343.890 95.105 344.060 95.275 ;
        RECT 345.070 95.085 345.240 95.255 ;
        RECT 363.885 95.425 364.055 95.595 ;
        RECT 371.340 96.155 371.510 96.325 ;
        RECT 369.480 95.720 369.650 95.890 ;
        RECT 343.870 94.290 344.040 94.460 ;
        RECT 345.000 94.300 345.170 94.470 ;
        RECT 371.885 95.730 372.055 95.900 ;
        RECT 348.365 91.445 348.535 91.615 ;
        RECT 355.820 92.175 355.990 92.345 ;
        RECT 353.960 91.740 354.130 91.910 ;
        RECT 356.330 91.715 356.500 91.885 ;
        RECT 381.465 89.875 381.635 90.045 ;
        RECT 388.920 90.605 389.090 90.775 ;
        RECT 387.060 90.170 387.230 90.340 ;
        RECT 389.455 90.175 389.625 90.345 ;
        RECT 348.035 83.425 348.205 83.595 ;
        RECT 355.490 84.155 355.660 84.325 ;
        RECT 353.630 83.720 353.800 83.890 ;
        RECT 356.035 83.730 356.205 83.900 ;
        RECT 343.720 80.685 343.890 80.855 ;
        RECT 344.900 80.665 345.070 80.835 ;
        RECT 363.715 81.005 363.885 81.175 ;
        RECT 371.170 81.735 371.340 81.905 ;
        RECT 369.310 81.300 369.480 81.470 ;
        RECT 343.700 79.870 343.870 80.040 ;
        RECT 344.830 79.880 345.000 80.050 ;
        RECT 317.510 78.120 317.680 78.290 ;
        RECT 319.930 78.115 320.100 78.285 ;
        RECT 371.715 81.310 371.885 81.480 ;
        RECT 348.195 77.025 348.365 77.195 ;
        RECT 355.650 77.755 355.820 77.925 ;
        RECT 353.790 77.320 353.960 77.490 ;
        RECT 356.160 77.295 356.330 77.465 ;
        RECT 413.225 77.635 413.395 77.805 ;
        RECT 420.680 78.365 420.850 78.535 ;
        RECT 246.575 68.185 246.745 68.355 ;
        RECT 254.030 68.915 254.200 69.085 ;
        RECT 252.170 68.480 252.340 68.650 ;
        RECT 254.575 68.490 254.745 68.660 ;
        RECT 242.260 65.445 242.430 65.615 ;
        RECT 243.440 65.425 243.610 65.595 ;
        RECT 262.255 65.765 262.425 65.935 ;
        RECT 269.710 66.495 269.880 66.665 ;
        RECT 267.850 66.060 268.020 66.230 ;
        RECT 242.240 64.630 242.410 64.800 ;
        RECT 243.370 64.640 243.540 64.810 ;
        RECT 270.255 66.070 270.425 66.240 ;
        RECT 418.820 77.930 418.990 78.100 ;
        RECT 421.240 77.925 421.410 78.095 ;
        RECT 347.885 67.995 348.055 68.165 ;
        RECT 355.340 68.725 355.510 68.895 ;
        RECT 353.480 68.290 353.650 68.460 ;
        RECT 355.885 68.300 356.055 68.470 ;
        RECT 246.735 61.785 246.905 61.955 ;
        RECT 254.190 62.515 254.360 62.685 ;
        RECT 252.330 62.080 252.500 62.250 ;
        RECT 254.700 62.055 254.870 62.225 ;
        RECT 279.835 60.215 280.005 60.385 ;
        RECT 287.290 60.945 287.460 61.115 ;
        RECT 285.430 60.510 285.600 60.680 ;
        RECT 287.825 60.515 287.995 60.685 ;
        RECT 246.405 53.765 246.575 53.935 ;
        RECT 253.860 54.495 254.030 54.665 ;
        RECT 252.000 54.060 252.170 54.230 ;
        RECT 254.405 54.070 254.575 54.240 ;
        RECT 242.090 51.025 242.260 51.195 ;
        RECT 243.270 51.005 243.440 51.175 ;
        RECT 262.085 51.345 262.255 51.515 ;
        RECT 269.540 52.075 269.710 52.245 ;
        RECT 267.680 51.640 267.850 51.810 ;
        RECT 242.070 50.210 242.240 50.380 ;
        RECT 243.200 50.220 243.370 50.390 ;
        RECT 270.085 51.650 270.255 51.820 ;
        RECT 246.565 47.365 246.735 47.535 ;
        RECT 254.020 48.095 254.190 48.265 ;
        RECT 252.160 47.660 252.330 47.830 ;
        RECT 254.530 47.635 254.700 47.805 ;
        RECT 343.570 65.255 343.740 65.425 ;
        RECT 344.750 65.235 344.920 65.405 ;
        RECT 363.565 65.575 363.735 65.745 ;
        RECT 371.020 66.305 371.190 66.475 ;
        RECT 369.160 65.870 369.330 66.040 ;
        RECT 343.550 64.440 343.720 64.610 ;
        RECT 344.680 64.450 344.850 64.620 ;
        RECT 371.565 65.880 371.735 66.050 ;
        RECT 348.045 61.595 348.215 61.765 ;
        RECT 355.500 62.325 355.670 62.495 ;
        RECT 353.640 61.890 353.810 62.060 ;
        RECT 356.010 61.865 356.180 62.035 ;
        RECT 381.145 60.025 381.315 60.195 ;
        RECT 388.600 60.755 388.770 60.925 ;
        RECT 386.740 60.320 386.910 60.490 ;
        RECT 389.135 60.325 389.305 60.495 ;
        RECT 347.715 53.575 347.885 53.745 ;
        RECT 355.170 54.305 355.340 54.475 ;
        RECT 353.310 53.870 353.480 54.040 ;
        RECT 355.715 53.880 355.885 54.050 ;
        RECT 343.400 50.835 343.570 51.005 ;
        RECT 344.580 50.815 344.750 50.985 ;
        RECT 363.395 51.155 363.565 51.325 ;
        RECT 370.850 51.885 371.020 52.055 ;
        RECT 368.990 51.450 369.160 51.620 ;
        RECT 343.380 50.020 343.550 50.190 ;
        RECT 344.510 50.030 344.680 50.200 ;
        RECT 371.395 51.460 371.565 51.630 ;
        RECT 297.365 44.195 297.535 44.365 ;
        RECT 304.820 44.925 304.990 45.095 ;
        RECT 347.875 47.175 348.045 47.345 ;
        RECT 355.330 47.905 355.500 48.075 ;
        RECT 353.470 47.470 353.640 47.640 ;
        RECT 355.840 47.445 356.010 47.615 ;
        RECT 302.960 44.490 303.130 44.660 ;
        RECT 305.380 44.490 305.550 44.660 ;
        RECT 398.675 44.005 398.845 44.175 ;
        RECT 406.130 44.735 406.300 44.905 ;
        RECT 404.270 44.300 404.440 44.470 ;
        RECT 406.690 44.300 406.860 44.470 ;
        RECT 246.545 38.115 246.715 38.285 ;
        RECT 254.000 38.845 254.170 39.015 ;
        RECT 252.140 38.410 252.310 38.580 ;
        RECT 254.545 38.420 254.715 38.590 ;
        RECT 242.230 35.375 242.400 35.545 ;
        RECT 243.410 35.355 243.580 35.525 ;
        RECT 262.225 35.695 262.395 35.865 ;
        RECT 269.680 36.425 269.850 36.595 ;
        RECT 267.820 35.990 267.990 36.160 ;
        RECT 242.210 34.560 242.380 34.730 ;
        RECT 243.340 34.570 243.510 34.740 ;
        RECT 270.225 36.000 270.395 36.170 ;
        RECT 246.705 31.715 246.875 31.885 ;
        RECT 254.160 32.445 254.330 32.615 ;
        RECT 252.300 32.010 252.470 32.180 ;
        RECT 254.670 31.985 254.840 32.155 ;
        RECT 279.805 30.145 279.975 30.315 ;
        RECT 287.260 30.875 287.430 31.045 ;
        RECT 285.400 30.440 285.570 30.610 ;
        RECT 347.855 37.925 348.025 38.095 ;
        RECT 355.310 38.655 355.480 38.825 ;
        RECT 353.450 38.220 353.620 38.390 ;
        RECT 355.855 38.230 356.025 38.400 ;
        RECT 343.540 35.185 343.710 35.355 ;
        RECT 344.720 35.165 344.890 35.335 ;
        RECT 363.535 35.505 363.705 35.675 ;
        RECT 370.990 36.235 371.160 36.405 ;
        RECT 369.130 35.800 369.300 35.970 ;
        RECT 343.520 34.370 343.690 34.540 ;
        RECT 344.650 34.380 344.820 34.550 ;
        RECT 371.535 35.810 371.705 35.980 ;
        RECT 348.015 31.525 348.185 31.695 ;
        RECT 355.470 32.255 355.640 32.425 ;
        RECT 353.610 31.820 353.780 31.990 ;
        RECT 355.980 31.795 356.150 31.965 ;
        RECT 287.795 30.445 287.965 30.615 ;
        RECT 381.115 29.955 381.285 30.125 ;
        RECT 388.570 30.685 388.740 30.855 ;
        RECT 386.710 30.250 386.880 30.420 ;
        RECT 389.105 30.255 389.275 30.425 ;
        RECT 246.375 23.695 246.545 23.865 ;
        RECT 253.830 24.425 254.000 24.595 ;
        RECT 251.970 23.990 252.140 24.160 ;
        RECT 254.375 24.000 254.545 24.170 ;
        RECT 242.060 20.955 242.230 21.125 ;
        RECT 243.240 20.935 243.410 21.105 ;
        RECT 262.055 21.275 262.225 21.445 ;
        RECT 269.510 22.005 269.680 22.175 ;
        RECT 347.685 23.505 347.855 23.675 ;
        RECT 355.140 24.235 355.310 24.405 ;
        RECT 353.280 23.800 353.450 23.970 ;
        RECT 355.685 23.810 355.855 23.980 ;
        RECT 267.650 21.570 267.820 21.740 ;
        RECT 242.040 20.140 242.210 20.310 ;
        RECT 243.170 20.150 243.340 20.320 ;
        RECT 270.055 21.580 270.225 21.750 ;
        RECT 343.370 20.765 343.540 20.935 ;
        RECT 344.550 20.745 344.720 20.915 ;
        RECT 363.365 21.085 363.535 21.255 ;
        RECT 370.820 21.815 370.990 21.985 ;
        RECT 368.960 21.380 369.130 21.550 ;
        RECT 343.350 19.950 343.520 20.120 ;
        RECT 246.535 17.295 246.705 17.465 ;
        RECT 253.990 18.025 254.160 18.195 ;
        RECT 344.480 19.960 344.650 20.130 ;
        RECT 252.130 17.590 252.300 17.760 ;
        RECT 254.500 17.565 254.670 17.735 ;
        RECT 371.365 21.390 371.535 21.560 ;
        RECT 347.845 17.105 348.015 17.275 ;
        RECT 355.300 17.835 355.470 18.005 ;
        RECT 353.440 17.400 353.610 17.570 ;
        RECT 355.810 17.375 355.980 17.545 ;
      LAYER met1 ;
        RECT 100.840 255.680 101.070 255.710 ;
        RECT 100.840 255.430 101.090 255.680 ;
        RECT 337.370 255.620 337.600 255.650 ;
        RECT 100.840 252.230 101.070 255.430 ;
        RECT 337.370 255.370 337.620 255.620 ;
        RECT 100.840 251.980 101.140 252.230 ;
        RECT 337.370 252.170 337.600 255.370 ;
        RECT 337.370 251.920 337.670 252.170 ;
        RECT 12.020 250.980 18.480 251.140 ;
        RECT 12.020 250.930 18.490 250.980 ;
        RECT 12.030 249.840 12.230 250.930 ;
        RECT 11.430 249.640 12.230 249.840 ;
        RECT 11.430 248.640 11.630 249.640 ;
        RECT 18.290 249.390 18.490 250.930 ;
        RECT 113.330 250.790 119.790 250.950 ;
        RECT 248.550 250.920 255.010 251.080 ;
        RECT 248.550 250.870 255.020 250.920 ;
        RECT 113.330 250.740 119.800 250.790 ;
        RECT 113.340 249.650 113.540 250.740 ;
        RECT 112.740 249.450 113.540 249.650 ;
        RECT 18.290 249.090 18.580 249.390 ;
        RECT 16.430 248.640 19.130 248.940 ;
        RECT 10.780 248.350 11.630 248.640 ;
        RECT 27.700 248.560 34.160 248.720 ;
        RECT 27.700 248.510 34.170 248.560 ;
        RECT 27.710 247.420 27.910 248.510 ;
        RECT 27.110 247.220 27.910 247.420 ;
        RECT 27.110 246.220 27.310 247.220 ;
        RECT 33.970 246.970 34.170 248.510 ;
        RECT 112.740 248.450 112.940 249.450 ;
        RECT 119.600 249.200 119.800 250.740 ;
        RECT 248.560 249.780 248.760 250.870 ;
        RECT 247.960 249.580 248.760 249.780 ;
        RECT 119.600 248.900 119.890 249.200 ;
        RECT 117.740 248.450 120.440 248.750 ;
        RECT 247.960 248.580 248.160 249.580 ;
        RECT 254.820 249.330 255.020 250.870 ;
        RECT 349.860 250.730 356.320 250.890 ;
        RECT 349.860 250.680 356.330 250.730 ;
        RECT 349.870 249.590 350.070 250.680 ;
        RECT 349.270 249.390 350.070 249.590 ;
        RECT 254.820 249.030 255.110 249.330 ;
        RECT 252.960 248.580 255.660 248.880 ;
        RECT 112.090 248.160 112.940 248.450 ;
        RECT 129.010 248.370 135.470 248.530 ;
        RECT 129.010 248.320 135.480 248.370 ;
        RECT 129.020 247.230 129.220 248.320 ;
        RECT 128.420 247.030 129.220 247.230 ;
        RECT 33.970 246.670 34.260 246.970 ;
        RECT 32.110 246.220 34.810 246.520 ;
        RECT 26.460 245.930 27.310 246.220 ;
        RECT 128.420 246.030 128.620 247.030 ;
        RECT 135.280 246.780 135.480 248.320 ;
        RECT 247.310 248.290 248.160 248.580 ;
        RECT 264.230 248.500 270.690 248.660 ;
        RECT 264.230 248.450 270.700 248.500 ;
        RECT 264.240 247.360 264.440 248.450 ;
        RECT 263.640 247.160 264.440 247.360 ;
        RECT 135.280 246.480 135.570 246.780 ;
        RECT 133.420 246.030 136.120 246.330 ;
        RECT 263.640 246.160 263.840 247.160 ;
        RECT 270.500 246.910 270.700 248.450 ;
        RECT 349.270 248.390 349.470 249.390 ;
        RECT 356.130 249.140 356.330 250.680 ;
        RECT 356.130 248.840 356.420 249.140 ;
        RECT 354.270 248.390 356.970 248.690 ;
        RECT 348.620 248.100 349.470 248.390 ;
        RECT 365.540 248.310 372.000 248.470 ;
        RECT 365.540 248.260 372.010 248.310 ;
        RECT 365.550 247.170 365.750 248.260 ;
        RECT 364.950 246.970 365.750 247.170 ;
        RECT 270.500 246.610 270.790 246.910 ;
        RECT 268.640 246.160 271.340 246.460 ;
        RECT 6.530 245.830 6.810 245.910 ;
        RECT 7.710 245.870 7.990 245.900 ;
        RECT 7.690 245.830 8.000 245.870 ;
        RECT 6.520 245.640 8.000 245.830 ;
        RECT 127.770 245.740 128.620 246.030 ;
        RECT 262.990 245.870 263.840 246.160 ;
        RECT 364.950 245.970 365.150 246.970 ;
        RECT 371.810 246.720 372.010 248.260 ;
        RECT 371.810 246.420 372.100 246.720 ;
        RECT 369.950 245.970 372.650 246.270 ;
        RECT 243.060 245.770 243.340 245.850 ;
        RECT 244.240 245.810 244.520 245.840 ;
        RECT 244.220 245.770 244.530 245.810 ;
        RECT 107.840 245.640 108.120 245.720 ;
        RECT 109.020 245.680 109.300 245.710 ;
        RECT 109.000 245.640 109.310 245.680 ;
        RECT 6.520 245.630 7.990 245.640 ;
        RECT 6.530 245.580 6.810 245.630 ;
        RECT 7.710 245.570 7.990 245.630 ;
        RECT 107.830 245.450 109.310 245.640 ;
        RECT 243.050 245.580 244.530 245.770 ;
        RECT 364.300 245.680 365.150 245.970 ;
        RECT 344.370 245.580 344.650 245.660 ;
        RECT 345.550 245.620 345.830 245.650 ;
        RECT 345.530 245.580 345.840 245.620 ;
        RECT 243.050 245.570 244.520 245.580 ;
        RECT 243.060 245.520 243.340 245.570 ;
        RECT 244.240 245.510 244.520 245.570 ;
        RECT 107.830 245.440 109.300 245.450 ;
        RECT 107.840 245.390 108.120 245.440 ;
        RECT 109.020 245.380 109.300 245.440 ;
        RECT 344.360 245.390 345.840 245.580 ;
        RECT 344.360 245.380 345.830 245.390 ;
        RECT 344.370 245.330 344.650 245.380 ;
        RECT 345.550 245.320 345.830 245.380 ;
        RECT 6.510 245.050 6.780 245.090 ;
        RECT 7.640 245.050 7.930 245.100 ;
        RECT 6.510 244.860 7.930 245.050 ;
        RECT 243.040 244.990 243.310 245.030 ;
        RECT 244.170 244.990 244.460 245.040 ;
        RECT 6.510 244.760 6.780 244.860 ;
        RECT 7.640 244.770 7.930 244.860 ;
        RECT 107.820 244.860 108.090 244.900 ;
        RECT 108.950 244.860 109.240 244.910 ;
        RECT 12.180 244.580 18.640 244.740 ;
        RECT 107.820 244.670 109.240 244.860 ;
        RECT 243.040 244.800 244.460 244.990 ;
        RECT 243.040 244.700 243.310 244.800 ;
        RECT 244.170 244.710 244.460 244.800 ;
        RECT 344.350 244.800 344.620 244.840 ;
        RECT 345.480 244.800 345.770 244.850 ;
        RECT 12.180 244.530 18.650 244.580 ;
        RECT 107.820 244.570 108.090 244.670 ;
        RECT 108.950 244.580 109.240 244.670 ;
        RECT 12.190 243.440 12.390 244.530 ;
        RECT 11.590 243.240 12.390 243.440 ;
        RECT 11.590 242.240 11.790 243.240 ;
        RECT 18.450 242.990 18.650 244.530 ;
        RECT 113.490 244.390 119.950 244.550 ;
        RECT 248.710 244.520 255.170 244.680 ;
        RECT 344.350 244.610 345.770 244.800 ;
        RECT 248.710 244.470 255.180 244.520 ;
        RECT 344.350 244.510 344.620 244.610 ;
        RECT 345.480 244.520 345.770 244.610 ;
        RECT 113.490 244.340 119.960 244.390 ;
        RECT 113.500 243.250 113.700 244.340 ;
        RECT 45.280 243.010 51.740 243.170 ;
        RECT 112.900 243.050 113.700 243.250 ;
        RECT 18.450 242.690 18.740 242.990 ;
        RECT 45.280 242.960 51.750 243.010 ;
        RECT 16.590 242.240 19.290 242.540 ;
        RECT 10.940 241.950 11.790 242.240 ;
        RECT 45.290 241.870 45.490 242.960 ;
        RECT 44.690 241.670 45.490 241.870 ;
        RECT 44.690 240.670 44.890 241.670 ;
        RECT 51.550 241.420 51.750 242.960 ;
        RECT 112.900 242.050 113.100 243.050 ;
        RECT 119.760 242.800 119.960 244.340 ;
        RECT 248.720 243.380 248.920 244.470 ;
        RECT 248.120 243.180 248.920 243.380 ;
        RECT 146.590 242.820 153.050 242.980 ;
        RECT 119.760 242.500 120.050 242.800 ;
        RECT 146.590 242.770 153.060 242.820 ;
        RECT 117.900 242.050 120.600 242.350 ;
        RECT 112.250 241.760 113.100 242.050 ;
        RECT 146.600 241.680 146.800 242.770 ;
        RECT 146.000 241.480 146.800 241.680 ;
        RECT 51.550 241.120 51.840 241.420 ;
        RECT 49.690 240.670 52.390 240.970 ;
        RECT 44.040 240.380 44.890 240.670 ;
        RECT 146.000 240.480 146.200 241.480 ;
        RECT 152.860 241.230 153.060 242.770 ;
        RECT 248.120 242.180 248.320 243.180 ;
        RECT 254.980 242.930 255.180 244.470 ;
        RECT 350.020 244.330 356.480 244.490 ;
        RECT 350.020 244.280 356.490 244.330 ;
        RECT 350.030 243.190 350.230 244.280 ;
        RECT 281.810 242.950 288.270 243.110 ;
        RECT 349.430 242.990 350.230 243.190 ;
        RECT 254.980 242.630 255.270 242.930 ;
        RECT 281.810 242.900 288.280 242.950 ;
        RECT 253.120 242.180 255.820 242.480 ;
        RECT 247.470 241.890 248.320 242.180 ;
        RECT 281.820 241.810 282.020 242.900 ;
        RECT 281.220 241.610 282.020 241.810 ;
        RECT 152.860 240.930 153.150 241.230 ;
        RECT 151.000 240.480 153.700 240.780 ;
        RECT 281.220 240.610 281.420 241.610 ;
        RECT 288.080 241.360 288.280 242.900 ;
        RECT 349.430 241.990 349.630 242.990 ;
        RECT 356.290 242.740 356.490 244.280 ;
        RECT 383.120 242.760 389.580 242.920 ;
        RECT 356.290 242.440 356.580 242.740 ;
        RECT 383.120 242.710 389.590 242.760 ;
        RECT 354.430 241.990 357.130 242.290 ;
        RECT 348.780 241.700 349.630 241.990 ;
        RECT 383.130 241.620 383.330 242.710 ;
        RECT 382.530 241.420 383.330 241.620 ;
        RECT 288.080 241.060 288.370 241.360 ;
        RECT 286.220 240.610 288.920 240.910 ;
        RECT 145.350 240.190 146.200 240.480 ;
        RECT 280.570 240.320 281.420 240.610 ;
        RECT 382.530 240.420 382.730 241.420 ;
        RECT 389.390 241.170 389.590 242.710 ;
        RECT 389.390 240.870 389.680 241.170 ;
        RECT 387.530 240.420 390.230 240.720 ;
        RECT 381.880 240.130 382.730 240.420 ;
        RECT 11.850 236.560 18.310 236.720 ;
        RECT 11.850 236.510 18.320 236.560 ;
        RECT 11.860 235.420 12.060 236.510 ;
        RECT 11.260 235.220 12.060 235.420 ;
        RECT 11.260 234.220 11.460 235.220 ;
        RECT 18.120 234.970 18.320 236.510 ;
        RECT 113.160 236.370 119.620 236.530 ;
        RECT 248.380 236.500 254.840 236.660 ;
        RECT 248.380 236.450 254.850 236.500 ;
        RECT 113.160 236.320 119.630 236.370 ;
        RECT 113.170 235.230 113.370 236.320 ;
        RECT 112.570 235.030 113.370 235.230 ;
        RECT 18.120 234.670 18.410 234.970 ;
        RECT 16.260 234.220 18.960 234.520 ;
        RECT 10.610 233.930 11.460 234.220 ;
        RECT 27.530 234.140 33.990 234.300 ;
        RECT 27.530 234.090 34.000 234.140 ;
        RECT 27.540 233.000 27.740 234.090 ;
        RECT 26.940 232.800 27.740 233.000 ;
        RECT 26.940 231.800 27.140 232.800 ;
        RECT 33.800 232.550 34.000 234.090 ;
        RECT 112.570 234.030 112.770 235.030 ;
        RECT 119.430 234.780 119.630 236.320 ;
        RECT 248.390 235.360 248.590 236.450 ;
        RECT 247.790 235.160 248.590 235.360 ;
        RECT 119.430 234.480 119.720 234.780 ;
        RECT 117.570 234.030 120.270 234.330 ;
        RECT 247.790 234.160 247.990 235.160 ;
        RECT 254.650 234.910 254.850 236.450 ;
        RECT 349.690 236.310 356.150 236.470 ;
        RECT 349.690 236.260 356.160 236.310 ;
        RECT 349.700 235.170 349.900 236.260 ;
        RECT 349.100 234.970 349.900 235.170 ;
        RECT 254.650 234.610 254.940 234.910 ;
        RECT 252.790 234.160 255.490 234.460 ;
        RECT 111.920 233.740 112.770 234.030 ;
        RECT 128.840 233.950 135.300 234.110 ;
        RECT 128.840 233.900 135.310 233.950 ;
        RECT 128.850 232.810 129.050 233.900 ;
        RECT 128.250 232.610 129.050 232.810 ;
        RECT 33.800 232.250 34.090 232.550 ;
        RECT 31.940 231.800 34.640 232.100 ;
        RECT 26.290 231.510 27.140 231.800 ;
        RECT 128.250 231.610 128.450 232.610 ;
        RECT 135.110 232.360 135.310 233.900 ;
        RECT 247.140 233.870 247.990 234.160 ;
        RECT 264.060 234.080 270.520 234.240 ;
        RECT 264.060 234.030 270.530 234.080 ;
        RECT 264.070 232.940 264.270 234.030 ;
        RECT 263.470 232.740 264.270 232.940 ;
        RECT 135.110 232.060 135.400 232.360 ;
        RECT 133.250 231.610 135.950 231.910 ;
        RECT 263.470 231.740 263.670 232.740 ;
        RECT 270.330 232.490 270.530 234.030 ;
        RECT 349.100 233.970 349.300 234.970 ;
        RECT 355.960 234.720 356.160 236.260 ;
        RECT 355.960 234.420 356.250 234.720 ;
        RECT 354.100 233.970 356.800 234.270 ;
        RECT 348.450 233.680 349.300 233.970 ;
        RECT 365.370 233.890 371.830 234.050 ;
        RECT 365.370 233.840 371.840 233.890 ;
        RECT 365.380 232.750 365.580 233.840 ;
        RECT 364.780 232.550 365.580 232.750 ;
        RECT 270.330 232.190 270.620 232.490 ;
        RECT 268.470 231.740 271.170 232.040 ;
        RECT 6.360 231.410 6.640 231.490 ;
        RECT 7.540 231.450 7.820 231.480 ;
        RECT 7.520 231.410 7.830 231.450 ;
        RECT 6.350 231.220 7.830 231.410 ;
        RECT 127.600 231.320 128.450 231.610 ;
        RECT 262.820 231.450 263.670 231.740 ;
        RECT 364.780 231.550 364.980 232.550 ;
        RECT 371.640 232.300 371.840 233.840 ;
        RECT 371.640 232.000 371.930 232.300 ;
        RECT 369.780 231.550 372.480 231.850 ;
        RECT 242.890 231.350 243.170 231.430 ;
        RECT 244.070 231.390 244.350 231.420 ;
        RECT 244.050 231.350 244.360 231.390 ;
        RECT 107.670 231.220 107.950 231.300 ;
        RECT 108.850 231.260 109.130 231.290 ;
        RECT 108.830 231.220 109.140 231.260 ;
        RECT 6.350 231.210 7.820 231.220 ;
        RECT 6.360 231.160 6.640 231.210 ;
        RECT 7.540 231.150 7.820 231.210 ;
        RECT 107.660 231.030 109.140 231.220 ;
        RECT 242.880 231.160 244.360 231.350 ;
        RECT 364.130 231.260 364.980 231.550 ;
        RECT 344.200 231.160 344.480 231.240 ;
        RECT 345.380 231.200 345.660 231.230 ;
        RECT 345.360 231.160 345.670 231.200 ;
        RECT 242.880 231.150 244.350 231.160 ;
        RECT 242.890 231.100 243.170 231.150 ;
        RECT 244.070 231.090 244.350 231.150 ;
        RECT 107.660 231.020 109.130 231.030 ;
        RECT 107.670 230.970 107.950 231.020 ;
        RECT 108.850 230.960 109.130 231.020 ;
        RECT 344.190 230.970 345.670 231.160 ;
        RECT 344.190 230.960 345.660 230.970 ;
        RECT 344.200 230.910 344.480 230.960 ;
        RECT 345.380 230.900 345.660 230.960 ;
        RECT 6.340 230.630 6.610 230.670 ;
        RECT 7.470 230.630 7.760 230.680 ;
        RECT 6.340 230.440 7.760 230.630 ;
        RECT 242.870 230.570 243.140 230.610 ;
        RECT 244.000 230.570 244.290 230.620 ;
        RECT 6.340 230.340 6.610 230.440 ;
        RECT 7.470 230.350 7.760 230.440 ;
        RECT 107.650 230.440 107.920 230.480 ;
        RECT 108.780 230.440 109.070 230.490 ;
        RECT 12.010 230.160 18.470 230.320 ;
        RECT 107.650 230.250 109.070 230.440 ;
        RECT 242.870 230.380 244.290 230.570 ;
        RECT 242.870 230.280 243.140 230.380 ;
        RECT 244.000 230.290 244.290 230.380 ;
        RECT 344.180 230.380 344.450 230.420 ;
        RECT 345.310 230.380 345.600 230.430 ;
        RECT 12.010 230.110 18.480 230.160 ;
        RECT 107.650 230.150 107.920 230.250 ;
        RECT 108.780 230.160 109.070 230.250 ;
        RECT 12.020 229.020 12.220 230.110 ;
        RECT 11.420 228.820 12.220 229.020 ;
        RECT 11.420 227.820 11.620 228.820 ;
        RECT 18.280 228.570 18.480 230.110 ;
        RECT 113.320 229.970 119.780 230.130 ;
        RECT 248.540 230.100 255.000 230.260 ;
        RECT 344.180 230.190 345.600 230.380 ;
        RECT 248.540 230.050 255.010 230.100 ;
        RECT 344.180 230.090 344.450 230.190 ;
        RECT 345.310 230.100 345.600 230.190 ;
        RECT 113.320 229.920 119.790 229.970 ;
        RECT 113.330 228.830 113.530 229.920 ;
        RECT 112.730 228.630 113.530 228.830 ;
        RECT 18.280 228.270 18.570 228.570 ;
        RECT 16.420 227.820 19.120 228.120 ;
        RECT 10.770 227.530 11.620 227.820 ;
        RECT 112.730 227.630 112.930 228.630 ;
        RECT 119.590 228.380 119.790 229.920 ;
        RECT 248.550 228.960 248.750 230.050 ;
        RECT 247.950 228.760 248.750 228.960 ;
        RECT 119.590 228.080 119.880 228.380 ;
        RECT 117.730 227.630 120.430 227.930 ;
        RECT 247.950 227.760 248.150 228.760 ;
        RECT 254.810 228.510 255.010 230.050 ;
        RECT 349.850 229.910 356.310 230.070 ;
        RECT 349.850 229.860 356.320 229.910 ;
        RECT 349.860 228.770 350.060 229.860 ;
        RECT 349.260 228.570 350.060 228.770 ;
        RECT 254.810 228.210 255.100 228.510 ;
        RECT 252.950 227.760 255.650 228.060 ;
        RECT 112.080 227.340 112.930 227.630 ;
        RECT 247.300 227.470 248.150 227.760 ;
        RECT 349.260 227.570 349.460 228.570 ;
        RECT 356.120 228.320 356.320 229.860 ;
        RECT 356.120 228.020 356.410 228.320 ;
        RECT 354.260 227.570 356.960 227.870 ;
        RECT 348.610 227.280 349.460 227.570 ;
        RECT 62.810 226.990 69.270 227.150 ;
        RECT 62.810 226.940 69.280 226.990 ;
        RECT 62.820 225.850 63.020 226.940 ;
        RECT 62.220 225.650 63.020 225.850 ;
        RECT 62.220 224.650 62.420 225.650 ;
        RECT 69.080 225.400 69.280 226.940 ;
        RECT 164.120 226.800 170.580 226.960 ;
        RECT 299.340 226.930 305.800 227.090 ;
        RECT 299.340 226.880 305.810 226.930 ;
        RECT 164.120 226.750 170.590 226.800 ;
        RECT 164.130 225.660 164.330 226.750 ;
        RECT 163.530 225.460 164.330 225.660 ;
        RECT 69.080 225.100 69.370 225.400 ;
        RECT 67.220 224.650 69.920 224.950 ;
        RECT 61.570 224.360 62.420 224.650 ;
        RECT 163.530 224.460 163.730 225.460 ;
        RECT 170.390 225.210 170.590 226.750 ;
        RECT 299.350 225.790 299.550 226.880 ;
        RECT 298.750 225.590 299.550 225.790 ;
        RECT 170.390 224.910 170.680 225.210 ;
        RECT 168.530 224.460 171.230 224.760 ;
        RECT 298.750 224.590 298.950 225.590 ;
        RECT 305.610 225.340 305.810 226.880 ;
        RECT 400.650 226.740 407.110 226.900 ;
        RECT 400.650 226.690 407.120 226.740 ;
        RECT 400.660 225.600 400.860 226.690 ;
        RECT 400.060 225.400 400.860 225.600 ;
        RECT 305.610 225.040 305.900 225.340 ;
        RECT 303.750 224.590 306.450 224.890 ;
        RECT 162.880 224.170 163.730 224.460 ;
        RECT 298.100 224.300 298.950 224.590 ;
        RECT 400.060 224.400 400.260 225.400 ;
        RECT 406.920 225.150 407.120 226.690 ;
        RECT 406.920 224.850 407.210 225.150 ;
        RECT 405.060 224.400 407.760 224.700 ;
        RECT 399.410 224.110 400.260 224.400 ;
        RECT 11.990 220.910 18.450 221.070 ;
        RECT 11.990 220.860 18.460 220.910 ;
        RECT 12.000 219.770 12.200 220.860 ;
        RECT 11.400 219.570 12.200 219.770 ;
        RECT 11.400 218.570 11.600 219.570 ;
        RECT 18.260 219.320 18.460 220.860 ;
        RECT 113.300 220.720 119.760 220.880 ;
        RECT 248.520 220.850 254.980 221.010 ;
        RECT 248.520 220.800 254.990 220.850 ;
        RECT 113.300 220.670 119.770 220.720 ;
        RECT 113.310 219.580 113.510 220.670 ;
        RECT 112.710 219.380 113.510 219.580 ;
        RECT 18.260 219.020 18.550 219.320 ;
        RECT 16.400 218.570 19.100 218.870 ;
        RECT 10.750 218.280 11.600 218.570 ;
        RECT 27.670 218.490 34.130 218.650 ;
        RECT 27.670 218.440 34.140 218.490 ;
        RECT 27.680 217.350 27.880 218.440 ;
        RECT 27.080 217.150 27.880 217.350 ;
        RECT 27.080 216.150 27.280 217.150 ;
        RECT 33.940 216.900 34.140 218.440 ;
        RECT 112.710 218.380 112.910 219.380 ;
        RECT 119.570 219.130 119.770 220.670 ;
        RECT 248.530 219.710 248.730 220.800 ;
        RECT 247.930 219.510 248.730 219.710 ;
        RECT 119.570 218.830 119.860 219.130 ;
        RECT 117.710 218.380 120.410 218.680 ;
        RECT 247.930 218.510 248.130 219.510 ;
        RECT 254.790 219.260 254.990 220.800 ;
        RECT 349.830 220.660 356.290 220.820 ;
        RECT 349.830 220.610 356.300 220.660 ;
        RECT 349.840 219.520 350.040 220.610 ;
        RECT 349.240 219.320 350.040 219.520 ;
        RECT 254.790 218.960 255.080 219.260 ;
        RECT 252.930 218.510 255.630 218.810 ;
        RECT 112.060 218.090 112.910 218.380 ;
        RECT 128.980 218.300 135.440 218.460 ;
        RECT 128.980 218.250 135.450 218.300 ;
        RECT 128.990 217.160 129.190 218.250 ;
        RECT 128.390 216.960 129.190 217.160 ;
        RECT 33.940 216.600 34.230 216.900 ;
        RECT 32.080 216.150 34.780 216.450 ;
        RECT 26.430 215.860 27.280 216.150 ;
        RECT 128.390 215.960 128.590 216.960 ;
        RECT 135.250 216.710 135.450 218.250 ;
        RECT 247.280 218.220 248.130 218.510 ;
        RECT 264.200 218.430 270.660 218.590 ;
        RECT 264.200 218.380 270.670 218.430 ;
        RECT 264.210 217.290 264.410 218.380 ;
        RECT 263.610 217.090 264.410 217.290 ;
        RECT 135.250 216.410 135.540 216.710 ;
        RECT 133.390 215.960 136.090 216.260 ;
        RECT 263.610 216.090 263.810 217.090 ;
        RECT 270.470 216.840 270.670 218.380 ;
        RECT 349.240 218.320 349.440 219.320 ;
        RECT 356.100 219.070 356.300 220.610 ;
        RECT 356.100 218.770 356.390 219.070 ;
        RECT 354.240 218.320 356.940 218.620 ;
        RECT 348.590 218.030 349.440 218.320 ;
        RECT 365.510 218.240 371.970 218.400 ;
        RECT 365.510 218.190 371.980 218.240 ;
        RECT 365.520 217.100 365.720 218.190 ;
        RECT 364.920 216.900 365.720 217.100 ;
        RECT 270.470 216.540 270.760 216.840 ;
        RECT 268.610 216.090 271.310 216.390 ;
        RECT 6.500 215.760 6.780 215.840 ;
        RECT 7.680 215.800 7.960 215.830 ;
        RECT 7.660 215.760 7.970 215.800 ;
        RECT 6.490 215.570 7.970 215.760 ;
        RECT 127.740 215.670 128.590 215.960 ;
        RECT 262.960 215.800 263.810 216.090 ;
        RECT 364.920 215.900 365.120 216.900 ;
        RECT 371.780 216.650 371.980 218.190 ;
        RECT 371.780 216.350 372.070 216.650 ;
        RECT 369.920 215.900 372.620 216.200 ;
        RECT 243.030 215.700 243.310 215.780 ;
        RECT 244.210 215.740 244.490 215.770 ;
        RECT 244.190 215.700 244.500 215.740 ;
        RECT 107.810 215.570 108.090 215.650 ;
        RECT 108.990 215.610 109.270 215.640 ;
        RECT 108.970 215.570 109.280 215.610 ;
        RECT 6.490 215.560 7.960 215.570 ;
        RECT 6.500 215.510 6.780 215.560 ;
        RECT 7.680 215.500 7.960 215.560 ;
        RECT 107.800 215.380 109.280 215.570 ;
        RECT 243.020 215.510 244.500 215.700 ;
        RECT 364.270 215.610 365.120 215.900 ;
        RECT 344.340 215.510 344.620 215.590 ;
        RECT 345.520 215.550 345.800 215.580 ;
        RECT 345.500 215.510 345.810 215.550 ;
        RECT 243.020 215.500 244.490 215.510 ;
        RECT 243.030 215.450 243.310 215.500 ;
        RECT 244.210 215.440 244.490 215.500 ;
        RECT 107.800 215.370 109.270 215.380 ;
        RECT 107.810 215.320 108.090 215.370 ;
        RECT 108.990 215.310 109.270 215.370 ;
        RECT 344.330 215.320 345.810 215.510 ;
        RECT 344.330 215.310 345.800 215.320 ;
        RECT 344.340 215.260 344.620 215.310 ;
        RECT 345.520 215.250 345.800 215.310 ;
        RECT 6.480 214.980 6.750 215.020 ;
        RECT 7.610 214.980 7.900 215.030 ;
        RECT 6.480 214.790 7.900 214.980 ;
        RECT 243.010 214.920 243.280 214.960 ;
        RECT 244.140 214.920 244.430 214.970 ;
        RECT 6.480 214.690 6.750 214.790 ;
        RECT 7.610 214.700 7.900 214.790 ;
        RECT 107.790 214.790 108.060 214.830 ;
        RECT 108.920 214.790 109.210 214.840 ;
        RECT 12.150 214.510 18.610 214.670 ;
        RECT 107.790 214.600 109.210 214.790 ;
        RECT 243.010 214.730 244.430 214.920 ;
        RECT 243.010 214.630 243.280 214.730 ;
        RECT 244.140 214.640 244.430 214.730 ;
        RECT 344.320 214.730 344.590 214.770 ;
        RECT 345.450 214.730 345.740 214.780 ;
        RECT 12.150 214.460 18.620 214.510 ;
        RECT 107.790 214.500 108.060 214.600 ;
        RECT 108.920 214.510 109.210 214.600 ;
        RECT 12.160 213.370 12.360 214.460 ;
        RECT 11.560 213.170 12.360 213.370 ;
        RECT 11.560 212.170 11.760 213.170 ;
        RECT 18.420 212.920 18.620 214.460 ;
        RECT 113.460 214.320 119.920 214.480 ;
        RECT 248.680 214.450 255.140 214.610 ;
        RECT 344.320 214.540 345.740 214.730 ;
        RECT 248.680 214.400 255.150 214.450 ;
        RECT 344.320 214.440 344.590 214.540 ;
        RECT 345.450 214.450 345.740 214.540 ;
        RECT 113.460 214.270 119.930 214.320 ;
        RECT 113.470 213.180 113.670 214.270 ;
        RECT 45.250 212.940 51.710 213.100 ;
        RECT 112.870 212.980 113.670 213.180 ;
        RECT 18.420 212.620 18.710 212.920 ;
        RECT 45.250 212.890 51.720 212.940 ;
        RECT 16.560 212.170 19.260 212.470 ;
        RECT 10.910 211.880 11.760 212.170 ;
        RECT 45.260 211.800 45.460 212.890 ;
        RECT 44.660 211.600 45.460 211.800 ;
        RECT 44.660 210.600 44.860 211.600 ;
        RECT 51.520 211.350 51.720 212.890 ;
        RECT 112.870 211.980 113.070 212.980 ;
        RECT 119.730 212.730 119.930 214.270 ;
        RECT 248.690 213.310 248.890 214.400 ;
        RECT 248.090 213.110 248.890 213.310 ;
        RECT 146.560 212.750 153.020 212.910 ;
        RECT 119.730 212.430 120.020 212.730 ;
        RECT 146.560 212.700 153.030 212.750 ;
        RECT 117.870 211.980 120.570 212.280 ;
        RECT 112.220 211.690 113.070 211.980 ;
        RECT 146.570 211.610 146.770 212.700 ;
        RECT 145.970 211.410 146.770 211.610 ;
        RECT 51.520 211.050 51.810 211.350 ;
        RECT 49.660 210.600 52.360 210.900 ;
        RECT 44.010 210.310 44.860 210.600 ;
        RECT 145.970 210.410 146.170 211.410 ;
        RECT 152.830 211.160 153.030 212.700 ;
        RECT 248.090 212.110 248.290 213.110 ;
        RECT 254.950 212.860 255.150 214.400 ;
        RECT 349.990 214.260 356.450 214.420 ;
        RECT 349.990 214.210 356.460 214.260 ;
        RECT 350.000 213.120 350.200 214.210 ;
        RECT 281.780 212.880 288.240 213.040 ;
        RECT 349.400 212.920 350.200 213.120 ;
        RECT 254.950 212.560 255.240 212.860 ;
        RECT 281.780 212.830 288.250 212.880 ;
        RECT 253.090 212.110 255.790 212.410 ;
        RECT 247.440 211.820 248.290 212.110 ;
        RECT 281.790 211.740 281.990 212.830 ;
        RECT 281.190 211.540 281.990 211.740 ;
        RECT 152.830 210.860 153.120 211.160 ;
        RECT 150.970 210.410 153.670 210.710 ;
        RECT 281.190 210.540 281.390 211.540 ;
        RECT 288.050 211.290 288.250 212.830 ;
        RECT 349.400 211.920 349.600 212.920 ;
        RECT 356.260 212.670 356.460 214.210 ;
        RECT 383.090 212.690 389.550 212.850 ;
        RECT 356.260 212.370 356.550 212.670 ;
        RECT 383.090 212.640 389.560 212.690 ;
        RECT 354.400 211.920 357.100 212.220 ;
        RECT 348.750 211.630 349.600 211.920 ;
        RECT 383.100 211.550 383.300 212.640 ;
        RECT 382.500 211.350 383.300 211.550 ;
        RECT 288.050 210.990 288.340 211.290 ;
        RECT 286.190 210.540 288.890 210.840 ;
        RECT 145.320 210.120 146.170 210.410 ;
        RECT 280.540 210.250 281.390 210.540 ;
        RECT 382.500 210.350 382.700 211.350 ;
        RECT 389.360 211.100 389.560 212.640 ;
        RECT 389.360 210.800 389.650 211.100 ;
        RECT 387.500 210.350 390.200 210.650 ;
        RECT 381.850 210.060 382.700 210.350 ;
        RECT 11.820 206.490 18.280 206.650 ;
        RECT 11.820 206.440 18.290 206.490 ;
        RECT 11.830 205.350 12.030 206.440 ;
        RECT 11.230 205.150 12.030 205.350 ;
        RECT 11.230 204.150 11.430 205.150 ;
        RECT 18.090 204.900 18.290 206.440 ;
        RECT 113.130 206.300 119.590 206.460 ;
        RECT 248.350 206.430 254.810 206.590 ;
        RECT 248.350 206.380 254.820 206.430 ;
        RECT 113.130 206.250 119.600 206.300 ;
        RECT 113.140 205.160 113.340 206.250 ;
        RECT 112.540 204.960 113.340 205.160 ;
        RECT 18.090 204.600 18.380 204.900 ;
        RECT 16.230 204.150 18.930 204.450 ;
        RECT 10.580 203.860 11.430 204.150 ;
        RECT 27.500 204.070 33.960 204.230 ;
        RECT 27.500 204.020 33.970 204.070 ;
        RECT 27.510 202.930 27.710 204.020 ;
        RECT 26.910 202.730 27.710 202.930 ;
        RECT 26.910 201.730 27.110 202.730 ;
        RECT 33.770 202.480 33.970 204.020 ;
        RECT 112.540 203.960 112.740 204.960 ;
        RECT 119.400 204.710 119.600 206.250 ;
        RECT 248.360 205.290 248.560 206.380 ;
        RECT 247.760 205.090 248.560 205.290 ;
        RECT 119.400 204.410 119.690 204.710 ;
        RECT 117.540 203.960 120.240 204.260 ;
        RECT 247.760 204.090 247.960 205.090 ;
        RECT 254.620 204.840 254.820 206.380 ;
        RECT 349.660 206.240 356.120 206.400 ;
        RECT 349.660 206.190 356.130 206.240 ;
        RECT 349.670 205.100 349.870 206.190 ;
        RECT 349.070 204.900 349.870 205.100 ;
        RECT 254.620 204.540 254.910 204.840 ;
        RECT 252.760 204.090 255.460 204.390 ;
        RECT 111.890 203.670 112.740 203.960 ;
        RECT 128.810 203.880 135.270 204.040 ;
        RECT 128.810 203.830 135.280 203.880 ;
        RECT 128.820 202.740 129.020 203.830 ;
        RECT 128.220 202.540 129.020 202.740 ;
        RECT 33.770 202.180 34.060 202.480 ;
        RECT 31.910 201.730 34.610 202.030 ;
        RECT 26.260 201.440 27.110 201.730 ;
        RECT 128.220 201.540 128.420 202.540 ;
        RECT 135.080 202.290 135.280 203.830 ;
        RECT 247.110 203.800 247.960 204.090 ;
        RECT 264.030 204.010 270.490 204.170 ;
        RECT 264.030 203.960 270.500 204.010 ;
        RECT 264.040 202.870 264.240 203.960 ;
        RECT 263.440 202.670 264.240 202.870 ;
        RECT 135.080 201.990 135.370 202.290 ;
        RECT 133.220 201.540 135.920 201.840 ;
        RECT 263.440 201.670 263.640 202.670 ;
        RECT 270.300 202.420 270.500 203.960 ;
        RECT 349.070 203.900 349.270 204.900 ;
        RECT 355.930 204.650 356.130 206.190 ;
        RECT 355.930 204.350 356.220 204.650 ;
        RECT 354.070 203.900 356.770 204.200 ;
        RECT 348.420 203.610 349.270 203.900 ;
        RECT 365.340 203.820 371.800 203.980 ;
        RECT 365.340 203.770 371.810 203.820 ;
        RECT 365.350 202.680 365.550 203.770 ;
        RECT 364.750 202.480 365.550 202.680 ;
        RECT 270.300 202.120 270.590 202.420 ;
        RECT 268.440 201.670 271.140 201.970 ;
        RECT 6.330 201.340 6.610 201.420 ;
        RECT 7.510 201.380 7.790 201.410 ;
        RECT 7.490 201.340 7.800 201.380 ;
        RECT 6.320 201.150 7.800 201.340 ;
        RECT 127.570 201.250 128.420 201.540 ;
        RECT 262.790 201.380 263.640 201.670 ;
        RECT 364.750 201.480 364.950 202.480 ;
        RECT 371.610 202.230 371.810 203.770 ;
        RECT 371.610 201.930 371.900 202.230 ;
        RECT 369.750 201.480 372.450 201.780 ;
        RECT 242.860 201.280 243.140 201.360 ;
        RECT 244.040 201.320 244.320 201.350 ;
        RECT 244.020 201.280 244.330 201.320 ;
        RECT 107.640 201.150 107.920 201.230 ;
        RECT 108.820 201.190 109.100 201.220 ;
        RECT 108.800 201.150 109.110 201.190 ;
        RECT 6.320 201.140 7.790 201.150 ;
        RECT 6.330 201.090 6.610 201.140 ;
        RECT 7.510 201.080 7.790 201.140 ;
        RECT 107.630 200.960 109.110 201.150 ;
        RECT 242.850 201.090 244.330 201.280 ;
        RECT 364.100 201.190 364.950 201.480 ;
        RECT 344.170 201.090 344.450 201.170 ;
        RECT 345.350 201.130 345.630 201.160 ;
        RECT 345.330 201.090 345.640 201.130 ;
        RECT 242.850 201.080 244.320 201.090 ;
        RECT 242.860 201.030 243.140 201.080 ;
        RECT 244.040 201.020 244.320 201.080 ;
        RECT 107.630 200.950 109.100 200.960 ;
        RECT 107.640 200.900 107.920 200.950 ;
        RECT 108.820 200.890 109.100 200.950 ;
        RECT 344.160 200.900 345.640 201.090 ;
        RECT 344.160 200.890 345.630 200.900 ;
        RECT 77.010 200.700 83.470 200.860 ;
        RECT 344.170 200.840 344.450 200.890 ;
        RECT 345.350 200.830 345.630 200.890 ;
        RECT 77.010 200.650 83.480 200.700 ;
        RECT 6.310 200.560 6.580 200.600 ;
        RECT 7.440 200.560 7.730 200.610 ;
        RECT 6.310 200.370 7.730 200.560 ;
        RECT 6.310 200.270 6.580 200.370 ;
        RECT 7.440 200.280 7.730 200.370 ;
        RECT 11.980 200.090 18.440 200.250 ;
        RECT 11.980 200.040 18.450 200.090 ;
        RECT 11.990 198.950 12.190 200.040 ;
        RECT 11.390 198.750 12.190 198.950 ;
        RECT 11.390 197.750 11.590 198.750 ;
        RECT 18.250 198.500 18.450 200.040 ;
        RECT 77.020 199.560 77.220 200.650 ;
        RECT 76.420 199.360 77.220 199.560 ;
        RECT 18.250 198.200 18.540 198.500 ;
        RECT 76.420 198.360 76.620 199.360 ;
        RECT 83.280 199.110 83.480 200.650 ;
        RECT 178.320 200.510 184.780 200.670 ;
        RECT 313.540 200.640 320.000 200.800 ;
        RECT 313.540 200.590 320.010 200.640 ;
        RECT 178.320 200.460 184.790 200.510 ;
        RECT 107.620 200.370 107.890 200.410 ;
        RECT 108.750 200.370 109.040 200.420 ;
        RECT 107.620 200.180 109.040 200.370 ;
        RECT 107.620 200.080 107.890 200.180 ;
        RECT 108.750 200.090 109.040 200.180 ;
        RECT 113.290 199.900 119.750 200.060 ;
        RECT 113.290 199.850 119.760 199.900 ;
        RECT 83.280 198.810 83.570 199.110 ;
        RECT 113.300 198.760 113.500 199.850 ;
        RECT 81.420 198.610 84.120 198.660 ;
        RECT 81.420 198.380 84.170 198.610 ;
        RECT 112.700 198.560 113.500 198.760 ;
        RECT 81.420 198.360 84.120 198.380 ;
        RECT 75.770 198.070 76.620 198.360 ;
        RECT 16.390 197.750 19.090 198.050 ;
        RECT 10.740 197.460 11.590 197.750 ;
        RECT 112.700 197.560 112.900 198.560 ;
        RECT 119.560 198.310 119.760 199.850 ;
        RECT 178.330 199.370 178.530 200.460 ;
        RECT 177.730 199.170 178.530 199.370 ;
        RECT 119.560 198.010 119.850 198.310 ;
        RECT 177.730 198.170 177.930 199.170 ;
        RECT 184.590 198.920 184.790 200.460 ;
        RECT 242.840 200.500 243.110 200.540 ;
        RECT 243.970 200.500 244.260 200.550 ;
        RECT 242.840 200.310 244.260 200.500 ;
        RECT 242.840 200.210 243.110 200.310 ;
        RECT 243.970 200.220 244.260 200.310 ;
        RECT 248.510 200.030 254.970 200.190 ;
        RECT 248.510 199.980 254.980 200.030 ;
        RECT 184.590 198.620 184.880 198.920 ;
        RECT 248.520 198.890 248.720 199.980 ;
        RECT 247.920 198.690 248.720 198.890 ;
        RECT 182.730 198.420 185.430 198.470 ;
        RECT 182.730 198.190 185.480 198.420 ;
        RECT 182.730 198.170 185.430 198.190 ;
        RECT 177.080 197.880 177.930 198.170 ;
        RECT 117.700 197.560 120.400 197.860 ;
        RECT 247.920 197.690 248.120 198.690 ;
        RECT 254.780 198.440 254.980 199.980 ;
        RECT 313.550 199.500 313.750 200.590 ;
        RECT 312.950 199.300 313.750 199.500 ;
        RECT 254.780 198.140 255.070 198.440 ;
        RECT 312.950 198.300 313.150 199.300 ;
        RECT 319.810 199.050 320.010 200.590 ;
        RECT 414.850 200.450 421.310 200.610 ;
        RECT 414.850 200.400 421.320 200.450 ;
        RECT 344.150 200.310 344.420 200.350 ;
        RECT 345.280 200.310 345.570 200.360 ;
        RECT 344.150 200.120 345.570 200.310 ;
        RECT 344.150 200.020 344.420 200.120 ;
        RECT 345.280 200.030 345.570 200.120 ;
        RECT 349.820 199.840 356.280 200.000 ;
        RECT 349.820 199.790 356.290 199.840 ;
        RECT 319.810 198.750 320.100 199.050 ;
        RECT 349.830 198.700 350.030 199.790 ;
        RECT 317.950 198.550 320.650 198.600 ;
        RECT 317.950 198.320 320.700 198.550 ;
        RECT 349.230 198.500 350.030 198.700 ;
        RECT 317.950 198.300 320.650 198.320 ;
        RECT 312.300 198.010 313.150 198.300 ;
        RECT 252.920 197.690 255.620 197.990 ;
        RECT 112.050 197.270 112.900 197.560 ;
        RECT 247.270 197.400 248.120 197.690 ;
        RECT 349.230 197.500 349.430 198.500 ;
        RECT 356.090 198.250 356.290 199.790 ;
        RECT 414.860 199.310 415.060 200.400 ;
        RECT 414.260 199.110 415.060 199.310 ;
        RECT 356.090 197.950 356.380 198.250 ;
        RECT 414.260 198.110 414.460 199.110 ;
        RECT 421.120 198.860 421.320 200.400 ;
        RECT 421.120 198.560 421.410 198.860 ;
        RECT 419.260 198.360 421.960 198.410 ;
        RECT 419.260 198.130 422.010 198.360 ;
        RECT 419.260 198.110 421.960 198.130 ;
        RECT 413.610 197.820 414.460 198.110 ;
        RECT 354.230 197.500 356.930 197.800 ;
        RECT 348.580 197.210 349.430 197.500 ;
        RECT 11.670 191.060 18.130 191.220 ;
        RECT 11.670 191.010 18.140 191.060 ;
        RECT 11.680 189.920 11.880 191.010 ;
        RECT 11.080 189.720 11.880 189.920 ;
        RECT 11.080 188.720 11.280 189.720 ;
        RECT 17.940 189.470 18.140 191.010 ;
        RECT 112.980 190.870 119.440 191.030 ;
        RECT 248.200 191.000 254.660 191.160 ;
        RECT 248.200 190.950 254.670 191.000 ;
        RECT 112.980 190.820 119.450 190.870 ;
        RECT 112.990 189.730 113.190 190.820 ;
        RECT 112.390 189.530 113.190 189.730 ;
        RECT 17.940 189.170 18.230 189.470 ;
        RECT 16.080 188.720 18.780 189.020 ;
        RECT 10.430 188.430 11.280 188.720 ;
        RECT 27.350 188.640 33.810 188.800 ;
        RECT 27.350 188.590 33.820 188.640 ;
        RECT 27.360 187.500 27.560 188.590 ;
        RECT 26.760 187.300 27.560 187.500 ;
        RECT 26.760 186.300 26.960 187.300 ;
        RECT 33.620 187.050 33.820 188.590 ;
        RECT 112.390 188.530 112.590 189.530 ;
        RECT 119.250 189.280 119.450 190.820 ;
        RECT 248.210 189.860 248.410 190.950 ;
        RECT 247.610 189.660 248.410 189.860 ;
        RECT 119.250 188.980 119.540 189.280 ;
        RECT 117.390 188.530 120.090 188.830 ;
        RECT 247.610 188.660 247.810 189.660 ;
        RECT 254.470 189.410 254.670 190.950 ;
        RECT 349.510 190.810 355.970 190.970 ;
        RECT 349.510 190.760 355.980 190.810 ;
        RECT 349.520 189.670 349.720 190.760 ;
        RECT 348.920 189.470 349.720 189.670 ;
        RECT 254.470 189.110 254.760 189.410 ;
        RECT 252.610 188.660 255.310 188.960 ;
        RECT 111.740 188.240 112.590 188.530 ;
        RECT 128.660 188.450 135.120 188.610 ;
        RECT 128.660 188.400 135.130 188.450 ;
        RECT 128.670 187.310 128.870 188.400 ;
        RECT 128.070 187.110 128.870 187.310 ;
        RECT 33.620 186.750 33.910 187.050 ;
        RECT 31.760 186.300 34.460 186.600 ;
        RECT 26.110 186.010 26.960 186.300 ;
        RECT 128.070 186.110 128.270 187.110 ;
        RECT 134.930 186.860 135.130 188.400 ;
        RECT 246.960 188.370 247.810 188.660 ;
        RECT 263.880 188.580 270.340 188.740 ;
        RECT 263.880 188.530 270.350 188.580 ;
        RECT 263.890 187.440 264.090 188.530 ;
        RECT 263.290 187.240 264.090 187.440 ;
        RECT 134.930 186.560 135.220 186.860 ;
        RECT 133.070 186.110 135.770 186.410 ;
        RECT 263.290 186.240 263.490 187.240 ;
        RECT 270.150 186.990 270.350 188.530 ;
        RECT 348.920 188.470 349.120 189.470 ;
        RECT 355.780 189.220 355.980 190.760 ;
        RECT 355.780 188.920 356.070 189.220 ;
        RECT 353.920 188.470 356.620 188.770 ;
        RECT 348.270 188.180 349.120 188.470 ;
        RECT 365.190 188.390 371.650 188.550 ;
        RECT 365.190 188.340 371.660 188.390 ;
        RECT 365.200 187.250 365.400 188.340 ;
        RECT 364.600 187.050 365.400 187.250 ;
        RECT 270.150 186.690 270.440 186.990 ;
        RECT 268.290 186.240 270.990 186.540 ;
        RECT 6.180 185.910 6.460 185.990 ;
        RECT 7.360 185.950 7.640 185.980 ;
        RECT 7.340 185.910 7.650 185.950 ;
        RECT 6.170 185.720 7.650 185.910 ;
        RECT 127.420 185.820 128.270 186.110 ;
        RECT 262.640 185.950 263.490 186.240 ;
        RECT 364.600 186.050 364.800 187.050 ;
        RECT 371.460 186.800 371.660 188.340 ;
        RECT 371.460 186.500 371.750 186.800 ;
        RECT 369.600 186.050 372.300 186.350 ;
        RECT 242.710 185.850 242.990 185.930 ;
        RECT 243.890 185.890 244.170 185.920 ;
        RECT 243.870 185.850 244.180 185.890 ;
        RECT 107.490 185.720 107.770 185.800 ;
        RECT 108.670 185.760 108.950 185.790 ;
        RECT 108.650 185.720 108.960 185.760 ;
        RECT 6.170 185.710 7.640 185.720 ;
        RECT 6.180 185.660 6.460 185.710 ;
        RECT 7.360 185.650 7.640 185.710 ;
        RECT 107.480 185.530 108.960 185.720 ;
        RECT 242.700 185.660 244.180 185.850 ;
        RECT 363.950 185.760 364.800 186.050 ;
        RECT 344.020 185.660 344.300 185.740 ;
        RECT 345.200 185.700 345.480 185.730 ;
        RECT 345.180 185.660 345.490 185.700 ;
        RECT 242.700 185.650 244.170 185.660 ;
        RECT 242.710 185.600 242.990 185.650 ;
        RECT 243.890 185.590 244.170 185.650 ;
        RECT 107.480 185.520 108.950 185.530 ;
        RECT 107.490 185.470 107.770 185.520 ;
        RECT 108.670 185.460 108.950 185.520 ;
        RECT 344.010 185.470 345.490 185.660 ;
        RECT 344.010 185.460 345.480 185.470 ;
        RECT 344.020 185.410 344.300 185.460 ;
        RECT 345.200 185.400 345.480 185.460 ;
        RECT 6.160 185.130 6.430 185.170 ;
        RECT 7.290 185.130 7.580 185.180 ;
        RECT 6.160 184.940 7.580 185.130 ;
        RECT 242.690 185.070 242.960 185.110 ;
        RECT 243.820 185.070 244.110 185.120 ;
        RECT 6.160 184.840 6.430 184.940 ;
        RECT 7.290 184.850 7.580 184.940 ;
        RECT 107.470 184.940 107.740 184.980 ;
        RECT 108.600 184.940 108.890 184.990 ;
        RECT 11.830 184.660 18.290 184.820 ;
        RECT 107.470 184.750 108.890 184.940 ;
        RECT 242.690 184.880 244.110 185.070 ;
        RECT 242.690 184.780 242.960 184.880 ;
        RECT 243.820 184.790 244.110 184.880 ;
        RECT 344.000 184.880 344.270 184.920 ;
        RECT 345.130 184.880 345.420 184.930 ;
        RECT 11.830 184.610 18.300 184.660 ;
        RECT 107.470 184.650 107.740 184.750 ;
        RECT 108.600 184.660 108.890 184.750 ;
        RECT 11.840 183.520 12.040 184.610 ;
        RECT 11.240 183.320 12.040 183.520 ;
        RECT 11.240 182.320 11.440 183.320 ;
        RECT 18.100 183.070 18.300 184.610 ;
        RECT 113.140 184.470 119.600 184.630 ;
        RECT 248.360 184.600 254.820 184.760 ;
        RECT 344.000 184.690 345.420 184.880 ;
        RECT 248.360 184.550 254.830 184.600 ;
        RECT 344.000 184.590 344.270 184.690 ;
        RECT 345.130 184.600 345.420 184.690 ;
        RECT 113.140 184.420 119.610 184.470 ;
        RECT 113.150 183.330 113.350 184.420 ;
        RECT 44.930 183.090 51.390 183.250 ;
        RECT 112.550 183.130 113.350 183.330 ;
        RECT 18.100 182.770 18.390 183.070 ;
        RECT 44.930 183.040 51.400 183.090 ;
        RECT 16.240 182.320 18.940 182.620 ;
        RECT 10.590 182.030 11.440 182.320 ;
        RECT 44.940 181.950 45.140 183.040 ;
        RECT 44.340 181.750 45.140 181.950 ;
        RECT 44.340 180.750 44.540 181.750 ;
        RECT 51.200 181.500 51.400 183.040 ;
        RECT 112.550 182.130 112.750 183.130 ;
        RECT 119.410 182.880 119.610 184.420 ;
        RECT 248.370 183.460 248.570 184.550 ;
        RECT 247.770 183.260 248.570 183.460 ;
        RECT 146.240 182.900 152.700 183.060 ;
        RECT 119.410 182.580 119.700 182.880 ;
        RECT 146.240 182.850 152.710 182.900 ;
        RECT 117.550 182.130 120.250 182.430 ;
        RECT 111.900 181.840 112.750 182.130 ;
        RECT 146.250 181.760 146.450 182.850 ;
        RECT 145.650 181.560 146.450 181.760 ;
        RECT 51.200 181.200 51.490 181.500 ;
        RECT 49.340 180.750 52.040 181.050 ;
        RECT 43.690 180.460 44.540 180.750 ;
        RECT 145.650 180.560 145.850 181.560 ;
        RECT 152.510 181.310 152.710 182.850 ;
        RECT 247.770 182.260 247.970 183.260 ;
        RECT 254.630 183.010 254.830 184.550 ;
        RECT 349.670 184.410 356.130 184.570 ;
        RECT 349.670 184.360 356.140 184.410 ;
        RECT 349.680 183.270 349.880 184.360 ;
        RECT 281.460 183.030 287.920 183.190 ;
        RECT 349.080 183.070 349.880 183.270 ;
        RECT 254.630 182.710 254.920 183.010 ;
        RECT 281.460 182.980 287.930 183.030 ;
        RECT 252.770 182.260 255.470 182.560 ;
        RECT 247.120 181.970 247.970 182.260 ;
        RECT 281.470 181.890 281.670 182.980 ;
        RECT 280.870 181.690 281.670 181.890 ;
        RECT 152.510 181.010 152.800 181.310 ;
        RECT 150.650 180.560 153.350 180.860 ;
        RECT 280.870 180.690 281.070 181.690 ;
        RECT 287.730 181.440 287.930 182.980 ;
        RECT 349.080 182.070 349.280 183.070 ;
        RECT 355.940 182.820 356.140 184.360 ;
        RECT 382.770 182.840 389.230 183.000 ;
        RECT 355.940 182.520 356.230 182.820 ;
        RECT 382.770 182.790 389.240 182.840 ;
        RECT 354.080 182.070 356.780 182.370 ;
        RECT 348.430 181.780 349.280 182.070 ;
        RECT 382.780 181.700 382.980 182.790 ;
        RECT 382.180 181.500 382.980 181.700 ;
        RECT 287.730 181.140 288.020 181.440 ;
        RECT 285.870 180.690 288.570 180.990 ;
        RECT 145.000 180.270 145.850 180.560 ;
        RECT 280.220 180.400 281.070 180.690 ;
        RECT 382.180 180.500 382.380 181.500 ;
        RECT 389.040 181.250 389.240 182.790 ;
        RECT 389.040 180.950 389.330 181.250 ;
        RECT 387.180 180.500 389.880 180.800 ;
        RECT 381.530 180.210 382.380 180.500 ;
        RECT 11.500 176.640 17.960 176.800 ;
        RECT 11.500 176.590 17.970 176.640 ;
        RECT 11.510 175.500 11.710 176.590 ;
        RECT 10.910 175.300 11.710 175.500 ;
        RECT 10.910 174.300 11.110 175.300 ;
        RECT 17.770 175.050 17.970 176.590 ;
        RECT 112.810 176.450 119.270 176.610 ;
        RECT 248.030 176.580 254.490 176.740 ;
        RECT 248.030 176.530 254.500 176.580 ;
        RECT 112.810 176.400 119.280 176.450 ;
        RECT 112.820 175.310 113.020 176.400 ;
        RECT 112.220 175.110 113.020 175.310 ;
        RECT 17.770 174.750 18.060 175.050 ;
        RECT 15.910 174.300 18.610 174.600 ;
        RECT 10.260 174.010 11.110 174.300 ;
        RECT 27.180 174.220 33.640 174.380 ;
        RECT 27.180 174.170 33.650 174.220 ;
        RECT 27.190 173.080 27.390 174.170 ;
        RECT 26.590 172.880 27.390 173.080 ;
        RECT 26.590 171.880 26.790 172.880 ;
        RECT 33.450 172.630 33.650 174.170 ;
        RECT 112.220 174.110 112.420 175.110 ;
        RECT 119.080 174.860 119.280 176.400 ;
        RECT 248.040 175.440 248.240 176.530 ;
        RECT 247.440 175.240 248.240 175.440 ;
        RECT 119.080 174.560 119.370 174.860 ;
        RECT 117.220 174.110 119.920 174.410 ;
        RECT 247.440 174.240 247.640 175.240 ;
        RECT 254.300 174.990 254.500 176.530 ;
        RECT 349.340 176.390 355.800 176.550 ;
        RECT 349.340 176.340 355.810 176.390 ;
        RECT 349.350 175.250 349.550 176.340 ;
        RECT 348.750 175.050 349.550 175.250 ;
        RECT 254.300 174.690 254.590 174.990 ;
        RECT 252.440 174.240 255.140 174.540 ;
        RECT 111.570 173.820 112.420 174.110 ;
        RECT 128.490 174.030 134.950 174.190 ;
        RECT 128.490 173.980 134.960 174.030 ;
        RECT 128.500 172.890 128.700 173.980 ;
        RECT 127.900 172.690 128.700 172.890 ;
        RECT 33.450 172.330 33.740 172.630 ;
        RECT 31.590 171.880 34.290 172.180 ;
        RECT 25.940 171.590 26.790 171.880 ;
        RECT 127.900 171.690 128.100 172.690 ;
        RECT 134.760 172.440 134.960 173.980 ;
        RECT 246.790 173.950 247.640 174.240 ;
        RECT 263.710 174.160 270.170 174.320 ;
        RECT 263.710 174.110 270.180 174.160 ;
        RECT 263.720 173.020 263.920 174.110 ;
        RECT 263.120 172.820 263.920 173.020 ;
        RECT 134.760 172.140 135.050 172.440 ;
        RECT 132.900 171.690 135.600 171.990 ;
        RECT 263.120 171.820 263.320 172.820 ;
        RECT 269.980 172.570 270.180 174.110 ;
        RECT 348.750 174.050 348.950 175.050 ;
        RECT 355.610 174.800 355.810 176.340 ;
        RECT 355.610 174.500 355.900 174.800 ;
        RECT 353.750 174.050 356.450 174.350 ;
        RECT 348.100 173.760 348.950 174.050 ;
        RECT 365.020 173.970 371.480 174.130 ;
        RECT 365.020 173.920 371.490 173.970 ;
        RECT 365.030 172.830 365.230 173.920 ;
        RECT 364.430 172.630 365.230 172.830 ;
        RECT 269.980 172.270 270.270 172.570 ;
        RECT 268.120 171.820 270.820 172.120 ;
        RECT 6.010 171.490 6.290 171.570 ;
        RECT 7.190 171.530 7.470 171.560 ;
        RECT 7.170 171.490 7.480 171.530 ;
        RECT 6.000 171.300 7.480 171.490 ;
        RECT 127.250 171.400 128.100 171.690 ;
        RECT 262.470 171.530 263.320 171.820 ;
        RECT 364.430 171.630 364.630 172.630 ;
        RECT 371.290 172.380 371.490 173.920 ;
        RECT 371.290 172.080 371.580 172.380 ;
        RECT 369.430 171.630 372.130 171.930 ;
        RECT 242.540 171.430 242.820 171.510 ;
        RECT 243.720 171.470 244.000 171.500 ;
        RECT 243.700 171.430 244.010 171.470 ;
        RECT 107.320 171.300 107.600 171.380 ;
        RECT 108.500 171.340 108.780 171.370 ;
        RECT 108.480 171.300 108.790 171.340 ;
        RECT 6.000 171.290 7.470 171.300 ;
        RECT 6.010 171.240 6.290 171.290 ;
        RECT 7.190 171.230 7.470 171.290 ;
        RECT 107.310 171.110 108.790 171.300 ;
        RECT 242.530 171.240 244.010 171.430 ;
        RECT 363.780 171.340 364.630 171.630 ;
        RECT 343.850 171.240 344.130 171.320 ;
        RECT 345.030 171.280 345.310 171.310 ;
        RECT 345.010 171.240 345.320 171.280 ;
        RECT 242.530 171.230 244.000 171.240 ;
        RECT 242.540 171.180 242.820 171.230 ;
        RECT 243.720 171.170 244.000 171.230 ;
        RECT 107.310 171.100 108.780 171.110 ;
        RECT 107.320 171.050 107.600 171.100 ;
        RECT 108.500 171.040 108.780 171.100 ;
        RECT 343.840 171.050 345.320 171.240 ;
        RECT 343.840 171.040 345.310 171.050 ;
        RECT 343.850 170.990 344.130 171.040 ;
        RECT 345.030 170.980 345.310 171.040 ;
        RECT 5.990 170.710 6.260 170.750 ;
        RECT 7.120 170.710 7.410 170.760 ;
        RECT 5.990 170.520 7.410 170.710 ;
        RECT 242.520 170.650 242.790 170.690 ;
        RECT 243.650 170.650 243.940 170.700 ;
        RECT 5.990 170.420 6.260 170.520 ;
        RECT 7.120 170.430 7.410 170.520 ;
        RECT 107.300 170.520 107.570 170.560 ;
        RECT 108.430 170.520 108.720 170.570 ;
        RECT 11.660 170.240 18.120 170.400 ;
        RECT 107.300 170.330 108.720 170.520 ;
        RECT 242.520 170.460 243.940 170.650 ;
        RECT 242.520 170.360 242.790 170.460 ;
        RECT 243.650 170.370 243.940 170.460 ;
        RECT 343.830 170.460 344.100 170.500 ;
        RECT 344.960 170.460 345.250 170.510 ;
        RECT 11.660 170.190 18.130 170.240 ;
        RECT 107.300 170.230 107.570 170.330 ;
        RECT 108.430 170.240 108.720 170.330 ;
        RECT 11.670 169.100 11.870 170.190 ;
        RECT 11.070 168.900 11.870 169.100 ;
        RECT 11.070 167.900 11.270 168.900 ;
        RECT 17.930 168.650 18.130 170.190 ;
        RECT 112.970 170.050 119.430 170.210 ;
        RECT 248.190 170.180 254.650 170.340 ;
        RECT 343.830 170.270 345.250 170.460 ;
        RECT 248.190 170.130 254.660 170.180 ;
        RECT 343.830 170.170 344.100 170.270 ;
        RECT 344.960 170.180 345.250 170.270 ;
        RECT 112.970 170.000 119.440 170.050 ;
        RECT 112.980 168.910 113.180 170.000 ;
        RECT 112.380 168.710 113.180 168.910 ;
        RECT 17.930 168.350 18.220 168.650 ;
        RECT 16.070 167.900 18.770 168.200 ;
        RECT 10.420 167.610 11.270 167.900 ;
        RECT 112.380 167.710 112.580 168.710 ;
        RECT 119.240 168.460 119.440 170.000 ;
        RECT 248.200 169.040 248.400 170.130 ;
        RECT 247.600 168.840 248.400 169.040 ;
        RECT 119.240 168.160 119.530 168.460 ;
        RECT 117.380 167.710 120.080 168.010 ;
        RECT 247.600 167.840 247.800 168.840 ;
        RECT 254.460 168.590 254.660 170.130 ;
        RECT 349.500 169.990 355.960 170.150 ;
        RECT 349.500 169.940 355.970 169.990 ;
        RECT 349.510 168.850 349.710 169.940 ;
        RECT 348.910 168.650 349.710 168.850 ;
        RECT 254.460 168.290 254.750 168.590 ;
        RECT 252.600 167.840 255.300 168.140 ;
        RECT 111.730 167.420 112.580 167.710 ;
        RECT 246.950 167.550 247.800 167.840 ;
        RECT 348.910 167.650 349.110 168.650 ;
        RECT 355.770 168.400 355.970 169.940 ;
        RECT 355.770 168.100 356.060 168.400 ;
        RECT 353.910 167.650 356.610 167.950 ;
        RECT 348.260 167.360 349.110 167.650 ;
        RECT 62.460 167.070 68.920 167.230 ;
        RECT 62.460 167.020 68.930 167.070 ;
        RECT 62.470 165.930 62.670 167.020 ;
        RECT 61.870 165.730 62.670 165.930 ;
        RECT 61.870 164.730 62.070 165.730 ;
        RECT 68.730 165.480 68.930 167.020 ;
        RECT 163.770 166.880 170.230 167.040 ;
        RECT 298.990 167.010 305.450 167.170 ;
        RECT 298.990 166.960 305.460 167.010 ;
        RECT 163.770 166.830 170.240 166.880 ;
        RECT 163.780 165.740 163.980 166.830 ;
        RECT 163.180 165.540 163.980 165.740 ;
        RECT 68.730 165.180 69.020 165.480 ;
        RECT 66.870 164.730 69.570 165.030 ;
        RECT 61.220 164.440 62.070 164.730 ;
        RECT 163.180 164.540 163.380 165.540 ;
        RECT 170.040 165.290 170.240 166.830 ;
        RECT 299.000 165.870 299.200 166.960 ;
        RECT 298.400 165.670 299.200 165.870 ;
        RECT 170.040 164.990 170.330 165.290 ;
        RECT 168.180 164.540 170.880 164.840 ;
        RECT 298.400 164.670 298.600 165.670 ;
        RECT 305.260 165.420 305.460 166.960 ;
        RECT 400.300 166.820 406.760 166.980 ;
        RECT 400.300 166.770 406.770 166.820 ;
        RECT 400.310 165.680 400.510 166.770 ;
        RECT 399.710 165.480 400.510 165.680 ;
        RECT 305.260 165.120 305.550 165.420 ;
        RECT 303.400 164.670 306.100 164.970 ;
        RECT 162.530 164.250 163.380 164.540 ;
        RECT 297.750 164.380 298.600 164.670 ;
        RECT 399.710 164.480 399.910 165.480 ;
        RECT 406.570 165.230 406.770 166.770 ;
        RECT 406.570 164.930 406.860 165.230 ;
        RECT 404.710 164.480 407.410 164.780 ;
        RECT 399.060 164.190 399.910 164.480 ;
        RECT 11.640 160.990 18.100 161.150 ;
        RECT 11.640 160.940 18.110 160.990 ;
        RECT 11.650 159.850 11.850 160.940 ;
        RECT 11.050 159.650 11.850 159.850 ;
        RECT 11.050 158.650 11.250 159.650 ;
        RECT 17.910 159.400 18.110 160.940 ;
        RECT 112.950 160.800 119.410 160.960 ;
        RECT 248.170 160.930 254.630 161.090 ;
        RECT 248.170 160.880 254.640 160.930 ;
        RECT 112.950 160.750 119.420 160.800 ;
        RECT 112.960 159.660 113.160 160.750 ;
        RECT 112.360 159.460 113.160 159.660 ;
        RECT 17.910 159.100 18.200 159.400 ;
        RECT 16.050 158.650 18.750 158.950 ;
        RECT 10.400 158.360 11.250 158.650 ;
        RECT 27.320 158.570 33.780 158.730 ;
        RECT 27.320 158.520 33.790 158.570 ;
        RECT 27.330 157.430 27.530 158.520 ;
        RECT 26.730 157.230 27.530 157.430 ;
        RECT 26.730 156.230 26.930 157.230 ;
        RECT 33.590 156.980 33.790 158.520 ;
        RECT 112.360 158.460 112.560 159.460 ;
        RECT 119.220 159.210 119.420 160.750 ;
        RECT 248.180 159.790 248.380 160.880 ;
        RECT 247.580 159.590 248.380 159.790 ;
        RECT 119.220 158.910 119.510 159.210 ;
        RECT 117.360 158.460 120.060 158.760 ;
        RECT 247.580 158.590 247.780 159.590 ;
        RECT 254.440 159.340 254.640 160.880 ;
        RECT 349.480 160.740 355.940 160.900 ;
        RECT 349.480 160.690 355.950 160.740 ;
        RECT 349.490 159.600 349.690 160.690 ;
        RECT 348.890 159.400 349.690 159.600 ;
        RECT 254.440 159.040 254.730 159.340 ;
        RECT 252.580 158.590 255.280 158.890 ;
        RECT 111.710 158.170 112.560 158.460 ;
        RECT 128.630 158.380 135.090 158.540 ;
        RECT 128.630 158.330 135.100 158.380 ;
        RECT 128.640 157.240 128.840 158.330 ;
        RECT 128.040 157.040 128.840 157.240 ;
        RECT 33.590 156.680 33.880 156.980 ;
        RECT 31.730 156.230 34.430 156.530 ;
        RECT 26.080 155.940 26.930 156.230 ;
        RECT 128.040 156.040 128.240 157.040 ;
        RECT 134.900 156.790 135.100 158.330 ;
        RECT 246.930 158.300 247.780 158.590 ;
        RECT 263.850 158.510 270.310 158.670 ;
        RECT 263.850 158.460 270.320 158.510 ;
        RECT 263.860 157.370 264.060 158.460 ;
        RECT 263.260 157.170 264.060 157.370 ;
        RECT 134.900 156.490 135.190 156.790 ;
        RECT 133.040 156.040 135.740 156.340 ;
        RECT 263.260 156.170 263.460 157.170 ;
        RECT 270.120 156.920 270.320 158.460 ;
        RECT 348.890 158.400 349.090 159.400 ;
        RECT 355.750 159.150 355.950 160.690 ;
        RECT 355.750 158.850 356.040 159.150 ;
        RECT 353.890 158.400 356.590 158.700 ;
        RECT 348.240 158.110 349.090 158.400 ;
        RECT 365.160 158.320 371.620 158.480 ;
        RECT 365.160 158.270 371.630 158.320 ;
        RECT 365.170 157.180 365.370 158.270 ;
        RECT 364.570 156.980 365.370 157.180 ;
        RECT 270.120 156.620 270.410 156.920 ;
        RECT 268.260 156.170 270.960 156.470 ;
        RECT 6.150 155.840 6.430 155.920 ;
        RECT 7.330 155.880 7.610 155.910 ;
        RECT 7.310 155.840 7.620 155.880 ;
        RECT 6.140 155.650 7.620 155.840 ;
        RECT 127.390 155.750 128.240 156.040 ;
        RECT 262.610 155.880 263.460 156.170 ;
        RECT 364.570 155.980 364.770 156.980 ;
        RECT 371.430 156.730 371.630 158.270 ;
        RECT 371.430 156.430 371.720 156.730 ;
        RECT 369.570 155.980 372.270 156.280 ;
        RECT 242.680 155.780 242.960 155.860 ;
        RECT 243.860 155.820 244.140 155.850 ;
        RECT 243.840 155.780 244.150 155.820 ;
        RECT 107.460 155.650 107.740 155.730 ;
        RECT 108.640 155.690 108.920 155.720 ;
        RECT 108.620 155.650 108.930 155.690 ;
        RECT 6.140 155.640 7.610 155.650 ;
        RECT 6.150 155.590 6.430 155.640 ;
        RECT 7.330 155.580 7.610 155.640 ;
        RECT 107.450 155.460 108.930 155.650 ;
        RECT 242.670 155.590 244.150 155.780 ;
        RECT 363.920 155.690 364.770 155.980 ;
        RECT 343.990 155.590 344.270 155.670 ;
        RECT 345.170 155.630 345.450 155.660 ;
        RECT 345.150 155.590 345.460 155.630 ;
        RECT 242.670 155.580 244.140 155.590 ;
        RECT 242.680 155.530 242.960 155.580 ;
        RECT 243.860 155.520 244.140 155.580 ;
        RECT 107.450 155.450 108.920 155.460 ;
        RECT 107.460 155.400 107.740 155.450 ;
        RECT 108.640 155.390 108.920 155.450 ;
        RECT 343.980 155.400 345.460 155.590 ;
        RECT 343.980 155.390 345.450 155.400 ;
        RECT 343.990 155.340 344.270 155.390 ;
        RECT 345.170 155.330 345.450 155.390 ;
        RECT 6.130 155.060 6.400 155.100 ;
        RECT 7.260 155.060 7.550 155.110 ;
        RECT 6.130 154.870 7.550 155.060 ;
        RECT 242.660 155.000 242.930 155.040 ;
        RECT 243.790 155.000 244.080 155.050 ;
        RECT 6.130 154.770 6.400 154.870 ;
        RECT 7.260 154.780 7.550 154.870 ;
        RECT 107.440 154.870 107.710 154.910 ;
        RECT 108.570 154.870 108.860 154.920 ;
        RECT 11.800 154.590 18.260 154.750 ;
        RECT 107.440 154.680 108.860 154.870 ;
        RECT 242.660 154.810 244.080 155.000 ;
        RECT 242.660 154.710 242.930 154.810 ;
        RECT 243.790 154.720 244.080 154.810 ;
        RECT 343.970 154.810 344.240 154.850 ;
        RECT 345.100 154.810 345.390 154.860 ;
        RECT 11.800 154.540 18.270 154.590 ;
        RECT 107.440 154.580 107.710 154.680 ;
        RECT 108.570 154.590 108.860 154.680 ;
        RECT 11.810 153.450 12.010 154.540 ;
        RECT 11.210 153.250 12.010 153.450 ;
        RECT 11.210 152.250 11.410 153.250 ;
        RECT 18.070 153.000 18.270 154.540 ;
        RECT 113.110 154.400 119.570 154.560 ;
        RECT 248.330 154.530 254.790 154.690 ;
        RECT 343.970 154.620 345.390 154.810 ;
        RECT 248.330 154.480 254.800 154.530 ;
        RECT 343.970 154.520 344.240 154.620 ;
        RECT 345.100 154.530 345.390 154.620 ;
        RECT 113.110 154.350 119.580 154.400 ;
        RECT 113.120 153.260 113.320 154.350 ;
        RECT 44.900 153.020 51.360 153.180 ;
        RECT 112.520 153.060 113.320 153.260 ;
        RECT 18.070 152.700 18.360 153.000 ;
        RECT 44.900 152.970 51.370 153.020 ;
        RECT 16.210 152.250 18.910 152.550 ;
        RECT 10.560 151.960 11.410 152.250 ;
        RECT 44.910 151.880 45.110 152.970 ;
        RECT 44.310 151.680 45.110 151.880 ;
        RECT 44.310 150.680 44.510 151.680 ;
        RECT 51.170 151.430 51.370 152.970 ;
        RECT 112.520 152.060 112.720 153.060 ;
        RECT 119.380 152.810 119.580 154.350 ;
        RECT 248.340 153.390 248.540 154.480 ;
        RECT 247.740 153.190 248.540 153.390 ;
        RECT 146.210 152.830 152.670 152.990 ;
        RECT 119.380 152.510 119.670 152.810 ;
        RECT 146.210 152.780 152.680 152.830 ;
        RECT 117.520 152.060 120.220 152.360 ;
        RECT 111.870 151.770 112.720 152.060 ;
        RECT 146.220 151.690 146.420 152.780 ;
        RECT 145.620 151.490 146.420 151.690 ;
        RECT 51.170 151.130 51.460 151.430 ;
        RECT 49.310 150.680 52.010 150.980 ;
        RECT 43.660 150.390 44.510 150.680 ;
        RECT 145.620 150.490 145.820 151.490 ;
        RECT 152.480 151.240 152.680 152.780 ;
        RECT 247.740 152.190 247.940 153.190 ;
        RECT 254.600 152.940 254.800 154.480 ;
        RECT 349.640 154.340 356.100 154.500 ;
        RECT 349.640 154.290 356.110 154.340 ;
        RECT 349.650 153.200 349.850 154.290 ;
        RECT 281.430 152.960 287.890 153.120 ;
        RECT 349.050 153.000 349.850 153.200 ;
        RECT 254.600 152.640 254.890 152.940 ;
        RECT 281.430 152.910 287.900 152.960 ;
        RECT 252.740 152.190 255.440 152.490 ;
        RECT 247.090 151.900 247.940 152.190 ;
        RECT 281.440 151.820 281.640 152.910 ;
        RECT 280.840 151.620 281.640 151.820 ;
        RECT 152.480 150.940 152.770 151.240 ;
        RECT 150.620 150.490 153.320 150.790 ;
        RECT 280.840 150.620 281.040 151.620 ;
        RECT 287.700 151.370 287.900 152.910 ;
        RECT 349.050 152.000 349.250 153.000 ;
        RECT 355.910 152.750 356.110 154.290 ;
        RECT 382.740 152.770 389.200 152.930 ;
        RECT 355.910 152.450 356.200 152.750 ;
        RECT 382.740 152.720 389.210 152.770 ;
        RECT 354.050 152.000 356.750 152.300 ;
        RECT 348.400 151.710 349.250 152.000 ;
        RECT 382.750 151.630 382.950 152.720 ;
        RECT 382.150 151.430 382.950 151.630 ;
        RECT 287.700 151.070 287.990 151.370 ;
        RECT 285.840 150.620 288.540 150.920 ;
        RECT 144.970 150.200 145.820 150.490 ;
        RECT 280.190 150.330 281.040 150.620 ;
        RECT 382.150 150.430 382.350 151.430 ;
        RECT 389.010 151.180 389.210 152.720 ;
        RECT 389.010 150.880 389.300 151.180 ;
        RECT 387.150 150.430 389.850 150.730 ;
        RECT 381.500 150.140 382.350 150.430 ;
        RECT 11.470 146.570 17.930 146.730 ;
        RECT 11.470 146.520 17.940 146.570 ;
        RECT 11.480 145.430 11.680 146.520 ;
        RECT 10.880 145.230 11.680 145.430 ;
        RECT 10.880 144.230 11.080 145.230 ;
        RECT 17.740 144.980 17.940 146.520 ;
        RECT 112.780 146.380 119.240 146.540 ;
        RECT 248.000 146.510 254.460 146.670 ;
        RECT 248.000 146.460 254.470 146.510 ;
        RECT 112.780 146.330 119.250 146.380 ;
        RECT 112.790 145.240 112.990 146.330 ;
        RECT 112.190 145.040 112.990 145.240 ;
        RECT 17.740 144.680 18.030 144.980 ;
        RECT 15.880 144.230 18.580 144.530 ;
        RECT 10.230 143.940 11.080 144.230 ;
        RECT 27.150 144.150 33.610 144.310 ;
        RECT 27.150 144.100 33.620 144.150 ;
        RECT 27.160 143.010 27.360 144.100 ;
        RECT 26.560 142.810 27.360 143.010 ;
        RECT 26.560 141.810 26.760 142.810 ;
        RECT 33.420 142.560 33.620 144.100 ;
        RECT 112.190 144.040 112.390 145.040 ;
        RECT 119.050 144.790 119.250 146.330 ;
        RECT 248.010 145.370 248.210 146.460 ;
        RECT 247.410 145.170 248.210 145.370 ;
        RECT 119.050 144.490 119.340 144.790 ;
        RECT 117.190 144.040 119.890 144.340 ;
        RECT 247.410 144.170 247.610 145.170 ;
        RECT 254.270 144.920 254.470 146.460 ;
        RECT 349.310 146.320 355.770 146.480 ;
        RECT 349.310 146.270 355.780 146.320 ;
        RECT 349.320 145.180 349.520 146.270 ;
        RECT 348.720 144.980 349.520 145.180 ;
        RECT 254.270 144.620 254.560 144.920 ;
        RECT 252.410 144.170 255.110 144.470 ;
        RECT 111.540 143.750 112.390 144.040 ;
        RECT 128.460 143.960 134.920 144.120 ;
        RECT 128.460 143.910 134.930 143.960 ;
        RECT 128.470 142.820 128.670 143.910 ;
        RECT 127.870 142.620 128.670 142.820 ;
        RECT 33.420 142.260 33.710 142.560 ;
        RECT 31.560 141.810 34.260 142.110 ;
        RECT 25.910 141.520 26.760 141.810 ;
        RECT 127.870 141.620 128.070 142.620 ;
        RECT 134.730 142.370 134.930 143.910 ;
        RECT 246.760 143.880 247.610 144.170 ;
        RECT 263.680 144.090 270.140 144.250 ;
        RECT 263.680 144.040 270.150 144.090 ;
        RECT 263.690 142.950 263.890 144.040 ;
        RECT 263.090 142.750 263.890 142.950 ;
        RECT 134.730 142.070 135.020 142.370 ;
        RECT 132.870 141.620 135.570 141.920 ;
        RECT 263.090 141.750 263.290 142.750 ;
        RECT 269.950 142.500 270.150 144.040 ;
        RECT 348.720 143.980 348.920 144.980 ;
        RECT 355.580 144.730 355.780 146.270 ;
        RECT 355.580 144.430 355.870 144.730 ;
        RECT 353.720 143.980 356.420 144.280 ;
        RECT 348.070 143.690 348.920 143.980 ;
        RECT 364.990 143.900 371.450 144.060 ;
        RECT 364.990 143.850 371.460 143.900 ;
        RECT 365.000 142.760 365.200 143.850 ;
        RECT 364.400 142.560 365.200 142.760 ;
        RECT 269.950 142.200 270.240 142.500 ;
        RECT 268.090 141.750 270.790 142.050 ;
        RECT 5.980 141.420 6.260 141.500 ;
        RECT 7.160 141.460 7.440 141.490 ;
        RECT 7.140 141.420 7.450 141.460 ;
        RECT 5.970 141.230 7.450 141.420 ;
        RECT 127.220 141.330 128.070 141.620 ;
        RECT 262.440 141.460 263.290 141.750 ;
        RECT 364.400 141.560 364.600 142.560 ;
        RECT 371.260 142.310 371.460 143.850 ;
        RECT 371.260 142.010 371.550 142.310 ;
        RECT 369.400 141.560 372.100 141.860 ;
        RECT 242.510 141.360 242.790 141.440 ;
        RECT 243.690 141.400 243.970 141.430 ;
        RECT 243.670 141.360 243.980 141.400 ;
        RECT 107.290 141.230 107.570 141.310 ;
        RECT 108.470 141.270 108.750 141.300 ;
        RECT 108.450 141.230 108.760 141.270 ;
        RECT 5.970 141.220 7.440 141.230 ;
        RECT 5.980 141.170 6.260 141.220 ;
        RECT 7.160 141.160 7.440 141.220 ;
        RECT 107.280 141.040 108.760 141.230 ;
        RECT 242.500 141.170 243.980 141.360 ;
        RECT 363.750 141.270 364.600 141.560 ;
        RECT 343.820 141.170 344.100 141.250 ;
        RECT 345.000 141.210 345.280 141.240 ;
        RECT 344.980 141.170 345.290 141.210 ;
        RECT 242.500 141.160 243.970 141.170 ;
        RECT 242.510 141.110 242.790 141.160 ;
        RECT 243.690 141.100 243.970 141.160 ;
        RECT 107.280 141.030 108.750 141.040 ;
        RECT 107.290 140.980 107.570 141.030 ;
        RECT 108.470 140.970 108.750 141.030 ;
        RECT 343.810 140.980 345.290 141.170 ;
        RECT 343.810 140.970 345.280 140.980 ;
        RECT 343.820 140.920 344.100 140.970 ;
        RECT 345.000 140.910 345.280 140.970 ;
        RECT 5.960 140.640 6.230 140.680 ;
        RECT 7.090 140.640 7.380 140.690 ;
        RECT 5.960 140.450 7.380 140.640 ;
        RECT 242.490 140.580 242.760 140.620 ;
        RECT 243.620 140.580 243.910 140.630 ;
        RECT 5.960 140.350 6.230 140.450 ;
        RECT 7.090 140.360 7.380 140.450 ;
        RECT 107.270 140.450 107.540 140.490 ;
        RECT 108.400 140.450 108.690 140.500 ;
        RECT 11.630 140.170 18.090 140.330 ;
        RECT 107.270 140.260 108.690 140.450 ;
        RECT 242.490 140.390 243.910 140.580 ;
        RECT 242.490 140.290 242.760 140.390 ;
        RECT 243.620 140.300 243.910 140.390 ;
        RECT 343.800 140.390 344.070 140.430 ;
        RECT 344.930 140.390 345.220 140.440 ;
        RECT 11.630 140.120 18.100 140.170 ;
        RECT 107.270 140.160 107.540 140.260 ;
        RECT 108.400 140.170 108.690 140.260 ;
        RECT 11.640 139.030 11.840 140.120 ;
        RECT 11.040 138.830 11.840 139.030 ;
        RECT 11.040 137.830 11.240 138.830 ;
        RECT 17.900 138.580 18.100 140.120 ;
        RECT 112.940 139.980 119.400 140.140 ;
        RECT 248.160 140.110 254.620 140.270 ;
        RECT 343.800 140.200 345.220 140.390 ;
        RECT 248.160 140.060 254.630 140.110 ;
        RECT 343.800 140.100 344.070 140.200 ;
        RECT 344.930 140.110 345.220 140.200 ;
        RECT 112.940 139.930 119.410 139.980 ;
        RECT 112.950 138.840 113.150 139.930 ;
        RECT 112.350 138.640 113.150 138.840 ;
        RECT 17.900 138.280 18.190 138.580 ;
        RECT 16.040 137.830 18.740 138.130 ;
        RECT 10.390 137.540 11.240 137.830 ;
        RECT 93.340 137.560 99.800 137.720 ;
        RECT 112.350 137.640 112.550 138.640 ;
        RECT 119.210 138.390 119.410 139.930 ;
        RECT 220.930 139.700 227.390 139.860 ;
        RECT 220.930 139.650 227.400 139.700 ;
        RECT 220.940 138.560 221.140 139.650 ;
        RECT 119.210 138.090 119.500 138.390 ;
        RECT 220.340 138.360 221.140 138.560 ;
        RECT 117.350 137.640 120.050 137.940 ;
        RECT 93.340 137.510 99.810 137.560 ;
        RECT 93.350 136.420 93.550 137.510 ;
        RECT 92.750 136.220 93.550 136.420 ;
        RECT 92.750 135.220 92.950 136.220 ;
        RECT 99.610 135.970 99.810 137.510 ;
        RECT 111.700 137.350 112.550 137.640 ;
        RECT 194.650 137.370 201.110 137.530 ;
        RECT 194.650 137.320 201.120 137.370 ;
        RECT 220.340 137.360 220.540 138.360 ;
        RECT 227.200 138.110 227.400 139.650 ;
        RECT 248.170 138.970 248.370 140.060 ;
        RECT 247.570 138.770 248.370 138.970 ;
        RECT 227.200 137.810 227.490 138.110 ;
        RECT 247.570 137.770 247.770 138.770 ;
        RECT 254.430 138.520 254.630 140.060 ;
        RECT 349.470 139.920 355.930 140.080 ;
        RECT 349.470 139.870 355.940 139.920 ;
        RECT 349.480 138.780 349.680 139.870 ;
        RECT 348.880 138.580 349.680 138.780 ;
        RECT 254.430 138.220 254.720 138.520 ;
        RECT 252.570 137.770 255.270 138.070 ;
        RECT 246.920 137.480 247.770 137.770 ;
        RECT 329.870 137.500 336.330 137.660 ;
        RECT 348.880 137.580 349.080 138.580 ;
        RECT 355.740 138.330 355.940 139.870 ;
        RECT 457.460 139.640 463.920 139.800 ;
        RECT 457.460 139.590 463.930 139.640 ;
        RECT 457.470 138.500 457.670 139.590 ;
        RECT 355.740 138.030 356.030 138.330 ;
        RECT 456.870 138.300 457.670 138.500 ;
        RECT 353.880 137.580 356.580 137.880 ;
        RECT 329.870 137.450 336.340 137.500 ;
        RECT 194.660 136.230 194.860 137.320 ;
        RECT 194.060 136.030 194.860 136.230 ;
        RECT 99.610 135.670 99.900 135.970 ;
        RECT 97.750 135.240 100.520 135.520 ;
        RECT 97.750 135.220 100.450 135.240 ;
        RECT 92.100 134.930 92.950 135.220 ;
        RECT 194.060 135.030 194.260 136.030 ;
        RECT 200.920 135.780 201.120 137.320 ;
        RECT 219.690 137.070 220.540 137.360 ;
        RECT 329.880 136.360 330.080 137.450 ;
        RECT 329.280 136.160 330.080 136.360 ;
        RECT 200.920 135.480 201.210 135.780 ;
        RECT 199.060 135.050 201.830 135.330 ;
        RECT 329.280 135.160 329.480 136.160 ;
        RECT 336.140 135.910 336.340 137.450 ;
        RECT 348.230 137.290 349.080 137.580 ;
        RECT 431.180 137.310 437.640 137.470 ;
        RECT 431.180 137.260 437.650 137.310 ;
        RECT 456.870 137.300 457.070 138.300 ;
        RECT 463.730 138.050 463.930 139.590 ;
        RECT 463.730 137.750 464.020 138.050 ;
        RECT 431.190 136.170 431.390 137.260 ;
        RECT 430.590 135.970 431.390 136.170 ;
        RECT 336.140 135.610 336.430 135.910 ;
        RECT 334.280 135.180 337.050 135.460 ;
        RECT 334.280 135.160 336.980 135.180 ;
        RECT 199.060 135.030 201.760 135.050 ;
        RECT 193.410 134.740 194.260 135.030 ;
        RECT 328.630 134.870 329.480 135.160 ;
        RECT 430.590 134.970 430.790 135.970 ;
        RECT 437.450 135.720 437.650 137.260 ;
        RECT 456.220 137.010 457.070 137.300 ;
        RECT 474.760 137.290 481.220 137.450 ;
        RECT 474.760 137.240 481.230 137.290 ;
        RECT 474.770 136.150 474.970 137.240 ;
        RECT 474.170 135.950 474.970 136.150 ;
        RECT 437.450 135.420 437.740 135.720 ;
        RECT 435.590 134.990 438.360 135.270 ;
        RECT 435.590 134.970 438.290 134.990 ;
        RECT 429.940 134.680 430.790 134.970 ;
        RECT 474.170 134.950 474.370 135.950 ;
        RECT 481.030 135.700 481.230 137.240 ;
        RECT 481.030 135.400 481.320 135.700 ;
        RECT 473.520 134.660 474.370 134.950 ;
        RECT 11.520 130.740 17.980 130.900 ;
        RECT 11.520 130.690 17.990 130.740 ;
        RECT 11.530 129.600 11.730 130.690 ;
        RECT 10.930 129.400 11.730 129.600 ;
        RECT 10.930 128.400 11.130 129.400 ;
        RECT 17.790 129.150 17.990 130.690 ;
        RECT 112.830 130.550 119.290 130.710 ;
        RECT 248.050 130.680 254.510 130.840 ;
        RECT 248.050 130.630 254.520 130.680 ;
        RECT 112.830 130.500 119.300 130.550 ;
        RECT 112.840 129.410 113.040 130.500 ;
        RECT 112.240 129.210 113.040 129.410 ;
        RECT 17.790 128.850 18.080 129.150 ;
        RECT 15.930 128.400 18.630 128.700 ;
        RECT 10.280 128.110 11.130 128.400 ;
        RECT 27.200 128.320 33.660 128.480 ;
        RECT 27.200 128.270 33.670 128.320 ;
        RECT 27.210 127.180 27.410 128.270 ;
        RECT 26.610 126.980 27.410 127.180 ;
        RECT 26.610 125.980 26.810 126.980 ;
        RECT 33.470 126.730 33.670 128.270 ;
        RECT 112.240 128.210 112.440 129.210 ;
        RECT 119.100 128.960 119.300 130.500 ;
        RECT 248.060 129.540 248.260 130.630 ;
        RECT 247.460 129.340 248.260 129.540 ;
        RECT 119.100 128.660 119.390 128.960 ;
        RECT 117.240 128.210 119.940 128.510 ;
        RECT 247.460 128.340 247.660 129.340 ;
        RECT 254.320 129.090 254.520 130.630 ;
        RECT 349.360 130.490 355.820 130.650 ;
        RECT 349.360 130.440 355.830 130.490 ;
        RECT 349.370 129.350 349.570 130.440 ;
        RECT 348.770 129.150 349.570 129.350 ;
        RECT 254.320 128.790 254.610 129.090 ;
        RECT 252.460 128.340 255.160 128.640 ;
        RECT 111.590 127.920 112.440 128.210 ;
        RECT 128.510 128.130 134.970 128.290 ;
        RECT 128.510 128.080 134.980 128.130 ;
        RECT 128.520 126.990 128.720 128.080 ;
        RECT 127.920 126.790 128.720 126.990 ;
        RECT 33.470 126.430 33.760 126.730 ;
        RECT 31.610 125.980 34.310 126.280 ;
        RECT 25.960 125.690 26.810 125.980 ;
        RECT 127.920 125.790 128.120 126.790 ;
        RECT 134.780 126.540 134.980 128.080 ;
        RECT 246.810 128.050 247.660 128.340 ;
        RECT 263.730 128.260 270.190 128.420 ;
        RECT 263.730 128.210 270.200 128.260 ;
        RECT 263.740 127.120 263.940 128.210 ;
        RECT 263.140 126.920 263.940 127.120 ;
        RECT 134.780 126.240 135.070 126.540 ;
        RECT 132.920 125.790 135.620 126.090 ;
        RECT 263.140 125.920 263.340 126.920 ;
        RECT 270.000 126.670 270.200 128.210 ;
        RECT 348.770 128.150 348.970 129.150 ;
        RECT 355.630 128.900 355.830 130.440 ;
        RECT 355.630 128.600 355.920 128.900 ;
        RECT 353.770 128.150 356.470 128.450 ;
        RECT 348.120 127.860 348.970 128.150 ;
        RECT 365.040 128.070 371.500 128.230 ;
        RECT 365.040 128.020 371.510 128.070 ;
        RECT 365.050 126.930 365.250 128.020 ;
        RECT 364.450 126.730 365.250 126.930 ;
        RECT 270.000 126.370 270.290 126.670 ;
        RECT 268.140 125.920 270.840 126.220 ;
        RECT 6.030 125.590 6.310 125.670 ;
        RECT 7.210 125.630 7.490 125.660 ;
        RECT 7.190 125.590 7.500 125.630 ;
        RECT 6.020 125.400 7.500 125.590 ;
        RECT 127.270 125.500 128.120 125.790 ;
        RECT 262.490 125.630 263.340 125.920 ;
        RECT 364.450 125.730 364.650 126.730 ;
        RECT 371.310 126.480 371.510 128.020 ;
        RECT 371.310 126.180 371.600 126.480 ;
        RECT 369.450 125.730 372.150 126.030 ;
        RECT 242.560 125.530 242.840 125.610 ;
        RECT 243.740 125.570 244.020 125.600 ;
        RECT 243.720 125.530 244.030 125.570 ;
        RECT 107.340 125.400 107.620 125.480 ;
        RECT 108.520 125.440 108.800 125.470 ;
        RECT 108.500 125.400 108.810 125.440 ;
        RECT 6.020 125.390 7.490 125.400 ;
        RECT 6.030 125.340 6.310 125.390 ;
        RECT 7.210 125.330 7.490 125.390 ;
        RECT 107.330 125.210 108.810 125.400 ;
        RECT 242.550 125.340 244.030 125.530 ;
        RECT 363.800 125.440 364.650 125.730 ;
        RECT 343.870 125.340 344.150 125.420 ;
        RECT 345.050 125.380 345.330 125.410 ;
        RECT 345.030 125.340 345.340 125.380 ;
        RECT 242.550 125.330 244.020 125.340 ;
        RECT 242.560 125.280 242.840 125.330 ;
        RECT 243.740 125.270 244.020 125.330 ;
        RECT 107.330 125.200 108.800 125.210 ;
        RECT 107.340 125.150 107.620 125.200 ;
        RECT 108.520 125.140 108.800 125.200 ;
        RECT 343.860 125.150 345.340 125.340 ;
        RECT 343.860 125.140 345.330 125.150 ;
        RECT 343.870 125.090 344.150 125.140 ;
        RECT 345.050 125.080 345.330 125.140 ;
        RECT 6.010 124.810 6.280 124.850 ;
        RECT 7.140 124.810 7.430 124.860 ;
        RECT 6.010 124.620 7.430 124.810 ;
        RECT 242.540 124.750 242.810 124.790 ;
        RECT 243.670 124.750 243.960 124.800 ;
        RECT 6.010 124.520 6.280 124.620 ;
        RECT 7.140 124.530 7.430 124.620 ;
        RECT 107.320 124.620 107.590 124.660 ;
        RECT 108.450 124.620 108.740 124.670 ;
        RECT 11.680 124.340 18.140 124.500 ;
        RECT 107.320 124.430 108.740 124.620 ;
        RECT 242.540 124.560 243.960 124.750 ;
        RECT 242.540 124.460 242.810 124.560 ;
        RECT 243.670 124.470 243.960 124.560 ;
        RECT 343.850 124.560 344.120 124.600 ;
        RECT 344.980 124.560 345.270 124.610 ;
        RECT 11.680 124.290 18.150 124.340 ;
        RECT 107.320 124.330 107.590 124.430 ;
        RECT 108.450 124.340 108.740 124.430 ;
        RECT 11.690 123.200 11.890 124.290 ;
        RECT 11.090 123.000 11.890 123.200 ;
        RECT 11.090 122.000 11.290 123.000 ;
        RECT 17.950 122.750 18.150 124.290 ;
        RECT 112.990 124.150 119.450 124.310 ;
        RECT 248.210 124.280 254.670 124.440 ;
        RECT 343.850 124.370 345.270 124.560 ;
        RECT 248.210 124.230 254.680 124.280 ;
        RECT 343.850 124.270 344.120 124.370 ;
        RECT 344.980 124.280 345.270 124.370 ;
        RECT 112.990 124.100 119.460 124.150 ;
        RECT 113.000 123.010 113.200 124.100 ;
        RECT 44.780 122.770 51.240 122.930 ;
        RECT 112.400 122.810 113.200 123.010 ;
        RECT 17.950 122.450 18.240 122.750 ;
        RECT 44.780 122.720 51.250 122.770 ;
        RECT 16.090 122.000 18.790 122.300 ;
        RECT 10.440 121.710 11.290 122.000 ;
        RECT 44.790 121.630 44.990 122.720 ;
        RECT 44.190 121.430 44.990 121.630 ;
        RECT 44.190 120.430 44.390 121.430 ;
        RECT 51.050 121.180 51.250 122.720 ;
        RECT 112.400 121.810 112.600 122.810 ;
        RECT 119.260 122.560 119.460 124.100 ;
        RECT 248.220 123.140 248.420 124.230 ;
        RECT 247.620 122.940 248.420 123.140 ;
        RECT 146.090 122.580 152.550 122.740 ;
        RECT 119.260 122.260 119.550 122.560 ;
        RECT 146.090 122.530 152.560 122.580 ;
        RECT 117.400 121.810 120.100 122.110 ;
        RECT 111.750 121.520 112.600 121.810 ;
        RECT 146.100 121.440 146.300 122.530 ;
        RECT 145.500 121.240 146.300 121.440 ;
        RECT 51.050 120.880 51.340 121.180 ;
        RECT 49.190 120.430 51.890 120.730 ;
        RECT 43.540 120.140 44.390 120.430 ;
        RECT 145.500 120.240 145.700 121.240 ;
        RECT 152.360 120.990 152.560 122.530 ;
        RECT 247.620 121.940 247.820 122.940 ;
        RECT 254.480 122.690 254.680 124.230 ;
        RECT 349.520 124.090 355.980 124.250 ;
        RECT 349.520 124.040 355.990 124.090 ;
        RECT 349.530 122.950 349.730 124.040 ;
        RECT 281.310 122.710 287.770 122.870 ;
        RECT 348.930 122.750 349.730 122.950 ;
        RECT 254.480 122.390 254.770 122.690 ;
        RECT 281.310 122.660 287.780 122.710 ;
        RECT 252.620 121.940 255.320 122.240 ;
        RECT 246.970 121.650 247.820 121.940 ;
        RECT 281.320 121.570 281.520 122.660 ;
        RECT 280.720 121.370 281.520 121.570 ;
        RECT 152.360 120.690 152.650 120.990 ;
        RECT 150.500 120.240 153.200 120.540 ;
        RECT 280.720 120.370 280.920 121.370 ;
        RECT 287.580 121.120 287.780 122.660 ;
        RECT 348.930 121.750 349.130 122.750 ;
        RECT 355.790 122.500 355.990 124.040 ;
        RECT 382.620 122.520 389.080 122.680 ;
        RECT 355.790 122.200 356.080 122.500 ;
        RECT 382.620 122.470 389.090 122.520 ;
        RECT 353.930 121.750 356.630 122.050 ;
        RECT 348.280 121.460 349.130 121.750 ;
        RECT 382.630 121.380 382.830 122.470 ;
        RECT 382.030 121.180 382.830 121.380 ;
        RECT 287.580 120.820 287.870 121.120 ;
        RECT 285.720 120.370 288.420 120.670 ;
        RECT 144.850 119.950 145.700 120.240 ;
        RECT 280.070 120.080 280.920 120.370 ;
        RECT 382.030 120.180 382.230 121.180 ;
        RECT 388.890 120.930 389.090 122.470 ;
        RECT 388.890 120.630 389.180 120.930 ;
        RECT 387.030 120.180 389.730 120.480 ;
        RECT 381.380 119.890 382.230 120.180 ;
        RECT 11.350 116.320 17.810 116.480 ;
        RECT 11.350 116.270 17.820 116.320 ;
        RECT 11.360 115.180 11.560 116.270 ;
        RECT 10.760 114.980 11.560 115.180 ;
        RECT 10.760 113.980 10.960 114.980 ;
        RECT 17.620 114.730 17.820 116.270 ;
        RECT 112.660 116.130 119.120 116.290 ;
        RECT 247.880 116.260 254.340 116.420 ;
        RECT 247.880 116.210 254.350 116.260 ;
        RECT 112.660 116.080 119.130 116.130 ;
        RECT 112.670 114.990 112.870 116.080 ;
        RECT 112.070 114.790 112.870 114.990 ;
        RECT 17.620 114.430 17.910 114.730 ;
        RECT 15.760 113.980 18.460 114.280 ;
        RECT 10.110 113.690 10.960 113.980 ;
        RECT 27.030 113.900 33.490 114.060 ;
        RECT 27.030 113.850 33.500 113.900 ;
        RECT 27.040 112.760 27.240 113.850 ;
        RECT 26.440 112.560 27.240 112.760 ;
        RECT 26.440 111.560 26.640 112.560 ;
        RECT 33.300 112.310 33.500 113.850 ;
        RECT 112.070 113.790 112.270 114.790 ;
        RECT 118.930 114.540 119.130 116.080 ;
        RECT 247.890 115.120 248.090 116.210 ;
        RECT 247.290 114.920 248.090 115.120 ;
        RECT 118.930 114.240 119.220 114.540 ;
        RECT 117.070 113.790 119.770 114.090 ;
        RECT 247.290 113.920 247.490 114.920 ;
        RECT 254.150 114.670 254.350 116.210 ;
        RECT 349.190 116.070 355.650 116.230 ;
        RECT 349.190 116.020 355.660 116.070 ;
        RECT 349.200 114.930 349.400 116.020 ;
        RECT 348.600 114.730 349.400 114.930 ;
        RECT 254.150 114.370 254.440 114.670 ;
        RECT 252.290 113.920 254.990 114.220 ;
        RECT 111.420 113.500 112.270 113.790 ;
        RECT 128.340 113.710 134.800 113.870 ;
        RECT 128.340 113.660 134.810 113.710 ;
        RECT 128.350 112.570 128.550 113.660 ;
        RECT 127.750 112.370 128.550 112.570 ;
        RECT 33.300 112.010 33.590 112.310 ;
        RECT 31.440 111.560 34.140 111.860 ;
        RECT 25.790 111.270 26.640 111.560 ;
        RECT 127.750 111.370 127.950 112.370 ;
        RECT 134.610 112.120 134.810 113.660 ;
        RECT 246.640 113.630 247.490 113.920 ;
        RECT 263.560 113.840 270.020 114.000 ;
        RECT 263.560 113.790 270.030 113.840 ;
        RECT 263.570 112.700 263.770 113.790 ;
        RECT 262.970 112.500 263.770 112.700 ;
        RECT 134.610 111.820 134.900 112.120 ;
        RECT 132.750 111.370 135.450 111.670 ;
        RECT 262.970 111.500 263.170 112.500 ;
        RECT 269.830 112.250 270.030 113.790 ;
        RECT 348.600 113.730 348.800 114.730 ;
        RECT 355.460 114.480 355.660 116.020 ;
        RECT 355.460 114.180 355.750 114.480 ;
        RECT 353.600 113.730 356.300 114.030 ;
        RECT 347.950 113.440 348.800 113.730 ;
        RECT 364.870 113.650 371.330 113.810 ;
        RECT 364.870 113.600 371.340 113.650 ;
        RECT 364.880 112.510 365.080 113.600 ;
        RECT 364.280 112.310 365.080 112.510 ;
        RECT 269.830 111.950 270.120 112.250 ;
        RECT 267.970 111.500 270.670 111.800 ;
        RECT 5.860 111.170 6.140 111.250 ;
        RECT 7.040 111.210 7.320 111.240 ;
        RECT 7.020 111.170 7.330 111.210 ;
        RECT 5.850 110.980 7.330 111.170 ;
        RECT 127.100 111.080 127.950 111.370 ;
        RECT 262.320 111.210 263.170 111.500 ;
        RECT 364.280 111.310 364.480 112.310 ;
        RECT 371.140 112.060 371.340 113.600 ;
        RECT 371.140 111.760 371.430 112.060 ;
        RECT 369.280 111.310 371.980 111.610 ;
        RECT 242.390 111.110 242.670 111.190 ;
        RECT 243.570 111.150 243.850 111.180 ;
        RECT 243.550 111.110 243.860 111.150 ;
        RECT 107.170 110.980 107.450 111.060 ;
        RECT 108.350 111.020 108.630 111.050 ;
        RECT 108.330 110.980 108.640 111.020 ;
        RECT 5.850 110.970 7.320 110.980 ;
        RECT 5.860 110.920 6.140 110.970 ;
        RECT 7.040 110.910 7.320 110.970 ;
        RECT 107.160 110.790 108.640 110.980 ;
        RECT 242.380 110.920 243.860 111.110 ;
        RECT 363.630 111.020 364.480 111.310 ;
        RECT 343.700 110.920 343.980 111.000 ;
        RECT 344.880 110.960 345.160 110.990 ;
        RECT 344.860 110.920 345.170 110.960 ;
        RECT 242.380 110.910 243.850 110.920 ;
        RECT 242.390 110.860 242.670 110.910 ;
        RECT 243.570 110.850 243.850 110.910 ;
        RECT 107.160 110.780 108.630 110.790 ;
        RECT 107.170 110.730 107.450 110.780 ;
        RECT 108.350 110.720 108.630 110.780 ;
        RECT 343.690 110.730 345.170 110.920 ;
        RECT 343.690 110.720 345.160 110.730 ;
        RECT 343.700 110.670 343.980 110.720 ;
        RECT 344.880 110.660 345.160 110.720 ;
        RECT 5.840 110.390 6.110 110.430 ;
        RECT 6.970 110.390 7.260 110.440 ;
        RECT 5.840 110.200 7.260 110.390 ;
        RECT 242.370 110.330 242.640 110.370 ;
        RECT 243.500 110.330 243.790 110.380 ;
        RECT 5.840 110.100 6.110 110.200 ;
        RECT 6.970 110.110 7.260 110.200 ;
        RECT 107.150 110.200 107.420 110.240 ;
        RECT 108.280 110.200 108.570 110.250 ;
        RECT 11.510 109.920 17.970 110.080 ;
        RECT 107.150 110.010 108.570 110.200 ;
        RECT 242.370 110.140 243.790 110.330 ;
        RECT 242.370 110.040 242.640 110.140 ;
        RECT 243.500 110.050 243.790 110.140 ;
        RECT 343.680 110.140 343.950 110.180 ;
        RECT 344.810 110.140 345.100 110.190 ;
        RECT 11.510 109.870 17.980 109.920 ;
        RECT 107.150 109.910 107.420 110.010 ;
        RECT 108.280 109.920 108.570 110.010 ;
        RECT 11.520 108.780 11.720 109.870 ;
        RECT 10.920 108.580 11.720 108.780 ;
        RECT 10.920 107.580 11.120 108.580 ;
        RECT 17.780 108.330 17.980 109.870 ;
        RECT 112.820 109.730 119.280 109.890 ;
        RECT 248.040 109.860 254.500 110.020 ;
        RECT 343.680 109.950 345.100 110.140 ;
        RECT 248.040 109.810 254.510 109.860 ;
        RECT 343.680 109.850 343.950 109.950 ;
        RECT 344.810 109.860 345.100 109.950 ;
        RECT 112.820 109.680 119.290 109.730 ;
        RECT 112.830 108.590 113.030 109.680 ;
        RECT 112.230 108.390 113.030 108.590 ;
        RECT 17.780 108.030 18.070 108.330 ;
        RECT 15.920 107.580 18.620 107.880 ;
        RECT 10.270 107.290 11.120 107.580 ;
        RECT 112.230 107.390 112.430 108.390 ;
        RECT 119.090 108.140 119.290 109.680 ;
        RECT 248.050 108.720 248.250 109.810 ;
        RECT 247.450 108.520 248.250 108.720 ;
        RECT 119.090 107.840 119.380 108.140 ;
        RECT 117.230 107.390 119.930 107.690 ;
        RECT 247.450 107.520 247.650 108.520 ;
        RECT 254.310 108.270 254.510 109.810 ;
        RECT 349.350 109.670 355.810 109.830 ;
        RECT 349.350 109.620 355.820 109.670 ;
        RECT 349.360 108.530 349.560 109.620 ;
        RECT 348.760 108.330 349.560 108.530 ;
        RECT 254.310 107.970 254.600 108.270 ;
        RECT 252.450 107.520 255.150 107.820 ;
        RECT 111.580 107.100 112.430 107.390 ;
        RECT 246.800 107.230 247.650 107.520 ;
        RECT 348.760 107.330 348.960 108.330 ;
        RECT 355.620 108.080 355.820 109.620 ;
        RECT 355.620 107.780 355.910 108.080 ;
        RECT 353.760 107.330 356.460 107.630 ;
        RECT 348.110 107.040 348.960 107.330 ;
        RECT 62.310 106.750 68.770 106.910 ;
        RECT 62.310 106.700 68.780 106.750 ;
        RECT 62.320 105.610 62.520 106.700 ;
        RECT 61.720 105.410 62.520 105.610 ;
        RECT 61.720 104.410 61.920 105.410 ;
        RECT 68.580 105.160 68.780 106.700 ;
        RECT 163.620 106.560 170.080 106.720 ;
        RECT 298.840 106.690 305.300 106.850 ;
        RECT 298.840 106.640 305.310 106.690 ;
        RECT 163.620 106.510 170.090 106.560 ;
        RECT 163.630 105.420 163.830 106.510 ;
        RECT 163.030 105.220 163.830 105.420 ;
        RECT 68.580 104.860 68.870 105.160 ;
        RECT 66.720 104.410 69.420 104.710 ;
        RECT 61.070 104.120 61.920 104.410 ;
        RECT 163.030 104.220 163.230 105.220 ;
        RECT 169.890 104.970 170.090 106.510 ;
        RECT 298.850 105.550 299.050 106.640 ;
        RECT 298.250 105.350 299.050 105.550 ;
        RECT 169.890 104.670 170.180 104.970 ;
        RECT 168.030 104.220 170.730 104.520 ;
        RECT 298.250 104.350 298.450 105.350 ;
        RECT 305.110 105.100 305.310 106.640 ;
        RECT 400.150 106.500 406.610 106.660 ;
        RECT 400.150 106.450 406.620 106.500 ;
        RECT 400.160 105.360 400.360 106.450 ;
        RECT 399.560 105.160 400.360 105.360 ;
        RECT 305.110 104.800 305.400 105.100 ;
        RECT 303.250 104.350 305.950 104.650 ;
        RECT 162.380 103.930 163.230 104.220 ;
        RECT 297.600 104.060 298.450 104.350 ;
        RECT 399.560 104.160 399.760 105.160 ;
        RECT 406.420 104.910 406.620 106.450 ;
        RECT 406.420 104.610 406.710 104.910 ;
        RECT 404.560 104.160 407.260 104.460 ;
        RECT 398.910 103.870 399.760 104.160 ;
        RECT 11.490 100.670 17.950 100.830 ;
        RECT 11.490 100.620 17.960 100.670 ;
        RECT 11.500 99.530 11.700 100.620 ;
        RECT 10.900 99.330 11.700 99.530 ;
        RECT 10.900 98.330 11.100 99.330 ;
        RECT 17.760 99.080 17.960 100.620 ;
        RECT 112.800 100.480 119.260 100.640 ;
        RECT 248.020 100.610 254.480 100.770 ;
        RECT 248.020 100.560 254.490 100.610 ;
        RECT 112.800 100.430 119.270 100.480 ;
        RECT 112.810 99.340 113.010 100.430 ;
        RECT 112.210 99.140 113.010 99.340 ;
        RECT 17.760 98.780 18.050 99.080 ;
        RECT 15.900 98.330 18.600 98.630 ;
        RECT 10.250 98.040 11.100 98.330 ;
        RECT 27.170 98.250 33.630 98.410 ;
        RECT 27.170 98.200 33.640 98.250 ;
        RECT 27.180 97.110 27.380 98.200 ;
        RECT 26.580 96.910 27.380 97.110 ;
        RECT 26.580 95.910 26.780 96.910 ;
        RECT 33.440 96.660 33.640 98.200 ;
        RECT 112.210 98.140 112.410 99.140 ;
        RECT 119.070 98.890 119.270 100.430 ;
        RECT 248.030 99.470 248.230 100.560 ;
        RECT 247.430 99.270 248.230 99.470 ;
        RECT 119.070 98.590 119.360 98.890 ;
        RECT 117.210 98.140 119.910 98.440 ;
        RECT 247.430 98.270 247.630 99.270 ;
        RECT 254.290 99.020 254.490 100.560 ;
        RECT 349.330 100.420 355.790 100.580 ;
        RECT 349.330 100.370 355.800 100.420 ;
        RECT 349.340 99.280 349.540 100.370 ;
        RECT 348.740 99.080 349.540 99.280 ;
        RECT 254.290 98.720 254.580 99.020 ;
        RECT 252.430 98.270 255.130 98.570 ;
        RECT 111.560 97.850 112.410 98.140 ;
        RECT 128.480 98.060 134.940 98.220 ;
        RECT 128.480 98.010 134.950 98.060 ;
        RECT 128.490 96.920 128.690 98.010 ;
        RECT 127.890 96.720 128.690 96.920 ;
        RECT 33.440 96.360 33.730 96.660 ;
        RECT 31.580 95.910 34.280 96.210 ;
        RECT 25.930 95.620 26.780 95.910 ;
        RECT 127.890 95.720 128.090 96.720 ;
        RECT 134.750 96.470 134.950 98.010 ;
        RECT 246.780 97.980 247.630 98.270 ;
        RECT 263.700 98.190 270.160 98.350 ;
        RECT 263.700 98.140 270.170 98.190 ;
        RECT 263.710 97.050 263.910 98.140 ;
        RECT 263.110 96.850 263.910 97.050 ;
        RECT 134.750 96.170 135.040 96.470 ;
        RECT 132.890 95.720 135.590 96.020 ;
        RECT 263.110 95.850 263.310 96.850 ;
        RECT 269.970 96.600 270.170 98.140 ;
        RECT 348.740 98.080 348.940 99.080 ;
        RECT 355.600 98.830 355.800 100.370 ;
        RECT 355.600 98.530 355.890 98.830 ;
        RECT 353.740 98.080 356.440 98.380 ;
        RECT 348.090 97.790 348.940 98.080 ;
        RECT 365.010 98.000 371.470 98.160 ;
        RECT 365.010 97.950 371.480 98.000 ;
        RECT 365.020 96.860 365.220 97.950 ;
        RECT 364.420 96.660 365.220 96.860 ;
        RECT 269.970 96.300 270.260 96.600 ;
        RECT 268.110 95.850 270.810 96.150 ;
        RECT 6.000 95.520 6.280 95.600 ;
        RECT 7.180 95.560 7.460 95.590 ;
        RECT 7.160 95.520 7.470 95.560 ;
        RECT 5.990 95.330 7.470 95.520 ;
        RECT 127.240 95.430 128.090 95.720 ;
        RECT 262.460 95.560 263.310 95.850 ;
        RECT 364.420 95.660 364.620 96.660 ;
        RECT 371.280 96.410 371.480 97.950 ;
        RECT 371.280 96.110 371.570 96.410 ;
        RECT 369.420 95.660 372.120 95.960 ;
        RECT 242.530 95.460 242.810 95.540 ;
        RECT 243.710 95.500 243.990 95.530 ;
        RECT 243.690 95.460 244.000 95.500 ;
        RECT 107.310 95.330 107.590 95.410 ;
        RECT 108.490 95.370 108.770 95.400 ;
        RECT 108.470 95.330 108.780 95.370 ;
        RECT 5.990 95.320 7.460 95.330 ;
        RECT 6.000 95.270 6.280 95.320 ;
        RECT 7.180 95.260 7.460 95.320 ;
        RECT 107.300 95.140 108.780 95.330 ;
        RECT 242.520 95.270 244.000 95.460 ;
        RECT 363.770 95.370 364.620 95.660 ;
        RECT 343.840 95.270 344.120 95.350 ;
        RECT 345.020 95.310 345.300 95.340 ;
        RECT 345.000 95.270 345.310 95.310 ;
        RECT 242.520 95.260 243.990 95.270 ;
        RECT 242.530 95.210 242.810 95.260 ;
        RECT 243.710 95.200 243.990 95.260 ;
        RECT 107.300 95.130 108.770 95.140 ;
        RECT 107.310 95.080 107.590 95.130 ;
        RECT 108.490 95.070 108.770 95.130 ;
        RECT 343.830 95.080 345.310 95.270 ;
        RECT 343.830 95.070 345.300 95.080 ;
        RECT 343.840 95.020 344.120 95.070 ;
        RECT 345.020 95.010 345.300 95.070 ;
        RECT 5.980 94.740 6.250 94.780 ;
        RECT 7.110 94.740 7.400 94.790 ;
        RECT 5.980 94.550 7.400 94.740 ;
        RECT 242.510 94.680 242.780 94.720 ;
        RECT 243.640 94.680 243.930 94.730 ;
        RECT 5.980 94.450 6.250 94.550 ;
        RECT 7.110 94.460 7.400 94.550 ;
        RECT 107.290 94.550 107.560 94.590 ;
        RECT 108.420 94.550 108.710 94.600 ;
        RECT 11.650 94.270 18.110 94.430 ;
        RECT 107.290 94.360 108.710 94.550 ;
        RECT 242.510 94.490 243.930 94.680 ;
        RECT 242.510 94.390 242.780 94.490 ;
        RECT 243.640 94.400 243.930 94.490 ;
        RECT 343.820 94.490 344.090 94.530 ;
        RECT 344.950 94.490 345.240 94.540 ;
        RECT 11.650 94.220 18.120 94.270 ;
        RECT 107.290 94.260 107.560 94.360 ;
        RECT 108.420 94.270 108.710 94.360 ;
        RECT 11.660 93.130 11.860 94.220 ;
        RECT 11.060 92.930 11.860 93.130 ;
        RECT 11.060 91.930 11.260 92.930 ;
        RECT 17.920 92.680 18.120 94.220 ;
        RECT 112.960 94.080 119.420 94.240 ;
        RECT 248.180 94.210 254.640 94.370 ;
        RECT 343.820 94.300 345.240 94.490 ;
        RECT 248.180 94.160 254.650 94.210 ;
        RECT 343.820 94.200 344.090 94.300 ;
        RECT 344.950 94.210 345.240 94.300 ;
        RECT 112.960 94.030 119.430 94.080 ;
        RECT 112.970 92.940 113.170 94.030 ;
        RECT 44.750 92.700 51.210 92.860 ;
        RECT 112.370 92.740 113.170 92.940 ;
        RECT 17.920 92.380 18.210 92.680 ;
        RECT 44.750 92.650 51.220 92.700 ;
        RECT 16.060 91.930 18.760 92.230 ;
        RECT 10.410 91.640 11.260 91.930 ;
        RECT 44.760 91.560 44.960 92.650 ;
        RECT 44.160 91.360 44.960 91.560 ;
        RECT 44.160 90.360 44.360 91.360 ;
        RECT 51.020 91.110 51.220 92.650 ;
        RECT 112.370 91.740 112.570 92.740 ;
        RECT 119.230 92.490 119.430 94.030 ;
        RECT 248.190 93.070 248.390 94.160 ;
        RECT 247.590 92.870 248.390 93.070 ;
        RECT 146.060 92.510 152.520 92.670 ;
        RECT 119.230 92.190 119.520 92.490 ;
        RECT 146.060 92.460 152.530 92.510 ;
        RECT 117.370 91.740 120.070 92.040 ;
        RECT 111.720 91.450 112.570 91.740 ;
        RECT 146.070 91.370 146.270 92.460 ;
        RECT 145.470 91.170 146.270 91.370 ;
        RECT 51.020 90.810 51.310 91.110 ;
        RECT 49.160 90.360 51.860 90.660 ;
        RECT 43.510 90.070 44.360 90.360 ;
        RECT 145.470 90.170 145.670 91.170 ;
        RECT 152.330 90.920 152.530 92.460 ;
        RECT 247.590 91.870 247.790 92.870 ;
        RECT 254.450 92.620 254.650 94.160 ;
        RECT 349.490 94.020 355.950 94.180 ;
        RECT 349.490 93.970 355.960 94.020 ;
        RECT 349.500 92.880 349.700 93.970 ;
        RECT 281.280 92.640 287.740 92.800 ;
        RECT 348.900 92.680 349.700 92.880 ;
        RECT 254.450 92.320 254.740 92.620 ;
        RECT 281.280 92.590 287.750 92.640 ;
        RECT 252.590 91.870 255.290 92.170 ;
        RECT 246.940 91.580 247.790 91.870 ;
        RECT 281.290 91.500 281.490 92.590 ;
        RECT 280.690 91.300 281.490 91.500 ;
        RECT 152.330 90.620 152.620 90.920 ;
        RECT 150.470 90.170 153.170 90.470 ;
        RECT 280.690 90.300 280.890 91.300 ;
        RECT 287.550 91.050 287.750 92.590 ;
        RECT 348.900 91.680 349.100 92.680 ;
        RECT 355.760 92.430 355.960 93.970 ;
        RECT 382.590 92.450 389.050 92.610 ;
        RECT 355.760 92.130 356.050 92.430 ;
        RECT 382.590 92.400 389.060 92.450 ;
        RECT 353.900 91.680 356.600 91.980 ;
        RECT 348.250 91.390 349.100 91.680 ;
        RECT 382.600 91.310 382.800 92.400 ;
        RECT 382.000 91.110 382.800 91.310 ;
        RECT 287.550 90.750 287.840 91.050 ;
        RECT 285.690 90.300 288.390 90.600 ;
        RECT 144.820 89.880 145.670 90.170 ;
        RECT 280.040 90.010 280.890 90.300 ;
        RECT 382.000 90.110 382.200 91.110 ;
        RECT 388.860 90.860 389.060 92.400 ;
        RECT 388.860 90.560 389.150 90.860 ;
        RECT 387.000 90.110 389.700 90.410 ;
        RECT 381.350 89.820 382.200 90.110 ;
        RECT 11.320 86.250 17.780 86.410 ;
        RECT 11.320 86.200 17.790 86.250 ;
        RECT 11.330 85.110 11.530 86.200 ;
        RECT 10.730 84.910 11.530 85.110 ;
        RECT 10.730 83.910 10.930 84.910 ;
        RECT 17.590 84.660 17.790 86.200 ;
        RECT 112.630 86.060 119.090 86.220 ;
        RECT 247.850 86.190 254.310 86.350 ;
        RECT 247.850 86.140 254.320 86.190 ;
        RECT 112.630 86.010 119.100 86.060 ;
        RECT 112.640 84.920 112.840 86.010 ;
        RECT 112.040 84.720 112.840 84.920 ;
        RECT 17.590 84.360 17.880 84.660 ;
        RECT 15.730 83.910 18.430 84.210 ;
        RECT 10.080 83.620 10.930 83.910 ;
        RECT 27.000 83.830 33.460 83.990 ;
        RECT 27.000 83.780 33.470 83.830 ;
        RECT 27.010 82.690 27.210 83.780 ;
        RECT 26.410 82.490 27.210 82.690 ;
        RECT 26.410 81.490 26.610 82.490 ;
        RECT 33.270 82.240 33.470 83.780 ;
        RECT 112.040 83.720 112.240 84.720 ;
        RECT 118.900 84.470 119.100 86.010 ;
        RECT 247.860 85.050 248.060 86.140 ;
        RECT 247.260 84.850 248.060 85.050 ;
        RECT 118.900 84.170 119.190 84.470 ;
        RECT 117.040 83.720 119.740 84.020 ;
        RECT 247.260 83.850 247.460 84.850 ;
        RECT 254.120 84.600 254.320 86.140 ;
        RECT 349.160 86.000 355.620 86.160 ;
        RECT 349.160 85.950 355.630 86.000 ;
        RECT 349.170 84.860 349.370 85.950 ;
        RECT 348.570 84.660 349.370 84.860 ;
        RECT 254.120 84.300 254.410 84.600 ;
        RECT 252.260 83.850 254.960 84.150 ;
        RECT 111.390 83.430 112.240 83.720 ;
        RECT 128.310 83.640 134.770 83.800 ;
        RECT 128.310 83.590 134.780 83.640 ;
        RECT 128.320 82.500 128.520 83.590 ;
        RECT 127.720 82.300 128.520 82.500 ;
        RECT 33.270 81.940 33.560 82.240 ;
        RECT 31.410 81.490 34.110 81.790 ;
        RECT 25.760 81.200 26.610 81.490 ;
        RECT 127.720 81.300 127.920 82.300 ;
        RECT 134.580 82.050 134.780 83.590 ;
        RECT 246.610 83.560 247.460 83.850 ;
        RECT 263.530 83.770 269.990 83.930 ;
        RECT 263.530 83.720 270.000 83.770 ;
        RECT 263.540 82.630 263.740 83.720 ;
        RECT 262.940 82.430 263.740 82.630 ;
        RECT 134.580 81.750 134.870 82.050 ;
        RECT 132.720 81.300 135.420 81.600 ;
        RECT 262.940 81.430 263.140 82.430 ;
        RECT 269.800 82.180 270.000 83.720 ;
        RECT 348.570 83.660 348.770 84.660 ;
        RECT 355.430 84.410 355.630 85.950 ;
        RECT 355.430 84.110 355.720 84.410 ;
        RECT 353.570 83.660 356.270 83.960 ;
        RECT 347.920 83.370 348.770 83.660 ;
        RECT 364.840 83.580 371.300 83.740 ;
        RECT 364.840 83.530 371.310 83.580 ;
        RECT 364.850 82.440 365.050 83.530 ;
        RECT 364.250 82.240 365.050 82.440 ;
        RECT 269.800 81.880 270.090 82.180 ;
        RECT 267.940 81.430 270.640 81.730 ;
        RECT 5.830 81.100 6.110 81.180 ;
        RECT 7.010 81.140 7.290 81.170 ;
        RECT 6.990 81.100 7.300 81.140 ;
        RECT 5.820 80.910 7.300 81.100 ;
        RECT 127.070 81.010 127.920 81.300 ;
        RECT 262.290 81.140 263.140 81.430 ;
        RECT 364.250 81.240 364.450 82.240 ;
        RECT 371.110 81.990 371.310 83.530 ;
        RECT 371.110 81.690 371.400 81.990 ;
        RECT 369.250 81.240 371.950 81.540 ;
        RECT 242.360 81.040 242.640 81.120 ;
        RECT 243.540 81.080 243.820 81.110 ;
        RECT 243.520 81.040 243.830 81.080 ;
        RECT 107.140 80.910 107.420 80.990 ;
        RECT 108.320 80.950 108.600 80.980 ;
        RECT 108.300 80.910 108.610 80.950 ;
        RECT 5.820 80.900 7.290 80.910 ;
        RECT 5.830 80.850 6.110 80.900 ;
        RECT 7.010 80.840 7.290 80.900 ;
        RECT 107.130 80.720 108.610 80.910 ;
        RECT 242.350 80.850 243.830 81.040 ;
        RECT 363.600 80.950 364.450 81.240 ;
        RECT 343.670 80.850 343.950 80.930 ;
        RECT 344.850 80.890 345.130 80.920 ;
        RECT 344.830 80.850 345.140 80.890 ;
        RECT 242.350 80.840 243.820 80.850 ;
        RECT 242.360 80.790 242.640 80.840 ;
        RECT 243.540 80.780 243.820 80.840 ;
        RECT 107.130 80.710 108.600 80.720 ;
        RECT 107.140 80.660 107.420 80.710 ;
        RECT 108.320 80.650 108.600 80.710 ;
        RECT 343.660 80.660 345.140 80.850 ;
        RECT 343.660 80.650 345.130 80.660 ;
        RECT 76.510 80.460 82.970 80.620 ;
        RECT 343.670 80.600 343.950 80.650 ;
        RECT 344.850 80.590 345.130 80.650 ;
        RECT 76.510 80.410 82.980 80.460 ;
        RECT 5.810 80.320 6.080 80.360 ;
        RECT 6.940 80.320 7.230 80.370 ;
        RECT 5.810 80.130 7.230 80.320 ;
        RECT 5.810 80.030 6.080 80.130 ;
        RECT 6.940 80.040 7.230 80.130 ;
        RECT 11.480 79.850 17.940 80.010 ;
        RECT 11.480 79.800 17.950 79.850 ;
        RECT 11.490 78.710 11.690 79.800 ;
        RECT 10.890 78.510 11.690 78.710 ;
        RECT 10.890 77.510 11.090 78.510 ;
        RECT 17.750 78.260 17.950 79.800 ;
        RECT 76.520 79.320 76.720 80.410 ;
        RECT 75.920 79.120 76.720 79.320 ;
        RECT 17.750 77.960 18.040 78.260 ;
        RECT 75.920 78.120 76.120 79.120 ;
        RECT 82.780 78.870 82.980 80.410 ;
        RECT 177.820 80.270 184.280 80.430 ;
        RECT 313.040 80.400 319.500 80.560 ;
        RECT 313.040 80.350 319.510 80.400 ;
        RECT 177.820 80.220 184.290 80.270 ;
        RECT 107.120 80.130 107.390 80.170 ;
        RECT 108.250 80.130 108.540 80.180 ;
        RECT 107.120 79.940 108.540 80.130 ;
        RECT 107.120 79.840 107.390 79.940 ;
        RECT 108.250 79.850 108.540 79.940 ;
        RECT 112.790 79.660 119.250 79.820 ;
        RECT 112.790 79.610 119.260 79.660 ;
        RECT 82.780 78.570 83.070 78.870 ;
        RECT 112.800 78.520 113.000 79.610 ;
        RECT 80.920 78.370 83.620 78.420 ;
        RECT 80.920 78.140 83.670 78.370 ;
        RECT 112.200 78.320 113.000 78.520 ;
        RECT 80.920 78.120 83.620 78.140 ;
        RECT 75.270 77.830 76.120 78.120 ;
        RECT 15.890 77.510 18.590 77.810 ;
        RECT 10.240 77.220 11.090 77.510 ;
        RECT 112.200 77.320 112.400 78.320 ;
        RECT 119.060 78.070 119.260 79.610 ;
        RECT 177.830 79.130 178.030 80.220 ;
        RECT 177.230 78.930 178.030 79.130 ;
        RECT 119.060 77.770 119.350 78.070 ;
        RECT 177.230 77.930 177.430 78.930 ;
        RECT 184.090 78.680 184.290 80.220 ;
        RECT 242.340 80.260 242.610 80.300 ;
        RECT 243.470 80.260 243.760 80.310 ;
        RECT 242.340 80.070 243.760 80.260 ;
        RECT 242.340 79.970 242.610 80.070 ;
        RECT 243.470 79.980 243.760 80.070 ;
        RECT 248.010 79.790 254.470 79.950 ;
        RECT 248.010 79.740 254.480 79.790 ;
        RECT 184.090 78.380 184.380 78.680 ;
        RECT 248.020 78.650 248.220 79.740 ;
        RECT 247.420 78.450 248.220 78.650 ;
        RECT 182.230 78.180 184.930 78.230 ;
        RECT 182.230 77.950 184.980 78.180 ;
        RECT 182.230 77.930 184.930 77.950 ;
        RECT 176.580 77.640 177.430 77.930 ;
        RECT 117.200 77.320 119.900 77.620 ;
        RECT 247.420 77.450 247.620 78.450 ;
        RECT 254.280 78.200 254.480 79.740 ;
        RECT 313.050 79.260 313.250 80.350 ;
        RECT 312.450 79.060 313.250 79.260 ;
        RECT 254.280 77.900 254.570 78.200 ;
        RECT 312.450 78.060 312.650 79.060 ;
        RECT 319.310 78.810 319.510 80.350 ;
        RECT 414.350 80.210 420.810 80.370 ;
        RECT 414.350 80.160 420.820 80.210 ;
        RECT 343.650 80.070 343.920 80.110 ;
        RECT 344.780 80.070 345.070 80.120 ;
        RECT 343.650 79.880 345.070 80.070 ;
        RECT 343.650 79.780 343.920 79.880 ;
        RECT 344.780 79.790 345.070 79.880 ;
        RECT 349.320 79.600 355.780 79.760 ;
        RECT 349.320 79.550 355.790 79.600 ;
        RECT 319.310 78.510 319.600 78.810 ;
        RECT 349.330 78.460 349.530 79.550 ;
        RECT 317.450 78.310 320.150 78.360 ;
        RECT 317.450 78.080 320.200 78.310 ;
        RECT 348.730 78.260 349.530 78.460 ;
        RECT 317.450 78.060 320.150 78.080 ;
        RECT 311.800 77.770 312.650 78.060 ;
        RECT 252.420 77.450 255.120 77.750 ;
        RECT 111.550 77.030 112.400 77.320 ;
        RECT 246.770 77.160 247.620 77.450 ;
        RECT 348.730 77.260 348.930 78.260 ;
        RECT 355.590 78.010 355.790 79.550 ;
        RECT 414.360 79.070 414.560 80.160 ;
        RECT 413.760 78.870 414.560 79.070 ;
        RECT 355.590 77.710 355.880 78.010 ;
        RECT 413.760 77.870 413.960 78.870 ;
        RECT 420.620 78.620 420.820 80.160 ;
        RECT 420.620 78.320 420.910 78.620 ;
        RECT 418.760 78.120 421.460 78.170 ;
        RECT 418.760 77.890 421.510 78.120 ;
        RECT 418.760 77.870 421.460 77.890 ;
        RECT 413.110 77.580 413.960 77.870 ;
        RECT 353.730 77.260 356.430 77.560 ;
        RECT 348.080 76.970 348.930 77.260 ;
        RECT 11.170 70.820 17.630 70.980 ;
        RECT 11.170 70.770 17.640 70.820 ;
        RECT 11.180 69.680 11.380 70.770 ;
        RECT 10.580 69.480 11.380 69.680 ;
        RECT 10.580 68.480 10.780 69.480 ;
        RECT 17.440 69.230 17.640 70.770 ;
        RECT 112.480 70.630 118.940 70.790 ;
        RECT 247.700 70.760 254.160 70.920 ;
        RECT 247.700 70.710 254.170 70.760 ;
        RECT 112.480 70.580 118.950 70.630 ;
        RECT 112.490 69.490 112.690 70.580 ;
        RECT 111.890 69.290 112.690 69.490 ;
        RECT 17.440 68.930 17.730 69.230 ;
        RECT 15.580 68.480 18.280 68.780 ;
        RECT 9.930 68.190 10.780 68.480 ;
        RECT 26.850 68.400 33.310 68.560 ;
        RECT 26.850 68.350 33.320 68.400 ;
        RECT 26.860 67.260 27.060 68.350 ;
        RECT 26.260 67.060 27.060 67.260 ;
        RECT 26.260 66.060 26.460 67.060 ;
        RECT 33.120 66.810 33.320 68.350 ;
        RECT 111.890 68.290 112.090 69.290 ;
        RECT 118.750 69.040 118.950 70.580 ;
        RECT 247.710 69.620 247.910 70.710 ;
        RECT 247.110 69.420 247.910 69.620 ;
        RECT 118.750 68.740 119.040 69.040 ;
        RECT 116.890 68.290 119.590 68.590 ;
        RECT 247.110 68.420 247.310 69.420 ;
        RECT 253.970 69.170 254.170 70.710 ;
        RECT 349.010 70.570 355.470 70.730 ;
        RECT 349.010 70.520 355.480 70.570 ;
        RECT 349.020 69.430 349.220 70.520 ;
        RECT 348.420 69.230 349.220 69.430 ;
        RECT 253.970 68.870 254.260 69.170 ;
        RECT 252.110 68.420 254.810 68.720 ;
        RECT 111.240 68.000 112.090 68.290 ;
        RECT 128.160 68.210 134.620 68.370 ;
        RECT 128.160 68.160 134.630 68.210 ;
        RECT 128.170 67.070 128.370 68.160 ;
        RECT 127.570 66.870 128.370 67.070 ;
        RECT 33.120 66.510 33.410 66.810 ;
        RECT 31.260 66.060 33.960 66.360 ;
        RECT 25.610 65.770 26.460 66.060 ;
        RECT 127.570 65.870 127.770 66.870 ;
        RECT 134.430 66.620 134.630 68.160 ;
        RECT 246.460 68.130 247.310 68.420 ;
        RECT 263.380 68.340 269.840 68.500 ;
        RECT 263.380 68.290 269.850 68.340 ;
        RECT 263.390 67.200 263.590 68.290 ;
        RECT 262.790 67.000 263.590 67.200 ;
        RECT 134.430 66.320 134.720 66.620 ;
        RECT 132.570 65.870 135.270 66.170 ;
        RECT 262.790 66.000 262.990 67.000 ;
        RECT 269.650 66.750 269.850 68.290 ;
        RECT 348.420 68.230 348.620 69.230 ;
        RECT 355.280 68.980 355.480 70.520 ;
        RECT 355.280 68.680 355.570 68.980 ;
        RECT 353.420 68.230 356.120 68.530 ;
        RECT 347.770 67.940 348.620 68.230 ;
        RECT 364.690 68.150 371.150 68.310 ;
        RECT 364.690 68.100 371.160 68.150 ;
        RECT 364.700 67.010 364.900 68.100 ;
        RECT 364.100 66.810 364.900 67.010 ;
        RECT 269.650 66.450 269.940 66.750 ;
        RECT 267.790 66.000 270.490 66.300 ;
        RECT 5.680 65.670 5.960 65.750 ;
        RECT 6.860 65.710 7.140 65.740 ;
        RECT 6.840 65.670 7.150 65.710 ;
        RECT 5.670 65.480 7.150 65.670 ;
        RECT 126.920 65.580 127.770 65.870 ;
        RECT 262.140 65.710 262.990 66.000 ;
        RECT 364.100 65.810 364.300 66.810 ;
        RECT 370.960 66.560 371.160 68.100 ;
        RECT 370.960 66.260 371.250 66.560 ;
        RECT 369.100 65.810 371.800 66.110 ;
        RECT 242.210 65.610 242.490 65.690 ;
        RECT 243.390 65.650 243.670 65.680 ;
        RECT 243.370 65.610 243.680 65.650 ;
        RECT 106.990 65.480 107.270 65.560 ;
        RECT 108.170 65.520 108.450 65.550 ;
        RECT 108.150 65.480 108.460 65.520 ;
        RECT 5.670 65.470 7.140 65.480 ;
        RECT 5.680 65.420 5.960 65.470 ;
        RECT 6.860 65.410 7.140 65.470 ;
        RECT 106.980 65.290 108.460 65.480 ;
        RECT 242.200 65.420 243.680 65.610 ;
        RECT 363.450 65.520 364.300 65.810 ;
        RECT 343.520 65.420 343.800 65.500 ;
        RECT 344.700 65.460 344.980 65.490 ;
        RECT 344.680 65.420 344.990 65.460 ;
        RECT 242.200 65.410 243.670 65.420 ;
        RECT 242.210 65.360 242.490 65.410 ;
        RECT 243.390 65.350 243.670 65.410 ;
        RECT 106.980 65.280 108.450 65.290 ;
        RECT 106.990 65.230 107.270 65.280 ;
        RECT 108.170 65.220 108.450 65.280 ;
        RECT 343.510 65.230 344.990 65.420 ;
        RECT 343.510 65.220 344.980 65.230 ;
        RECT 343.520 65.170 343.800 65.220 ;
        RECT 344.700 65.160 344.980 65.220 ;
        RECT 5.660 64.890 5.930 64.930 ;
        RECT 6.790 64.890 7.080 64.940 ;
        RECT 5.660 64.700 7.080 64.890 ;
        RECT 242.190 64.830 242.460 64.870 ;
        RECT 243.320 64.830 243.610 64.880 ;
        RECT 5.660 64.600 5.930 64.700 ;
        RECT 6.790 64.610 7.080 64.700 ;
        RECT 106.970 64.700 107.240 64.740 ;
        RECT 108.100 64.700 108.390 64.750 ;
        RECT 11.330 64.420 17.790 64.580 ;
        RECT 106.970 64.510 108.390 64.700 ;
        RECT 242.190 64.640 243.610 64.830 ;
        RECT 242.190 64.540 242.460 64.640 ;
        RECT 243.320 64.550 243.610 64.640 ;
        RECT 343.500 64.640 343.770 64.680 ;
        RECT 344.630 64.640 344.920 64.690 ;
        RECT 11.330 64.370 17.800 64.420 ;
        RECT 106.970 64.410 107.240 64.510 ;
        RECT 108.100 64.420 108.390 64.510 ;
        RECT 11.340 63.280 11.540 64.370 ;
        RECT 10.740 63.080 11.540 63.280 ;
        RECT 10.740 62.080 10.940 63.080 ;
        RECT 17.600 62.830 17.800 64.370 ;
        RECT 112.640 64.230 119.100 64.390 ;
        RECT 247.860 64.360 254.320 64.520 ;
        RECT 343.500 64.450 344.920 64.640 ;
        RECT 247.860 64.310 254.330 64.360 ;
        RECT 343.500 64.350 343.770 64.450 ;
        RECT 344.630 64.360 344.920 64.450 ;
        RECT 112.640 64.180 119.110 64.230 ;
        RECT 112.650 63.090 112.850 64.180 ;
        RECT 44.430 62.850 50.890 63.010 ;
        RECT 112.050 62.890 112.850 63.090 ;
        RECT 17.600 62.530 17.890 62.830 ;
        RECT 44.430 62.800 50.900 62.850 ;
        RECT 15.740 62.080 18.440 62.380 ;
        RECT 10.090 61.790 10.940 62.080 ;
        RECT 44.440 61.710 44.640 62.800 ;
        RECT 43.840 61.510 44.640 61.710 ;
        RECT 43.840 60.510 44.040 61.510 ;
        RECT 50.700 61.260 50.900 62.800 ;
        RECT 112.050 61.890 112.250 62.890 ;
        RECT 118.910 62.640 119.110 64.180 ;
        RECT 247.870 63.220 248.070 64.310 ;
        RECT 247.270 63.020 248.070 63.220 ;
        RECT 145.740 62.660 152.200 62.820 ;
        RECT 118.910 62.340 119.200 62.640 ;
        RECT 145.740 62.610 152.210 62.660 ;
        RECT 117.050 61.890 119.750 62.190 ;
        RECT 111.400 61.600 112.250 61.890 ;
        RECT 145.750 61.520 145.950 62.610 ;
        RECT 145.150 61.320 145.950 61.520 ;
        RECT 50.700 60.960 50.990 61.260 ;
        RECT 48.840 60.510 51.540 60.810 ;
        RECT 43.190 60.220 44.040 60.510 ;
        RECT 145.150 60.320 145.350 61.320 ;
        RECT 152.010 61.070 152.210 62.610 ;
        RECT 247.270 62.020 247.470 63.020 ;
        RECT 254.130 62.770 254.330 64.310 ;
        RECT 349.170 64.170 355.630 64.330 ;
        RECT 349.170 64.120 355.640 64.170 ;
        RECT 349.180 63.030 349.380 64.120 ;
        RECT 280.960 62.790 287.420 62.950 ;
        RECT 348.580 62.830 349.380 63.030 ;
        RECT 254.130 62.470 254.420 62.770 ;
        RECT 280.960 62.740 287.430 62.790 ;
        RECT 252.270 62.020 254.970 62.320 ;
        RECT 246.620 61.730 247.470 62.020 ;
        RECT 280.970 61.650 281.170 62.740 ;
        RECT 280.370 61.450 281.170 61.650 ;
        RECT 152.010 60.770 152.300 61.070 ;
        RECT 150.150 60.320 152.850 60.620 ;
        RECT 280.370 60.450 280.570 61.450 ;
        RECT 287.230 61.200 287.430 62.740 ;
        RECT 348.580 61.830 348.780 62.830 ;
        RECT 355.440 62.580 355.640 64.120 ;
        RECT 382.270 62.600 388.730 62.760 ;
        RECT 355.440 62.280 355.730 62.580 ;
        RECT 382.270 62.550 388.740 62.600 ;
        RECT 353.580 61.830 356.280 62.130 ;
        RECT 347.930 61.540 348.780 61.830 ;
        RECT 382.280 61.460 382.480 62.550 ;
        RECT 381.680 61.260 382.480 61.460 ;
        RECT 287.230 60.900 287.520 61.200 ;
        RECT 285.370 60.450 288.070 60.750 ;
        RECT 144.500 60.030 145.350 60.320 ;
        RECT 279.720 60.160 280.570 60.450 ;
        RECT 381.680 60.260 381.880 61.260 ;
        RECT 388.540 61.010 388.740 62.550 ;
        RECT 388.540 60.710 388.830 61.010 ;
        RECT 386.680 60.260 389.380 60.560 ;
        RECT 381.030 59.970 381.880 60.260 ;
        RECT 11.000 56.400 17.460 56.560 ;
        RECT 11.000 56.350 17.470 56.400 ;
        RECT 11.010 55.260 11.210 56.350 ;
        RECT 10.410 55.060 11.210 55.260 ;
        RECT 10.410 54.060 10.610 55.060 ;
        RECT 17.270 54.810 17.470 56.350 ;
        RECT 112.310 56.210 118.770 56.370 ;
        RECT 247.530 56.340 253.990 56.500 ;
        RECT 247.530 56.290 254.000 56.340 ;
        RECT 112.310 56.160 118.780 56.210 ;
        RECT 112.320 55.070 112.520 56.160 ;
        RECT 111.720 54.870 112.520 55.070 ;
        RECT 17.270 54.510 17.560 54.810 ;
        RECT 15.410 54.060 18.110 54.360 ;
        RECT 9.760 53.770 10.610 54.060 ;
        RECT 26.680 53.980 33.140 54.140 ;
        RECT 26.680 53.930 33.150 53.980 ;
        RECT 26.690 52.840 26.890 53.930 ;
        RECT 26.090 52.640 26.890 52.840 ;
        RECT 26.090 51.640 26.290 52.640 ;
        RECT 32.950 52.390 33.150 53.930 ;
        RECT 111.720 53.870 111.920 54.870 ;
        RECT 118.580 54.620 118.780 56.160 ;
        RECT 247.540 55.200 247.740 56.290 ;
        RECT 246.940 55.000 247.740 55.200 ;
        RECT 118.580 54.320 118.870 54.620 ;
        RECT 116.720 53.870 119.420 54.170 ;
        RECT 246.940 54.000 247.140 55.000 ;
        RECT 253.800 54.750 254.000 56.290 ;
        RECT 348.840 56.150 355.300 56.310 ;
        RECT 348.840 56.100 355.310 56.150 ;
        RECT 348.850 55.010 349.050 56.100 ;
        RECT 348.250 54.810 349.050 55.010 ;
        RECT 253.800 54.450 254.090 54.750 ;
        RECT 251.940 54.000 254.640 54.300 ;
        RECT 111.070 53.580 111.920 53.870 ;
        RECT 127.990 53.790 134.450 53.950 ;
        RECT 127.990 53.740 134.460 53.790 ;
        RECT 128.000 52.650 128.200 53.740 ;
        RECT 127.400 52.450 128.200 52.650 ;
        RECT 32.950 52.090 33.240 52.390 ;
        RECT 31.090 51.640 33.790 51.940 ;
        RECT 25.440 51.350 26.290 51.640 ;
        RECT 127.400 51.450 127.600 52.450 ;
        RECT 134.260 52.200 134.460 53.740 ;
        RECT 246.290 53.710 247.140 54.000 ;
        RECT 263.210 53.920 269.670 54.080 ;
        RECT 263.210 53.870 269.680 53.920 ;
        RECT 263.220 52.780 263.420 53.870 ;
        RECT 262.620 52.580 263.420 52.780 ;
        RECT 134.260 51.900 134.550 52.200 ;
        RECT 132.400 51.450 135.100 51.750 ;
        RECT 262.620 51.580 262.820 52.580 ;
        RECT 269.480 52.330 269.680 53.870 ;
        RECT 348.250 53.810 348.450 54.810 ;
        RECT 355.110 54.560 355.310 56.100 ;
        RECT 355.110 54.260 355.400 54.560 ;
        RECT 353.250 53.810 355.950 54.110 ;
        RECT 347.600 53.520 348.450 53.810 ;
        RECT 364.520 53.730 370.980 53.890 ;
        RECT 364.520 53.680 370.990 53.730 ;
        RECT 364.530 52.590 364.730 53.680 ;
        RECT 363.930 52.390 364.730 52.590 ;
        RECT 269.480 52.030 269.770 52.330 ;
        RECT 267.620 51.580 270.320 51.880 ;
        RECT 5.510 51.250 5.790 51.330 ;
        RECT 6.690 51.290 6.970 51.320 ;
        RECT 6.670 51.250 6.980 51.290 ;
        RECT 5.500 51.060 6.980 51.250 ;
        RECT 126.750 51.160 127.600 51.450 ;
        RECT 261.970 51.290 262.820 51.580 ;
        RECT 363.930 51.390 364.130 52.390 ;
        RECT 370.790 52.140 370.990 53.680 ;
        RECT 370.790 51.840 371.080 52.140 ;
        RECT 368.930 51.390 371.630 51.690 ;
        RECT 242.040 51.190 242.320 51.270 ;
        RECT 243.220 51.230 243.500 51.260 ;
        RECT 243.200 51.190 243.510 51.230 ;
        RECT 106.820 51.060 107.100 51.140 ;
        RECT 108.000 51.100 108.280 51.130 ;
        RECT 107.980 51.060 108.290 51.100 ;
        RECT 5.500 51.050 6.970 51.060 ;
        RECT 5.510 51.000 5.790 51.050 ;
        RECT 6.690 50.990 6.970 51.050 ;
        RECT 106.810 50.870 108.290 51.060 ;
        RECT 242.030 51.000 243.510 51.190 ;
        RECT 363.280 51.100 364.130 51.390 ;
        RECT 343.350 51.000 343.630 51.080 ;
        RECT 344.530 51.040 344.810 51.070 ;
        RECT 344.510 51.000 344.820 51.040 ;
        RECT 242.030 50.990 243.500 51.000 ;
        RECT 242.040 50.940 242.320 50.990 ;
        RECT 243.220 50.930 243.500 50.990 ;
        RECT 106.810 50.860 108.280 50.870 ;
        RECT 106.820 50.810 107.100 50.860 ;
        RECT 108.000 50.800 108.280 50.860 ;
        RECT 343.340 50.810 344.820 51.000 ;
        RECT 343.340 50.800 344.810 50.810 ;
        RECT 343.350 50.750 343.630 50.800 ;
        RECT 344.530 50.740 344.810 50.800 ;
        RECT 5.490 50.470 5.760 50.510 ;
        RECT 6.620 50.470 6.910 50.520 ;
        RECT 5.490 50.280 6.910 50.470 ;
        RECT 242.020 50.410 242.290 50.450 ;
        RECT 243.150 50.410 243.440 50.460 ;
        RECT 5.490 50.180 5.760 50.280 ;
        RECT 6.620 50.190 6.910 50.280 ;
        RECT 106.800 50.280 107.070 50.320 ;
        RECT 107.930 50.280 108.220 50.330 ;
        RECT 11.160 50.000 17.620 50.160 ;
        RECT 106.800 50.090 108.220 50.280 ;
        RECT 242.020 50.220 243.440 50.410 ;
        RECT 242.020 50.120 242.290 50.220 ;
        RECT 243.150 50.130 243.440 50.220 ;
        RECT 343.330 50.220 343.600 50.260 ;
        RECT 344.460 50.220 344.750 50.270 ;
        RECT 11.160 49.950 17.630 50.000 ;
        RECT 106.800 49.990 107.070 50.090 ;
        RECT 107.930 50.000 108.220 50.090 ;
        RECT 11.170 48.860 11.370 49.950 ;
        RECT 10.570 48.660 11.370 48.860 ;
        RECT 10.570 47.660 10.770 48.660 ;
        RECT 17.430 48.410 17.630 49.950 ;
        RECT 112.470 49.810 118.930 49.970 ;
        RECT 247.690 49.940 254.150 50.100 ;
        RECT 343.330 50.030 344.750 50.220 ;
        RECT 247.690 49.890 254.160 49.940 ;
        RECT 343.330 49.930 343.600 50.030 ;
        RECT 344.460 49.940 344.750 50.030 ;
        RECT 112.470 49.760 118.940 49.810 ;
        RECT 112.480 48.670 112.680 49.760 ;
        RECT 111.880 48.470 112.680 48.670 ;
        RECT 17.430 48.110 17.720 48.410 ;
        RECT 15.570 47.660 18.270 47.960 ;
        RECT 9.920 47.370 10.770 47.660 ;
        RECT 111.880 47.470 112.080 48.470 ;
        RECT 118.740 48.220 118.940 49.760 ;
        RECT 247.700 48.800 247.900 49.890 ;
        RECT 247.100 48.600 247.900 48.800 ;
        RECT 118.740 47.920 119.030 48.220 ;
        RECT 116.880 47.470 119.580 47.770 ;
        RECT 247.100 47.600 247.300 48.600 ;
        RECT 253.960 48.350 254.160 49.890 ;
        RECT 349.000 49.750 355.460 49.910 ;
        RECT 349.000 49.700 355.470 49.750 ;
        RECT 349.010 48.610 349.210 49.700 ;
        RECT 348.410 48.410 349.210 48.610 ;
        RECT 253.960 48.050 254.250 48.350 ;
        RECT 252.100 47.600 254.800 47.900 ;
        RECT 111.230 47.180 112.080 47.470 ;
        RECT 246.450 47.310 247.300 47.600 ;
        RECT 348.410 47.410 348.610 48.410 ;
        RECT 355.270 48.160 355.470 49.700 ;
        RECT 355.270 47.860 355.560 48.160 ;
        RECT 353.410 47.410 356.110 47.710 ;
        RECT 347.760 47.120 348.610 47.410 ;
        RECT 61.960 46.830 68.420 46.990 ;
        RECT 61.960 46.780 68.430 46.830 ;
        RECT 61.970 45.690 62.170 46.780 ;
        RECT 61.370 45.490 62.170 45.690 ;
        RECT 61.370 44.490 61.570 45.490 ;
        RECT 68.230 45.240 68.430 46.780 ;
        RECT 163.270 46.640 169.730 46.800 ;
        RECT 298.490 46.770 304.950 46.930 ;
        RECT 298.490 46.720 304.960 46.770 ;
        RECT 163.270 46.590 169.740 46.640 ;
        RECT 163.280 45.500 163.480 46.590 ;
        RECT 162.680 45.300 163.480 45.500 ;
        RECT 68.230 44.940 68.520 45.240 ;
        RECT 66.370 44.490 69.070 44.790 ;
        RECT 60.720 44.200 61.570 44.490 ;
        RECT 162.680 44.300 162.880 45.300 ;
        RECT 169.540 45.050 169.740 46.590 ;
        RECT 298.500 45.630 298.700 46.720 ;
        RECT 297.900 45.430 298.700 45.630 ;
        RECT 169.540 44.750 169.830 45.050 ;
        RECT 167.680 44.300 170.380 44.600 ;
        RECT 297.900 44.430 298.100 45.430 ;
        RECT 304.760 45.180 304.960 46.720 ;
        RECT 399.800 46.580 406.260 46.740 ;
        RECT 399.800 46.530 406.270 46.580 ;
        RECT 399.810 45.440 400.010 46.530 ;
        RECT 399.210 45.240 400.010 45.440 ;
        RECT 304.760 44.880 305.050 45.180 ;
        RECT 302.900 44.430 305.600 44.730 ;
        RECT 162.030 44.010 162.880 44.300 ;
        RECT 297.250 44.140 298.100 44.430 ;
        RECT 399.210 44.240 399.410 45.240 ;
        RECT 406.070 44.990 406.270 46.530 ;
        RECT 406.070 44.690 406.360 44.990 ;
        RECT 404.210 44.240 406.910 44.540 ;
        RECT 398.560 43.950 399.410 44.240 ;
        RECT 11.140 40.750 17.600 40.910 ;
        RECT 11.140 40.700 17.610 40.750 ;
        RECT 11.150 39.610 11.350 40.700 ;
        RECT 10.550 39.410 11.350 39.610 ;
        RECT 10.550 38.410 10.750 39.410 ;
        RECT 17.410 39.160 17.610 40.700 ;
        RECT 112.450 40.560 118.910 40.720 ;
        RECT 247.670 40.690 254.130 40.850 ;
        RECT 247.670 40.640 254.140 40.690 ;
        RECT 112.450 40.510 118.920 40.560 ;
        RECT 112.460 39.420 112.660 40.510 ;
        RECT 111.860 39.220 112.660 39.420 ;
        RECT 17.410 38.860 17.700 39.160 ;
        RECT 15.550 38.410 18.250 38.710 ;
        RECT 9.900 38.120 10.750 38.410 ;
        RECT 26.820 38.330 33.280 38.490 ;
        RECT 26.820 38.280 33.290 38.330 ;
        RECT 26.830 37.190 27.030 38.280 ;
        RECT 26.230 36.990 27.030 37.190 ;
        RECT 26.230 35.990 26.430 36.990 ;
        RECT 33.090 36.740 33.290 38.280 ;
        RECT 111.860 38.220 112.060 39.220 ;
        RECT 118.720 38.970 118.920 40.510 ;
        RECT 247.680 39.550 247.880 40.640 ;
        RECT 247.080 39.350 247.880 39.550 ;
        RECT 118.720 38.670 119.010 38.970 ;
        RECT 116.860 38.220 119.560 38.520 ;
        RECT 247.080 38.350 247.280 39.350 ;
        RECT 253.940 39.100 254.140 40.640 ;
        RECT 348.980 40.500 355.440 40.660 ;
        RECT 348.980 40.450 355.450 40.500 ;
        RECT 348.990 39.360 349.190 40.450 ;
        RECT 348.390 39.160 349.190 39.360 ;
        RECT 253.940 38.800 254.230 39.100 ;
        RECT 252.080 38.350 254.780 38.650 ;
        RECT 111.210 37.930 112.060 38.220 ;
        RECT 128.130 38.140 134.590 38.300 ;
        RECT 128.130 38.090 134.600 38.140 ;
        RECT 128.140 37.000 128.340 38.090 ;
        RECT 127.540 36.800 128.340 37.000 ;
        RECT 33.090 36.440 33.380 36.740 ;
        RECT 31.230 35.990 33.930 36.290 ;
        RECT 25.580 35.700 26.430 35.990 ;
        RECT 127.540 35.800 127.740 36.800 ;
        RECT 134.400 36.550 134.600 38.090 ;
        RECT 246.430 38.060 247.280 38.350 ;
        RECT 263.350 38.270 269.810 38.430 ;
        RECT 263.350 38.220 269.820 38.270 ;
        RECT 263.360 37.130 263.560 38.220 ;
        RECT 262.760 36.930 263.560 37.130 ;
        RECT 134.400 36.250 134.690 36.550 ;
        RECT 132.540 35.800 135.240 36.100 ;
        RECT 262.760 35.930 262.960 36.930 ;
        RECT 269.620 36.680 269.820 38.220 ;
        RECT 348.390 38.160 348.590 39.160 ;
        RECT 355.250 38.910 355.450 40.450 ;
        RECT 355.250 38.610 355.540 38.910 ;
        RECT 353.390 38.160 356.090 38.460 ;
        RECT 347.740 37.870 348.590 38.160 ;
        RECT 364.660 38.080 371.120 38.240 ;
        RECT 364.660 38.030 371.130 38.080 ;
        RECT 364.670 36.940 364.870 38.030 ;
        RECT 364.070 36.740 364.870 36.940 ;
        RECT 269.620 36.380 269.910 36.680 ;
        RECT 267.760 35.930 270.460 36.230 ;
        RECT 5.650 35.600 5.930 35.680 ;
        RECT 6.830 35.640 7.110 35.670 ;
        RECT 6.810 35.600 7.120 35.640 ;
        RECT 5.640 35.410 7.120 35.600 ;
        RECT 126.890 35.510 127.740 35.800 ;
        RECT 262.110 35.640 262.960 35.930 ;
        RECT 364.070 35.740 364.270 36.740 ;
        RECT 370.930 36.490 371.130 38.030 ;
        RECT 370.930 36.190 371.220 36.490 ;
        RECT 369.070 35.740 371.770 36.040 ;
        RECT 242.180 35.540 242.460 35.620 ;
        RECT 243.360 35.580 243.640 35.610 ;
        RECT 243.340 35.540 243.650 35.580 ;
        RECT 106.960 35.410 107.240 35.490 ;
        RECT 108.140 35.450 108.420 35.480 ;
        RECT 108.120 35.410 108.430 35.450 ;
        RECT 5.640 35.400 7.110 35.410 ;
        RECT 5.650 35.350 5.930 35.400 ;
        RECT 6.830 35.340 7.110 35.400 ;
        RECT 106.950 35.220 108.430 35.410 ;
        RECT 242.170 35.350 243.650 35.540 ;
        RECT 363.420 35.450 364.270 35.740 ;
        RECT 343.490 35.350 343.770 35.430 ;
        RECT 344.670 35.390 344.950 35.420 ;
        RECT 344.650 35.350 344.960 35.390 ;
        RECT 242.170 35.340 243.640 35.350 ;
        RECT 242.180 35.290 242.460 35.340 ;
        RECT 243.360 35.280 243.640 35.340 ;
        RECT 106.950 35.210 108.420 35.220 ;
        RECT 106.960 35.160 107.240 35.210 ;
        RECT 108.140 35.150 108.420 35.210 ;
        RECT 343.480 35.160 344.960 35.350 ;
        RECT 343.480 35.150 344.950 35.160 ;
        RECT 343.490 35.100 343.770 35.150 ;
        RECT 344.670 35.090 344.950 35.150 ;
        RECT 5.630 34.820 5.900 34.860 ;
        RECT 6.760 34.820 7.050 34.870 ;
        RECT 5.630 34.630 7.050 34.820 ;
        RECT 242.160 34.760 242.430 34.800 ;
        RECT 243.290 34.760 243.580 34.810 ;
        RECT 5.630 34.530 5.900 34.630 ;
        RECT 6.760 34.540 7.050 34.630 ;
        RECT 106.940 34.630 107.210 34.670 ;
        RECT 108.070 34.630 108.360 34.680 ;
        RECT 11.300 34.350 17.760 34.510 ;
        RECT 106.940 34.440 108.360 34.630 ;
        RECT 242.160 34.570 243.580 34.760 ;
        RECT 242.160 34.470 242.430 34.570 ;
        RECT 243.290 34.480 243.580 34.570 ;
        RECT 343.470 34.570 343.740 34.610 ;
        RECT 344.600 34.570 344.890 34.620 ;
        RECT 11.300 34.300 17.770 34.350 ;
        RECT 106.940 34.340 107.210 34.440 ;
        RECT 108.070 34.350 108.360 34.440 ;
        RECT 11.310 33.210 11.510 34.300 ;
        RECT 10.710 33.010 11.510 33.210 ;
        RECT 10.710 32.010 10.910 33.010 ;
        RECT 17.570 32.760 17.770 34.300 ;
        RECT 112.610 34.160 119.070 34.320 ;
        RECT 247.830 34.290 254.290 34.450 ;
        RECT 343.470 34.380 344.890 34.570 ;
        RECT 247.830 34.240 254.300 34.290 ;
        RECT 343.470 34.280 343.740 34.380 ;
        RECT 344.600 34.290 344.890 34.380 ;
        RECT 112.610 34.110 119.080 34.160 ;
        RECT 112.620 33.020 112.820 34.110 ;
        RECT 44.400 32.780 50.860 32.940 ;
        RECT 112.020 32.820 112.820 33.020 ;
        RECT 17.570 32.460 17.860 32.760 ;
        RECT 44.400 32.730 50.870 32.780 ;
        RECT 15.710 32.010 18.410 32.310 ;
        RECT 10.060 31.720 10.910 32.010 ;
        RECT 44.410 31.640 44.610 32.730 ;
        RECT 43.810 31.440 44.610 31.640 ;
        RECT 43.810 30.440 44.010 31.440 ;
        RECT 50.670 31.190 50.870 32.730 ;
        RECT 112.020 31.820 112.220 32.820 ;
        RECT 118.880 32.570 119.080 34.110 ;
        RECT 247.840 33.150 248.040 34.240 ;
        RECT 247.240 32.950 248.040 33.150 ;
        RECT 145.710 32.590 152.170 32.750 ;
        RECT 118.880 32.270 119.170 32.570 ;
        RECT 145.710 32.540 152.180 32.590 ;
        RECT 117.020 31.820 119.720 32.120 ;
        RECT 111.370 31.530 112.220 31.820 ;
        RECT 145.720 31.450 145.920 32.540 ;
        RECT 145.120 31.250 145.920 31.450 ;
        RECT 50.670 30.890 50.960 31.190 ;
        RECT 48.810 30.440 51.510 30.740 ;
        RECT 43.160 30.150 44.010 30.440 ;
        RECT 145.120 30.250 145.320 31.250 ;
        RECT 151.980 31.000 152.180 32.540 ;
        RECT 247.240 31.950 247.440 32.950 ;
        RECT 254.100 32.700 254.300 34.240 ;
        RECT 349.140 34.100 355.600 34.260 ;
        RECT 349.140 34.050 355.610 34.100 ;
        RECT 349.150 32.960 349.350 34.050 ;
        RECT 280.930 32.720 287.390 32.880 ;
        RECT 348.550 32.760 349.350 32.960 ;
        RECT 254.100 32.400 254.390 32.700 ;
        RECT 280.930 32.670 287.400 32.720 ;
        RECT 252.240 31.950 254.940 32.250 ;
        RECT 246.590 31.660 247.440 31.950 ;
        RECT 280.940 31.580 281.140 32.670 ;
        RECT 280.340 31.380 281.140 31.580 ;
        RECT 151.980 30.700 152.270 31.000 ;
        RECT 150.120 30.250 152.820 30.550 ;
        RECT 280.340 30.380 280.540 31.380 ;
        RECT 287.200 31.130 287.400 32.670 ;
        RECT 348.550 31.760 348.750 32.760 ;
        RECT 355.410 32.510 355.610 34.050 ;
        RECT 382.240 32.530 388.700 32.690 ;
        RECT 355.410 32.210 355.700 32.510 ;
        RECT 382.240 32.480 388.710 32.530 ;
        RECT 353.550 31.760 356.250 32.060 ;
        RECT 347.900 31.470 348.750 31.760 ;
        RECT 382.250 31.390 382.450 32.480 ;
        RECT 381.650 31.190 382.450 31.390 ;
        RECT 287.200 30.830 287.490 31.130 ;
        RECT 285.340 30.380 288.040 30.680 ;
        RECT 144.470 29.960 145.320 30.250 ;
        RECT 279.690 30.090 280.540 30.380 ;
        RECT 381.650 30.190 381.850 31.190 ;
        RECT 388.510 30.940 388.710 32.480 ;
        RECT 388.510 30.640 388.800 30.940 ;
        RECT 386.650 30.190 389.350 30.490 ;
        RECT 381.000 29.900 381.850 30.190 ;
        RECT 10.970 26.330 17.430 26.490 ;
        RECT 10.970 26.280 17.440 26.330 ;
        RECT 10.980 25.190 11.180 26.280 ;
        RECT 10.380 24.990 11.180 25.190 ;
        RECT 10.380 23.990 10.580 24.990 ;
        RECT 17.240 24.740 17.440 26.280 ;
        RECT 112.280 26.140 118.740 26.300 ;
        RECT 247.500 26.270 253.960 26.430 ;
        RECT 247.500 26.220 253.970 26.270 ;
        RECT 112.280 26.090 118.750 26.140 ;
        RECT 112.290 25.000 112.490 26.090 ;
        RECT 111.690 24.800 112.490 25.000 ;
        RECT 17.240 24.440 17.530 24.740 ;
        RECT 15.380 23.990 18.080 24.290 ;
        RECT 9.730 23.700 10.580 23.990 ;
        RECT 26.650 23.910 33.110 24.070 ;
        RECT 26.650 23.860 33.120 23.910 ;
        RECT 26.660 22.770 26.860 23.860 ;
        RECT 26.060 22.570 26.860 22.770 ;
        RECT 26.060 21.570 26.260 22.570 ;
        RECT 32.920 22.320 33.120 23.860 ;
        RECT 111.690 23.800 111.890 24.800 ;
        RECT 118.550 24.550 118.750 26.090 ;
        RECT 247.510 25.130 247.710 26.220 ;
        RECT 246.910 24.930 247.710 25.130 ;
        RECT 118.550 24.250 118.840 24.550 ;
        RECT 116.690 23.800 119.390 24.100 ;
        RECT 246.910 23.930 247.110 24.930 ;
        RECT 253.770 24.680 253.970 26.220 ;
        RECT 348.810 26.080 355.270 26.240 ;
        RECT 348.810 26.030 355.280 26.080 ;
        RECT 348.820 24.940 349.020 26.030 ;
        RECT 348.220 24.740 349.020 24.940 ;
        RECT 253.770 24.380 254.060 24.680 ;
        RECT 251.910 23.930 254.610 24.230 ;
        RECT 111.040 23.510 111.890 23.800 ;
        RECT 127.960 23.720 134.420 23.880 ;
        RECT 127.960 23.670 134.430 23.720 ;
        RECT 127.970 22.580 128.170 23.670 ;
        RECT 127.370 22.380 128.170 22.580 ;
        RECT 32.920 22.020 33.210 22.320 ;
        RECT 31.060 21.570 33.760 21.870 ;
        RECT 25.410 21.280 26.260 21.570 ;
        RECT 127.370 21.380 127.570 22.380 ;
        RECT 134.230 22.130 134.430 23.670 ;
        RECT 246.260 23.640 247.110 23.930 ;
        RECT 263.180 23.850 269.640 24.010 ;
        RECT 263.180 23.800 269.650 23.850 ;
        RECT 263.190 22.710 263.390 23.800 ;
        RECT 262.590 22.510 263.390 22.710 ;
        RECT 134.230 21.830 134.520 22.130 ;
        RECT 132.370 21.380 135.070 21.680 ;
        RECT 262.590 21.510 262.790 22.510 ;
        RECT 269.450 22.260 269.650 23.800 ;
        RECT 348.220 23.740 348.420 24.740 ;
        RECT 355.080 24.490 355.280 26.030 ;
        RECT 355.080 24.190 355.370 24.490 ;
        RECT 353.220 23.740 355.920 24.040 ;
        RECT 347.570 23.450 348.420 23.740 ;
        RECT 364.490 23.660 370.950 23.820 ;
        RECT 364.490 23.610 370.960 23.660 ;
        RECT 364.500 22.520 364.700 23.610 ;
        RECT 363.900 22.320 364.700 22.520 ;
        RECT 269.450 21.960 269.740 22.260 ;
        RECT 267.590 21.510 270.290 21.810 ;
        RECT 5.480 21.180 5.760 21.260 ;
        RECT 6.660 21.220 6.940 21.250 ;
        RECT 6.640 21.180 6.950 21.220 ;
        RECT 5.470 20.990 6.950 21.180 ;
        RECT 126.720 21.090 127.570 21.380 ;
        RECT 261.940 21.220 262.790 21.510 ;
        RECT 363.900 21.320 364.100 22.320 ;
        RECT 370.760 22.070 370.960 23.610 ;
        RECT 370.760 21.770 371.050 22.070 ;
        RECT 368.900 21.320 371.600 21.620 ;
        RECT 242.010 21.120 242.290 21.200 ;
        RECT 243.190 21.160 243.470 21.190 ;
        RECT 243.170 21.120 243.480 21.160 ;
        RECT 106.790 20.990 107.070 21.070 ;
        RECT 107.970 21.030 108.250 21.060 ;
        RECT 107.950 20.990 108.260 21.030 ;
        RECT 5.470 20.980 6.940 20.990 ;
        RECT 5.480 20.930 5.760 20.980 ;
        RECT 6.660 20.920 6.940 20.980 ;
        RECT 106.780 20.800 108.260 20.990 ;
        RECT 242.000 20.930 243.480 21.120 ;
        RECT 363.250 21.030 364.100 21.320 ;
        RECT 343.320 20.930 343.600 21.010 ;
        RECT 344.500 20.970 344.780 21.000 ;
        RECT 344.480 20.930 344.790 20.970 ;
        RECT 242.000 20.920 243.470 20.930 ;
        RECT 242.010 20.870 242.290 20.920 ;
        RECT 243.190 20.860 243.470 20.920 ;
        RECT 106.780 20.790 108.250 20.800 ;
        RECT 106.790 20.740 107.070 20.790 ;
        RECT 107.970 20.730 108.250 20.790 ;
        RECT 343.310 20.740 344.790 20.930 ;
        RECT 343.310 20.730 344.780 20.740 ;
        RECT 343.320 20.680 343.600 20.730 ;
        RECT 344.500 20.670 344.780 20.730 ;
        RECT 5.460 20.400 5.730 20.440 ;
        RECT 6.590 20.400 6.880 20.450 ;
        RECT 5.460 20.210 6.880 20.400 ;
        RECT 241.990 20.340 242.260 20.380 ;
        RECT 243.120 20.340 243.410 20.390 ;
        RECT 5.460 20.110 5.730 20.210 ;
        RECT 6.590 20.120 6.880 20.210 ;
        RECT 106.770 20.210 107.040 20.250 ;
        RECT 107.900 20.210 108.190 20.260 ;
        RECT 11.130 19.930 17.590 20.090 ;
        RECT 106.770 20.020 108.190 20.210 ;
        RECT 241.990 20.150 243.410 20.340 ;
        RECT 241.990 20.050 242.260 20.150 ;
        RECT 243.120 20.060 243.410 20.150 ;
        RECT 343.300 20.150 343.570 20.190 ;
        RECT 344.430 20.150 344.720 20.200 ;
        RECT 11.130 19.880 17.600 19.930 ;
        RECT 106.770 19.920 107.040 20.020 ;
        RECT 107.900 19.930 108.190 20.020 ;
        RECT 11.140 18.790 11.340 19.880 ;
        RECT 10.540 18.590 11.340 18.790 ;
        RECT 10.540 17.590 10.740 18.590 ;
        RECT 17.400 18.340 17.600 19.880 ;
        RECT 112.440 19.740 118.900 19.900 ;
        RECT 247.660 19.870 254.120 20.030 ;
        RECT 343.300 19.960 344.720 20.150 ;
        RECT 247.660 19.820 254.130 19.870 ;
        RECT 343.300 19.860 343.570 19.960 ;
        RECT 344.430 19.870 344.720 19.960 ;
        RECT 112.440 19.690 118.910 19.740 ;
        RECT 112.450 18.600 112.650 19.690 ;
        RECT 111.850 18.400 112.650 18.600 ;
        RECT 17.400 18.040 17.690 18.340 ;
        RECT 15.540 17.590 18.240 17.890 ;
        RECT 9.890 17.300 10.740 17.590 ;
        RECT 111.850 17.400 112.050 18.400 ;
        RECT 118.710 18.150 118.910 19.690 ;
        RECT 247.670 18.730 247.870 19.820 ;
        RECT 247.070 18.530 247.870 18.730 ;
        RECT 118.710 17.850 119.000 18.150 ;
        RECT 116.850 17.400 119.550 17.700 ;
        RECT 247.070 17.530 247.270 18.530 ;
        RECT 253.930 18.280 254.130 19.820 ;
        RECT 348.970 19.680 355.430 19.840 ;
        RECT 348.970 19.630 355.440 19.680 ;
        RECT 348.980 18.540 349.180 19.630 ;
        RECT 348.380 18.340 349.180 18.540 ;
        RECT 253.930 17.980 254.220 18.280 ;
        RECT 252.070 17.530 254.770 17.830 ;
        RECT 111.200 17.110 112.050 17.400 ;
        RECT 246.420 17.240 247.270 17.530 ;
        RECT 348.380 17.340 348.580 18.340 ;
        RECT 355.240 18.090 355.440 19.630 ;
        RECT 355.240 17.790 355.530 18.090 ;
        RECT 353.380 17.340 356.080 17.640 ;
        RECT 347.730 17.050 348.580 17.340 ;
  END
END 8bitdac_layout
END LIBRARY

