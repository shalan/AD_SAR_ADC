VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC_8BIT
  CLASS BLOCK ;
  FOREIGN DAC_8BIT ;
  ORIGIN 0.000 0.000 ;
  SIZE 499.220 BY 320.560 ;
  PIN d0
    PORT
      LAYER li1 ;
        RECT 106.460 19.395 106.760 25.600 ;
    END
    PORT
      LAYER met2 ;
        RECT 106.710 0.000 107.290 4.000 ;
    END
  END d0
  PIN d1
    PORT
      LAYER li1 ;
        RECT 121.850 19.960 122.150 26.270 ;
    END
    PORT
      LAYER met2 ;
        RECT 124.095 0.000 124.675 4.000 ;
    END
  END d1
  PIN d2
    PORT
      LAYER li1 ;
        RECT 138.550 20.880 138.850 27.510 ;
    END
    PORT
      LAYER met2 ;
        RECT 139.380 0.000 139.960 10.345 ;
    END
  END d2
  PIN d3
    PORT
      LAYER li1 ;
        RECT 155.520 21.790 155.820 28.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 157.775 0.000 158.355 10.345 ;
    END
  END d3
  PIN d4
    PORT
      LAYER li1 ;
        RECT 171.730 23.100 172.030 30.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 175.845 0.000 176.425 10.340 ;
    END
  END d4
  PIN d5
    PORT
      LAYER li1 ;
        RECT 189.040 23.410 189.340 48.150 ;
    END
    PORT
      LAYER met2 ;
        RECT 193.520 0.000 194.100 10.340 ;
    END
  END d5
  PIN d6
    PORT
      LAYER li1 ;
        RECT 215.460 24.380 215.790 31.770 ;
    END
    PORT
      LAYER met2 ;
        RECT 220.960 0.000 221.540 10.345 ;
    END
  END d6
  PIN x2_out_v
    PORT
      LAYER li1 ;
        RECT 480.860 155.910 481.070 158.160 ;
    END
  END x2_out_v
  PIN x1_out_v
    PORT
      LAYER li1 ;
        RECT 480.750 161.920 480.980 163.420 ;
    END
  END x1_out_v
  PIN out_v
    PORT
      LAYER li1 ;
        RECT 481.825 160.250 482.600 160.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 484.820 160.105 499.220 160.705 ;
    END
  END out_v
  PIN d7
    PORT
      LAYER li1 ;
        RECT 469.650 159.460 469.835 159.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 467.920 149.270 499.220 150.070 ;
    END
  END d7
  PIN inp1
    PORT
      LAYER li1 ;
        RECT 3.980 278.435 4.270 278.670 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.995 280.105 4.885 320.560 ;
    END
  END inp1
  PIN x2_vref1
    PORT
      LAYER li1 ;
        RECT 103.880 34.250 104.390 35.180 ;
    END
  END x2_vref1
  PIN x1_vref5
    PORT
      LAYER li1 ;
        RECT 103.000 36.230 103.510 37.100 ;
    END
  END x1_vref5
  PIN inp2
    PORT
      LAYER met2 ;
        RECT 339.785 0.000 340.365 10.275 ;
    END
  END inp2

  PIN gnd
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 55.030 281.005 60.350 320.560 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.185 279.130 19.505 320.560 ;
    END
  END vdd
  OBS
      LAYER li1 ;
        RECT 0.000 278.840 481.825 283.120 ;
        RECT 0.000 278.265 3.810 278.840 ;
        RECT 4.440 278.265 481.825 278.840 ;
        RECT 0.000 163.590 481.825 278.265 ;
        RECT 0.000 161.750 480.580 163.590 ;
        RECT 481.150 161.750 481.825 163.590 ;
        RECT 0.000 160.740 481.825 161.750 ;
        RECT 0.000 160.090 481.655 160.740 ;
        RECT 0.000 159.290 469.480 160.090 ;
        RECT 470.005 160.080 481.655 160.090 ;
        RECT 470.005 159.290 481.825 160.080 ;
        RECT 0.000 158.330 481.825 159.290 ;
        RECT 0.000 155.740 480.690 158.330 ;
        RECT 481.240 155.740 481.825 158.330 ;
        RECT 0.000 48.320 481.825 155.740 ;
        RECT 0.000 37.270 188.870 48.320 ;
        RECT 0.000 36.060 102.830 37.270 ;
        RECT 103.680 36.060 188.870 37.270 ;
        RECT 0.000 35.350 188.870 36.060 ;
        RECT 0.000 34.080 103.710 35.350 ;
        RECT 104.560 34.080 188.870 35.350 ;
        RECT 0.000 30.580 188.870 34.080 ;
        RECT 0.000 29.150 171.560 30.580 ;
        RECT 0.000 27.680 155.350 29.150 ;
        RECT 0.000 26.440 138.380 27.680 ;
        RECT 0.000 25.770 121.680 26.440 ;
        RECT 0.000 19.225 106.290 25.770 ;
        RECT 106.930 19.790 121.680 25.770 ;
        RECT 122.320 20.710 138.380 26.440 ;
        RECT 139.020 21.620 155.350 27.680 ;
        RECT 155.990 22.930 171.560 29.150 ;
        RECT 172.200 23.240 188.870 30.580 ;
        RECT 189.510 31.940 481.825 48.320 ;
        RECT 189.510 24.210 215.290 31.940 ;
        RECT 215.960 24.210 481.825 31.940 ;
        RECT 189.510 23.240 481.825 24.210 ;
        RECT 172.200 22.930 481.825 23.240 ;
        RECT 155.990 21.620 481.825 22.930 ;
        RECT 139.020 20.710 481.825 21.620 ;
        RECT 122.320 19.790 481.825 20.710 ;
        RECT 106.930 19.225 481.825 19.790 ;
        RECT 0.000 19.150 481.825 19.225 ;
      LAYER met1 ;
        RECT 3.125 10.265 483.290 282.230 ;
      LAYER met2 ;
        RECT 3.125 279.825 3.715 318.560 ;
        RECT 5.165 279.825 485.000 318.560 ;
        RECT 3.125 158.550 485.000 279.825 ;
        RECT 3.125 157.530 469.390 158.550 ;
        RECT 470.645 157.530 485.000 158.550 ;
        RECT 3.125 10.625 485.000 157.530 ;
        RECT 3.125 4.280 139.100 10.625 ;
        RECT 3.125 4.000 106.430 4.280 ;
        RECT 107.570 4.000 123.815 4.280 ;
        RECT 124.955 4.000 139.100 4.280 ;
        RECT 140.240 4.000 157.495 10.625 ;
        RECT 158.635 10.620 220.680 10.625 ;
        RECT 158.635 4.000 175.565 10.620 ;
        RECT 176.705 4.000 193.240 10.620 ;
        RECT 194.380 4.000 220.680 10.620 ;
        RECT 221.820 10.555 485.000 10.625 ;
        RECT 221.820 4.000 339.505 10.555 ;
        RECT 340.645 4.000 485.000 10.555 ;
      LAYER met3 ;
        RECT 10.220 161.105 497.080 282.315 ;
        RECT 10.220 159.705 484.420 161.105 ;
        RECT 10.220 150.470 497.080 159.705 ;
        RECT 10.220 148.870 467.520 150.470 ;
        RECT 10.220 44.630 497.080 148.870 ;
      LAYER met4 ;
        RECT 10.230 278.730 13.785 282.810 ;
        RECT 19.905 280.605 54.630 282.810 ;
        RECT 60.750 280.605 474.450 282.810 ;
        RECT 19.905 278.730 474.450 280.605 ;
        RECT 10.230 166.410 474.450 278.730 ;
        RECT 10.230 162.560 473.680 166.410 ;
        RECT 10.230 45.490 474.450 162.560 ;
  END
END DAC_8BIT
END LIBRARY

