(* blackbox *)
module sky130_fd_sc_hvl__inv_1 (
    A   ,
    VGND   ,
    VNB    ,
    VPB    ,
    VPWR   ,
    Y   
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
endmodule

(* blackbox *)
module sky130_fd_sc_hvl__inv_4 (
    A   ,
    VGND   ,
    VNB    ,
    VPB    ,
    VPWR   ,
    Y   
);

    output Y   ;
    input  A   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
endmodule



(* blackbox *)
module sky130_fd_sc_hvl__nand3_1 (

    A   ,
    B   ,
    C   ,
    VGND   ,
    VNB    ,
    VPB    ,
    VPWR   ,
    Y 
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
endmodule


(* blackbox *)
module sky130_fd_sc_hvl__nor3_1 (
    A   ,
    B   ,
    C   ,
    VGND   ,
    VNB    ,
    VPB    ,
    VPWR   ,
    Y
);

    output Y   ;
    input  A   ;
    input  B   ;
    input  C   ;
    input  VPWR;
    input  VGND;
    input  VPB ;
    input  VNB ;
endmodule

