magic
tech sky130A
magscale 1 2
timestamp 1626434083
<< locali >>
rect 236469 335971 236503 336617
rect 314577 336583 314611 336685
rect 316417 336379 316451 336617
rect 354873 336583 354907 336685
rect 380909 336039 380943 336141
rect 425529 7123 425563 7837
rect 162593 4981 162961 5015
rect 162593 4811 162627 4981
rect 162685 4811 162719 4913
rect 171793 3451 171827 4165
rect 269865 3995 269899 4165
rect 272475 4097 272717 4131
rect 272567 4029 272659 4063
rect 269957 3791 269991 3961
rect 272625 3927 272659 4029
rect 275937 3961 276305 3995
rect 271797 3519 271831 3757
rect 272441 3655 272475 3893
rect 271797 3485 271889 3519
rect 110429 3043 110463 3145
rect 117973 2907 118007 3009
rect 258181 2907 258215 3485
rect 272533 3383 272567 3825
rect 274925 3587 274959 3689
rect 275937 3587 275971 3961
rect 272625 3383 272659 3485
rect 277317 3383 277351 3485
rect 277259 3349 277351 3383
rect 278053 3315 278087 3621
rect 278145 3247 278179 3893
rect 325525 3587 325559 3825
rect 325617 3723 325651 4097
<< viali >>
rect 314577 336685 314611 336719
rect 236469 336617 236503 336651
rect 354873 336685 354907 336719
rect 314577 336549 314611 336583
rect 316417 336617 316451 336651
rect 354873 336549 354907 336583
rect 316417 336345 316451 336379
rect 380909 336141 380943 336175
rect 380909 336005 380943 336039
rect 236469 335937 236503 335971
rect 425529 7837 425563 7871
rect 425529 7089 425563 7123
rect 162961 4981 162995 5015
rect 162593 4777 162627 4811
rect 162685 4913 162719 4947
rect 162685 4777 162719 4811
rect 171793 4165 171827 4199
rect 269865 4165 269899 4199
rect 272441 4097 272475 4131
rect 272717 4097 272751 4131
rect 325617 4097 325651 4131
rect 272533 4029 272567 4063
rect 269865 3961 269899 3995
rect 269957 3961 269991 3995
rect 272441 3893 272475 3927
rect 272625 3893 272659 3927
rect 276305 3961 276339 3995
rect 269957 3757 269991 3791
rect 271797 3757 271831 3791
rect 272441 3621 272475 3655
rect 272533 3825 272567 3859
rect 171793 3417 171827 3451
rect 258181 3485 258215 3519
rect 271889 3485 271923 3519
rect 110429 3145 110463 3179
rect 110429 3009 110463 3043
rect 117973 3009 118007 3043
rect 117973 2873 118007 2907
rect 274925 3689 274959 3723
rect 274925 3553 274959 3587
rect 278145 3893 278179 3927
rect 275937 3553 275971 3587
rect 278053 3621 278087 3655
rect 272533 3349 272567 3383
rect 272625 3485 272659 3519
rect 277317 3485 277351 3519
rect 272625 3349 272659 3383
rect 277225 3349 277259 3383
rect 278053 3281 278087 3315
rect 325525 3825 325559 3859
rect 325617 3689 325651 3723
rect 325525 3553 325559 3587
rect 278145 3213 278179 3247
rect 258181 2873 258215 2907
<< metal1 >>
rect 360102 700884 360108 700936
rect 360160 700924 360166 700936
rect 429838 700924 429844 700936
rect 360160 700896 429844 700924
rect 360160 700884 360166 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 367002 700816 367008 700868
rect 367060 700856 367066 700868
rect 446122 700856 446128 700868
rect 367060 700828 446128 700856
rect 367060 700816 367066 700828
rect 446122 700816 446128 700828
rect 446180 700816 446186 700868
rect 373902 700748 373908 700800
rect 373960 700788 373966 700800
rect 462314 700788 462320 700800
rect 373960 700760 462320 700788
rect 373960 700748 373966 700760
rect 462314 700748 462320 700760
rect 462372 700748 462378 700800
rect 382182 700680 382188 700732
rect 382240 700720 382246 700732
rect 478506 700720 478512 700732
rect 382240 700692 478512 700720
rect 382240 700680 382246 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 389082 700612 389088 700664
rect 389140 700652 389146 700664
rect 494790 700652 494796 700664
rect 389140 700624 494796 700652
rect 389140 700612 389146 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 395982 700544 395988 700596
rect 396040 700584 396046 700596
rect 510982 700584 510988 700596
rect 396040 700556 510988 700584
rect 396040 700544 396046 700556
rect 510982 700544 510988 700556
rect 511040 700544 511046 700596
rect 331122 700476 331128 700528
rect 331180 700516 331186 700528
rect 364978 700516 364984 700528
rect 331180 700488 364984 700516
rect 331180 700476 331186 700488
rect 364978 700476 364984 700488
rect 365036 700476 365042 700528
rect 402882 700476 402888 700528
rect 402940 700516 402946 700528
rect 527174 700516 527180 700528
rect 402940 700488 527180 700516
rect 402940 700476 402946 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 338022 700408 338028 700460
rect 338080 700448 338086 700460
rect 381170 700448 381176 700460
rect 338080 700420 381176 700448
rect 338080 700408 338086 700420
rect 381170 700408 381176 700420
rect 381228 700408 381234 700460
rect 411162 700408 411168 700460
rect 411220 700448 411226 700460
rect 543458 700448 543464 700460
rect 411220 700420 543464 700448
rect 411220 700408 411226 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 235902 700380 235908 700392
rect 235224 700352 235908 700380
rect 235224 700340 235230 700352
rect 235902 700340 235908 700352
rect 235960 700340 235966 700392
rect 317322 700340 317328 700392
rect 317380 700380 317386 700392
rect 332502 700380 332508 700392
rect 317380 700352 332508 700380
rect 317380 700340 317386 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 344922 700340 344928 700392
rect 344980 700380 344986 700392
rect 397454 700380 397460 700392
rect 344980 700352 397460 700380
rect 344980 700340 344986 700352
rect 397454 700340 397460 700352
rect 397512 700340 397518 700392
rect 418062 700340 418068 700392
rect 418120 700380 418126 700392
rect 559650 700380 559656 700392
rect 418120 700352 559656 700380
rect 418120 700340 418126 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 324222 700272 324228 700324
rect 324280 700312 324286 700324
rect 348786 700312 348792 700324
rect 324280 700284 348792 700312
rect 324280 700272 324286 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 353202 700272 353208 700324
rect 353260 700312 353266 700324
rect 413646 700312 413652 700324
rect 353260 700284 413652 700312
rect 353260 700272 353266 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 424962 700272 424968 700324
rect 425020 700312 425026 700324
rect 575842 700312 575848 700324
rect 425020 700284 575848 700312
rect 425020 700272 425026 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 56778 700136 56784 700188
rect 56836 700176 56842 700188
rect 57882 700176 57888 700188
rect 56836 700148 57888 700176
rect 56836 700136 56842 700148
rect 57882 700136 57888 700148
rect 57940 700136 57946 700188
rect 186498 700136 186504 700188
rect 186556 700176 186562 700188
rect 187602 700176 187608 700188
rect 186556 700148 187608 700176
rect 186556 700136 186562 700148
rect 187602 700136 187608 700148
rect 187660 700136 187666 700188
rect 251450 700068 251456 700120
rect 251508 700108 251514 700120
rect 252462 700108 252468 700120
rect 251508 700080 252468 700108
rect 251508 700068 251514 700080
rect 252462 700068 252468 700080
rect 252520 700068 252526 700120
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 122742 699700 122748 699712
rect 121696 699672 122748 699700
rect 121696 699660 121702 699672
rect 122742 699660 122748 699672
rect 122800 699660 122806 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 309778 699660 309784 699712
rect 309836 699700 309842 699712
rect 316310 699700 316316 699712
rect 309836 699672 316316 699700
rect 309836 699660 309842 699672
rect 316310 699660 316316 699672
rect 316368 699660 316374 699712
rect 429838 696940 429844 696992
rect 429896 696980 429902 696992
rect 580166 696980 580172 696992
rect 429896 696952 580172 696980
rect 429896 696940 429902 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429930 683136 429936 683188
rect 429988 683176 429994 683188
rect 580166 683176 580172 683188
rect 429988 683148 580172 683176
rect 429988 683136 429994 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 430022 670692 430028 670744
rect 430080 670732 430086 670744
rect 580166 670732 580172 670744
rect 430080 670704 580172 670732
rect 430080 670692 430086 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 430114 643084 430120 643136
rect 430172 643124 430178 643136
rect 580166 643124 580172 643136
rect 430172 643096 580172 643124
rect 430172 643084 430178 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 430206 630640 430212 630692
rect 430264 630680 430270 630692
rect 579982 630680 579988 630692
rect 430264 630652 579988 630680
rect 430264 630640 430270 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 430298 616836 430304 616888
rect 430356 616876 430362 616888
rect 580166 616876 580172 616888
rect 430356 616848 580172 616876
rect 430356 616836 430362 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 430390 590656 430396 590708
rect 430448 590696 430454 590708
rect 579614 590696 579620 590708
rect 430448 590668 579620 590696
rect 430448 590656 430454 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 430482 576852 430488 576904
rect 430540 576892 430546 576904
rect 579614 576892 579620 576904
rect 430540 576864 579620 576892
rect 430540 576852 430546 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 429746 563048 429752 563100
rect 429804 563088 429810 563100
rect 579890 563088 579896 563100
rect 429804 563060 579896 563088
rect 429804 563048 429810 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 429654 536800 429660 536852
rect 429712 536840 429718 536852
rect 580166 536840 580172 536852
rect 429712 536812 580172 536840
rect 429712 536800 429718 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 429562 524424 429568 524476
rect 429620 524464 429626 524476
rect 580166 524464 580172 524476
rect 429620 524436 580172 524464
rect 429620 524424 429626 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 171042 500896 171048 500948
rect 171100 500936 171106 500948
rect 243814 500936 243820 500948
rect 171100 500908 243820 500936
rect 171100 500896 171106 500908
rect 243814 500896 243820 500908
rect 243872 500896 243878 500948
rect 300762 500896 300768 500948
rect 300820 500936 300826 500948
rect 301590 500936 301596 500948
rect 300820 500908 301596 500936
rect 300820 500896 300826 500908
rect 301590 500896 301596 500908
rect 301648 500896 301654 500948
rect 308766 500896 308772 500948
rect 308824 500936 308830 500948
rect 309778 500936 309784 500948
rect 308824 500908 309784 500936
rect 308824 500896 308830 500908
rect 309778 500896 309784 500908
rect 309836 500896 309842 500948
rect 359366 500896 359372 500948
rect 359424 500936 359430 500948
rect 360102 500936 360108 500948
rect 359424 500908 360108 500936
rect 359424 500896 359430 500908
rect 360102 500896 360108 500908
rect 360160 500896 360166 500948
rect 380986 500896 380992 500948
rect 381044 500936 381050 500948
rect 382182 500936 382188 500948
rect 381044 500908 382188 500936
rect 381044 500896 381050 500908
rect 382182 500896 382188 500908
rect 382240 500896 382246 500948
rect 388254 500896 388260 500948
rect 388312 500936 388318 500948
rect 389082 500936 389088 500948
rect 388312 500908 389088 500936
rect 388312 500896 388318 500908
rect 389082 500896 389088 500908
rect 389140 500896 389146 500948
rect 417142 500896 417148 500948
rect 417200 500936 417206 500948
rect 418062 500936 418068 500948
rect 417200 500908 418068 500936
rect 417200 500896 417206 500908
rect 418062 500896 418068 500908
rect 418120 500896 418126 500948
rect 154482 500828 154488 500880
rect 154540 500868 154546 500880
rect 236546 500868 236552 500880
rect 154540 500840 236552 500868
rect 154540 500828 154546 500840
rect 236546 500828 236552 500840
rect 236604 500828 236610 500880
rect 137922 500760 137928 500812
rect 137980 500800 137986 500812
rect 229370 500800 229376 500812
rect 137980 500772 229376 500800
rect 137980 500760 137986 500772
rect 229370 500760 229376 500772
rect 229428 500760 229434 500812
rect 122742 500692 122748 500744
rect 122800 500732 122806 500744
rect 222102 500732 222108 500744
rect 122800 500704 222108 500732
rect 122800 500692 122806 500704
rect 222102 500692 222108 500704
rect 222160 500692 222166 500744
rect 106182 500624 106188 500676
rect 106240 500664 106246 500676
rect 214926 500664 214932 500676
rect 106240 500636 214932 500664
rect 106240 500624 106246 500636
rect 214926 500624 214932 500636
rect 214984 500624 214990 500676
rect 89622 500556 89628 500608
rect 89680 500596 89686 500608
rect 207658 500596 207664 500608
rect 89680 500568 207664 500596
rect 89680 500556 89686 500568
rect 207658 500556 207664 500568
rect 207716 500556 207722 500608
rect 316034 500556 316040 500608
rect 316092 500596 316098 500608
rect 317322 500596 317328 500608
rect 316092 500568 317328 500596
rect 316092 500556 316098 500568
rect 317322 500556 317328 500568
rect 317380 500556 317386 500608
rect 409874 500556 409880 500608
rect 409932 500596 409938 500608
rect 411162 500596 411168 500608
rect 409932 500568 411168 500596
rect 409932 500556 409938 500568
rect 411162 500556 411168 500568
rect 411220 500556 411226 500608
rect 73062 500488 73068 500540
rect 73120 500528 73126 500540
rect 200482 500528 200488 500540
rect 73120 500500 200488 500528
rect 73120 500488 73126 500500
rect 200482 500488 200488 500500
rect 200540 500488 200546 500540
rect 323210 500488 323216 500540
rect 323268 500528 323274 500540
rect 324222 500528 324228 500540
rect 323268 500500 324228 500528
rect 323268 500488 323274 500500
rect 324222 500488 324228 500500
rect 324280 500488 324286 500540
rect 57882 500420 57888 500472
rect 57940 500460 57946 500472
rect 193214 500460 193220 500472
rect 57940 500432 193220 500460
rect 57940 500420 57946 500432
rect 193214 500420 193220 500432
rect 193272 500420 193278 500472
rect 235902 500420 235908 500472
rect 235960 500460 235966 500472
rect 272702 500460 272708 500472
rect 235960 500432 272708 500460
rect 235960 500420 235966 500432
rect 272702 500420 272708 500432
rect 272760 500420 272766 500472
rect 352098 500420 352104 500472
rect 352156 500460 352162 500472
rect 353202 500460 353208 500472
rect 352156 500432 353208 500460
rect 352156 500420 352162 500432
rect 353202 500420 353208 500432
rect 353260 500420 353266 500472
rect 41322 500352 41328 500404
rect 41380 500392 41386 500404
rect 186038 500392 186044 500404
rect 41380 500364 186044 500392
rect 41380 500352 41386 500364
rect 186038 500352 186044 500364
rect 186096 500352 186102 500404
rect 219342 500352 219348 500404
rect 219400 500392 219406 500404
rect 265434 500392 265440 500404
rect 219400 500364 265440 500392
rect 219400 500352 219406 500364
rect 265434 500352 265440 500364
rect 265492 500352 265498 500404
rect 24762 500284 24768 500336
rect 24820 500324 24826 500336
rect 178770 500324 178776 500336
rect 24820 500296 178776 500324
rect 24820 500284 24826 500296
rect 178770 500284 178776 500296
rect 178828 500284 178834 500336
rect 202782 500284 202788 500336
rect 202840 500324 202846 500336
rect 258258 500324 258264 500336
rect 202840 500296 258264 500324
rect 202840 500284 202846 500296
rect 258258 500284 258264 500296
rect 258316 500284 258322 500336
rect 267642 500284 267648 500336
rect 267700 500324 267706 500336
rect 287146 500324 287152 500336
rect 267700 500296 287152 500324
rect 267700 500284 267706 500296
rect 287146 500284 287152 500296
rect 287204 500284 287210 500336
rect 8202 500216 8208 500268
rect 8260 500256 8266 500268
rect 171594 500256 171600 500268
rect 8260 500228 171600 500256
rect 8260 500216 8266 500228
rect 171594 500216 171600 500228
rect 171652 500216 171658 500268
rect 187602 500216 187608 500268
rect 187660 500256 187666 500268
rect 250990 500256 250996 500268
rect 187660 500228 250996 500256
rect 187660 500216 187666 500228
rect 250990 500216 250996 500228
rect 251048 500216 251054 500268
rect 252462 500216 252468 500268
rect 252520 500256 252526 500268
rect 279878 500256 279884 500268
rect 252520 500228 279884 500256
rect 252520 500216 252526 500228
rect 279878 500216 279884 500228
rect 279936 500216 279942 500268
rect 284202 500216 284208 500268
rect 284260 500256 284266 500268
rect 294322 500256 294328 500268
rect 284260 500228 294328 500256
rect 284260 500216 284266 500228
rect 294322 500216 294328 500228
rect 294380 500216 294386 500268
rect 3418 493960 3424 494012
rect 3476 494000 3482 494012
rect 165614 494000 165620 494012
rect 3476 493972 165620 494000
rect 3476 493960 3482 493972
rect 165614 493960 165620 493972
rect 165672 493960 165678 494012
rect 3510 491240 3516 491292
rect 3568 491280 3574 491292
rect 165614 491280 165620 491292
rect 3568 491252 165620 491280
rect 3568 491240 3574 491252
rect 165614 491240 165620 491252
rect 165672 491240 165678 491292
rect 3602 488452 3608 488504
rect 3660 488492 3666 488504
rect 165614 488492 165620 488504
rect 3660 488464 165620 488492
rect 3660 488452 3666 488464
rect 165614 488452 165620 488464
rect 165672 488452 165678 488504
rect 429378 488452 429384 488504
rect 429436 488492 429442 488504
rect 580258 488492 580264 488504
rect 429436 488464 580264 488492
rect 429436 488452 429442 488464
rect 580258 488452 580264 488464
rect 580316 488452 580322 488504
rect 3694 485732 3700 485784
rect 3752 485772 3758 485784
rect 165614 485772 165620 485784
rect 3752 485744 165620 485772
rect 3752 485732 3758 485744
rect 165614 485732 165620 485744
rect 165672 485732 165678 485784
rect 429838 484372 429844 484424
rect 429896 484412 429902 484424
rect 579614 484412 579620 484424
rect 429896 484384 579620 484412
rect 429896 484372 429902 484384
rect 579614 484372 579620 484384
rect 579672 484372 579678 484424
rect 3786 481584 3792 481636
rect 3844 481624 3850 481636
rect 165614 481624 165620 481636
rect 3844 481596 165620 481624
rect 3844 481584 3850 481596
rect 165614 481584 165620 481596
rect 165672 481584 165678 481636
rect 3878 478796 3884 478848
rect 3936 478836 3942 478848
rect 165614 478836 165620 478848
rect 3936 478808 165620 478836
rect 3936 478796 3942 478808
rect 165614 478796 165620 478808
rect 165672 478796 165678 478848
rect 3970 476008 3976 476060
rect 4028 476048 4034 476060
rect 165614 476048 165620 476060
rect 4028 476020 165620 476048
rect 4028 476008 4034 476020
rect 165614 476008 165620 476020
rect 165672 476008 165678 476060
rect 429470 476008 429476 476060
rect 429528 476048 429534 476060
rect 580350 476048 580356 476060
rect 429528 476020 580356 476048
rect 429528 476008 429534 476020
rect 580350 476008 580356 476020
rect 580408 476008 580414 476060
rect 4062 473288 4068 473340
rect 4120 473328 4126 473340
rect 165614 473328 165620 473340
rect 4120 473300 165620 473328
rect 4120 473288 4126 473300
rect 165614 473288 165620 473300
rect 165672 473288 165678 473340
rect 429930 470568 429936 470620
rect 429988 470608 429994 470620
rect 579614 470608 579620 470620
rect 429988 470580 579620 470608
rect 429988 470568 429994 470580
rect 579614 470568 579620 470580
rect 579672 470568 579678 470620
rect 3326 470500 3332 470552
rect 3384 470540 3390 470552
rect 165614 470540 165620 470552
rect 3384 470512 165620 470540
rect 3384 470500 3390 470512
rect 165614 470500 165620 470512
rect 165672 470500 165678 470552
rect 3234 467780 3240 467832
rect 3292 467820 3298 467832
rect 165614 467820 165620 467832
rect 3292 467792 165620 467820
rect 3292 467780 3298 467792
rect 165614 467780 165620 467792
rect 165672 467780 165678 467832
rect 3142 464992 3148 465044
rect 3200 465032 3206 465044
rect 165614 465032 165620 465044
rect 3200 465004 165620 465032
rect 3200 464992 3206 465004
rect 165614 464992 165620 465004
rect 165672 464992 165678 465044
rect 429194 463632 429200 463684
rect 429252 463672 429258 463684
rect 580442 463672 580448 463684
rect 429252 463644 580448 463672
rect 429252 463632 429258 463644
rect 580442 463632 580448 463644
rect 580500 463632 580506 463684
rect 3050 460844 3056 460896
rect 3108 460884 3114 460896
rect 165614 460884 165620 460896
rect 3108 460856 165620 460884
rect 3108 460844 3114 460856
rect 165614 460844 165620 460856
rect 165672 460844 165678 460896
rect 2958 458124 2964 458176
rect 3016 458164 3022 458176
rect 165614 458164 165620 458176
rect 3016 458136 165620 458164
rect 3016 458124 3022 458136
rect 165614 458124 165620 458136
rect 165672 458124 165678 458176
rect 430022 456764 430028 456816
rect 430080 456804 430086 456816
rect 580166 456804 580172 456816
rect 430080 456776 580172 456804
rect 430080 456764 430086 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 2866 455336 2872 455388
rect 2924 455376 2930 455388
rect 165614 455376 165620 455388
rect 2924 455348 165620 455376
rect 2924 455336 2930 455348
rect 165614 455336 165620 455348
rect 165672 455336 165678 455388
rect 429194 455336 429200 455388
rect 429252 455376 429258 455388
rect 580534 455376 580540 455388
rect 429252 455348 580540 455376
rect 429252 455336 429258 455348
rect 580534 455336 580540 455348
rect 580592 455336 580598 455388
rect 2774 452548 2780 452600
rect 2832 452588 2838 452600
rect 165614 452588 165620 452600
rect 2832 452560 165620 452588
rect 2832 452548 2838 452560
rect 165614 452548 165620 452560
rect 165672 452548 165678 452600
rect 429562 451188 429568 451240
rect 429620 451228 429626 451240
rect 580626 451228 580632 451240
rect 429620 451200 580632 451228
rect 429620 451188 429626 451200
rect 580626 451188 580632 451200
rect 580684 451188 580690 451240
rect 3418 449828 3424 449880
rect 3476 449868 3482 449880
rect 165614 449868 165620 449880
rect 3476 449840 165620 449868
rect 3476 449828 3482 449840
rect 165614 449828 165620 449840
rect 165672 449828 165678 449880
rect 3510 447040 3516 447092
rect 3568 447080 3574 447092
rect 165614 447080 165620 447092
rect 3568 447052 165620 447080
rect 3568 447040 3574 447052
rect 165614 447040 165620 447052
rect 165672 447040 165678 447092
rect 429838 444388 429844 444440
rect 429896 444428 429902 444440
rect 580166 444428 580172 444440
rect 429896 444400 580172 444428
rect 429896 444388 429902 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 3602 444320 3608 444372
rect 3660 444360 3666 444372
rect 165614 444360 165620 444372
rect 3660 444332 165620 444360
rect 3660 444320 3666 444332
rect 165614 444320 165620 444332
rect 165672 444320 165678 444372
rect 3694 440172 3700 440224
rect 3752 440212 3758 440224
rect 165614 440212 165620 440224
rect 3752 440184 165620 440212
rect 3752 440172 3758 440184
rect 165614 440172 165620 440184
rect 165672 440172 165678 440224
rect 3418 436704 3424 436756
rect 3476 436744 3482 436756
rect 165614 436744 165620 436756
rect 3476 436716 165620 436744
rect 3476 436704 3482 436716
rect 165614 436704 165620 436716
rect 165672 436704 165678 436756
rect 3418 433304 3424 433356
rect 3476 433344 3482 433356
rect 165614 433344 165620 433356
rect 3476 433316 165620 433344
rect 3476 433304 3482 433316
rect 165614 433304 165620 433316
rect 165672 433304 165678 433356
rect 429930 431876 429936 431928
rect 429988 431916 429994 431928
rect 579798 431916 579804 431928
rect 429988 431888 579804 431916
rect 429988 431876 429994 431888
rect 579798 431876 579804 431888
rect 579856 431876 579862 431928
rect 3786 430584 3792 430636
rect 3844 430624 3850 430636
rect 165614 430624 165620 430636
rect 3844 430596 165620 430624
rect 3844 430584 3850 430596
rect 165614 430584 165620 430596
rect 165672 430584 165678 430636
rect 3694 427796 3700 427848
rect 3752 427836 3758 427848
rect 165614 427836 165620 427848
rect 3752 427808 165620 427836
rect 3752 427796 3758 427808
rect 165614 427796 165620 427808
rect 165672 427796 165678 427848
rect 3602 420928 3608 420980
rect 3660 420968 3666 420980
rect 165614 420968 165620 420980
rect 3660 420940 165620 420968
rect 3660 420928 3666 420940
rect 165614 420928 165620 420940
rect 165672 420928 165678 420980
rect 429838 419432 429844 419484
rect 429896 419472 429902 419484
rect 580166 419472 580172 419484
rect 429896 419444 580172 419472
rect 429896 419432 429902 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 3510 418140 3516 418192
rect 3568 418180 3574 418192
rect 165614 418180 165620 418192
rect 3568 418152 165620 418180
rect 3568 418140 3574 418152
rect 165614 418140 165620 418152
rect 165672 418140 165678 418192
rect 3418 415420 3424 415472
rect 3476 415460 3482 415472
rect 165614 415460 165620 415472
rect 3476 415432 165620 415460
rect 3476 415420 3482 415432
rect 165614 415420 165620 415432
rect 165672 415420 165678 415472
rect 429562 414808 429568 414860
rect 429620 414848 429626 414860
rect 433978 414848 433984 414860
rect 429620 414820 433984 414848
rect 429620 414808 429626 414820
rect 433978 414808 433984 414820
rect 434036 414808 434042 414860
rect 429562 411272 429568 411324
rect 429620 411312 429626 411324
rect 435358 411312 435364 411324
rect 429620 411284 435364 411312
rect 429620 411272 429626 411284
rect 435358 411272 435364 411284
rect 435416 411272 435422 411324
rect 429470 408484 429476 408536
rect 429528 408524 429534 408536
rect 461578 408524 461584 408536
rect 429528 408496 461584 408524
rect 429528 408484 429534 408496
rect 461578 408484 461584 408496
rect 461636 408484 461642 408536
rect 3142 407124 3148 407176
rect 3200 407164 3206 407176
rect 165614 407164 165620 407176
rect 3200 407136 165620 407164
rect 3200 407124 3206 407136
rect 165614 407124 165620 407136
rect 165672 407124 165678 407176
rect 430206 405628 430212 405680
rect 430264 405668 430270 405680
rect 580166 405668 580172 405680
rect 430264 405640 580172 405668
rect 430264 405628 430270 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 3234 404336 3240 404388
rect 3292 404376 3298 404388
rect 165614 404376 165620 404388
rect 3292 404348 165620 404376
rect 3292 404336 3298 404348
rect 165614 404336 165620 404348
rect 165672 404336 165678 404388
rect 429562 402704 429568 402756
rect 429620 402744 429626 402756
rect 432598 402744 432604 402756
rect 429620 402716 432604 402744
rect 429620 402704 429626 402716
rect 432598 402704 432604 402716
rect 432656 402704 432662 402756
rect 22738 394680 22744 394732
rect 22796 394720 22802 394732
rect 165614 394720 165620 394732
rect 22796 394692 165620 394720
rect 22796 394680 22802 394692
rect 165614 394680 165620 394692
rect 165672 394680 165678 394732
rect 7558 391960 7564 392012
rect 7616 392000 7622 392012
rect 165614 392000 165620 392012
rect 7616 391972 165620 392000
rect 7616 391960 7622 391972
rect 165614 391960 165620 391972
rect 165672 391960 165678 392012
rect 430114 391892 430120 391944
rect 430172 391932 430178 391944
rect 580166 391932 580172 391944
rect 430172 391904 580172 391932
rect 430172 391892 430178 391904
rect 580166 391892 580172 391904
rect 580224 391892 580230 391944
rect 429562 390736 429568 390788
rect 429620 390776 429626 390788
rect 431218 390776 431224 390788
rect 429620 390748 431224 390776
rect 429620 390736 429626 390748
rect 431218 390736 431224 390748
rect 431276 390736 431282 390788
rect 429562 387812 429568 387864
rect 429620 387852 429626 387864
rect 454678 387852 454684 387864
rect 429620 387824 454684 387852
rect 429620 387812 429626 387824
rect 454678 387812 454684 387824
rect 454736 387812 454742 387864
rect 3326 384956 3332 385008
rect 3384 384996 3390 385008
rect 166258 384996 166264 385008
rect 3384 384968 166264 384996
rect 3384 384956 3390 384968
rect 166258 384956 166264 384968
rect 166316 384956 166322 385008
rect 3326 383664 3332 383716
rect 3384 383704 3390 383716
rect 165614 383704 165620 383716
rect 3384 383676 165620 383704
rect 3384 383664 3390 383676
rect 165614 383664 165620 383676
rect 165672 383664 165678 383716
rect 14458 379516 14464 379568
rect 14516 379556 14522 379568
rect 165614 379556 165620 379568
rect 14516 379528 165620 379556
rect 14516 379516 14522 379528
rect 165614 379516 165620 379528
rect 165672 379516 165678 379568
rect 430022 379448 430028 379500
rect 430080 379488 430086 379500
rect 580166 379488 580172 379500
rect 430080 379460 580172 379488
rect 430080 379448 430086 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 4062 374008 4068 374060
rect 4120 374048 4126 374060
rect 165614 374048 165620 374060
rect 4120 374020 165620 374048
rect 4120 374008 4126 374020
rect 165614 374008 165620 374020
rect 165672 374008 165678 374060
rect 25498 371220 25504 371272
rect 25556 371260 25562 371272
rect 165614 371260 165620 371272
rect 25556 371232 165620 371260
rect 25556 371220 25562 371232
rect 165614 371220 165620 371232
rect 165672 371220 165678 371272
rect 3970 368500 3976 368552
rect 4028 368540 4034 368552
rect 165614 368540 165620 368552
rect 4028 368512 165620 368540
rect 4028 368500 4034 368512
rect 165614 368500 165620 368512
rect 165672 368500 165678 368552
rect 429930 368500 429936 368552
rect 429988 368540 429994 368552
rect 447778 368540 447784 368552
rect 429988 368512 447784 368540
rect 429988 368500 429994 368512
rect 447778 368500 447784 368512
rect 447836 368500 447842 368552
rect 430022 365644 430028 365696
rect 430080 365684 430086 365696
rect 580166 365684 580172 365696
rect 430080 365656 580172 365684
rect 430080 365644 430086 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3878 362924 3884 362976
rect 3936 362964 3942 362976
rect 165614 362964 165620 362976
rect 3936 362936 165620 362964
rect 3936 362924 3942 362936
rect 165614 362924 165620 362936
rect 165672 362924 165678 362976
rect 3786 358776 3792 358828
rect 3844 358816 3850 358828
rect 165614 358816 165620 358828
rect 3844 358788 165620 358816
rect 3844 358776 3850 358788
rect 165614 358776 165620 358788
rect 165672 358776 165678 358828
rect 15838 356056 15844 356108
rect 15896 356096 15902 356108
rect 165614 356096 165620 356108
rect 15896 356068 165620 356096
rect 15896 356056 15902 356068
rect 165614 356056 165620 356068
rect 165672 356056 165678 356108
rect 3694 353268 3700 353320
rect 3752 353308 3758 353320
rect 165614 353308 165620 353320
rect 3752 353280 165620 353308
rect 3752 353268 3758 353280
rect 165614 353268 165620 353280
rect 165672 353268 165678 353320
rect 429930 353200 429936 353252
rect 429988 353240 429994 353252
rect 580166 353240 580172 353252
rect 429988 353212 580172 353240
rect 429988 353200 429994 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 32398 350548 32404 350600
rect 32456 350588 32462 350600
rect 165614 350588 165620 350600
rect 32456 350560 165620 350588
rect 32456 350548 32462 350560
rect 165614 350548 165620 350560
rect 165672 350548 165678 350600
rect 429838 350548 429844 350600
rect 429896 350588 429902 350600
rect 442258 350588 442264 350600
rect 429896 350560 442264 350588
rect 429896 350548 429902 350560
rect 442258 350548 442264 350560
rect 442316 350548 442322 350600
rect 3602 347760 3608 347812
rect 3660 347800 3666 347812
rect 165614 347800 165620 347812
rect 3660 347772 165620 347800
rect 3660 347760 3666 347772
rect 165614 347760 165620 347772
rect 165672 347760 165678 347812
rect 429838 347760 429844 347812
rect 429896 347800 429902 347812
rect 439498 347800 439504 347812
rect 429896 347772 439504 347800
rect 429896 347760 429902 347772
rect 439498 347760 439504 347772
rect 439556 347760 439562 347812
rect 3510 345040 3516 345092
rect 3568 345080 3574 345092
rect 165614 345080 165620 345092
rect 3568 345052 165620 345080
rect 3568 345040 3574 345052
rect 165614 345040 165620 345052
rect 165672 345040 165678 345092
rect 3418 342252 3424 342304
rect 3476 342292 3482 342304
rect 165614 342292 165620 342304
rect 3476 342264 165620 342292
rect 3476 342252 3482 342264
rect 165614 342252 165620 342264
rect 165672 342252 165678 342304
rect 429102 339464 429108 339516
rect 429160 339504 429166 339516
rect 489178 339504 489184 339516
rect 429160 339476 489184 339504
rect 429160 339464 429166 339476
rect 489178 339464 489184 339476
rect 489236 339464 489242 339516
rect 433978 339396 433984 339448
rect 434036 339436 434042 339448
rect 579982 339436 579988 339448
rect 434036 339408 579988 339436
rect 434036 339396 434042 339408
rect 579982 339396 579988 339408
rect 580040 339396 580046 339448
rect 17218 338104 17224 338156
rect 17276 338144 17282 338156
rect 165614 338144 165620 338156
rect 17276 338116 165620 338144
rect 17276 338104 17282 338116
rect 165614 338104 165620 338116
rect 165672 338104 165678 338156
rect 178034 336676 178040 336728
rect 178092 336716 178098 336728
rect 178310 336716 178316 336728
rect 178092 336688 178316 336716
rect 178092 336676 178098 336688
rect 178310 336676 178316 336688
rect 178368 336676 178374 336728
rect 188338 336676 188344 336728
rect 188396 336716 188402 336728
rect 190270 336716 190276 336728
rect 188396 336688 190276 336716
rect 188396 336676 188402 336688
rect 190270 336676 190276 336688
rect 190328 336676 190334 336728
rect 191834 336676 191840 336728
rect 191892 336716 191898 336728
rect 192110 336716 192116 336728
rect 191892 336688 192116 336716
rect 191892 336676 191898 336688
rect 192110 336676 192116 336688
rect 192168 336676 192174 336728
rect 235994 336676 236000 336728
rect 236052 336716 236058 336728
rect 236270 336716 236276 336728
rect 236052 336688 236276 336716
rect 236052 336676 236058 336688
rect 236270 336676 236276 336688
rect 236328 336676 236334 336728
rect 270494 336716 270500 336728
rect 236380 336688 270500 336716
rect 231762 336608 231768 336660
rect 231820 336648 231826 336660
rect 236380 336648 236408 336688
rect 270494 336676 270500 336688
rect 270552 336676 270558 336728
rect 270678 336676 270684 336728
rect 270736 336716 270742 336728
rect 271414 336716 271420 336728
rect 270736 336688 271420 336716
rect 270736 336676 270742 336688
rect 271414 336676 271420 336688
rect 271472 336676 271478 336728
rect 286962 336676 286968 336728
rect 287020 336716 287026 336728
rect 295518 336716 295524 336728
rect 287020 336688 295524 336716
rect 287020 336676 287026 336688
rect 295518 336676 295524 336688
rect 295576 336676 295582 336728
rect 303890 336676 303896 336728
rect 303948 336716 303954 336728
rect 304902 336716 304908 336728
rect 303948 336688 304908 336716
rect 303948 336676 303954 336688
rect 304902 336676 304908 336688
rect 304960 336676 304966 336728
rect 306558 336676 306564 336728
rect 306616 336716 306622 336728
rect 307662 336716 307668 336728
rect 306616 336688 307668 336716
rect 306616 336676 306622 336688
rect 307662 336676 307668 336688
rect 307720 336676 307726 336728
rect 308674 336676 308680 336728
rect 308732 336716 308738 336728
rect 309778 336716 309784 336728
rect 308732 336688 309784 336716
rect 308732 336676 308738 336688
rect 309778 336676 309784 336688
rect 309836 336676 309842 336728
rect 312906 336676 312912 336728
rect 312964 336716 312970 336728
rect 314565 336719 314623 336725
rect 312964 336688 314516 336716
rect 312964 336676 312970 336688
rect 231820 336620 236408 336648
rect 236457 336651 236515 336657
rect 231820 336608 231826 336620
rect 236457 336617 236469 336651
rect 236503 336648 236515 336651
rect 270218 336648 270224 336660
rect 236503 336620 270224 336648
rect 236503 336617 236515 336620
rect 236457 336611 236515 336617
rect 270218 336608 270224 336620
rect 270276 336608 270282 336660
rect 285582 336608 285588 336660
rect 285640 336648 285646 336660
rect 294966 336648 294972 336660
rect 285640 336620 294972 336648
rect 285640 336608 285646 336620
rect 294966 336608 294972 336620
rect 295024 336608 295030 336660
rect 308122 336608 308128 336660
rect 308180 336648 308186 336660
rect 311158 336648 311164 336660
rect 308180 336620 311164 336648
rect 308180 336608 308186 336620
rect 311158 336608 311164 336620
rect 311216 336608 311222 336660
rect 312354 336608 312360 336660
rect 312412 336648 312418 336660
rect 313182 336648 313188 336660
rect 312412 336620 313188 336648
rect 312412 336608 312418 336620
rect 313182 336608 313188 336620
rect 313240 336608 313246 336660
rect 314488 336648 314516 336688
rect 314565 336685 314577 336719
rect 314611 336716 314623 336719
rect 314611 336688 316540 336716
rect 314611 336685 314623 336688
rect 314565 336679 314623 336685
rect 316405 336651 316463 336657
rect 316405 336648 316417 336651
rect 314488 336620 316417 336648
rect 316405 336617 316417 336620
rect 316451 336617 316463 336651
rect 316512 336648 316540 336688
rect 316586 336676 316592 336728
rect 316644 336716 316650 336728
rect 317322 336716 317328 336728
rect 316644 336688 317328 336716
rect 316644 336676 316650 336688
rect 317322 336676 317328 336688
rect 317380 336676 317386 336728
rect 318702 336676 318708 336728
rect 318760 336716 318766 336728
rect 319438 336716 319444 336728
rect 318760 336688 319444 336716
rect 318760 336676 318766 336688
rect 319438 336676 319444 336688
rect 319496 336676 319502 336728
rect 320266 336676 320272 336728
rect 320324 336716 320330 336728
rect 321370 336716 321376 336728
rect 320324 336688 321376 336716
rect 320324 336676 320330 336688
rect 321370 336676 321376 336688
rect 321428 336676 321434 336728
rect 321830 336676 321836 336728
rect 321888 336716 321894 336728
rect 322658 336716 322664 336728
rect 321888 336688 322664 336716
rect 321888 336676 321894 336688
rect 322658 336676 322664 336688
rect 322716 336676 322722 336728
rect 326062 336676 326068 336728
rect 326120 336716 326126 336728
rect 326982 336716 326988 336728
rect 326120 336688 326988 336716
rect 326120 336676 326126 336688
rect 326982 336676 326988 336688
rect 327040 336676 327046 336728
rect 327074 336676 327080 336728
rect 327132 336716 327138 336728
rect 328270 336716 328276 336728
rect 327132 336688 328276 336716
rect 327132 336676 327138 336688
rect 328270 336676 328276 336688
rect 328328 336676 328334 336728
rect 332870 336676 332876 336728
rect 332928 336716 332934 336728
rect 333882 336716 333888 336728
rect 332928 336688 333888 336716
rect 332928 336676 332934 336688
rect 333882 336676 333888 336688
rect 333940 336676 333946 336728
rect 334434 336676 334440 336728
rect 334492 336716 334498 336728
rect 335170 336716 335176 336728
rect 334492 336688 335176 336716
rect 334492 336676 334498 336688
rect 335170 336676 335176 336688
rect 335228 336676 335234 336728
rect 335538 336676 335544 336728
rect 335596 336716 335602 336728
rect 336642 336716 336648 336728
rect 335596 336688 336648 336716
rect 335596 336676 335602 336688
rect 336642 336676 336648 336688
rect 336700 336676 336706 336728
rect 337102 336676 337108 336728
rect 337160 336716 337166 336728
rect 338022 336716 338028 336728
rect 337160 336688 338028 336716
rect 337160 336676 337166 336688
rect 338022 336676 338028 336688
rect 338080 336676 338086 336728
rect 338114 336676 338120 336728
rect 338172 336716 338178 336728
rect 339218 336716 339224 336728
rect 338172 336688 339224 336716
rect 338172 336676 338178 336688
rect 339218 336676 339224 336688
rect 339276 336676 339282 336728
rect 339678 336676 339684 336728
rect 339736 336716 339742 336728
rect 340598 336716 340604 336728
rect 339736 336688 340604 336716
rect 339736 336676 339742 336688
rect 340598 336676 340604 336688
rect 340656 336676 340662 336728
rect 341334 336676 341340 336728
rect 341392 336716 341398 336728
rect 342070 336716 342076 336728
rect 341392 336688 342076 336716
rect 341392 336676 341398 336688
rect 342070 336676 342076 336688
rect 342128 336676 342134 336728
rect 342346 336676 342352 336728
rect 342404 336716 342410 336728
rect 343450 336716 343456 336728
rect 342404 336688 343456 336716
rect 342404 336676 342410 336688
rect 343450 336676 343456 336688
rect 343508 336676 343514 336728
rect 343910 336676 343916 336728
rect 343968 336716 343974 336728
rect 344922 336716 344928 336728
rect 343968 336688 344928 336716
rect 343968 336676 343974 336688
rect 344922 336676 344928 336688
rect 344980 336676 344986 336728
rect 345474 336676 345480 336728
rect 345532 336716 345538 336728
rect 346210 336716 346216 336728
rect 345532 336688 346216 336716
rect 345532 336676 345538 336688
rect 346210 336676 346216 336688
rect 346268 336676 346274 336728
rect 347130 336676 347136 336728
rect 347188 336716 347194 336728
rect 347590 336716 347596 336728
rect 347188 336688 347596 336716
rect 347188 336676 347194 336688
rect 347590 336676 347596 336688
rect 347648 336676 347654 336728
rect 348142 336676 348148 336728
rect 348200 336716 348206 336728
rect 349062 336716 349068 336728
rect 348200 336688 349068 336716
rect 348200 336676 348206 336688
rect 349062 336676 349068 336688
rect 349120 336676 349126 336728
rect 352374 336676 352380 336728
rect 352432 336716 352438 336728
rect 353202 336716 353208 336728
rect 352432 336688 353208 336716
rect 352432 336676 352438 336688
rect 353202 336676 353208 336688
rect 353260 336676 353266 336728
rect 353386 336676 353392 336728
rect 353444 336716 353450 336728
rect 354490 336716 354496 336728
rect 353444 336688 354496 336716
rect 353444 336676 353450 336688
rect 354490 336676 354496 336688
rect 354548 336676 354554 336728
rect 354861 336719 354919 336725
rect 354861 336716 354873 336719
rect 354646 336688 354873 336716
rect 320450 336648 320456 336660
rect 316512 336620 320456 336648
rect 316405 336611 316463 336617
rect 320450 336608 320456 336620
rect 320508 336608 320514 336660
rect 333974 336608 333980 336660
rect 334032 336648 334038 336660
rect 335262 336648 335268 336660
rect 334032 336620 335268 336648
rect 334032 336608 334038 336620
rect 335262 336608 335268 336620
rect 335320 336608 335326 336660
rect 338666 336608 338672 336660
rect 338724 336648 338730 336660
rect 339402 336648 339408 336660
rect 338724 336620 339408 336648
rect 338724 336608 338730 336620
rect 339402 336608 339408 336620
rect 339460 336608 339466 336660
rect 349706 336608 349712 336660
rect 349764 336648 349770 336660
rect 349764 336620 352236 336648
rect 349764 336608 349770 336620
rect 224862 336540 224868 336592
rect 224920 336580 224926 336592
rect 267642 336580 267648 336592
rect 224920 336552 267648 336580
rect 224920 336540 224926 336552
rect 267642 336540 267648 336552
rect 267700 336540 267706 336592
rect 282822 336540 282828 336592
rect 282880 336580 282886 336592
rect 293402 336580 293408 336592
rect 282880 336552 293408 336580
rect 282880 336540 282886 336552
rect 293402 336540 293408 336552
rect 293460 336540 293466 336592
rect 310790 336540 310796 336592
rect 310848 336580 310854 336592
rect 314565 336583 314623 336589
rect 314565 336580 314577 336583
rect 310848 336552 314577 336580
rect 310848 336540 310854 336552
rect 314565 336549 314577 336552
rect 314611 336549 314623 336583
rect 314565 336543 314623 336549
rect 316034 336540 316040 336592
rect 316092 336580 316098 336592
rect 317230 336580 317236 336592
rect 316092 336552 317236 336580
rect 316092 336540 316098 336552
rect 317230 336540 317236 336552
rect 317288 336540 317294 336592
rect 317598 336540 317604 336592
rect 317656 336580 317662 336592
rect 318702 336580 318708 336592
rect 317656 336552 318708 336580
rect 317656 336540 317662 336552
rect 318702 336540 318708 336552
rect 318760 336540 318766 336592
rect 329190 336540 329196 336592
rect 329248 336580 329254 336592
rect 329742 336580 329748 336592
rect 329248 336552 329748 336580
rect 329248 336540 329254 336552
rect 329742 336540 329748 336552
rect 329800 336540 329806 336592
rect 335998 336540 336004 336592
rect 336056 336580 336062 336592
rect 336550 336580 336556 336592
rect 336056 336552 336556 336580
rect 336056 336540 336062 336552
rect 336550 336540 336556 336552
rect 336608 336540 336614 336592
rect 351270 336540 351276 336592
rect 351328 336580 351334 336592
rect 351822 336580 351828 336592
rect 351328 336552 351828 336580
rect 351328 336540 351334 336552
rect 351822 336540 351828 336552
rect 351880 336540 351886 336592
rect 352208 336580 352236 336620
rect 352834 336608 352840 336660
rect 352892 336648 352898 336660
rect 354646 336648 354674 336688
rect 354861 336685 354873 336688
rect 354907 336685 354919 336719
rect 354861 336679 354919 336685
rect 354950 336676 354956 336728
rect 355008 336716 355014 336728
rect 355962 336716 355968 336728
rect 355008 336688 355968 336716
rect 355008 336676 355014 336688
rect 355962 336676 355968 336688
rect 356020 336676 356026 336728
rect 356514 336676 356520 336728
rect 356572 336716 356578 336728
rect 357342 336716 357348 336728
rect 356572 336688 357348 336716
rect 356572 336676 356578 336688
rect 357342 336676 357348 336688
rect 357400 336676 357406 336728
rect 357618 336676 357624 336728
rect 357676 336716 357682 336728
rect 358722 336716 358728 336728
rect 357676 336688 358728 336716
rect 357676 336676 357682 336688
rect 358722 336676 358728 336688
rect 358780 336676 358786 336728
rect 359182 336676 359188 336728
rect 359240 336716 359246 336728
rect 360102 336716 360108 336728
rect 359240 336688 360108 336716
rect 359240 336676 359246 336688
rect 360102 336676 360108 336688
rect 360160 336676 360166 336728
rect 360746 336676 360752 336728
rect 360804 336716 360810 336728
rect 361482 336716 361488 336728
rect 360804 336688 361488 336716
rect 360804 336676 360810 336688
rect 361482 336676 361488 336688
rect 361540 336676 361546 336728
rect 361850 336676 361856 336728
rect 361908 336716 361914 336728
rect 362862 336716 362868 336728
rect 361908 336688 362868 336716
rect 361908 336676 361914 336688
rect 362862 336676 362868 336688
rect 362920 336676 362926 336728
rect 363414 336676 363420 336728
rect 363472 336716 363478 336728
rect 364150 336716 364156 336728
rect 363472 336688 364156 336716
rect 363472 336676 363478 336688
rect 364150 336676 364156 336688
rect 364208 336676 364214 336728
rect 364426 336676 364432 336728
rect 364484 336716 364490 336728
rect 365622 336716 365628 336728
rect 364484 336688 365628 336716
rect 364484 336676 364490 336688
rect 365622 336676 365628 336688
rect 365680 336676 365686 336728
rect 365990 336676 365996 336728
rect 366048 336716 366054 336728
rect 367002 336716 367008 336728
rect 366048 336688 367008 336716
rect 366048 336676 366054 336688
rect 367002 336676 367008 336688
rect 367060 336676 367066 336728
rect 367094 336676 367100 336728
rect 367152 336716 367158 336728
rect 368382 336716 368388 336728
rect 367152 336688 368388 336716
rect 367152 336676 367158 336688
rect 368382 336676 368388 336688
rect 368440 336676 368446 336728
rect 370222 336676 370228 336728
rect 370280 336716 370286 336728
rect 371142 336716 371148 336728
rect 370280 336688 371148 336716
rect 370280 336676 370286 336688
rect 371142 336676 371148 336688
rect 371200 336676 371206 336728
rect 371326 336676 371332 336728
rect 371384 336716 371390 336728
rect 372430 336716 372436 336728
rect 371384 336688 372436 336716
rect 371384 336676 371390 336688
rect 372430 336676 372436 336688
rect 372488 336676 372494 336728
rect 374454 336676 374460 336728
rect 374512 336716 374518 336728
rect 375282 336716 375288 336728
rect 374512 336688 375288 336716
rect 374512 336676 374518 336688
rect 375282 336676 375288 336688
rect 375340 336676 375346 336728
rect 375466 336676 375472 336728
rect 375524 336716 375530 336728
rect 376570 336716 376576 336728
rect 375524 336688 376576 336716
rect 375524 336676 375530 336688
rect 376570 336676 376576 336688
rect 376628 336676 376634 336728
rect 377122 336676 377128 336728
rect 377180 336716 377186 336728
rect 378042 336716 378048 336728
rect 377180 336688 378048 336716
rect 377180 336676 377186 336688
rect 378042 336676 378048 336688
rect 378100 336676 378106 336728
rect 378686 336676 378692 336728
rect 378744 336716 378750 336728
rect 379422 336716 379428 336728
rect 378744 336688 379428 336716
rect 378744 336676 378750 336688
rect 379422 336676 379428 336688
rect 379480 336676 379486 336728
rect 380618 336676 380624 336728
rect 380676 336716 380682 336728
rect 380802 336716 380808 336728
rect 380676 336688 380808 336716
rect 380676 336676 380682 336688
rect 380802 336676 380808 336688
rect 380860 336676 380866 336728
rect 382366 336676 382372 336728
rect 382424 336716 382430 336728
rect 383562 336716 383568 336728
rect 382424 336688 383568 336716
rect 382424 336676 382430 336688
rect 383562 336676 383568 336688
rect 383620 336676 383626 336728
rect 384942 336676 384948 336728
rect 385000 336716 385006 336728
rect 385678 336716 385684 336728
rect 385000 336688 385684 336716
rect 385000 336676 385006 336688
rect 385678 336676 385684 336688
rect 385736 336676 385742 336728
rect 388162 336676 388168 336728
rect 388220 336716 388226 336728
rect 388990 336716 388996 336728
rect 388220 336688 388996 336716
rect 388220 336676 388226 336688
rect 388990 336676 388996 336688
rect 389048 336676 389054 336728
rect 390738 336676 390744 336728
rect 390796 336716 390802 336728
rect 391750 336716 391756 336728
rect 390796 336688 391756 336716
rect 390796 336676 390802 336688
rect 391750 336676 391756 336688
rect 391808 336676 391814 336728
rect 392302 336676 392308 336728
rect 392360 336716 392366 336728
rect 393130 336716 393136 336728
rect 392360 336688 393136 336716
rect 392360 336676 392366 336688
rect 393130 336676 393136 336688
rect 393188 336676 393194 336728
rect 394970 336676 394976 336728
rect 395028 336716 395034 336728
rect 395982 336716 395988 336728
rect 395028 336688 395988 336716
rect 395028 336676 395034 336688
rect 395982 336676 395988 336688
rect 396040 336676 396046 336728
rect 396534 336676 396540 336728
rect 396592 336716 396598 336728
rect 397270 336716 397276 336728
rect 396592 336688 397276 336716
rect 396592 336676 396598 336688
rect 397270 336676 397276 336688
rect 397328 336676 397334 336728
rect 398098 336676 398104 336728
rect 398156 336716 398162 336728
rect 398650 336716 398656 336728
rect 398156 336688 398656 336716
rect 398156 336676 398162 336688
rect 398650 336676 398656 336688
rect 398708 336676 398714 336728
rect 399202 336676 399208 336728
rect 399260 336716 399266 336728
rect 400122 336716 400128 336728
rect 399260 336688 400128 336716
rect 399260 336676 399266 336688
rect 400122 336676 400128 336688
rect 400180 336676 400186 336728
rect 400214 336676 400220 336728
rect 400272 336716 400278 336728
rect 401318 336716 401324 336728
rect 400272 336688 401324 336716
rect 400272 336676 400278 336688
rect 401318 336676 401324 336688
rect 401376 336676 401382 336728
rect 402330 336676 402336 336728
rect 402388 336716 402394 336728
rect 402882 336716 402888 336728
rect 402388 336688 402888 336716
rect 402388 336676 402394 336688
rect 402882 336676 402888 336688
rect 402940 336676 402946 336728
rect 404446 336676 404452 336728
rect 404504 336716 404510 336728
rect 405550 336716 405556 336728
rect 404504 336688 405556 336716
rect 404504 336676 404510 336688
rect 405550 336676 405556 336688
rect 405608 336676 405614 336728
rect 406010 336676 406016 336728
rect 406068 336716 406074 336728
rect 407022 336716 407028 336728
rect 406068 336688 407028 336716
rect 406068 336676 406074 336688
rect 407022 336676 407028 336688
rect 407080 336676 407086 336728
rect 407114 336676 407120 336728
rect 407172 336716 407178 336728
rect 408310 336716 408316 336728
rect 407172 336688 408316 336716
rect 407172 336676 407178 336688
rect 408310 336676 408316 336688
rect 408368 336676 408374 336728
rect 408678 336676 408684 336728
rect 408736 336716 408742 336728
rect 409690 336716 409696 336728
rect 408736 336688 409696 336716
rect 408736 336676 408742 336688
rect 409690 336676 409696 336688
rect 409748 336676 409754 336728
rect 410242 336676 410248 336728
rect 410300 336716 410306 336728
rect 411162 336716 411168 336728
rect 410300 336688 411168 336716
rect 410300 336676 410306 336688
rect 411162 336676 411168 336688
rect 411220 336676 411226 336728
rect 411806 336676 411812 336728
rect 411864 336716 411870 336728
rect 412450 336716 412456 336728
rect 411864 336688 412456 336716
rect 411864 336676 411870 336688
rect 412450 336676 412456 336688
rect 412508 336676 412514 336728
rect 413370 336676 413376 336728
rect 413428 336716 413434 336728
rect 413830 336716 413836 336728
rect 413428 336688 413836 336716
rect 413428 336676 413434 336688
rect 413830 336676 413836 336688
rect 413888 336676 413894 336728
rect 414474 336676 414480 336728
rect 414532 336716 414538 336728
rect 415302 336716 415308 336728
rect 414532 336688 415308 336716
rect 414532 336676 414538 336688
rect 415302 336676 415308 336688
rect 415360 336676 415366 336728
rect 415486 336676 415492 336728
rect 415544 336716 415550 336728
rect 416498 336716 416504 336728
rect 415544 336688 416504 336716
rect 415544 336676 415550 336688
rect 416498 336676 416504 336688
rect 416556 336676 416562 336728
rect 418154 336676 418160 336728
rect 418212 336716 418218 336728
rect 419350 336716 419356 336728
rect 418212 336688 419356 336716
rect 418212 336676 418218 336688
rect 419350 336676 419356 336688
rect 419408 336676 419414 336728
rect 419718 336676 419724 336728
rect 419776 336716 419782 336728
rect 420730 336716 420736 336728
rect 419776 336688 420736 336716
rect 419776 336676 419782 336688
rect 420730 336676 420736 336688
rect 420788 336676 420794 336728
rect 422846 336676 422852 336728
rect 422904 336716 422910 336728
rect 423490 336716 423496 336728
rect 422904 336688 423496 336716
rect 422904 336676 422910 336688
rect 423490 336676 423496 336688
rect 423548 336676 423554 336728
rect 424410 336676 424416 336728
rect 424468 336716 424474 336728
rect 424870 336716 424876 336728
rect 424468 336688 424876 336716
rect 424468 336676 424474 336688
rect 424870 336676 424876 336688
rect 424928 336676 424934 336728
rect 407390 336648 407396 336660
rect 352892 336620 354674 336648
rect 354784 336620 407396 336648
rect 352892 336608 352898 336620
rect 352208 336552 354674 336580
rect 159358 336472 159364 336524
rect 159416 336512 159422 336524
rect 203978 336512 203984 336524
rect 159416 336484 203984 336512
rect 159416 336472 159422 336484
rect 203978 336472 203984 336484
rect 204036 336472 204042 336524
rect 227622 336472 227628 336524
rect 227680 336512 227686 336524
rect 268654 336512 268660 336524
rect 227680 336484 268660 336512
rect 227680 336472 227686 336484
rect 268654 336472 268660 336484
rect 268712 336472 268718 336524
rect 280890 336472 280896 336524
rect 280948 336512 280954 336524
rect 291470 336512 291476 336524
rect 280948 336484 291476 336512
rect 280948 336472 280954 336484
rect 291470 336472 291476 336484
rect 291528 336472 291534 336524
rect 311802 336472 311808 336524
rect 311860 336512 311866 336524
rect 323118 336512 323124 336524
rect 311860 336484 323124 336512
rect 311860 336472 311866 336484
rect 323118 336472 323124 336484
rect 323176 336472 323182 336524
rect 354646 336512 354674 336552
rect 354784 336512 354812 336620
rect 407390 336608 407396 336620
rect 407448 336608 407454 336660
rect 416038 336608 416044 336660
rect 416096 336648 416102 336660
rect 416682 336648 416688 336660
rect 416096 336620 416688 336648
rect 416096 336608 416102 336620
rect 416682 336608 416688 336620
rect 416740 336608 416746 336660
rect 417050 336608 417056 336660
rect 417108 336648 417114 336660
rect 417970 336648 417976 336660
rect 417108 336620 417976 336648
rect 417108 336608 417114 336620
rect 417970 336608 417976 336620
rect 418028 336608 418034 336660
rect 421282 336608 421288 336660
rect 421340 336648 421346 336660
rect 422202 336648 422208 336660
rect 421340 336620 422208 336648
rect 421340 336608 421346 336620
rect 422202 336608 422208 336620
rect 422260 336608 422266 336660
rect 422386 336608 422392 336660
rect 422444 336648 422450 336660
rect 423582 336648 423588 336660
rect 422444 336620 423588 336648
rect 422444 336608 422450 336620
rect 423582 336608 423588 336620
rect 423640 336608 423646 336660
rect 354861 336583 354919 336589
rect 354861 336549 354873 336583
rect 354907 336580 354919 336583
rect 415670 336580 415676 336592
rect 354907 336552 415676 336580
rect 354907 336549 354919 336552
rect 354861 336543 354919 336549
rect 415670 336540 415676 336552
rect 415728 336540 415734 336592
rect 426526 336540 426532 336592
rect 426584 336580 426590 336592
rect 427538 336580 427544 336592
rect 426584 336552 427544 336580
rect 426584 336540 426590 336552
rect 427538 336540 427544 336552
rect 427596 336540 427602 336592
rect 422570 336512 422576 336524
rect 354646 336484 354812 336512
rect 360212 336484 422576 336512
rect 125502 336404 125508 336456
rect 125560 336444 125566 336456
rect 223390 336444 223396 336456
rect 125560 336416 223396 336444
rect 125560 336404 125566 336416
rect 223390 336404 223396 336416
rect 223448 336404 223454 336456
rect 223482 336404 223488 336456
rect 223540 336444 223546 336456
rect 267090 336444 267096 336456
rect 223540 336416 267096 336444
rect 223540 336404 223546 336416
rect 267090 336404 267096 336416
rect 267148 336404 267154 336456
rect 278038 336404 278044 336456
rect 278096 336444 278102 336456
rect 290274 336444 290280 336456
rect 278096 336416 290280 336444
rect 278096 336404 278102 336416
rect 290274 336404 290280 336416
rect 290332 336404 290338 336456
rect 313366 336404 313372 336456
rect 313424 336444 313430 336456
rect 318058 336444 318064 336456
rect 313424 336416 318064 336444
rect 313424 336404 313430 336416
rect 318058 336404 318064 336416
rect 318116 336404 318122 336456
rect 319162 336404 319168 336456
rect 319220 336444 319226 336456
rect 320082 336444 320088 336456
rect 319220 336416 320088 336444
rect 319220 336404 319226 336416
rect 320082 336404 320088 336416
rect 320140 336404 320146 336456
rect 356054 336404 356060 336456
rect 356112 336444 356118 336456
rect 360212 336444 360240 336484
rect 422570 336472 422576 336484
rect 422628 336472 422634 336524
rect 356112 336416 360240 336444
rect 356112 336404 356118 336416
rect 362310 336404 362316 336456
rect 362368 336444 362374 336456
rect 436094 336444 436100 336456
rect 362368 336416 436100 336444
rect 362368 336404 362374 336416
rect 436094 336404 436100 336416
rect 436152 336404 436158 336456
rect 114462 336336 114468 336388
rect 114520 336376 114526 336388
rect 218698 336376 218704 336388
rect 114520 336348 218704 336376
rect 114520 336336 114526 336348
rect 218698 336336 218704 336348
rect 218756 336336 218762 336388
rect 220722 336336 220728 336388
rect 220780 336376 220786 336388
rect 266078 336376 266084 336388
rect 220780 336348 266084 336376
rect 220780 336336 220786 336348
rect 266078 336336 266084 336348
rect 266136 336336 266142 336388
rect 281442 336336 281448 336388
rect 281500 336376 281506 336388
rect 292850 336376 292856 336388
rect 281500 336348 292856 336376
rect 281500 336336 281506 336348
rect 292850 336336 292856 336348
rect 292908 336336 292914 336388
rect 294598 336336 294604 336388
rect 294656 336376 294662 336388
rect 298646 336376 298652 336388
rect 294656 336348 298652 336376
rect 294656 336336 294662 336348
rect 298646 336336 298652 336348
rect 298704 336336 298710 336388
rect 306006 336336 306012 336388
rect 306064 336376 306070 336388
rect 309318 336376 309324 336388
rect 306064 336348 309324 336376
rect 306064 336336 306070 336348
rect 309318 336336 309324 336348
rect 309376 336336 309382 336388
rect 310238 336336 310244 336388
rect 310296 336376 310302 336388
rect 313918 336376 313924 336388
rect 310296 336348 313924 336376
rect 310296 336336 310302 336348
rect 313918 336336 313924 336348
rect 313976 336336 313982 336388
rect 316405 336379 316463 336385
rect 316405 336345 316417 336379
rect 316451 336376 316463 336379
rect 324406 336376 324412 336388
rect 316451 336348 324412 336376
rect 316451 336345 316463 336348
rect 316405 336339 316463 336345
rect 324406 336336 324412 336348
rect 324464 336336 324470 336388
rect 369210 336336 369216 336388
rect 369268 336376 369274 336388
rect 370498 336376 370504 336388
rect 369268 336348 370504 336376
rect 369268 336336 369274 336348
rect 370498 336336 370504 336348
rect 370556 336336 370562 336388
rect 442994 336376 443000 336388
rect 370608 336348 443000 336376
rect 35158 336268 35164 336320
rect 35216 336308 35222 336320
rect 180794 336308 180800 336320
rect 35216 336280 180800 336308
rect 35216 336268 35222 336280
rect 180794 336268 180800 336280
rect 180852 336268 180858 336320
rect 217962 336268 217968 336320
rect 218020 336308 218026 336320
rect 264422 336308 264428 336320
rect 218020 336280 264428 336308
rect 218020 336268 218026 336280
rect 264422 336268 264428 336280
rect 264480 336268 264486 336320
rect 277210 336268 277216 336320
rect 277268 336308 277274 336320
rect 290734 336308 290740 336320
rect 277268 336280 290740 336308
rect 277268 336268 277274 336280
rect 290734 336268 290740 336280
rect 290792 336268 290798 336320
rect 311342 336268 311348 336320
rect 311400 336308 311406 336320
rect 321830 336308 321836 336320
rect 311400 336280 321836 336308
rect 311400 336268 311406 336280
rect 321830 336268 321836 336280
rect 321888 336268 321894 336320
rect 330202 336268 330208 336320
rect 330260 336308 330266 336320
rect 352558 336308 352564 336320
rect 330260 336280 352564 336308
rect 330260 336268 330266 336280
rect 352558 336268 352564 336280
rect 352616 336268 352622 336320
rect 29638 336200 29644 336252
rect 29696 336240 29702 336252
rect 176562 336240 176568 336252
rect 29696 336212 176568 336240
rect 29696 336200 29702 336212
rect 176562 336200 176568 336212
rect 176620 336200 176626 336252
rect 219250 336200 219256 336252
rect 219308 336240 219314 336252
rect 265526 336240 265532 336252
rect 219308 336212 265532 336240
rect 219308 336200 219314 336212
rect 265526 336200 265532 336212
rect 265584 336200 265590 336252
rect 277302 336200 277308 336252
rect 277360 336240 277366 336252
rect 291286 336240 291292 336252
rect 277360 336212 291292 336240
rect 277360 336200 277366 336212
rect 291286 336200 291292 336212
rect 291344 336200 291350 336252
rect 307570 336200 307576 336252
rect 307628 336240 307634 336252
rect 313366 336240 313372 336252
rect 307628 336212 313372 336240
rect 307628 336200 307634 336212
rect 313366 336200 313372 336212
rect 313424 336200 313430 336252
rect 314470 336200 314476 336252
rect 314528 336240 314534 336252
rect 327718 336240 327724 336252
rect 314528 336212 327724 336240
rect 314528 336200 314534 336212
rect 327718 336200 327724 336212
rect 327776 336200 327782 336252
rect 328638 336200 328644 336252
rect 328696 336240 328702 336252
rect 349798 336240 349804 336252
rect 328696 336212 349804 336240
rect 328696 336200 328702 336212
rect 349798 336200 349804 336212
rect 349856 336200 349862 336252
rect 365530 336200 365536 336252
rect 365588 336240 365594 336252
rect 370608 336240 370636 336348
rect 442994 336336 443000 336348
rect 443052 336336 443058 336388
rect 449894 336308 449900 336320
rect 365588 336212 370636 336240
rect 371344 336280 449900 336308
rect 365588 336200 365594 336212
rect 28258 336132 28264 336184
rect 28316 336172 28322 336184
rect 177114 336172 177120 336184
rect 28316 336144 177120 336172
rect 28316 336132 28322 336144
rect 177114 336132 177120 336144
rect 177172 336132 177178 336184
rect 213822 336132 213828 336184
rect 213880 336172 213886 336184
rect 262858 336172 262864 336184
rect 213880 336144 262864 336172
rect 213880 336132 213886 336144
rect 262858 336132 262864 336144
rect 262916 336132 262922 336184
rect 271782 336132 271788 336184
rect 271840 336172 271846 336184
rect 288710 336172 288716 336184
rect 271840 336144 288716 336172
rect 271840 336132 271846 336144
rect 288710 336132 288716 336144
rect 288768 336132 288774 336184
rect 292482 336132 292488 336184
rect 292540 336172 292546 336184
rect 297634 336172 297640 336184
rect 292540 336144 297640 336172
rect 292540 336132 292546 336144
rect 297634 336132 297640 336144
rect 297692 336132 297698 336184
rect 304994 336132 305000 336184
rect 305052 336172 305058 336184
rect 306190 336172 306196 336184
rect 305052 336144 306196 336172
rect 305052 336132 305058 336144
rect 306190 336132 306196 336144
rect 306248 336132 306254 336184
rect 319714 336132 319720 336184
rect 319772 336172 319778 336184
rect 341058 336172 341064 336184
rect 319772 336144 341064 336172
rect 319772 336132 319778 336144
rect 341058 336132 341064 336144
rect 341116 336132 341122 336184
rect 344462 336132 344468 336184
rect 344520 336172 344526 336184
rect 358078 336172 358084 336184
rect 344520 336144 358084 336172
rect 344520 336132 344526 336144
rect 358078 336132 358084 336144
rect 358136 336132 358142 336184
rect 368658 336132 368664 336184
rect 368716 336172 368722 336184
rect 371344 336172 371372 336280
rect 449894 336268 449900 336280
rect 449952 336268 449958 336320
rect 371786 336200 371792 336252
rect 371844 336240 371850 336252
rect 456794 336240 456800 336252
rect 371844 336212 456800 336240
rect 371844 336200 371850 336212
rect 456794 336200 456800 336212
rect 456852 336200 456858 336252
rect 368716 336144 371372 336172
rect 368716 336132 368722 336144
rect 379698 336132 379704 336184
rect 379756 336172 379762 336184
rect 380802 336172 380808 336184
rect 379756 336144 380808 336172
rect 379756 336132 379762 336144
rect 380802 336132 380808 336144
rect 380860 336132 380866 336184
rect 380897 336175 380955 336181
rect 380897 336141 380909 336175
rect 380943 336172 380955 336175
rect 465074 336172 465080 336184
rect 380943 336144 465080 336172
rect 380943 336141 380955 336144
rect 380897 336135 380955 336141
rect 465074 336132 465080 336144
rect 465132 336132 465138 336184
rect 18598 336064 18604 336116
rect 18656 336104 18662 336116
rect 172882 336104 172888 336116
rect 18656 336076 172888 336104
rect 18656 336064 18662 336076
rect 172882 336064 172888 336076
rect 172940 336064 172946 336116
rect 191098 336064 191104 336116
rect 191156 336104 191162 336116
rect 216214 336104 216220 336116
rect 191156 336076 216220 336104
rect 191156 336064 191162 336076
rect 216214 336064 216220 336076
rect 216272 336064 216278 336116
rect 216582 336064 216588 336116
rect 216640 336104 216646 336116
rect 263962 336104 263968 336116
rect 216640 336076 263968 336104
rect 216640 336064 216646 336076
rect 263962 336064 263968 336076
rect 264020 336064 264026 336116
rect 269022 336064 269028 336116
rect 269080 336104 269086 336116
rect 287054 336104 287060 336116
rect 269080 336076 287060 336104
rect 269080 336064 269086 336076
rect 287054 336064 287060 336076
rect 287112 336064 287118 336116
rect 289722 336064 289728 336116
rect 289780 336104 289786 336116
rect 296530 336104 296536 336116
rect 289780 336076 296536 336104
rect 289780 336064 289786 336076
rect 296530 336064 296536 336076
rect 296588 336064 296594 336116
rect 296622 336064 296628 336116
rect 296680 336104 296686 336116
rect 299750 336104 299756 336116
rect 296680 336076 299756 336104
rect 296680 336064 296686 336076
rect 299750 336064 299756 336076
rect 299808 336064 299814 336116
rect 315022 336064 315028 336116
rect 315080 336104 315086 336116
rect 330018 336104 330024 336116
rect 315080 336076 330024 336104
rect 315080 336064 315086 336076
rect 330018 336064 330024 336076
rect 330076 336064 330082 336116
rect 349154 336064 349160 336116
rect 349212 336104 349218 336116
rect 350350 336104 350356 336116
rect 349212 336076 350356 336104
rect 349212 336064 349218 336076
rect 350350 336064 350356 336076
rect 350408 336064 350414 336116
rect 378134 336064 378140 336116
rect 378192 336104 378198 336116
rect 471974 336104 471980 336116
rect 378192 336076 471980 336104
rect 378192 336064 378198 336076
rect 471974 336064 471980 336076
rect 472032 336064 472038 336116
rect 10318 335996 10324 336048
rect 10376 336036 10382 336048
rect 170214 336036 170220 336048
rect 10376 336008 170220 336036
rect 10376 335996 10382 336008
rect 170214 335996 170220 336008
rect 170272 335996 170278 336048
rect 212442 335996 212448 336048
rect 212500 336036 212506 336048
rect 262306 336036 262312 336048
rect 212500 336008 262312 336036
rect 212500 335996 212506 336008
rect 262306 335996 262312 336008
rect 262364 335996 262370 336048
rect 264882 335996 264888 336048
rect 264940 336036 264946 336048
rect 285214 336036 285220 336048
rect 264940 336008 285220 336036
rect 264940 335996 264946 336008
rect 285214 335996 285220 336008
rect 285272 335996 285278 336048
rect 285490 335996 285496 336048
rect 285548 336036 285554 336048
rect 294414 336036 294420 336048
rect 285548 336008 294420 336036
rect 285548 335996 285554 336008
rect 294414 335996 294420 336008
rect 294472 335996 294478 336048
rect 326522 335996 326528 336048
rect 326580 336036 326586 336048
rect 326580 336008 335354 336036
rect 326580 335996 326586 336008
rect 230382 335928 230388 335980
rect 230440 335968 230446 335980
rect 236457 335971 236515 335977
rect 236457 335968 236469 335971
rect 230440 335940 236469 335968
rect 230440 335928 230446 335940
rect 236457 335937 236469 335940
rect 236503 335937 236515 335971
rect 236457 335931 236515 335937
rect 242802 335928 242808 335980
rect 242860 335968 242866 335980
rect 275554 335968 275560 335980
rect 242860 335940 275560 335968
rect 242860 335928 242866 335940
rect 275554 335928 275560 335940
rect 275612 335928 275618 335980
rect 309686 335928 309692 335980
rect 309744 335968 309750 335980
rect 317506 335968 317512 335980
rect 309744 335940 317512 335968
rect 309744 335928 309750 335940
rect 317506 335928 317512 335940
rect 317564 335928 317570 335980
rect 324498 335928 324504 335980
rect 324556 335968 324562 335980
rect 325418 335968 325424 335980
rect 324556 335940 325424 335968
rect 324556 335928 324562 335940
rect 325418 335928 325424 335940
rect 325476 335928 325482 335980
rect 335326 335968 335354 336008
rect 358170 335996 358176 336048
rect 358228 336036 358234 336048
rect 374638 336036 374644 336048
rect 358228 336008 374644 336036
rect 358228 335996 358234 336008
rect 374638 335996 374644 336008
rect 374696 335996 374702 336048
rect 375006 335996 375012 336048
rect 375064 336036 375070 336048
rect 380897 336039 380955 336045
rect 380897 336036 380909 336039
rect 375064 336008 380909 336036
rect 375064 335996 375070 336008
rect 380897 336005 380909 336008
rect 380943 336005 380955 336039
rect 380897 335999 380955 336005
rect 381262 335996 381268 336048
rect 381320 336036 381326 336048
rect 478874 336036 478880 336048
rect 381320 336008 478880 336036
rect 381320 335996 381326 336008
rect 478874 335996 478880 336008
rect 478932 335996 478938 336048
rect 356146 335968 356152 335980
rect 335326 335940 356152 335968
rect 356146 335928 356152 335940
rect 356204 335928 356210 335980
rect 385494 335928 385500 335980
rect 385552 335968 385558 335980
rect 386322 335968 386328 335980
rect 385552 335940 386328 335968
rect 385552 335928 385558 335940
rect 386322 335928 386328 335940
rect 386380 335928 386386 335980
rect 389174 335928 389180 335980
rect 389232 335968 389238 335980
rect 390278 335968 390284 335980
rect 389232 335940 390284 335968
rect 389232 335928 389238 335940
rect 390278 335928 390284 335940
rect 390336 335928 390342 335980
rect 393406 335928 393412 335980
rect 393464 335968 393470 335980
rect 394418 335968 394424 335980
rect 393464 335940 394424 335968
rect 393464 335928 393470 335940
rect 394418 335928 394424 335940
rect 394476 335928 394482 335980
rect 396074 335928 396080 335980
rect 396132 335968 396138 335980
rect 397362 335968 397368 335980
rect 396132 335940 397368 335968
rect 396132 335928 396138 335940
rect 397362 335928 397368 335940
rect 397420 335928 397426 335980
rect 397638 335928 397644 335980
rect 397696 335968 397702 335980
rect 398742 335968 398748 335980
rect 397696 335940 398748 335968
rect 397696 335928 397702 335940
rect 398742 335928 398748 335940
rect 398800 335928 398806 335980
rect 400766 335928 400772 335980
rect 400824 335968 400830 335980
rect 401502 335968 401508 335980
rect 400824 335940 401508 335968
rect 400824 335928 400830 335940
rect 401502 335928 401508 335940
rect 401560 335928 401566 335980
rect 240778 335860 240784 335912
rect 240836 335900 240842 335912
rect 243446 335900 243452 335912
rect 240836 335872 243452 335900
rect 240836 335860 240842 335872
rect 243446 335860 243452 335872
rect 243504 335860 243510 335912
rect 251082 335860 251088 335912
rect 251140 335900 251146 335912
rect 279234 335900 279240 335912
rect 251140 335872 279240 335900
rect 251140 335860 251146 335872
rect 279234 335860 279240 335872
rect 279292 335860 279298 335912
rect 345014 335860 345020 335912
rect 345072 335900 345078 335912
rect 346302 335900 346308 335912
rect 345072 335872 346308 335900
rect 345072 335860 345078 335872
rect 346302 335860 346308 335872
rect 346360 335860 346366 335912
rect 253842 335792 253848 335844
rect 253900 335832 253906 335844
rect 280798 335832 280804 335844
rect 253900 335804 280804 335832
rect 253900 335792 253906 335804
rect 280798 335792 280804 335804
rect 280856 335792 280862 335844
rect 259362 335724 259368 335776
rect 259420 335764 259426 335776
rect 282914 335764 282920 335776
rect 259420 335736 282920 335764
rect 259420 335724 259426 335736
rect 282914 335724 282920 335736
rect 282972 335724 282978 335776
rect 331306 335724 331312 335776
rect 331364 335764 331370 335776
rect 332410 335764 332416 335776
rect 331364 335736 332416 335764
rect 331364 335724 331370 335736
rect 332410 335724 332416 335736
rect 332468 335724 332474 335776
rect 210510 335656 210516 335708
rect 210568 335696 210574 335708
rect 211798 335696 211804 335708
rect 210568 335668 211804 335696
rect 210568 335656 210574 335668
rect 211798 335656 211804 335668
rect 211856 335656 211862 335708
rect 304442 335656 304448 335708
rect 304500 335696 304506 335708
rect 306650 335696 306656 335708
rect 304500 335668 306656 335696
rect 304500 335656 304506 335668
rect 306650 335656 306656 335668
rect 306708 335656 306714 335708
rect 340230 335656 340236 335708
rect 340288 335696 340294 335708
rect 340782 335696 340788 335708
rect 340288 335668 340788 335696
rect 340288 335656 340294 335668
rect 340782 335656 340788 335668
rect 340840 335656 340846 335708
rect 260742 335588 260748 335640
rect 260800 335628 260806 335640
rect 283926 335628 283932 335640
rect 260800 335600 283932 335628
rect 260800 335588 260806 335600
rect 283926 335588 283932 335600
rect 283984 335588 283990 335640
rect 291838 335588 291844 335640
rect 291896 335628 291902 335640
rect 297082 335628 297088 335640
rect 291896 335600 297088 335628
rect 291896 335588 291902 335600
rect 297082 335588 297088 335600
rect 297140 335588 297146 335640
rect 299382 335588 299388 335640
rect 299440 335628 299446 335640
rect 300762 335628 300768 335640
rect 299440 335600 300768 335628
rect 299440 335588 299446 335600
rect 300762 335588 300768 335600
rect 300820 335588 300826 335640
rect 360286 335588 360292 335640
rect 360344 335628 360350 335640
rect 361390 335628 361396 335640
rect 360344 335600 361396 335628
rect 360344 335588 360350 335600
rect 361390 335588 361396 335600
rect 361448 335588 361454 335640
rect 309226 335520 309232 335572
rect 309284 335560 309290 335572
rect 310422 335560 310428 335572
rect 309284 335532 310428 335560
rect 309284 335520 309290 335532
rect 310422 335520 310428 335532
rect 310480 335520 310486 335572
rect 346578 335520 346584 335572
rect 346636 335560 346642 335572
rect 347682 335560 347688 335572
rect 346636 335532 347688 335560
rect 346636 335520 346642 335532
rect 347682 335520 347688 335532
rect 347740 335520 347746 335572
rect 411254 335520 411260 335572
rect 411312 335560 411318 335572
rect 412542 335560 412548 335572
rect 411312 335532 412548 335560
rect 411312 335520 411318 335532
rect 412542 335520 412548 335532
rect 412600 335520 412606 335572
rect 307110 335452 307116 335504
rect 307168 335492 307174 335504
rect 312078 335492 312084 335504
rect 307168 335464 312084 335492
rect 307168 335452 307174 335464
rect 312078 335452 312084 335464
rect 312136 335452 312142 335504
rect 283558 335316 283564 335368
rect 283616 335356 283622 335368
rect 289170 335356 289176 335368
rect 283616 335328 289176 335356
rect 283616 335316 283622 335328
rect 289170 335316 289176 335328
rect 289228 335316 289234 335368
rect 383930 335316 383936 335368
rect 383988 335356 383994 335368
rect 383988 335328 384896 335356
rect 383988 335316 383994 335328
rect 384868 335220 384896 335328
rect 412910 335316 412916 335368
rect 412968 335356 412974 335368
rect 412968 335328 413692 335356
rect 412968 335316 412974 335328
rect 384942 335220 384948 335232
rect 384868 335192 384948 335220
rect 384942 335180 384948 335192
rect 385000 335180 385006 335232
rect 413664 335220 413692 335328
rect 423950 335316 423956 335368
rect 424008 335356 424014 335368
rect 424008 335328 424732 335356
rect 424008 335316 424014 335328
rect 413922 335220 413928 335232
rect 413664 335192 413928 335220
rect 413922 335180 413928 335192
rect 413980 335180 413986 335232
rect 424704 335220 424732 335328
rect 424962 335220 424968 335232
rect 424704 335192 424968 335220
rect 424962 335180 424968 335192
rect 425020 335180 425026 335232
rect 126882 334636 126888 334688
rect 126940 334676 126946 334688
rect 223942 334676 223948 334688
rect 126940 334648 223948 334676
rect 126940 334636 126946 334648
rect 223942 334636 223948 334648
rect 224000 334636 224006 334688
rect 386598 334636 386604 334688
rect 386656 334676 386662 334688
rect 489914 334676 489920 334688
rect 386656 334648 489920 334676
rect 386656 334636 386662 334648
rect 489914 334636 489920 334648
rect 489972 334636 489978 334688
rect 39298 334568 39304 334620
rect 39356 334608 39362 334620
rect 183370 334608 183376 334620
rect 39356 334580 183376 334608
rect 39356 334568 39362 334580
rect 183370 334568 183376 334580
rect 183428 334568 183434 334620
rect 202782 334568 202788 334620
rect 202840 334608 202846 334620
rect 258166 334608 258172 334620
rect 202840 334580 258172 334608
rect 202840 334568 202846 334580
rect 258166 334568 258172 334580
rect 258224 334568 258230 334620
rect 324958 334568 324964 334620
rect 325016 334608 325022 334620
rect 351914 334608 351920 334620
rect 325016 334580 351920 334608
rect 325016 334568 325022 334580
rect 351914 334568 351920 334580
rect 351972 334568 351978 334620
rect 404998 334568 405004 334620
rect 405056 334608 405062 334620
rect 531314 334608 531320 334620
rect 405056 334580 531320 334608
rect 405056 334568 405062 334580
rect 531314 334568 531320 334580
rect 531372 334568 531378 334620
rect 206922 333344 206928 333396
rect 206980 333384 206986 333396
rect 259730 333384 259736 333396
rect 206980 333356 259736 333384
rect 206980 333344 206986 333356
rect 259730 333344 259736 333356
rect 259788 333344 259794 333396
rect 161382 333276 161388 333328
rect 161440 333316 161446 333328
rect 161440 333288 219434 333316
rect 161440 333276 161446 333288
rect 95142 333208 95148 333260
rect 95200 333248 95206 333260
rect 95200 333220 200114 333248
rect 95200 333208 95206 333220
rect 200086 333180 200114 333220
rect 210234 333180 210240 333192
rect 200086 333152 210240 333180
rect 210234 333140 210240 333152
rect 210292 333140 210298 333192
rect 219406 333180 219434 333288
rect 372890 333276 372896 333328
rect 372948 333316 372954 333328
rect 459554 333316 459560 333328
rect 372948 333288 459560 333316
rect 372948 333276 372954 333288
rect 459554 333276 459560 333288
rect 459612 333276 459618 333328
rect 328178 333208 328184 333260
rect 328236 333248 328242 333260
rect 358814 333248 358820 333260
rect 328236 333220 358820 333248
rect 328236 333208 328242 333220
rect 358814 333208 358820 333220
rect 358872 333208 358878 333260
rect 394602 333208 394608 333260
rect 394660 333248 394666 333260
rect 507854 333248 507860 333260
rect 394660 333220 507860 333248
rect 394660 333208 394666 333220
rect 507854 333208 507860 333220
rect 507912 333208 507918 333260
rect 239766 333180 239772 333192
rect 219406 333152 239772 333180
rect 239766 333140 239772 333152
rect 239824 333140 239830 333192
rect 3050 332528 3056 332580
rect 3108 332568 3114 332580
rect 166902 332568 166908 332580
rect 3108 332540 166908 332568
rect 3108 332528 3114 332540
rect 166902 332528 166908 332540
rect 166960 332528 166966 332580
rect 195882 331916 195888 331968
rect 195940 331956 195946 331968
rect 254946 331956 254952 331968
rect 195940 331928 254952 331956
rect 195940 331916 195946 331928
rect 254946 331916 254952 331928
rect 255004 331916 255010 331968
rect 383378 331916 383384 331968
rect 383436 331956 383442 331968
rect 483014 331956 483020 331968
rect 383436 331928 483020 331956
rect 383436 331916 383442 331928
rect 483014 331916 483020 331928
rect 483072 331916 483078 331968
rect 140682 331848 140688 331900
rect 140740 331888 140746 331900
rect 230290 331888 230296 331900
rect 140740 331860 230296 331888
rect 140740 331848 140746 331860
rect 230290 331848 230296 331860
rect 230348 331848 230354 331900
rect 401778 331848 401784 331900
rect 401836 331888 401842 331900
rect 524414 331888 524420 331900
rect 401836 331860 524420 331888
rect 401836 331848 401842 331860
rect 524414 331848 524420 331860
rect 524472 331848 524478 331900
rect 193398 331168 193404 331220
rect 193456 331208 193462 331220
rect 193582 331208 193588 331220
rect 193456 331180 193588 331208
rect 193456 331168 193462 331180
rect 193582 331168 193588 331180
rect 193640 331168 193646 331220
rect 214190 331168 214196 331220
rect 214248 331208 214254 331220
rect 214374 331208 214380 331220
rect 214248 331180 214380 331208
rect 214248 331168 214254 331180
rect 214374 331168 214380 331180
rect 214432 331168 214438 331220
rect 232038 331168 232044 331220
rect 232096 331208 232102 331220
rect 232222 331208 232228 331220
rect 232096 331180 232228 331208
rect 232096 331168 232102 331180
rect 232222 331168 232228 331180
rect 232280 331168 232286 331220
rect 276198 330760 276204 330812
rect 276256 330760 276262 330812
rect 276216 330608 276244 330760
rect 165522 330556 165528 330608
rect 165580 330596 165586 330608
rect 241330 330596 241336 330608
rect 165580 330568 241336 330596
rect 165580 330556 165586 330568
rect 241330 330556 241336 330568
rect 241388 330556 241394 330608
rect 276198 330556 276204 330608
rect 276256 330556 276262 330608
rect 350810 330556 350816 330608
rect 350868 330596 350874 330608
rect 409874 330596 409880 330608
rect 350868 330568 409880 330596
rect 350868 330556 350874 330568
rect 409874 330556 409880 330568
rect 409932 330556 409938 330608
rect 21358 330488 21364 330540
rect 21416 330528 21422 330540
rect 173894 330528 173900 330540
rect 21416 330500 173900 330528
rect 21416 330488 21422 330500
rect 173894 330488 173900 330500
rect 173952 330488 173958 330540
rect 175366 330488 175372 330540
rect 175424 330528 175430 330540
rect 175642 330528 175648 330540
rect 175424 330500 175648 330528
rect 175424 330488 175430 330500
rect 175642 330488 175648 330500
rect 175700 330488 175706 330540
rect 197354 330488 197360 330540
rect 197412 330528 197418 330540
rect 198366 330528 198372 330540
rect 197412 330500 198372 330528
rect 197412 330488 197418 330500
rect 198366 330488 198372 330500
rect 198424 330488 198430 330540
rect 200114 330488 200120 330540
rect 200172 330528 200178 330540
rect 200942 330528 200948 330540
rect 200172 330500 200948 330528
rect 200172 330488 200178 330500
rect 200942 330488 200948 330500
rect 201000 330488 201006 330540
rect 202966 330488 202972 330540
rect 203024 330528 203030 330540
rect 203150 330528 203156 330540
rect 203024 330500 203156 330528
rect 203024 330488 203030 330500
rect 203150 330488 203156 330500
rect 203208 330488 203214 330540
rect 269206 330488 269212 330540
rect 269264 330528 269270 330540
rect 269390 330528 269396 330540
rect 269264 330500 269396 330528
rect 269264 330488 269270 330500
rect 269390 330488 269396 330500
rect 269448 330488 269454 330540
rect 270586 330488 270592 330540
rect 270644 330528 270650 330540
rect 271046 330528 271052 330540
rect 270644 330500 271052 330528
rect 270644 330488 270650 330500
rect 271046 330488 271052 330500
rect 271104 330488 271110 330540
rect 276106 330488 276112 330540
rect 276164 330528 276170 330540
rect 276750 330528 276756 330540
rect 276164 330500 276756 330528
rect 276164 330488 276170 330500
rect 276750 330488 276756 330500
rect 276808 330488 276814 330540
rect 277394 330488 277400 330540
rect 277452 330528 277458 330540
rect 278406 330528 278412 330540
rect 277452 330500 278412 330528
rect 277452 330488 277458 330500
rect 278406 330488 278412 330500
rect 278464 330488 278470 330540
rect 280246 330488 280252 330540
rect 280304 330528 280310 330540
rect 280982 330528 280988 330540
rect 280304 330500 280988 330528
rect 280304 330488 280310 330500
rect 280982 330488 280988 330500
rect 281040 330488 281046 330540
rect 281626 330488 281632 330540
rect 281684 330528 281690 330540
rect 282086 330528 282092 330540
rect 281684 330500 282092 330528
rect 281684 330488 281690 330500
rect 282086 330488 282092 330500
rect 282144 330488 282150 330540
rect 284478 330488 284484 330540
rect 284536 330528 284542 330540
rect 284662 330528 284668 330540
rect 284536 330500 284668 330528
rect 284536 330488 284542 330500
rect 284662 330488 284668 330500
rect 284720 330488 284726 330540
rect 300854 330488 300860 330540
rect 300912 330528 300918 330540
rect 301590 330528 301596 330540
rect 300912 330500 301596 330528
rect 300912 330488 300918 330500
rect 301590 330488 301596 330500
rect 301648 330488 301654 330540
rect 391290 330488 391296 330540
rect 391348 330528 391354 330540
rect 500954 330528 500960 330540
rect 391348 330500 500960 330528
rect 391348 330488 391354 330500
rect 500954 330488 500960 330500
rect 501012 330488 501018 330540
rect 168374 330420 168380 330472
rect 168432 330460 168438 330472
rect 168926 330460 168932 330472
rect 168432 330432 168932 330460
rect 168432 330420 168438 330432
rect 168926 330420 168932 330432
rect 168984 330420 168990 330472
rect 195974 329536 195980 329588
rect 196032 329576 196038 329588
rect 196710 329576 196716 329588
rect 196032 329548 196716 329576
rect 196032 329536 196038 329548
rect 196710 329536 196716 329548
rect 196768 329536 196774 329588
rect 129642 329128 129648 329180
rect 129700 329168 129706 329180
rect 225506 329168 225512 329180
rect 129700 329140 225512 329168
rect 129700 329128 129706 329140
rect 225506 329128 225512 329140
rect 225564 329128 225570 329180
rect 362770 329128 362776 329180
rect 362828 329168 362834 329180
rect 437474 329168 437480 329180
rect 362828 329140 437480 329168
rect 362828 329128 362834 329140
rect 437474 329128 437480 329140
rect 437532 329128 437538 329180
rect 119982 329060 119988 329112
rect 120040 329100 120046 329112
rect 221274 329100 221280 329112
rect 120040 329072 221280 329100
rect 120040 329060 120046 329072
rect 221274 329060 221280 329072
rect 221332 329060 221338 329112
rect 235902 329060 235908 329112
rect 235960 329100 235966 329112
rect 272886 329100 272892 329112
rect 235960 329072 272892 329100
rect 235960 329060 235966 329072
rect 272886 329060 272892 329072
rect 272944 329060 272950 329112
rect 380618 329060 380624 329112
rect 380676 329100 380682 329112
rect 477494 329100 477500 329112
rect 380676 329072 477500 329100
rect 380676 329060 380682 329072
rect 477494 329060 477500 329072
rect 477552 329060 477558 329112
rect 198734 328040 198740 328092
rect 198792 328080 198798 328092
rect 199470 328080 199476 328092
rect 198792 328052 199476 328080
rect 198792 328040 198798 328052
rect 199470 328040 199476 328052
rect 199528 328040 199534 328092
rect 131022 327768 131028 327820
rect 131080 327808 131086 327820
rect 225690 327808 225696 327820
rect 131080 327780 225696 327808
rect 131080 327768 131086 327780
rect 225690 327768 225696 327780
rect 225748 327768 225754 327820
rect 368014 327768 368020 327820
rect 368072 327808 368078 327820
rect 448514 327808 448520 327820
rect 368072 327780 448520 327808
rect 368072 327768 368078 327780
rect 448514 327768 448520 327780
rect 448572 327768 448578 327820
rect 11698 327700 11704 327752
rect 11756 327740 11762 327752
rect 172054 327740 172060 327752
rect 11756 327712 172060 327740
rect 11756 327700 11762 327712
rect 172054 327700 172060 327712
rect 172112 327700 172118 327752
rect 176562 327700 176568 327752
rect 176620 327740 176626 327752
rect 245746 327740 245752 327752
rect 176620 327712 245752 327740
rect 176620 327700 176626 327712
rect 245746 327700 245752 327712
rect 245804 327700 245810 327752
rect 398558 327700 398564 327752
rect 398616 327740 398622 327752
rect 517514 327740 517520 327752
rect 398616 327712 517520 327740
rect 398616 327700 398622 327712
rect 517514 327700 517520 327712
rect 517572 327700 517578 327752
rect 248598 326816 248604 326868
rect 248656 326816 248662 326868
rect 248616 326664 248644 326816
rect 248598 326612 248604 326664
rect 248656 326612 248662 326664
rect 169662 326408 169668 326460
rect 169720 326448 169726 326460
rect 242986 326448 242992 326460
rect 169720 326420 242992 326448
rect 169720 326408 169726 326420
rect 242986 326408 242992 326420
rect 243044 326408 243050 326460
rect 247126 326408 247132 326460
rect 247184 326408 247190 326460
rect 362862 326408 362868 326460
rect 362920 326448 362926 326460
rect 434714 326448 434720 326460
rect 362920 326420 434720 326448
rect 362920 326408 362926 326420
rect 434714 326408 434720 326420
rect 434772 326408 434778 326460
rect 88242 326340 88248 326392
rect 88300 326380 88306 326392
rect 88300 326352 205634 326380
rect 88300 326340 88306 326352
rect 186314 326272 186320 326324
rect 186372 326312 186378 326324
rect 186774 326312 186780 326324
rect 186372 326284 186780 326312
rect 186372 326272 186378 326284
rect 186774 326272 186780 326284
rect 186832 326272 186838 326324
rect 187694 326272 187700 326324
rect 187752 326312 187758 326324
rect 188430 326312 188436 326324
rect 187752 326284 188436 326312
rect 187752 326272 187758 326284
rect 188430 326272 188436 326284
rect 188488 326272 188494 326324
rect 189166 326272 189172 326324
rect 189224 326312 189230 326324
rect 189350 326312 189356 326324
rect 189224 326284 189356 326312
rect 189224 326272 189230 326284
rect 189350 326272 189356 326284
rect 189408 326272 189414 326324
rect 193306 326272 193312 326324
rect 193364 326312 193370 326324
rect 194134 326312 194140 326324
rect 193364 326284 194140 326312
rect 193364 326272 193370 326284
rect 194134 326272 194140 326284
rect 194192 326272 194198 326324
rect 194594 326272 194600 326324
rect 194652 326312 194658 326324
rect 195238 326312 195244 326324
rect 194652 326284 195244 326312
rect 194652 326272 194658 326284
rect 195238 326272 195244 326284
rect 195296 326272 195302 326324
rect 205606 326312 205634 326352
rect 207106 326340 207112 326392
rect 207164 326380 207170 326392
rect 207750 326380 207756 326392
rect 207164 326352 207756 326380
rect 207164 326340 207170 326352
rect 207750 326340 207756 326352
rect 207808 326340 207814 326392
rect 208486 326340 208492 326392
rect 208544 326380 208550 326392
rect 209406 326380 209412 326392
rect 208544 326352 209412 326380
rect 208544 326340 208550 326352
rect 209406 326340 209412 326352
rect 209464 326340 209470 326392
rect 214098 326340 214104 326392
rect 214156 326380 214162 326392
rect 214742 326380 214748 326392
rect 214156 326352 214748 326380
rect 214156 326340 214162 326352
rect 214742 326340 214748 326352
rect 214800 326340 214806 326392
rect 216766 326340 216772 326392
rect 216824 326380 216830 326392
rect 217318 326380 217324 326392
rect 216824 326352 217324 326380
rect 216824 326340 216830 326352
rect 217318 326340 217324 326352
rect 217376 326340 217382 326392
rect 222286 326340 222292 326392
rect 222344 326380 222350 326392
rect 222470 326380 222476 326392
rect 222344 326352 222476 326380
rect 222344 326340 222350 326352
rect 222470 326340 222476 326352
rect 222528 326340 222534 326392
rect 230474 326340 230480 326392
rect 230532 326380 230538 326392
rect 230934 326380 230940 326392
rect 230532 326352 230940 326380
rect 230532 326340 230538 326352
rect 230934 326340 230940 326352
rect 230992 326340 230998 326392
rect 231946 326340 231952 326392
rect 232004 326380 232010 326392
rect 232590 326380 232596 326392
rect 232004 326352 232596 326380
rect 232004 326340 232010 326352
rect 232590 326340 232596 326352
rect 232648 326340 232654 326392
rect 237374 326340 237380 326392
rect 237432 326380 237438 326392
rect 237650 326380 237656 326392
rect 237432 326352 237656 326380
rect 237432 326340 237438 326352
rect 237650 326340 237656 326352
rect 237708 326340 237714 326392
rect 241514 326340 241520 326392
rect 241572 326380 241578 326392
rect 241974 326380 241980 326392
rect 241572 326352 241980 326380
rect 241572 326340 241578 326352
rect 241974 326340 241980 326352
rect 242032 326340 242038 326392
rect 244274 326340 244280 326392
rect 244332 326380 244338 326392
rect 245102 326380 245108 326392
rect 244332 326352 245108 326380
rect 244332 326340 244338 326352
rect 245102 326340 245108 326352
rect 245160 326340 245166 326392
rect 207198 326312 207204 326324
rect 205606 326284 207204 326312
rect 207198 326272 207204 326284
rect 207256 326272 207262 326324
rect 247144 326256 247172 326408
rect 248506 326340 248512 326392
rect 248564 326380 248570 326392
rect 249334 326380 249340 326392
rect 248564 326352 249340 326380
rect 248564 326340 248570 326352
rect 249334 326340 249340 326352
rect 249392 326340 249398 326392
rect 258166 326340 258172 326392
rect 258224 326380 258230 326392
rect 258902 326380 258908 326392
rect 258224 326352 258908 326380
rect 258224 326340 258230 326352
rect 258902 326340 258908 326352
rect 258960 326340 258966 326392
rect 259546 326340 259552 326392
rect 259604 326380 259610 326392
rect 260374 326380 260380 326392
rect 259604 326352 260380 326380
rect 259604 326340 259610 326352
rect 260374 326340 260380 326352
rect 260432 326340 260438 326392
rect 333790 326340 333796 326392
rect 333848 326380 333854 326392
rect 371234 326380 371240 326392
rect 333848 326352 371240 326380
rect 333848 326340 333854 326352
rect 371234 326340 371240 326352
rect 371292 326340 371298 326392
rect 387610 326340 387616 326392
rect 387668 326380 387674 326392
rect 492674 326380 492680 326392
rect 387668 326352 492680 326380
rect 387668 326340 387674 326352
rect 492674 326340 492680 326352
rect 492732 326340 492738 326392
rect 237466 326204 237472 326256
rect 237524 326244 237530 326256
rect 238294 326244 238300 326256
rect 237524 326216 238300 326244
rect 237524 326204 237530 326216
rect 238294 326204 238300 326216
rect 238352 326204 238358 326256
rect 247126 326204 247132 326256
rect 247184 326204 247190 326256
rect 435358 325592 435364 325644
rect 435416 325632 435422 325644
rect 580166 325632 580172 325644
rect 435416 325604 580172 325632
rect 435416 325592 435422 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 133782 324980 133788 325032
rect 133840 325020 133846 325032
rect 226610 325020 226616 325032
rect 133840 324992 226616 325020
rect 133840 324980 133846 324992
rect 226610 324980 226616 324992
rect 226668 324980 226674 325032
rect 40678 324912 40684 324964
rect 40736 324952 40742 324964
rect 185118 324952 185124 324964
rect 40736 324924 185124 324952
rect 40736 324912 40742 324924
rect 185118 324912 185124 324924
rect 185176 324912 185182 324964
rect 347498 324912 347504 324964
rect 347556 324952 347562 324964
rect 402974 324952 402980 324964
rect 347556 324924 402980 324952
rect 347556 324912 347562 324924
rect 402974 324912 402980 324924
rect 403032 324912 403038 324964
rect 186406 324572 186412 324624
rect 186464 324612 186470 324624
rect 187326 324612 187332 324624
rect 186464 324584 187332 324612
rect 186464 324572 186470 324584
rect 187326 324572 187332 324584
rect 187384 324572 187390 324624
rect 178126 324368 178132 324420
rect 178184 324408 178190 324420
rect 178862 324408 178868 324420
rect 178184 324380 178868 324408
rect 178184 324368 178190 324380
rect 178862 324368 178868 324380
rect 178920 324368 178926 324420
rect 180886 324368 180892 324420
rect 180944 324408 180950 324420
rect 181438 324408 181444 324420
rect 180944 324380 181444 324408
rect 180944 324368 180950 324380
rect 181438 324368 181444 324380
rect 181496 324368 181502 324420
rect 236086 324368 236092 324420
rect 236144 324408 236150 324420
rect 236822 324408 236828 324420
rect 236144 324380 236828 324408
rect 236144 324368 236150 324380
rect 236822 324368 236828 324380
rect 236880 324368 236886 324420
rect 136542 323620 136548 323672
rect 136600 323660 136606 323672
rect 228266 323660 228272 323672
rect 136600 323632 228272 323660
rect 136600 323620 136606 323632
rect 228266 323620 228272 323632
rect 228324 323620 228330 323672
rect 355870 323620 355876 323672
rect 355928 323660 355934 323672
rect 420914 323660 420920 323672
rect 355928 323632 420920 323660
rect 355928 323620 355934 323632
rect 420914 323620 420920 323632
rect 420972 323620 420978 323672
rect 53742 323552 53748 323604
rect 53800 323592 53806 323604
rect 192018 323592 192024 323604
rect 53800 323564 192024 323592
rect 53800 323552 53806 323564
rect 192018 323552 192024 323564
rect 192076 323552 192082 323604
rect 248414 323552 248420 323604
rect 248472 323592 248478 323604
rect 248690 323592 248696 323604
rect 248472 323564 248696 323592
rect 248472 323552 248478 323564
rect 248690 323552 248696 323564
rect 248748 323552 248754 323604
rect 391750 323552 391756 323604
rect 391808 323592 391814 323604
rect 499574 323592 499580 323604
rect 391808 323564 499580 323592
rect 391808 323552 391814 323564
rect 499574 323552 499580 323564
rect 499632 323552 499638 323604
rect 182266 323484 182272 323536
rect 182324 323524 182330 323536
rect 182450 323524 182456 323536
rect 182324 323496 182456 323524
rect 182324 323484 182330 323496
rect 182450 323484 182456 323496
rect 182508 323484 182514 323536
rect 251174 323416 251180 323468
rect 251232 323456 251238 323468
rect 252094 323456 252100 323468
rect 251232 323428 252100 323456
rect 251232 323416 251238 323428
rect 252094 323416 252100 323428
rect 252152 323416 252158 323468
rect 147582 322192 147588 322244
rect 147640 322232 147646 322244
rect 233418 322232 233424 322244
rect 147640 322204 233424 322232
rect 147640 322192 147646 322204
rect 233418 322192 233424 322204
rect 233476 322192 233482 322244
rect 366910 322192 366916 322244
rect 366968 322232 366974 322244
rect 445754 322232 445760 322244
rect 366968 322204 445760 322232
rect 366968 322192 366974 322204
rect 445754 322192 445760 322204
rect 445812 322192 445818 322244
rect 247034 321648 247040 321700
rect 247092 321688 247098 321700
rect 247218 321688 247224 321700
rect 247092 321660 247224 321688
rect 247092 321648 247098 321660
rect 247218 321648 247224 321660
rect 247276 321648 247282 321700
rect 215386 321308 215392 321360
rect 215444 321348 215450 321360
rect 215570 321348 215576 321360
rect 215444 321320 215576 321348
rect 215444 321308 215450 321320
rect 215570 321308 215576 321320
rect 215628 321308 215634 321360
rect 144822 320832 144828 320884
rect 144880 320872 144886 320884
rect 232222 320872 232228 320884
rect 144880 320844 232228 320872
rect 144880 320832 144886 320844
rect 232222 320832 232228 320844
rect 232280 320832 232286 320884
rect 369762 320832 369768 320884
rect 369820 320872 369826 320884
rect 452654 320872 452660 320884
rect 369820 320844 452660 320872
rect 369820 320832 369826 320844
rect 452654 320832 452660 320844
rect 452712 320832 452718 320884
rect 3050 320084 3056 320136
rect 3108 320124 3114 320136
rect 166810 320124 166816 320136
rect 3108 320096 166816 320124
rect 3108 320084 3114 320096
rect 166810 320084 166816 320096
rect 166868 320084 166874 320136
rect 254026 319472 254032 319524
rect 254084 319512 254090 319524
rect 254210 319512 254216 319524
rect 254084 319484 254216 319512
rect 254084 319472 254090 319484
rect 254210 319472 254216 319484
rect 254268 319472 254274 319524
rect 375282 319404 375288 319456
rect 375340 319444 375346 319456
rect 463694 319444 463700 319456
rect 375340 319416 463700 319444
rect 375340 319404 375346 319416
rect 463694 319404 463700 319416
rect 463752 319404 463758 319456
rect 180702 318112 180708 318164
rect 180760 318152 180766 318164
rect 247770 318152 247776 318164
rect 180760 318124 247776 318152
rect 180760 318112 180766 318124
rect 247770 318112 247776 318124
rect 247828 318112 247834 318164
rect 113082 318044 113088 318096
rect 113140 318084 113146 318096
rect 218146 318084 218152 318096
rect 113140 318056 218152 318084
rect 113140 318044 113146 318056
rect 218146 318044 218152 318056
rect 218204 318044 218210 318096
rect 377950 318044 377956 318096
rect 378008 318084 378014 318096
rect 470594 318084 470600 318096
rect 378008 318056 470600 318084
rect 378008 318044 378014 318056
rect 470594 318044 470600 318056
rect 470652 318044 470658 318096
rect 137922 316684 137928 316736
rect 137980 316724 137986 316736
rect 229186 316724 229192 316736
rect 137980 316696 229192 316724
rect 137980 316684 137986 316696
rect 229186 316684 229192 316696
rect 229244 316684 229250 316736
rect 376478 316684 376484 316736
rect 376536 316724 376542 316736
rect 466454 316724 466460 316736
rect 376536 316696 466460 316724
rect 376536 316684 376542 316696
rect 466454 316684 466460 316696
rect 466512 316684 466518 316736
rect 162762 315256 162768 315308
rect 162820 315296 162826 315308
rect 240226 315296 240232 315308
rect 162820 315268 240232 315296
rect 162820 315256 162826 315268
rect 240226 315256 240232 315268
rect 240284 315256 240290 315308
rect 383470 315256 383476 315308
rect 383528 315296 383534 315308
rect 481634 315296 481640 315308
rect 383528 315268 481640 315296
rect 383528 315256 383534 315268
rect 481634 315256 481640 315268
rect 481692 315256 481698 315308
rect 142062 313896 142068 313948
rect 142120 313936 142126 313948
rect 230566 313936 230572 313948
rect 142120 313908 230572 313936
rect 142120 313896 142126 313908
rect 230566 313896 230572 313908
rect 230624 313896 230630 313948
rect 390278 313896 390284 313948
rect 390336 313936 390342 313948
rect 496814 313936 496820 313948
rect 390336 313908 496820 313936
rect 390336 313896 390342 313908
rect 496814 313896 496820 313908
rect 496872 313896 496878 313948
rect 461578 313216 461584 313268
rect 461636 313256 461642 313268
rect 580166 313256 580172 313268
rect 461636 313228 580172 313256
rect 461636 313216 461642 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 143442 312536 143448 312588
rect 143500 312576 143506 312588
rect 230474 312576 230480 312588
rect 143500 312548 230480 312576
rect 143500 312536 143506 312548
rect 230474 312536 230480 312548
rect 230532 312536 230538 312588
rect 99282 311108 99288 311160
rect 99340 311148 99346 311160
rect 210418 311148 210424 311160
rect 99340 311120 210424 311148
rect 99340 311108 99346 311120
rect 210418 311108 210424 311120
rect 210476 311108 210482 311160
rect 384850 311108 384856 311160
rect 384908 311148 384914 311160
rect 485774 311148 485780 311160
rect 384908 311120 485780 311148
rect 384908 311108 384914 311120
rect 485774 311108 485780 311120
rect 485832 311108 485838 311160
rect 33778 309748 33784 309800
rect 33836 309788 33842 309800
rect 179506 309788 179512 309800
rect 33836 309760 179512 309788
rect 33836 309748 33842 309760
rect 179506 309748 179512 309760
rect 179564 309748 179570 309800
rect 393130 309748 393136 309800
rect 393188 309788 393194 309800
rect 503714 309788 503720 309800
rect 393188 309760 503720 309788
rect 393188 309748 393194 309760
rect 503714 309748 503720 309760
rect 503772 309748 503778 309800
rect 124122 308388 124128 308440
rect 124180 308428 124186 308440
rect 222286 308428 222292 308440
rect 124180 308400 222292 308428
rect 124180 308388 124186 308400
rect 222286 308388 222292 308400
rect 222344 308388 222350 308440
rect 395890 308388 395896 308440
rect 395948 308428 395954 308440
rect 510614 308428 510620 308440
rect 395948 308400 510620 308428
rect 395948 308388 395954 308400
rect 510614 308388 510620 308400
rect 510672 308388 510678 308440
rect 106182 307028 106188 307080
rect 106240 307068 106246 307080
rect 214098 307068 214104 307080
rect 106240 307040 214104 307068
rect 106240 307028 106246 307040
rect 214098 307028 214104 307040
rect 214156 307028 214162 307080
rect 394510 307028 394516 307080
rect 394568 307068 394574 307080
rect 506474 307068 506480 307080
rect 394568 307040 506480 307068
rect 394568 307028 394574 307040
rect 506474 307028 506480 307040
rect 506532 307028 506538 307080
rect 43438 305600 43444 305652
rect 43496 305640 43502 305652
rect 186498 305640 186504 305652
rect 43496 305612 186504 305640
rect 43496 305600 43502 305612
rect 186498 305600 186504 305612
rect 186556 305600 186562 305652
rect 397178 305600 397184 305652
rect 397236 305640 397242 305652
rect 514754 305640 514760 305652
rect 397236 305612 514760 305640
rect 397236 305600 397242 305612
rect 514754 305600 514760 305612
rect 514812 305600 514818 305652
rect 36538 304240 36544 304292
rect 36596 304280 36602 304292
rect 180886 304280 180892 304292
rect 36596 304252 180892 304280
rect 36596 304240 36602 304252
rect 180886 304240 180892 304252
rect 180944 304240 180950 304292
rect 406930 304240 406936 304292
rect 406988 304280 406994 304292
rect 535454 304280 535460 304292
rect 406988 304252 535460 304280
rect 406988 304240 406994 304252
rect 535454 304240 535460 304252
rect 535512 304240 535518 304292
rect 57882 302880 57888 302932
rect 57940 302920 57946 302932
rect 193398 302920 193404 302932
rect 57940 302892 193404 302920
rect 57940 302880 57946 302892
rect 193398 302880 193404 302892
rect 193456 302880 193462 302932
rect 401318 302880 401324 302932
rect 401376 302920 401382 302932
rect 521654 302920 521660 302932
rect 401376 302892 521660 302920
rect 401376 302880 401382 302892
rect 521654 302880 521660 302892
rect 521712 302880 521718 302932
rect 50982 301452 50988 301504
rect 51040 301492 51046 301504
rect 188338 301492 188344 301504
rect 51040 301464 188344 301492
rect 51040 301452 51046 301464
rect 188338 301452 188344 301464
rect 188396 301452 188402 301504
rect 404170 301452 404176 301504
rect 404228 301492 404234 301504
rect 528554 301492 528560 301504
rect 404228 301464 528560 301492
rect 404228 301452 404234 301464
rect 528554 301452 528560 301464
rect 528612 301452 528618 301504
rect 46198 300092 46204 300144
rect 46256 300132 46262 300144
rect 187786 300132 187792 300144
rect 46256 300104 187792 300132
rect 46256 300092 46262 300104
rect 187786 300092 187792 300104
rect 187844 300092 187850 300144
rect 429194 299412 429200 299464
rect 429252 299452 429258 299464
rect 580166 299452 580172 299464
rect 429252 299424 580172 299452
rect 429252 299412 429258 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 61930 298732 61936 298784
rect 61988 298772 61994 298784
rect 194686 298772 194692 298784
rect 61988 298744 194692 298772
rect 61988 298732 61994 298744
rect 194686 298732 194692 298744
rect 194744 298732 194750 298784
rect 64782 297372 64788 297424
rect 64840 297412 64846 297424
rect 196158 297412 196164 297424
rect 64840 297384 196164 297412
rect 64840 297372 64846 297384
rect 196158 297372 196164 297384
rect 196216 297372 196222 297424
rect 68922 294584 68928 294636
rect 68980 294624 68986 294636
rect 197538 294624 197544 294636
rect 68980 294596 197544 294624
rect 68980 294584 68986 294596
rect 197538 294584 197544 294596
rect 197596 294584 197602 294636
rect 177942 290436 177948 290488
rect 178000 290476 178006 290488
rect 245654 290476 245660 290488
rect 178000 290448 245660 290476
rect 178000 290436 178006 290448
rect 245654 290436 245660 290448
rect 245712 290436 245718 290488
rect 173802 286288 173808 286340
rect 173860 286328 173866 286340
rect 244458 286328 244464 286340
rect 173860 286300 244464 286328
rect 173860 286288 173866 286300
rect 244458 286288 244464 286300
rect 244516 286288 244522 286340
rect 432598 285608 432604 285660
rect 432656 285648 432662 285660
rect 580166 285648 580172 285660
rect 432656 285620 580172 285648
rect 432656 285608 432662 285620
rect 580166 285608 580172 285620
rect 580224 285608 580230 285660
rect 3234 280100 3240 280152
rect 3292 280140 3298 280152
rect 166718 280140 166724 280152
rect 3292 280112 166724 280140
rect 3292 280100 3298 280112
rect 166718 280100 166724 280112
rect 166776 280100 166782 280152
rect 429286 273164 429292 273216
rect 429344 273204 429350 273216
rect 580166 273204 580172 273216
rect 429344 273176 580172 273204
rect 429344 273164 429350 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 135162 268336 135168 268388
rect 135220 268376 135226 268388
rect 226426 268376 226432 268388
rect 135220 268348 226432 268376
rect 135220 268336 135226 268348
rect 226426 268336 226432 268348
rect 226484 268336 226490 268388
rect 3050 267656 3056 267708
rect 3108 267696 3114 267708
rect 166626 267696 166632 267708
rect 3108 267668 166632 267696
rect 3108 267656 3114 267668
rect 166626 267656 166632 267668
rect 166684 267656 166690 267708
rect 429378 259360 429384 259412
rect 429436 259400 429442 259412
rect 580166 259400 580172 259412
rect 429436 259372 580172 259400
rect 429436 259360 429442 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 117222 255960 117228 256012
rect 117280 256000 117286 256012
rect 219526 256000 219532 256012
rect 117280 255972 219532 256000
rect 117280 255960 117286 255972
rect 219526 255960 219532 255972
rect 219584 255960 219590 256012
rect 3234 255212 3240 255264
rect 3292 255252 3298 255264
rect 22738 255252 22744 255264
rect 3292 255224 22744 255252
rect 3292 255212 3298 255224
rect 22738 255212 22744 255224
rect 22796 255212 22802 255264
rect 22738 253172 22744 253224
rect 22796 253212 22802 253224
rect 175366 253212 175372 253224
rect 22796 253184 175372 253212
rect 22796 253172 22802 253184
rect 175366 253172 175372 253184
rect 175424 253172 175430 253224
rect 386230 251812 386236 251864
rect 386288 251852 386294 251864
rect 490006 251852 490012 251864
rect 386288 251824 490012 251852
rect 386288 251812 386294 251824
rect 490006 251812 490012 251824
rect 490064 251812 490070 251864
rect 429470 245556 429476 245608
rect 429528 245596 429534 245608
rect 580166 245596 580172 245608
rect 429528 245568 580172 245596
rect 429528 245556 429534 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3234 241204 3240 241256
rect 3292 241244 3298 241256
rect 7558 241244 7564 241256
rect 3292 241216 7564 241244
rect 3292 241204 3298 241216
rect 7558 241204 7564 241216
rect 7616 241204 7622 241256
rect 431218 233180 431224 233232
rect 431276 233220 431282 233232
rect 579982 233220 579988 233232
rect 431276 233192 579988 233220
rect 431276 233180 431282 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 360010 232500 360016 232552
rect 360068 232540 360074 232552
rect 430574 232540 430580 232552
rect 360068 232512 430580 232540
rect 360068 232500 360074 232512
rect 430574 232500 430580 232512
rect 430632 232500 430638 232552
rect 3234 229032 3240 229084
rect 3292 229072 3298 229084
rect 166534 229072 166540 229084
rect 3292 229044 166540 229072
rect 3292 229032 3298 229044
rect 166534 229032 166540 229044
rect 166592 229032 166598 229084
rect 454678 219376 454684 219428
rect 454736 219416 454742 219428
rect 580166 219416 580172 219428
rect 454736 219388 580172 219416
rect 454736 219376 454742 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3234 215228 3240 215280
rect 3292 215268 3298 215280
rect 166442 215268 166448 215280
rect 3292 215240 166448 215268
rect 3292 215228 3298 215240
rect 166442 215228 166448 215240
rect 166500 215228 166506 215280
rect 429562 206932 429568 206984
rect 429620 206972 429626 206984
rect 579798 206972 579804 206984
rect 429620 206944 579804 206972
rect 429620 206932 429626 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 429654 193128 429660 193180
rect 429712 193168 429718 193180
rect 580166 193168 580172 193180
rect 429712 193140 580172 193168
rect 429712 193128 429718 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 14458 189020 14464 189032
rect 3384 188992 14464 189020
rect 3384 188980 3390 188992
rect 14458 188980 14464 188992
rect 14516 188980 14522 189032
rect 429746 179324 429752 179376
rect 429804 179364 429810 179376
rect 580166 179364 580172 179376
rect 429804 179336 580172 179364
rect 429804 179324 429810 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 25590 177284 25596 177336
rect 25648 177324 25654 177336
rect 178218 177324 178224 177336
rect 25648 177296 178224 177324
rect 25648 177284 25654 177296
rect 178218 177284 178224 177296
rect 178276 177284 178282 177336
rect 3326 176604 3332 176656
rect 3384 176644 3390 176656
rect 166350 176644 166356 176656
rect 3384 176616 166356 176644
rect 3384 176604 3390 176616
rect 166350 176604 166356 176616
rect 166408 176604 166414 176656
rect 372430 175924 372436 175976
rect 372488 175964 372494 175976
rect 456886 175964 456892 175976
rect 372488 175936 456892 175964
rect 372488 175924 372494 175936
rect 456886 175924 456892 175936
rect 456944 175924 456950 175976
rect 166902 174496 166908 174548
rect 166960 174536 166966 174548
rect 241606 174536 241612 174548
rect 166960 174508 241612 174536
rect 166960 174496 166966 174508
rect 241606 174496 241612 174508
rect 241664 174496 241670 174548
rect 365530 174496 365536 174548
rect 365588 174536 365594 174548
rect 441614 174536 441620 174548
rect 365588 174508 441620 174536
rect 365588 174496 365594 174508
rect 441614 174496 441620 174508
rect 441672 174496 441678 174548
rect 430482 166948 430488 167000
rect 430540 166988 430546 167000
rect 580166 166988 580172 167000
rect 430540 166960 580172 166988
rect 430540 166948 430546 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 430390 153144 430396 153196
rect 430448 153184 430454 153196
rect 580166 153184 580172 153196
rect 430448 153156 580172 153184
rect 430448 153144 430454 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 25498 150396 25504 150408
rect 3384 150368 25504 150396
rect 3384 150356 3390 150368
rect 25498 150356 25504 150368
rect 25556 150356 25562 150408
rect 447778 139340 447784 139392
rect 447836 139380 447842 139392
rect 580166 139380 580172 139392
rect 447836 139352 580172 139380
rect 447836 139340 447842 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 430298 126896 430304 126948
rect 430356 126936 430362 126948
rect 580166 126936 580172 126948
rect 430356 126908 580172 126936
rect 430356 126896 430362 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3142 124108 3148 124160
rect 3200 124148 3206 124160
rect 166258 124148 166264 124160
rect 3200 124120 166264 124148
rect 3200 124108 3206 124120
rect 166258 124108 166264 124120
rect 166316 124108 166322 124160
rect 430206 113092 430212 113144
rect 430264 113132 430270 113144
rect 579798 113132 579804 113144
rect 430264 113104 579804 113132
rect 430264 113092 430270 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 430114 100648 430120 100700
rect 430172 100688 430178 100700
rect 580166 100688 580172 100700
rect 430172 100660 580172 100688
rect 430172 100648 430178 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 430022 86912 430028 86964
rect 430080 86952 430086 86964
rect 580166 86952 580172 86964
rect 430080 86924 580172 86952
rect 430080 86912 430086 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 15838 85524 15844 85536
rect 3200 85496 15844 85524
rect 3200 85484 3206 85496
rect 15838 85484 15844 85496
rect 15896 85484 15902 85536
rect 429930 73108 429936 73160
rect 429988 73148 429994 73160
rect 580166 73148 580172 73160
rect 429988 73120 580172 73148
rect 429988 73108 429994 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 442258 60664 442264 60716
rect 442316 60704 442322 60716
rect 580166 60704 580172 60716
rect 442316 60676 580172 60704
rect 442316 60664 442322 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 2866 59304 2872 59356
rect 2924 59344 2930 59356
rect 32398 59344 32404 59356
rect 2924 59316 32404 59344
rect 2924 59304 2930 59316
rect 32398 59304 32404 59316
rect 32456 59304 32462 59356
rect 439498 46860 439504 46912
rect 439556 46900 439562 46912
rect 580166 46900 580172 46912
rect 439556 46872 580172 46900
rect 439556 46860 439562 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 364150 44820 364156 44872
rect 364208 44860 364214 44872
rect 438854 44860 438860 44872
rect 364208 44832 438860 44860
rect 364208 44820 364214 44832
rect 438854 44820 438860 44832
rect 438912 44820 438918 44872
rect 136450 35164 136456 35216
rect 136508 35204 136514 35216
rect 227714 35204 227720 35216
rect 136508 35176 227720 35204
rect 136508 35164 136514 35176
rect 227714 35164 227720 35176
rect 227772 35164 227778 35216
rect 368290 35164 368296 35216
rect 368348 35204 368354 35216
rect 448606 35204 448612 35216
rect 368348 35176 448612 35204
rect 368348 35164 368354 35176
rect 448606 35164 448612 35176
rect 448664 35164 448670 35216
rect 429838 33056 429844 33108
rect 429896 33096 429902 33108
rect 580166 33096 580172 33108
rect 429896 33068 580172 33096
rect 429896 33056 429902 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 209682 31016 209688 31068
rect 209740 31056 209746 31068
rect 259546 31056 259552 31068
rect 209740 31028 259552 31056
rect 209740 31016 209746 31028
rect 259546 31016 259552 31028
rect 259604 31016 259610 31068
rect 354398 31016 354404 31068
rect 354456 31056 354462 31068
rect 416774 31056 416780 31068
rect 354456 31028 416780 31056
rect 354456 31016 354462 31028
rect 416774 31016 416780 31028
rect 416832 31016 416838 31068
rect 346118 29588 346124 29640
rect 346176 29628 346182 29640
rect 398834 29628 398840 29640
rect 346176 29600 398840 29628
rect 346176 29588 346182 29600
rect 398834 29588 398840 29600
rect 398892 29588 398898 29640
rect 92382 28228 92388 28280
rect 92440 28268 92446 28280
rect 208578 28268 208584 28280
rect 92440 28240 208584 28268
rect 92440 28228 92446 28240
rect 208578 28228 208584 28240
rect 208636 28228 208642 28280
rect 353202 28228 353208 28280
rect 353260 28268 353266 28280
rect 414014 28268 414020 28280
rect 353260 28240 414020 28268
rect 353260 28228 353266 28240
rect 414014 28228 414020 28240
rect 414072 28228 414078 28280
rect 146202 26868 146208 26920
rect 146260 26908 146266 26920
rect 231946 26908 231952 26920
rect 146260 26880 231952 26908
rect 146260 26868 146266 26880
rect 231946 26868 231952 26880
rect 232004 26868 232010 26920
rect 358078 26868 358084 26920
rect 358136 26908 358142 26920
rect 396074 26908 396080 26920
rect 358136 26880 396080 26908
rect 358136 26868 358142 26880
rect 396074 26868 396080 26880
rect 396132 26868 396138 26920
rect 343358 25576 343364 25628
rect 343416 25616 343422 25628
rect 391934 25616 391940 25628
rect 343416 25588 391940 25616
rect 343416 25576 343422 25588
rect 391934 25576 391940 25588
rect 391992 25576 391998 25628
rect 139302 25508 139308 25560
rect 139360 25548 139366 25560
rect 229278 25548 229284 25560
rect 139360 25520 229284 25548
rect 139360 25508 139366 25520
rect 229278 25508 229284 25520
rect 229336 25508 229342 25560
rect 379330 25508 379336 25560
rect 379388 25548 379394 25560
rect 473354 25548 473360 25560
rect 379388 25520 473360 25548
rect 379388 25508 379394 25520
rect 473354 25508 473360 25520
rect 473412 25508 473418 25560
rect 200022 24080 200028 24132
rect 200080 24120 200086 24132
rect 255498 24120 255504 24132
rect 200080 24092 255504 24120
rect 200080 24080 200086 24092
rect 255498 24080 255504 24092
rect 255556 24080 255562 24132
rect 372522 24080 372528 24132
rect 372580 24120 372586 24132
rect 458174 24120 458180 24132
rect 372580 24092 458180 24120
rect 372580 24080 372586 24092
rect 458174 24080 458180 24092
rect 458232 24080 458238 24132
rect 177850 22720 177856 22772
rect 177908 22760 177914 22772
rect 247126 22760 247132 22772
rect 177908 22732 247132 22760
rect 177908 22720 177914 22732
rect 247126 22720 247132 22732
rect 247184 22720 247190 22772
rect 371050 22720 371056 22772
rect 371108 22760 371114 22772
rect 455414 22760 455420 22772
rect 371108 22732 455420 22760
rect 371108 22720 371114 22732
rect 455414 22720 455420 22732
rect 455472 22720 455478 22772
rect 188982 21360 188988 21412
rect 189040 21400 189046 21412
rect 251358 21400 251364 21412
rect 189040 21372 251364 21400
rect 189040 21360 189046 21372
rect 251358 21360 251364 21372
rect 251416 21360 251422 21412
rect 370498 21360 370504 21412
rect 370556 21400 370562 21412
rect 451274 21400 451280 21412
rect 370556 21372 451280 21400
rect 370556 21360 370562 21372
rect 451274 21360 451280 21372
rect 451332 21360 451338 21412
rect 336458 20000 336464 20052
rect 336516 20040 336522 20052
rect 378134 20040 378140 20052
rect 336516 20012 378140 20040
rect 336516 20000 336522 20012
rect 378134 20000 378140 20012
rect 378192 20000 378198 20052
rect 182082 19932 182088 19984
rect 182140 19972 182146 19984
rect 248598 19972 248604 19984
rect 182140 19944 248604 19972
rect 182140 19932 182146 19944
rect 248598 19932 248604 19944
rect 248656 19932 248662 19984
rect 357250 19932 357256 19984
rect 357308 19972 357314 19984
rect 423674 19972 423680 19984
rect 357308 19944 423680 19972
rect 357308 19932 357314 19944
rect 423674 19932 423680 19944
rect 423732 19932 423738 19984
rect 187602 18640 187608 18692
rect 187660 18680 187666 18692
rect 251266 18680 251272 18692
rect 187660 18652 251272 18680
rect 187660 18640 187666 18652
rect 251266 18640 251272 18652
rect 251324 18640 251330 18692
rect 332318 18640 332324 18692
rect 332376 18680 332382 18692
rect 367094 18680 367100 18692
rect 332376 18652 367100 18680
rect 332376 18640 332382 18652
rect 367094 18640 367100 18652
rect 367152 18640 367158 18692
rect 103422 18572 103428 18624
rect 103480 18612 103486 18624
rect 212626 18612 212632 18624
rect 103480 18584 212632 18612
rect 103480 18572 103486 18584
rect 212626 18572 212632 18584
rect 212684 18572 212690 18624
rect 367002 18572 367008 18624
rect 367060 18612 367066 18624
rect 444374 18612 444380 18624
rect 367060 18584 444380 18612
rect 367060 18572 367066 18584
rect 444374 18572 444380 18584
rect 444432 18572 444438 18624
rect 184842 17280 184848 17332
rect 184900 17320 184906 17332
rect 248506 17320 248512 17332
rect 184900 17292 248512 17320
rect 184900 17280 184906 17292
rect 248506 17280 248512 17292
rect 248564 17280 248570 17332
rect 85482 17212 85488 17264
rect 85540 17252 85546 17264
rect 204438 17252 204444 17264
rect 85540 17224 204444 17252
rect 85540 17212 85546 17224
rect 204438 17212 204444 17224
rect 204496 17212 204502 17264
rect 328270 17212 328276 17264
rect 328328 17252 328334 17264
rect 357526 17252 357532 17264
rect 328328 17224 357532 17252
rect 328328 17212 328334 17224
rect 357526 17212 357532 17224
rect 357584 17212 357590 17264
rect 365622 17212 365628 17264
rect 365680 17252 365686 17264
rect 440326 17252 440332 17264
rect 365680 17224 440332 17252
rect 365680 17212 365686 17224
rect 440326 17212 440332 17224
rect 440384 17212 440390 17264
rect 169570 15852 169576 15904
rect 169628 15892 169634 15904
rect 240778 15892 240784 15904
rect 169628 15864 240784 15892
rect 169628 15852 169634 15864
rect 240778 15852 240784 15864
rect 240836 15852 240842 15904
rect 324130 15852 324136 15904
rect 324188 15892 324194 15904
rect 349246 15892 349252 15904
rect 324188 15864 349252 15892
rect 324188 15852 324194 15864
rect 349246 15852 349252 15864
rect 349304 15852 349310 15904
rect 349798 15852 349804 15904
rect 349856 15892 349862 15904
rect 361114 15892 361120 15904
rect 349856 15864 361120 15892
rect 349856 15852 349862 15864
rect 361114 15852 361120 15864
rect 361172 15852 361178 15904
rect 361298 15852 361304 15904
rect 361356 15892 361362 15904
rect 434438 15892 434444 15904
rect 361356 15864 434444 15892
rect 361356 15852 361362 15864
rect 434438 15852 434444 15864
rect 434496 15852 434502 15904
rect 128262 14424 128268 14476
rect 128320 14464 128326 14476
rect 223666 14464 223672 14476
rect 128320 14436 223672 14464
rect 128320 14424 128326 14436
rect 223666 14424 223672 14436
rect 223724 14424 223730 14476
rect 233142 14424 233148 14476
rect 233200 14464 233206 14476
rect 270586 14464 270592 14476
rect 233200 14436 270592 14464
rect 233200 14424 233206 14436
rect 270586 14424 270592 14436
rect 270644 14424 270650 14476
rect 320082 14424 320088 14476
rect 320140 14464 320146 14476
rect 339862 14464 339868 14476
rect 320140 14436 339868 14464
rect 320140 14424 320146 14436
rect 339862 14424 339868 14436
rect 339920 14424 339926 14476
rect 340598 14424 340604 14476
rect 340656 14464 340662 14476
rect 385954 14464 385960 14476
rect 340656 14436 385960 14464
rect 340656 14424 340662 14436
rect 385954 14424 385960 14436
rect 386012 14424 386018 14476
rect 390370 14424 390376 14476
rect 390428 14464 390434 14476
rect 498194 14464 498200 14476
rect 390428 14436 498200 14464
rect 390428 14424 390434 14436
rect 498194 14424 498200 14436
rect 498252 14424 498258 14476
rect 183462 13132 183468 13184
rect 183520 13172 183526 13184
rect 248414 13172 248420 13184
rect 183520 13144 248420 13172
rect 183520 13132 183526 13144
rect 248414 13132 248420 13144
rect 248472 13132 248478 13184
rect 342070 13132 342076 13184
rect 342128 13172 342134 13184
rect 389450 13172 389456 13184
rect 342128 13144 389456 13172
rect 342128 13132 342134 13144
rect 389450 13132 389456 13144
rect 389508 13132 389514 13184
rect 131758 13064 131764 13116
rect 131816 13104 131822 13116
rect 226334 13104 226340 13116
rect 131816 13076 226340 13104
rect 131816 13064 131822 13076
rect 226334 13064 226340 13076
rect 226392 13064 226398 13116
rect 321278 13064 321284 13116
rect 321336 13104 321342 13116
rect 343358 13104 343364 13116
rect 321336 13076 343364 13104
rect 321336 13064 321342 13076
rect 343358 13064 343364 13076
rect 343416 13064 343422 13116
rect 388990 13064 388996 13116
rect 389048 13104 389054 13116
rect 494698 13104 494704 13116
rect 389048 13076 494704 13104
rect 389048 13064 389054 13076
rect 494698 13064 494704 13076
rect 494756 13064 494762 13116
rect 179046 11772 179052 11824
rect 179104 11812 179110 11824
rect 247034 11812 247040 11824
rect 179104 11784 247040 11812
rect 179104 11772 179110 11784
rect 247034 11772 247040 11784
rect 247092 11772 247098 11824
rect 322658 11772 322664 11824
rect 322716 11812 322722 11824
rect 345750 11812 345756 11824
rect 322716 11784 345756 11812
rect 322716 11772 322722 11784
rect 345750 11772 345756 11784
rect 345808 11772 345814 11824
rect 489178 11772 489184 11824
rect 489236 11812 489242 11824
rect 580258 11812 580264 11824
rect 489236 11784 580264 11812
rect 489236 11772 489242 11784
rect 580258 11772 580264 11784
rect 580316 11772 580322 11824
rect 110322 11704 110328 11756
rect 110380 11744 110386 11756
rect 191098 11744 191104 11756
rect 110380 11716 191104 11744
rect 110380 11704 110386 11716
rect 191098 11704 191104 11716
rect 191156 11704 191162 11756
rect 193122 11704 193128 11756
rect 193180 11744 193186 11756
rect 252646 11744 252652 11756
rect 193180 11716 252652 11744
rect 193180 11704 193186 11716
rect 252646 11704 252652 11716
rect 252704 11704 252710 11756
rect 339218 11704 339224 11756
rect 339276 11744 339282 11756
rect 382366 11744 382372 11756
rect 339276 11716 382372 11744
rect 339276 11704 339282 11716
rect 382366 11704 382372 11716
rect 382424 11704 382430 11756
rect 393222 11704 393228 11756
rect 393280 11744 393286 11756
rect 505370 11744 505376 11756
rect 393280 11716 505376 11744
rect 393280 11704 393286 11716
rect 505370 11704 505376 11716
rect 505428 11704 505434 11756
rect 186130 10344 186136 10396
rect 186188 10384 186194 10396
rect 249886 10384 249892 10396
rect 186188 10356 249892 10384
rect 186188 10344 186194 10356
rect 249886 10344 249892 10356
rect 249944 10344 249950 10396
rect 319438 10344 319444 10396
rect 319496 10384 319502 10396
rect 338666 10384 338672 10396
rect 319496 10356 338672 10384
rect 319496 10344 319502 10356
rect 338666 10344 338672 10356
rect 338724 10344 338730 10396
rect 350350 10344 350356 10396
rect 350408 10384 350414 10396
rect 407206 10384 407212 10396
rect 350408 10356 407212 10384
rect 350408 10344 350414 10356
rect 407206 10344 407212 10356
rect 407264 10344 407270 10396
rect 81342 10276 81348 10328
rect 81400 10316 81406 10328
rect 159358 10316 159364 10328
rect 81400 10288 159364 10316
rect 81400 10276 81406 10288
rect 159358 10276 159364 10288
rect 159416 10276 159422 10328
rect 172422 10276 172428 10328
rect 172480 10316 172486 10328
rect 244366 10316 244372 10328
rect 172480 10288 244372 10316
rect 172480 10276 172486 10288
rect 244366 10276 244372 10288
rect 244424 10276 244430 10328
rect 335078 10276 335084 10328
rect 335136 10316 335142 10328
rect 373994 10316 374000 10328
rect 335136 10288 374000 10316
rect 335136 10276 335142 10288
rect 373994 10276 374000 10288
rect 374052 10276 374058 10328
rect 385678 10276 385684 10328
rect 385736 10316 385742 10328
rect 487614 10316 487620 10328
rect 385736 10288 487620 10316
rect 385736 10276 385742 10288
rect 487614 10276 487620 10288
rect 487672 10276 487678 10328
rect 185118 9188 185124 9240
rect 185176 9228 185182 9240
rect 249794 9228 249800 9240
rect 185176 9200 249800 9228
rect 185176 9188 185182 9200
rect 249794 9188 249800 9200
rect 249852 9188 249858 9240
rect 77386 9120 77392 9172
rect 77444 9160 77450 9172
rect 201586 9160 201592 9172
rect 77444 9132 201592 9160
rect 77444 9120 77450 9132
rect 201586 9120 201592 9132
rect 201644 9120 201650 9172
rect 73798 9052 73804 9104
rect 73856 9092 73862 9104
rect 200298 9092 200304 9104
rect 73856 9064 200304 9092
rect 73856 9052 73862 9064
rect 200298 9052 200304 9064
rect 200356 9052 200362 9104
rect 70302 8984 70308 9036
rect 70360 9024 70366 9036
rect 198826 9024 198832 9036
rect 70360 8996 198832 9024
rect 70360 8984 70366 8996
rect 198826 8984 198832 8996
rect 198884 8984 198890 9036
rect 321370 8984 321376 9036
rect 321428 9024 321434 9036
rect 342162 9024 342168 9036
rect 321428 8996 342168 9024
rect 321428 8984 321434 8996
rect 342162 8984 342168 8996
rect 342220 8984 342226 9036
rect 374638 8984 374644 9036
rect 374696 9024 374702 9036
rect 427262 9024 427268 9036
rect 374696 8996 427268 9024
rect 374696 8984 374702 8996
rect 427262 8984 427268 8996
rect 427320 8984 427326 9036
rect 66714 8916 66720 8968
rect 66772 8956 66778 8968
rect 197446 8956 197452 8968
rect 66772 8928 197452 8956
rect 66772 8916 66778 8928
rect 197446 8916 197452 8928
rect 197504 8916 197510 8968
rect 228726 8916 228732 8968
rect 228784 8956 228790 8968
rect 269206 8956 269212 8968
rect 228784 8928 269212 8956
rect 228784 8916 228790 8928
rect 269206 8916 269212 8928
rect 269264 8916 269270 8968
rect 325510 8916 325516 8968
rect 325568 8956 325574 8968
rect 354030 8956 354036 8968
rect 325568 8928 354036 8956
rect 325568 8916 325574 8928
rect 354030 8916 354036 8928
rect 354088 8916 354094 8968
rect 382182 8916 382188 8968
rect 382240 8956 382246 8968
rect 480530 8956 480536 8968
rect 382240 8928 480536 8956
rect 382240 8916 382246 8928
rect 480530 8916 480536 8928
rect 480588 8916 480594 8968
rect 424686 8304 424692 8356
rect 424744 8344 424750 8356
rect 424962 8344 424968 8356
rect 424744 8316 424968 8344
rect 424744 8304 424750 8316
rect 424962 8304 424968 8316
rect 425020 8304 425026 8356
rect 108114 8236 108120 8288
rect 108172 8276 108178 8288
rect 215386 8276 215392 8288
rect 108172 8248 215392 8276
rect 108172 8236 108178 8248
rect 215386 8236 215392 8248
rect 215444 8236 215450 8288
rect 409598 8236 409604 8288
rect 409656 8276 409662 8288
rect 541986 8276 541992 8288
rect 409656 8248 541992 8276
rect 409656 8236 409662 8248
rect 541986 8236 541992 8248
rect 542044 8236 542050 8288
rect 104526 8168 104532 8220
rect 104584 8208 104590 8220
rect 214006 8208 214012 8220
rect 104584 8180 214012 8208
rect 104584 8168 104590 8180
rect 214006 8168 214012 8180
rect 214064 8168 214070 8220
rect 411070 8168 411076 8220
rect 411128 8208 411134 8220
rect 545482 8208 545488 8220
rect 411128 8180 545488 8208
rect 411128 8168 411134 8180
rect 545482 8168 545488 8180
rect 545540 8168 545546 8220
rect 101030 8100 101036 8152
rect 101088 8140 101094 8152
rect 212534 8140 212540 8152
rect 101088 8112 212540 8140
rect 101088 8100 101094 8112
rect 212534 8100 212540 8112
rect 212592 8100 212598 8152
rect 412358 8100 412364 8152
rect 412416 8140 412422 8152
rect 549070 8140 549076 8152
rect 412416 8112 549076 8140
rect 412416 8100 412422 8112
rect 549070 8100 549076 8112
rect 549128 8100 549134 8152
rect 97442 8032 97448 8084
rect 97500 8072 97506 8084
rect 211246 8072 211252 8084
rect 97500 8044 211252 8072
rect 97500 8032 97506 8044
rect 211246 8032 211252 8044
rect 211304 8032 211310 8084
rect 413738 8032 413744 8084
rect 413796 8072 413802 8084
rect 552658 8072 552664 8084
rect 413796 8044 552664 8072
rect 413796 8032 413802 8044
rect 552658 8032 552664 8044
rect 552716 8032 552722 8084
rect 93946 7964 93952 8016
rect 94004 8004 94010 8016
rect 208486 8004 208492 8016
rect 94004 7976 208492 8004
rect 94004 7964 94010 7976
rect 208486 7964 208492 7976
rect 208544 7964 208550 8016
rect 416498 7964 416504 8016
rect 416556 8004 416562 8016
rect 556154 8004 556160 8016
rect 416556 7976 556160 8004
rect 416556 7964 416562 7976
rect 556154 7964 556160 7976
rect 556212 7964 556218 8016
rect 90358 7896 90364 7948
rect 90416 7936 90422 7948
rect 207106 7936 207112 7948
rect 90416 7908 207112 7936
rect 90416 7896 90422 7908
rect 207106 7896 207112 7908
rect 207164 7896 207170 7948
rect 417970 7896 417976 7948
rect 418028 7936 418034 7948
rect 559742 7936 559748 7948
rect 418028 7908 559748 7936
rect 418028 7896 418034 7908
rect 559742 7896 559748 7908
rect 559800 7896 559806 7948
rect 86862 7828 86868 7880
rect 86920 7868 86926 7880
rect 205726 7868 205732 7880
rect 86920 7840 205732 7868
rect 86920 7828 86926 7840
rect 205726 7828 205732 7840
rect 205784 7828 205790 7880
rect 420638 7828 420644 7880
rect 420696 7868 420702 7880
rect 425517 7871 425575 7877
rect 420696 7840 425468 7868
rect 420696 7828 420702 7840
rect 63218 7760 63224 7812
rect 63276 7800 63282 7812
rect 196066 7800 196072 7812
rect 63276 7772 196072 7800
rect 63276 7760 63282 7772
rect 196066 7760 196072 7772
rect 196124 7760 196130 7812
rect 422110 7760 422116 7812
rect 422168 7800 422174 7812
rect 425440 7800 425468 7840
rect 425517 7837 425529 7871
rect 425563 7868 425575 7871
rect 563238 7868 563244 7880
rect 425563 7840 563244 7868
rect 425563 7837 425575 7840
rect 425517 7831 425575 7837
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 566826 7800 566832 7812
rect 422168 7772 425376 7800
rect 425440 7772 566832 7800
rect 422168 7760 422174 7772
rect 59630 7692 59636 7744
rect 59688 7732 59694 7744
rect 193306 7732 193312 7744
rect 59688 7704 193312 7732
rect 59688 7692 59694 7704
rect 193306 7692 193312 7704
rect 193364 7692 193370 7744
rect 423398 7692 423404 7744
rect 423456 7732 423462 7744
rect 425348 7732 425376 7772
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 570322 7732 570328 7744
rect 423456 7704 425284 7732
rect 425348 7704 570328 7732
rect 423456 7692 423462 7704
rect 56042 7624 56048 7676
rect 56100 7664 56106 7676
rect 191926 7664 191932 7676
rect 56100 7636 191932 7664
rect 56100 7624 56106 7636
rect 191926 7624 191932 7636
rect 191984 7624 191990 7676
rect 317138 7624 317144 7676
rect 317196 7664 317202 7676
rect 335078 7664 335084 7676
rect 317196 7636 335084 7664
rect 317196 7624 317202 7636
rect 335078 7624 335084 7636
rect 335136 7624 335142 7676
rect 424778 7624 424784 7676
rect 424836 7664 424842 7676
rect 425256 7664 425284 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 573910 7664 573916 7676
rect 424836 7636 425100 7664
rect 425256 7636 573916 7664
rect 424836 7624 424842 7636
rect 52546 7556 52552 7608
rect 52604 7596 52610 7608
rect 190546 7596 190552 7608
rect 52604 7568 190552 7596
rect 52604 7556 52610 7568
rect 190546 7556 190552 7568
rect 190604 7556 190610 7608
rect 239306 7556 239312 7608
rect 239364 7596 239370 7608
rect 273438 7596 273444 7608
rect 239364 7568 273444 7596
rect 239364 7556 239370 7568
rect 273438 7556 273444 7568
rect 273496 7556 273502 7608
rect 324222 7556 324228 7608
rect 324280 7596 324286 7608
rect 350350 7596 350356 7608
rect 324280 7568 350356 7596
rect 324280 7556 324286 7568
rect 350350 7556 350356 7568
rect 350408 7556 350414 7608
rect 423674 7556 423680 7608
rect 423732 7596 423738 7608
rect 424962 7596 424968 7608
rect 423732 7568 424968 7596
rect 423732 7556 423738 7568
rect 424962 7556 424968 7568
rect 425020 7556 425026 7608
rect 425072 7596 425100 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 577406 7596 577412 7608
rect 425072 7568 577412 7596
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 111610 7488 111616 7540
rect 111668 7528 111674 7540
rect 216766 7528 216772 7540
rect 111668 7500 216772 7528
rect 111668 7488 111674 7500
rect 216766 7488 216772 7500
rect 216824 7488 216830 7540
rect 408218 7488 408224 7540
rect 408276 7528 408282 7540
rect 538398 7528 538404 7540
rect 408276 7500 538404 7528
rect 408276 7488 408282 7500
rect 538398 7488 538404 7500
rect 538456 7488 538462 7540
rect 115198 7420 115204 7472
rect 115256 7460 115262 7472
rect 218238 7460 218244 7472
rect 115256 7432 218244 7460
rect 115256 7420 115262 7432
rect 218238 7420 218244 7432
rect 218296 7420 218302 7472
rect 407022 7420 407028 7472
rect 407080 7460 407086 7472
rect 534902 7460 534908 7472
rect 407080 7432 534908 7460
rect 407080 7420 407086 7432
rect 534902 7420 534908 7432
rect 534960 7420 534966 7472
rect 118786 7352 118792 7404
rect 118844 7392 118850 7404
rect 220906 7392 220912 7404
rect 118844 7364 220912 7392
rect 118844 7352 118850 7364
rect 220906 7352 220912 7364
rect 220964 7352 220970 7404
rect 405550 7352 405556 7404
rect 405608 7392 405614 7404
rect 531406 7392 531412 7404
rect 405608 7364 531412 7392
rect 405608 7352 405614 7364
rect 531406 7352 531412 7364
rect 531464 7352 531470 7404
rect 122282 7284 122288 7336
rect 122340 7324 122346 7336
rect 222378 7324 222384 7336
rect 122340 7296 222384 7324
rect 122340 7284 122346 7296
rect 222378 7284 222384 7296
rect 222436 7284 222442 7336
rect 402790 7284 402796 7336
rect 402848 7324 402854 7336
rect 527818 7324 527824 7336
rect 402848 7296 527824 7324
rect 402848 7284 402854 7296
rect 527818 7284 527824 7296
rect 527876 7284 527882 7336
rect 153010 7216 153016 7268
rect 153068 7256 153074 7268
rect 236178 7256 236184 7268
rect 153068 7228 236184 7256
rect 153068 7216 153074 7228
rect 236178 7216 236184 7228
rect 236236 7216 236242 7268
rect 361390 7216 361396 7268
rect 361448 7256 361454 7268
rect 432046 7256 432052 7268
rect 361448 7228 432052 7256
rect 361448 7216 361454 7228
rect 432046 7216 432052 7228
rect 432104 7216 432110 7268
rect 149514 7148 149520 7200
rect 149572 7188 149578 7200
rect 233326 7188 233332 7200
rect 149572 7160 233332 7188
rect 149572 7148 149578 7160
rect 233326 7148 233332 7160
rect 233384 7148 233390 7200
rect 358630 7148 358636 7200
rect 358688 7188 358694 7200
rect 428458 7188 428464 7200
rect 358688 7160 428464 7188
rect 358688 7148 358694 7160
rect 428458 7148 428464 7160
rect 428516 7148 428522 7200
rect 156598 7080 156604 7132
rect 156656 7120 156662 7132
rect 237558 7120 237564 7132
rect 156656 7092 237564 7120
rect 156656 7080 156662 7092
rect 237558 7080 237564 7092
rect 237616 7080 237622 7132
rect 419258 7080 419264 7132
rect 419316 7120 419322 7132
rect 425517 7123 425575 7129
rect 425517 7120 425529 7123
rect 419316 7092 425529 7120
rect 419316 7080 419322 7092
rect 425517 7089 425529 7092
rect 425563 7089 425575 7123
rect 425517 7083 425575 7089
rect 160094 7012 160100 7064
rect 160152 7052 160158 7064
rect 238754 7052 238760 7064
rect 160152 7024 238760 7052
rect 160152 7012 160158 7024
rect 238754 7012 238760 7024
rect 238812 7012 238818 7064
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 17218 6848 17224 6860
rect 3476 6820 17224 6848
rect 3476 6808 3482 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 83274 6808 83280 6860
rect 83332 6848 83338 6860
rect 204346 6848 204352 6860
rect 83332 6820 204352 6848
rect 83332 6808 83338 6820
rect 204346 6808 204352 6820
rect 204404 6808 204410 6860
rect 386322 6808 386328 6860
rect 386380 6848 386386 6860
rect 488810 6848 488816 6860
rect 386380 6820 488816 6848
rect 386380 6808 386386 6820
rect 488810 6808 488816 6820
rect 488868 6808 488874 6860
rect 48958 6740 48964 6792
rect 49016 6780 49022 6792
rect 189166 6780 189172 6792
rect 49016 6752 189172 6780
rect 49016 6740 49022 6752
rect 189166 6740 189172 6752
rect 189224 6740 189230 6792
rect 387518 6740 387524 6792
rect 387576 6780 387582 6792
rect 492306 6780 492312 6792
rect 387576 6752 492312 6780
rect 387576 6740 387582 6752
rect 492306 6740 492312 6752
rect 492364 6740 492370 6792
rect 44266 6672 44272 6724
rect 44324 6712 44330 6724
rect 186406 6712 186412 6724
rect 44324 6684 186412 6712
rect 44324 6672 44330 6684
rect 186406 6672 186412 6684
rect 186464 6672 186470 6724
rect 389082 6672 389088 6724
rect 389140 6712 389146 6724
rect 495894 6712 495900 6724
rect 389140 6684 495900 6712
rect 389140 6672 389146 6684
rect 495894 6672 495900 6684
rect 495952 6672 495958 6724
rect 40770 6604 40776 6656
rect 40828 6644 40834 6656
rect 185026 6644 185032 6656
rect 40828 6616 185032 6644
rect 40828 6604 40834 6616
rect 185026 6604 185032 6616
rect 185084 6604 185090 6656
rect 390462 6604 390468 6656
rect 390520 6644 390526 6656
rect 499390 6644 499396 6656
rect 390520 6616 499396 6644
rect 390520 6604 390526 6616
rect 499390 6604 499396 6616
rect 499448 6604 499454 6656
rect 37182 6536 37188 6588
rect 37240 6576 37246 6588
rect 183646 6576 183652 6588
rect 37240 6548 183652 6576
rect 37240 6536 37246 6548
rect 183646 6536 183652 6548
rect 183704 6536 183710 6588
rect 205082 6536 205088 6588
rect 205140 6576 205146 6588
rect 258166 6576 258172 6588
rect 205140 6548 258172 6576
rect 205140 6536 205146 6548
rect 258166 6536 258172 6548
rect 258224 6536 258230 6588
rect 391842 6536 391848 6588
rect 391900 6576 391906 6588
rect 502978 6576 502984 6588
rect 391900 6548 502984 6576
rect 391900 6536 391906 6548
rect 502978 6536 502984 6548
rect 503036 6536 503042 6588
rect 33594 6468 33600 6520
rect 33652 6508 33658 6520
rect 182266 6508 182272 6520
rect 33652 6480 182272 6508
rect 33652 6468 33658 6480
rect 182266 6468 182272 6480
rect 182324 6468 182330 6520
rect 201586 6468 201592 6520
rect 201644 6508 201650 6520
rect 256786 6508 256792 6520
rect 201644 6480 256792 6508
rect 201644 6468 201650 6480
rect 256786 6468 256792 6480
rect 256844 6468 256850 6520
rect 394418 6468 394424 6520
rect 394476 6508 394482 6520
rect 506566 6508 506572 6520
rect 394476 6480 506572 6508
rect 394476 6468 394482 6480
rect 506566 6468 506572 6480
rect 506624 6468 506630 6520
rect 30098 6400 30104 6452
rect 30156 6440 30162 6452
rect 180978 6440 180984 6452
rect 30156 6412 180984 6440
rect 30156 6400 30162 6412
rect 180978 6400 180984 6412
rect 181036 6400 181042 6452
rect 197906 6400 197912 6452
rect 197964 6440 197970 6452
rect 255406 6440 255412 6452
rect 197964 6412 255412 6440
rect 197964 6400 197970 6412
rect 255406 6400 255412 6412
rect 255464 6400 255470 6452
rect 395982 6400 395988 6452
rect 396040 6440 396046 6452
rect 510062 6440 510068 6452
rect 396040 6412 510068 6440
rect 396040 6400 396046 6412
rect 510062 6400 510068 6412
rect 510120 6400 510126 6452
rect 26510 6332 26516 6384
rect 26568 6372 26574 6384
rect 179414 6372 179420 6384
rect 26568 6344 179420 6372
rect 26568 6332 26574 6344
rect 179414 6332 179420 6344
rect 179472 6332 179478 6384
rect 194410 6332 194416 6384
rect 194468 6372 194474 6384
rect 254026 6372 254032 6384
rect 194468 6344 254032 6372
rect 194468 6332 194474 6344
rect 254026 6332 254032 6344
rect 254084 6332 254090 6384
rect 397270 6332 397276 6384
rect 397328 6372 397334 6384
rect 513558 6372 513564 6384
rect 397328 6344 513564 6372
rect 397328 6332 397334 6344
rect 513558 6332 513564 6344
rect 513616 6332 513622 6384
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 176746 6304 176752 6316
rect 21876 6276 176752 6304
rect 21876 6264 21882 6276
rect 176746 6264 176752 6276
rect 176804 6264 176810 6316
rect 190822 6264 190828 6316
rect 190880 6304 190886 6316
rect 252554 6304 252560 6316
rect 190880 6276 252560 6304
rect 190880 6264 190886 6276
rect 252554 6264 252560 6276
rect 252612 6264 252618 6316
rect 398650 6264 398656 6316
rect 398708 6304 398714 6316
rect 517146 6304 517152 6316
rect 398708 6276 517152 6304
rect 398708 6264 398714 6276
rect 517146 6264 517152 6276
rect 517204 6264 517210 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 171226 6236 171232 6248
rect 8812 6208 171232 6236
rect 8812 6196 8818 6208
rect 171226 6196 171232 6208
rect 171284 6196 171290 6248
rect 174262 6196 174268 6248
rect 174320 6236 174326 6248
rect 244274 6236 244280 6248
rect 174320 6208 244280 6236
rect 174320 6196 174326 6208
rect 244274 6196 244280 6208
rect 244332 6196 244338 6248
rect 315942 6196 315948 6248
rect 316000 6236 316006 6248
rect 331582 6236 331588 6248
rect 316000 6208 331588 6236
rect 316000 6196 316006 6208
rect 331582 6196 331588 6208
rect 331640 6196 331646 6248
rect 400030 6196 400036 6248
rect 400088 6236 400094 6248
rect 520734 6236 520740 6248
rect 400088 6208 520740 6236
rect 400088 6196 400094 6208
rect 520734 6196 520740 6208
rect 520792 6196 520798 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 169846 6168 169852 6180
rect 4120 6140 169852 6168
rect 4120 6128 4126 6140
rect 169846 6128 169852 6140
rect 169904 6128 169910 6180
rect 170766 6128 170772 6180
rect 170824 6168 170830 6180
rect 243078 6168 243084 6180
rect 170824 6140 243084 6168
rect 170824 6128 170830 6140
rect 243078 6128 243084 6140
rect 243136 6128 243142 6180
rect 322750 6128 322756 6180
rect 322808 6168 322814 6180
rect 346946 6168 346952 6180
rect 322808 6140 346952 6168
rect 322808 6128 322814 6140
rect 346946 6128 346952 6140
rect 347004 6128 347010 6180
rect 352558 6128 352564 6180
rect 352616 6168 352622 6180
rect 364610 6168 364616 6180
rect 352616 6140 364616 6168
rect 352616 6128 352622 6140
rect 364610 6128 364616 6140
rect 364668 6128 364674 6180
rect 401410 6128 401416 6180
rect 401468 6168 401474 6180
rect 524230 6168 524236 6180
rect 401468 6140 524236 6168
rect 401468 6128 401474 6140
rect 524230 6128 524236 6140
rect 524288 6128 524294 6180
rect 128170 6060 128176 6112
rect 128228 6100 128234 6112
rect 224954 6100 224960 6112
rect 128228 6072 224960 6100
rect 128228 6060 128234 6072
rect 224954 6060 224960 6072
rect 225012 6060 225018 6112
rect 384942 6060 384948 6112
rect 385000 6100 385006 6112
rect 485222 6100 485228 6112
rect 385000 6072 485228 6100
rect 385000 6060 385006 6072
rect 485222 6060 485228 6072
rect 485280 6060 485286 6112
rect 144730 5992 144736 6044
rect 144788 6032 144794 6044
rect 231854 6032 231860 6044
rect 144788 6004 231860 6032
rect 144788 5992 144794 6004
rect 231854 5992 231860 6004
rect 231912 5992 231918 6044
rect 383562 5992 383568 6044
rect 383620 6032 383626 6044
rect 481726 6032 481732 6044
rect 383620 6004 481732 6032
rect 383620 5992 383626 6004
rect 481726 5992 481732 6004
rect 481784 5992 481790 6044
rect 148318 5924 148324 5976
rect 148376 5964 148382 5976
rect 233234 5964 233240 5976
rect 148376 5936 233240 5964
rect 148376 5924 148382 5936
rect 233234 5924 233240 5936
rect 233292 5924 233298 5976
rect 380710 5924 380716 5976
rect 380768 5964 380774 5976
rect 476942 5964 476948 5976
rect 380768 5936 476948 5964
rect 380768 5924 380774 5936
rect 476942 5924 476948 5936
rect 477000 5924 477006 5976
rect 151814 5856 151820 5908
rect 151872 5896 151878 5908
rect 234706 5896 234712 5908
rect 151872 5868 234712 5896
rect 151872 5856 151878 5868
rect 234706 5856 234712 5868
rect 234764 5856 234770 5908
rect 379422 5856 379428 5908
rect 379480 5896 379486 5908
rect 473446 5896 473452 5908
rect 379480 5868 473452 5896
rect 379480 5856 379486 5868
rect 473446 5856 473452 5868
rect 473504 5856 473510 5908
rect 155402 5788 155408 5840
rect 155460 5828 155466 5840
rect 236086 5828 236092 5840
rect 155460 5800 236092 5828
rect 155460 5788 155466 5800
rect 236086 5788 236092 5800
rect 236144 5788 236150 5840
rect 378042 5788 378048 5840
rect 378100 5828 378106 5840
rect 469858 5828 469864 5840
rect 378100 5800 469864 5828
rect 378100 5788 378106 5800
rect 469858 5788 469864 5800
rect 469916 5788 469922 5840
rect 158898 5720 158904 5772
rect 158956 5760 158962 5772
rect 237466 5760 237472 5772
rect 158956 5732 237472 5760
rect 158956 5720 158962 5732
rect 237466 5720 237472 5732
rect 237524 5720 237530 5772
rect 376570 5720 376576 5772
rect 376628 5760 376634 5772
rect 466270 5760 466276 5772
rect 376628 5732 466276 5760
rect 376628 5720 376634 5732
rect 466270 5720 466276 5732
rect 466328 5720 466334 5772
rect 163682 5652 163688 5704
rect 163740 5692 163746 5704
rect 240318 5692 240324 5704
rect 163740 5664 240324 5692
rect 163740 5652 163746 5664
rect 240318 5652 240324 5664
rect 240376 5652 240382 5704
rect 373810 5652 373816 5704
rect 373868 5692 373874 5704
rect 462774 5692 462780 5704
rect 373868 5664 462780 5692
rect 373868 5652 373874 5664
rect 462774 5652 462780 5664
rect 462832 5652 462838 5704
rect 167178 5584 167184 5636
rect 167236 5624 167242 5636
rect 241514 5624 241520 5636
rect 167236 5596 241520 5624
rect 167236 5584 167242 5596
rect 241514 5584 241520 5596
rect 241572 5584 241578 5636
rect 62022 5448 62028 5500
rect 62080 5488 62086 5500
rect 194594 5488 194600 5500
rect 62080 5460 194600 5488
rect 62080 5448 62086 5460
rect 194594 5448 194600 5460
rect 194652 5448 194658 5500
rect 225138 5448 225144 5500
rect 225196 5488 225202 5500
rect 267826 5488 267832 5500
rect 225196 5460 267832 5488
rect 225196 5448 225202 5460
rect 267826 5448 267832 5460
rect 267884 5448 267890 5500
rect 343450 5448 343456 5500
rect 343508 5488 343514 5500
rect 391842 5488 391848 5500
rect 343508 5460 391848 5488
rect 343508 5448 343514 5460
rect 391842 5448 391848 5460
rect 391900 5448 391906 5500
rect 409690 5448 409696 5500
rect 409748 5488 409754 5500
rect 540790 5488 540796 5500
rect 409748 5460 540796 5488
rect 409748 5448 409754 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 58434 5380 58440 5432
rect 58492 5420 58498 5432
rect 193214 5420 193220 5432
rect 58492 5392 193220 5420
rect 58492 5380 58498 5392
rect 193214 5380 193220 5392
rect 193272 5380 193278 5432
rect 221550 5380 221556 5432
rect 221608 5420 221614 5432
rect 266446 5420 266452 5432
rect 221608 5392 266452 5420
rect 221608 5380 221614 5392
rect 266446 5380 266452 5392
rect 266504 5380 266510 5432
rect 340690 5380 340696 5432
rect 340748 5420 340754 5432
rect 388254 5420 388260 5432
rect 340748 5392 388260 5420
rect 340748 5380 340754 5392
rect 388254 5380 388260 5392
rect 388312 5380 388318 5432
rect 411162 5380 411168 5432
rect 411220 5420 411226 5432
rect 544378 5420 544384 5432
rect 411220 5392 544384 5420
rect 411220 5380 411226 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 54938 5312 54944 5364
rect 54996 5352 55002 5364
rect 191834 5352 191840 5364
rect 54996 5324 191840 5352
rect 54996 5312 55002 5324
rect 191834 5312 191840 5324
rect 191892 5312 191898 5364
rect 218054 5312 218060 5364
rect 218112 5352 218118 5364
rect 265066 5352 265072 5364
rect 218112 5324 265072 5352
rect 218112 5312 218118 5324
rect 265066 5312 265072 5324
rect 265124 5312 265130 5364
rect 344922 5312 344928 5364
rect 344980 5352 344986 5364
rect 395338 5352 395344 5364
rect 344980 5324 395344 5352
rect 344980 5312 344986 5324
rect 395338 5312 395344 5324
rect 395396 5312 395402 5364
rect 412450 5312 412456 5364
rect 412508 5352 412514 5364
rect 547874 5352 547880 5364
rect 412508 5324 547880 5352
rect 412508 5312 412514 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 51350 5244 51356 5296
rect 51408 5284 51414 5296
rect 190454 5284 190460 5296
rect 51408 5256 190460 5284
rect 51408 5244 51414 5256
rect 190454 5244 190460 5256
rect 190512 5244 190518 5296
rect 214466 5244 214472 5296
rect 214524 5284 214530 5296
rect 262306 5284 262312 5296
rect 214524 5256 262312 5284
rect 214524 5244 214530 5256
rect 262306 5244 262312 5256
rect 262364 5244 262370 5296
rect 346210 5244 346216 5296
rect 346268 5284 346274 5296
rect 398926 5284 398932 5296
rect 346268 5256 398932 5284
rect 346268 5244 346274 5256
rect 398926 5244 398932 5256
rect 398984 5244 398990 5296
rect 413830 5244 413836 5296
rect 413888 5284 413894 5296
rect 551462 5284 551468 5296
rect 413888 5256 551468 5284
rect 413888 5244 413894 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 47854 5176 47860 5228
rect 47912 5216 47918 5228
rect 189258 5216 189264 5228
rect 47912 5188 189264 5216
rect 47912 5176 47918 5188
rect 189258 5176 189264 5188
rect 189316 5176 189322 5228
rect 210970 5176 210976 5228
rect 211028 5216 211034 5228
rect 260926 5216 260932 5228
rect 211028 5188 260932 5216
rect 211028 5176 211034 5188
rect 260926 5176 260932 5188
rect 260984 5176 260990 5228
rect 347590 5176 347596 5228
rect 347648 5216 347654 5228
rect 402514 5216 402520 5228
rect 347648 5188 402520 5216
rect 347648 5176 347654 5188
rect 402514 5176 402520 5188
rect 402572 5176 402578 5228
rect 415210 5176 415216 5228
rect 415268 5216 415274 5228
rect 554958 5216 554964 5228
rect 415268 5188 554964 5216
rect 415268 5176 415274 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 175458 5148 175464 5160
rect 17092 5120 175464 5148
rect 17092 5108 17098 5120
rect 175458 5108 175464 5120
rect 175516 5108 175522 5160
rect 207382 5108 207388 5160
rect 207440 5148 207446 5160
rect 259638 5148 259644 5160
rect 207440 5120 259644 5148
rect 207440 5108 207446 5120
rect 259638 5108 259644 5120
rect 259696 5108 259702 5160
rect 348970 5108 348976 5160
rect 349028 5148 349034 5160
rect 406010 5148 406016 5160
rect 349028 5120 406016 5148
rect 349028 5108 349034 5120
rect 406010 5108 406016 5120
rect 406068 5108 406074 5160
rect 416590 5108 416596 5160
rect 416648 5148 416654 5160
rect 558546 5148 558552 5160
rect 416648 5120 558552 5148
rect 416648 5108 416654 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 162762 5080 162768 5092
rect 12400 5052 162768 5080
rect 12400 5040 12406 5052
rect 162762 5040 162768 5052
rect 162820 5040 162826 5092
rect 171134 5080 171140 5092
rect 162872 5052 171140 5080
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 162872 5012 162900 5052
rect 171134 5040 171140 5052
rect 171192 5040 171198 5092
rect 203886 5040 203892 5092
rect 203944 5080 203950 5092
rect 258258 5080 258264 5092
rect 203944 5052 258264 5080
rect 203944 5040 203950 5052
rect 258258 5040 258264 5052
rect 258316 5040 258322 5092
rect 350442 5040 350448 5092
rect 350500 5080 350506 5092
rect 409598 5080 409604 5092
rect 350500 5052 409604 5080
rect 350500 5040 350506 5052
rect 409598 5040 409604 5052
rect 409656 5040 409662 5092
rect 419350 5040 419356 5092
rect 419408 5080 419414 5092
rect 562042 5080 562048 5092
rect 419408 5052 562048 5080
rect 419408 5040 419414 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 7708 4984 162900 5012
rect 162949 5015 163007 5021
rect 7708 4972 7714 4984
rect 162949 4981 162961 5015
rect 162995 5012 163007 5015
rect 168466 5012 168472 5024
rect 162995 4984 168472 5012
rect 162995 4981 163007 4984
rect 162949 4975 163007 4981
rect 168466 4972 168472 4984
rect 168524 4972 168530 5024
rect 172606 5012 172612 5024
rect 171106 4984 172612 5012
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 162673 4947 162731 4953
rect 162673 4944 162685 4947
rect 2924 4916 162685 4944
rect 2924 4904 2930 4916
rect 162673 4913 162685 4916
rect 162719 4913 162731 4947
rect 162673 4907 162731 4913
rect 162762 4904 162768 4956
rect 162820 4944 162826 4956
rect 171106 4944 171134 4984
rect 172606 4972 172612 4984
rect 172664 4972 172670 5024
rect 200298 4972 200304 5024
rect 200356 5012 200362 5024
rect 256694 5012 256700 5024
rect 200356 4984 256700 5012
rect 200356 4972 200362 4984
rect 256694 4972 256700 4984
rect 256752 4972 256758 5024
rect 351730 4972 351736 5024
rect 351788 5012 351794 5024
rect 413094 5012 413100 5024
rect 351788 4984 413100 5012
rect 351788 4972 351794 4984
rect 413094 4972 413100 4984
rect 413152 4972 413158 5024
rect 420730 4972 420736 5024
rect 420788 5012 420794 5024
rect 565630 5012 565636 5024
rect 420788 4984 565636 5012
rect 420788 4972 420794 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 162820 4916 171134 4944
rect 162820 4904 162826 4916
rect 196802 4904 196808 4956
rect 196860 4944 196866 4956
rect 255314 4944 255320 4956
rect 196860 4916 255320 4944
rect 196860 4904 196866 4916
rect 255314 4904 255320 4916
rect 255372 4904 255378 4956
rect 354490 4904 354496 4956
rect 354548 4944 354554 4956
rect 416498 4944 416504 4956
rect 354548 4916 416504 4944
rect 354548 4904 354554 4916
rect 416498 4904 416504 4916
rect 416556 4904 416562 4956
rect 422202 4904 422208 4956
rect 422260 4944 422266 4956
rect 569126 4944 569132 4956
rect 422260 4916 569132 4944
rect 422260 4904 422266 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 166994 4876 167000 4888
rect 624 4848 167000 4876
rect 624 4836 630 4848
rect 166994 4836 167000 4848
rect 167052 4836 167058 4888
rect 193214 4836 193220 4888
rect 193272 4876 193278 4888
rect 254118 4876 254124 4888
rect 193272 4848 254124 4876
rect 193272 4836 193278 4848
rect 254118 4836 254124 4848
rect 254176 4836 254182 4888
rect 355962 4836 355968 4888
rect 356020 4876 356026 4888
rect 420178 4876 420184 4888
rect 356020 4848 420184 4876
rect 356020 4836 356026 4848
rect 420178 4836 420184 4848
rect 420236 4836 420242 4888
rect 423490 4836 423496 4888
rect 423548 4876 423554 4888
rect 572714 4876 572720 4888
rect 423548 4848 572720 4876
rect 423548 4836 423554 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 162581 4811 162639 4817
rect 162581 4808 162593 4811
rect 1728 4780 162593 4808
rect 1728 4768 1734 4780
rect 162581 4777 162593 4780
rect 162627 4777 162639 4811
rect 162581 4771 162639 4777
rect 162673 4811 162731 4817
rect 162673 4777 162685 4811
rect 162719 4808 162731 4811
rect 168374 4808 168380 4820
rect 162719 4780 168380 4808
rect 162719 4777 162731 4780
rect 162673 4771 162731 4777
rect 168374 4768 168380 4780
rect 168432 4768 168438 4820
rect 189718 4768 189724 4820
rect 189776 4808 189782 4820
rect 251174 4808 251180 4820
rect 189776 4780 251180 4808
rect 189776 4768 189782 4780
rect 251174 4768 251180 4780
rect 251232 4768 251238 4820
rect 357342 4768 357348 4820
rect 357400 4808 357406 4820
rect 423766 4808 423772 4820
rect 357400 4780 423772 4808
rect 357400 4768 357406 4780
rect 423766 4768 423772 4780
rect 423824 4768 423830 4820
rect 424870 4768 424876 4820
rect 424928 4808 424934 4820
rect 576302 4808 576308 4820
rect 424928 4780 576308 4808
rect 424928 4768 424934 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 65518 4700 65524 4752
rect 65576 4740 65582 4752
rect 195974 4740 195980 4752
rect 65576 4712 195980 4740
rect 65576 4700 65582 4712
rect 195974 4700 195980 4712
rect 196032 4700 196038 4752
rect 339310 4700 339316 4752
rect 339368 4740 339374 4752
rect 384758 4740 384764 4752
rect 339368 4712 384764 4740
rect 339368 4700 339374 4712
rect 384758 4700 384764 4712
rect 384816 4700 384822 4752
rect 408310 4700 408316 4752
rect 408368 4740 408374 4752
rect 537202 4740 537208 4752
rect 408368 4712 537208 4740
rect 408368 4700 408374 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 72602 4632 72608 4684
rect 72660 4672 72666 4684
rect 200206 4672 200212 4684
rect 72660 4644 200212 4672
rect 72660 4632 72666 4644
rect 200206 4632 200212 4644
rect 200264 4632 200270 4684
rect 337930 4632 337936 4684
rect 337988 4672 337994 4684
rect 381170 4672 381176 4684
rect 337988 4644 381176 4672
rect 337988 4632 337994 4644
rect 381170 4632 381176 4644
rect 381228 4632 381234 4684
rect 405458 4632 405464 4684
rect 405516 4672 405522 4684
rect 533706 4672 533712 4684
rect 405516 4644 533712 4672
rect 405516 4632 405522 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 69106 4564 69112 4616
rect 69164 4604 69170 4616
rect 197354 4604 197360 4616
rect 69164 4576 197360 4604
rect 69164 4564 69170 4576
rect 197354 4564 197360 4576
rect 197412 4564 197418 4616
rect 336550 4564 336556 4616
rect 336608 4604 336614 4616
rect 377674 4604 377680 4616
rect 336608 4576 377680 4604
rect 336608 4564 336614 4576
rect 377674 4564 377680 4576
rect 377732 4564 377738 4616
rect 404262 4564 404268 4616
rect 404320 4604 404326 4616
rect 530118 4604 530124 4616
rect 404320 4576 530124 4604
rect 404320 4564 404326 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 76190 4496 76196 4548
rect 76248 4536 76254 4548
rect 201494 4536 201500 4548
rect 76248 4508 201500 4536
rect 76248 4496 76254 4508
rect 201494 4496 201500 4508
rect 201552 4496 201558 4548
rect 335170 4496 335176 4548
rect 335228 4536 335234 4548
rect 335228 4508 369164 4536
rect 335228 4496 335234 4508
rect 79686 4428 79692 4480
rect 79744 4468 79750 4480
rect 202966 4468 202972 4480
rect 79744 4440 202972 4468
rect 79744 4428 79750 4440
rect 202966 4428 202972 4440
rect 203024 4428 203030 4480
rect 333882 4428 333888 4480
rect 333940 4468 333946 4480
rect 369136 4468 369164 4508
rect 402882 4496 402888 4548
rect 402940 4536 402946 4548
rect 526622 4536 526628 4548
rect 402940 4508 526628 4536
rect 402940 4496 402946 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 374086 4468 374092 4480
rect 333940 4440 369072 4468
rect 369136 4440 374092 4468
rect 333940 4428 333946 4440
rect 150618 4360 150624 4412
rect 150676 4400 150682 4412
rect 234614 4400 234620 4412
rect 150676 4372 234620 4400
rect 150676 4360 150682 4372
rect 234614 4360 234620 4372
rect 234672 4360 234678 4412
rect 332410 4360 332416 4412
rect 332468 4400 332474 4412
rect 367002 4400 367008 4412
rect 332468 4372 367008 4400
rect 332468 4360 332474 4372
rect 367002 4360 367008 4372
rect 367060 4360 367066 4412
rect 369044 4400 369072 4440
rect 374086 4428 374092 4440
rect 374144 4428 374150 4480
rect 401502 4428 401508 4480
rect 401560 4468 401566 4480
rect 523034 4468 523040 4480
rect 401560 4440 523040 4468
rect 401560 4428 401566 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 370590 4400 370596 4412
rect 369044 4372 370596 4400
rect 370590 4360 370596 4372
rect 370648 4360 370654 4412
rect 400122 4360 400128 4412
rect 400180 4400 400186 4412
rect 519538 4400 519544 4412
rect 400180 4372 519544 4400
rect 400180 4360 400186 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 154206 4292 154212 4344
rect 154264 4332 154270 4344
rect 235994 4332 236000 4344
rect 154264 4304 236000 4332
rect 154264 4292 154270 4304
rect 235994 4292 236000 4304
rect 236052 4292 236058 4344
rect 329650 4292 329656 4344
rect 329708 4332 329714 4344
rect 363506 4332 363512 4344
rect 329708 4304 363512 4332
rect 329708 4292 329714 4304
rect 363506 4292 363512 4304
rect 363564 4292 363570 4344
rect 398742 4292 398748 4344
rect 398800 4332 398806 4344
rect 515950 4332 515956 4344
rect 398800 4304 515956 4332
rect 398800 4292 398806 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 157794 4224 157800 4276
rect 157852 4264 157858 4276
rect 237374 4264 237380 4276
rect 157852 4236 237380 4264
rect 157852 4224 157858 4236
rect 237374 4224 237380 4236
rect 237432 4224 237438 4276
rect 397362 4224 397368 4276
rect 397420 4264 397426 4276
rect 512454 4264 512460 4276
rect 397420 4236 512460 4264
rect 397420 4224 397426 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 126974 4156 126980 4208
rect 127032 4196 127038 4208
rect 128262 4196 128268 4208
rect 127032 4168 128268 4196
rect 127032 4156 127038 4168
rect 128262 4156 128268 4168
rect 128320 4156 128326 4208
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 144822 4196 144828 4208
rect 143592 4168 144828 4196
rect 143592 4156 143598 4168
rect 144822 4156 144828 4168
rect 144880 4156 144886 4208
rect 168374 4156 168380 4208
rect 168432 4196 168438 4208
rect 169662 4196 169668 4208
rect 168432 4168 169668 4196
rect 168432 4156 168438 4168
rect 169662 4156 169668 4168
rect 169720 4156 169726 4208
rect 171781 4199 171839 4205
rect 171781 4165 171793 4199
rect 171827 4196 171839 4199
rect 178126 4196 178132 4208
rect 171827 4168 178132 4196
rect 171827 4165 171839 4168
rect 171781 4159 171839 4165
rect 178126 4156 178132 4168
rect 178184 4156 178190 4208
rect 269853 4199 269911 4205
rect 269853 4165 269865 4199
rect 269899 4196 269911 4199
rect 269899 4168 272564 4196
rect 269899 4165 269911 4168
rect 269853 4159 269911 4165
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 28258 4128 28264 4140
rect 20680 4100 28264 4128
rect 20680 4088 20686 4100
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 46198 4128 46204 4140
rect 45520 4100 46204 4128
rect 45520 4088 45526 4100
rect 46198 4088 46204 4100
rect 46256 4088 46262 4140
rect 85666 4088 85672 4140
rect 85724 4128 85730 4140
rect 205634 4128 205640 4140
rect 85724 4100 205640 4128
rect 85724 4088 85730 4100
rect 205634 4088 205640 4100
rect 205692 4088 205698 4140
rect 252370 4088 252376 4140
rect 252428 4128 252434 4140
rect 272429 4131 272487 4137
rect 272429 4128 272441 4131
rect 252428 4100 272441 4128
rect 252428 4088 252434 4100
rect 272429 4097 272441 4100
rect 272475 4097 272487 4131
rect 272536 4128 272564 4168
rect 448606 4156 448612 4208
rect 448664 4196 448670 4208
rect 449802 4196 449808 4208
rect 448664 4168 449808 4196
rect 448664 4156 448670 4168
rect 449802 4156 449808 4168
rect 449860 4156 449866 4208
rect 272705 4131 272763 4137
rect 272536 4100 272656 4128
rect 272429 4091 272487 4097
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 204254 4060 204260 4072
rect 82136 4032 204260 4060
rect 82136 4020 82142 4032
rect 204254 4020 204260 4032
rect 204312 4020 204318 4072
rect 248782 4020 248788 4072
rect 248840 4060 248846 4072
rect 272521 4063 272579 4069
rect 272521 4060 272533 4063
rect 248840 4032 272533 4060
rect 248840 4020 248846 4032
rect 272521 4029 272533 4032
rect 272567 4029 272579 4063
rect 272628 4060 272656 4100
rect 272705 4097 272717 4131
rect 272751 4128 272763 4131
rect 280338 4128 280344 4140
rect 272751 4100 280344 4128
rect 272751 4097 272763 4100
rect 272705 4091 272763 4097
rect 280338 4088 280344 4100
rect 280396 4088 280402 4140
rect 306282 4088 306288 4140
rect 306340 4128 306346 4140
rect 309042 4128 309048 4140
rect 306340 4100 309048 4128
rect 306340 4088 306346 4100
rect 309042 4088 309048 4100
rect 309100 4088 309106 4140
rect 309778 4088 309784 4140
rect 309836 4128 309842 4140
rect 310330 4128 310336 4140
rect 309836 4100 310336 4128
rect 309836 4088 309842 4100
rect 310330 4088 310336 4100
rect 310388 4088 310394 4140
rect 318610 4088 318616 4140
rect 318668 4128 318674 4140
rect 325605 4131 325663 4137
rect 325605 4128 325617 4131
rect 318668 4100 325617 4128
rect 318668 4088 318674 4100
rect 325605 4097 325617 4100
rect 325651 4097 325663 4131
rect 325605 4091 325663 4097
rect 338022 4088 338028 4140
rect 338080 4128 338086 4140
rect 379974 4128 379980 4140
rect 338080 4100 379980 4128
rect 338080 4088 338086 4100
rect 379974 4088 379980 4100
rect 380032 4088 380038 4140
rect 409782 4088 409788 4140
rect 409840 4128 409846 4140
rect 543182 4128 543188 4140
rect 409840 4100 543188 4128
rect 409840 4088 409846 4100
rect 543182 4088 543188 4100
rect 543240 4088 543246 4140
rect 277210 4060 277216 4072
rect 272628 4032 277216 4060
rect 272521 4023 272579 4029
rect 277210 4020 277216 4032
rect 277268 4020 277274 4072
rect 294874 4020 294880 4072
rect 294932 4060 294938 4072
rect 298278 4060 298284 4072
rect 294932 4032 298284 4060
rect 294932 4020 294938 4032
rect 298278 4020 298284 4032
rect 298336 4020 298342 4072
rect 317230 4020 317236 4072
rect 317288 4060 317294 4072
rect 325510 4060 325516 4072
rect 317288 4032 325516 4060
rect 317288 4020 317294 4032
rect 325510 4020 325516 4032
rect 325568 4020 325574 4072
rect 339402 4020 339408 4072
rect 339460 4060 339466 4072
rect 383562 4060 383568 4072
rect 339460 4032 383568 4060
rect 339460 4020 339466 4032
rect 383562 4020 383568 4032
rect 383620 4020 383626 4072
rect 412542 4020 412548 4072
rect 412600 4060 412606 4072
rect 546678 4060 546684 4072
rect 412600 4032 546684 4060
rect 412600 4020 412606 4032
rect 546678 4020 546684 4032
rect 546736 4020 546742 4072
rect 78582 3952 78588 4004
rect 78640 3992 78646 4004
rect 203058 3992 203064 4004
rect 78640 3964 203064 3992
rect 78640 3952 78646 3964
rect 203058 3952 203064 3964
rect 203116 3952 203122 4004
rect 247586 3952 247592 4004
rect 247644 3992 247650 4004
rect 269853 3995 269911 4001
rect 269853 3992 269865 3995
rect 247644 3964 269865 3992
rect 247644 3952 247650 3964
rect 269853 3961 269865 3964
rect 269899 3961 269911 3995
rect 269853 3955 269911 3961
rect 269945 3995 270003 4001
rect 269945 3961 269957 3995
rect 269991 3992 270003 3995
rect 276198 3992 276204 4004
rect 269991 3964 276204 3992
rect 269991 3961 270003 3964
rect 269945 3955 270003 3961
rect 276198 3952 276204 3964
rect 276256 3952 276262 4004
rect 276293 3995 276351 4001
rect 276293 3961 276305 3995
rect 276339 3992 276351 3995
rect 278038 3992 278044 4004
rect 276339 3964 278044 3992
rect 276339 3961 276351 3964
rect 276293 3955 276351 3961
rect 278038 3952 278044 3964
rect 278096 3952 278102 4004
rect 317322 3952 317328 4004
rect 317380 3992 317386 4004
rect 333882 3992 333888 4004
rect 317380 3964 333888 3992
rect 317380 3952 317386 3964
rect 333882 3952 333888 3964
rect 333940 3952 333946 4004
rect 340782 3952 340788 4004
rect 340840 3992 340846 4004
rect 387150 3992 387156 4004
rect 340840 3964 387156 3992
rect 340840 3952 340846 3964
rect 387150 3952 387156 3964
rect 387208 3952 387214 4004
rect 413922 3952 413928 4004
rect 413980 3992 413986 4004
rect 550266 3992 550272 4004
rect 413980 3964 550272 3992
rect 413980 3952 413986 3964
rect 550266 3952 550272 3964
rect 550324 3952 550330 4004
rect 74994 3884 75000 3936
rect 75052 3924 75058 3936
rect 200114 3924 200120 3936
rect 75052 3896 200120 3924
rect 75052 3884 75058 3896
rect 200114 3884 200120 3896
rect 200172 3884 200178 3936
rect 246390 3884 246396 3936
rect 246448 3924 246454 3936
rect 272429 3927 272487 3933
rect 272429 3924 272441 3927
rect 246448 3896 272441 3924
rect 246448 3884 246454 3896
rect 272429 3893 272441 3896
rect 272475 3893 272487 3927
rect 272429 3887 272487 3893
rect 272613 3927 272671 3933
rect 272613 3893 272625 3927
rect 272659 3924 272671 3927
rect 277394 3924 277400 3936
rect 272659 3896 277400 3924
rect 272659 3893 272671 3896
rect 272613 3887 272671 3893
rect 277394 3884 277400 3896
rect 277452 3884 277458 3936
rect 278133 3927 278191 3933
rect 278133 3893 278145 3927
rect 278179 3924 278191 3927
rect 281718 3924 281724 3936
rect 278179 3896 281724 3924
rect 278179 3893 278191 3896
rect 278133 3887 278191 3893
rect 281718 3884 281724 3896
rect 281776 3884 281782 3936
rect 318058 3884 318064 3936
rect 318116 3924 318122 3936
rect 326798 3924 326804 3936
rect 318116 3896 326804 3924
rect 318116 3884 318122 3896
rect 326798 3884 326804 3896
rect 326856 3884 326862 3936
rect 342070 3884 342076 3936
rect 342128 3924 342134 3936
rect 390646 3924 390652 3936
rect 342128 3896 390652 3924
rect 342128 3884 342134 3896
rect 390646 3884 390652 3896
rect 390704 3884 390710 3936
rect 415302 3884 415308 3936
rect 415360 3924 415366 3936
rect 553762 3924 553768 3936
rect 415360 3896 553768 3924
rect 415360 3884 415366 3896
rect 553762 3884 553768 3896
rect 553820 3884 553826 3936
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 198734 3856 198740 3868
rect 71556 3828 198740 3856
rect 71556 3816 71562 3828
rect 198734 3816 198740 3828
rect 198792 3816 198798 3868
rect 245194 3816 245200 3868
rect 245252 3856 245258 3868
rect 272521 3859 272579 3865
rect 245252 3828 271920 3856
rect 245252 3816 245258 3828
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 39298 3788 39304 3800
rect 34848 3760 39304 3788
rect 34848 3748 34854 3760
rect 39298 3748 39304 3760
rect 39356 3748 39362 3800
rect 46658 3748 46664 3800
rect 46716 3788 46722 3800
rect 187694 3788 187700 3800
rect 46716 3760 187700 3788
rect 46716 3748 46722 3760
rect 187694 3748 187700 3760
rect 187752 3748 187758 3800
rect 242894 3748 242900 3800
rect 242952 3788 242958 3800
rect 269945 3791 270003 3797
rect 269945 3788 269957 3791
rect 242952 3760 269957 3788
rect 242952 3748 242958 3760
rect 269945 3757 269957 3760
rect 269991 3757 270003 3791
rect 269945 3751 270003 3757
rect 270034 3748 270040 3800
rect 270092 3788 270098 3800
rect 271785 3791 271843 3797
rect 271785 3788 271797 3791
rect 270092 3760 271797 3788
rect 270092 3748 270098 3760
rect 271785 3757 271797 3760
rect 271831 3757 271843 3791
rect 271892 3788 271920 3828
rect 272521 3825 272533 3859
rect 272567 3856 272579 3859
rect 278958 3856 278964 3868
rect 272567 3828 278964 3856
rect 272567 3825 272579 3828
rect 272521 3819 272579 3825
rect 278958 3816 278964 3828
rect 279016 3816 279022 3868
rect 283558 3856 283564 3868
rect 279436 3828 283564 3856
rect 276106 3788 276112 3800
rect 271892 3760 276112 3788
rect 271785 3751 271843 3757
rect 276106 3748 276112 3760
rect 276164 3748 276170 3800
rect 277026 3748 277032 3800
rect 277084 3788 277090 3800
rect 277302 3788 277308 3800
rect 277084 3760 277308 3788
rect 277084 3748 277090 3760
rect 277302 3748 277308 3760
rect 277360 3748 277366 3800
rect 43070 3680 43076 3732
rect 43128 3720 43134 3732
rect 186314 3720 186320 3732
rect 43128 3692 186320 3720
rect 43128 3680 43134 3692
rect 186314 3680 186320 3692
rect 186372 3680 186378 3732
rect 240502 3680 240508 3732
rect 240560 3720 240566 3732
rect 274818 3720 274824 3732
rect 240560 3692 274824 3720
rect 240560 3680 240566 3692
rect 274818 3680 274824 3692
rect 274876 3680 274882 3732
rect 274913 3723 274971 3729
rect 274913 3689 274925 3723
rect 274959 3720 274971 3723
rect 279436 3720 279464 3828
rect 283558 3816 283564 3828
rect 283616 3816 283622 3868
rect 322842 3816 322848 3868
rect 322900 3856 322906 3868
rect 325513 3859 325571 3865
rect 325513 3856 325525 3859
rect 322900 3828 325525 3856
rect 322900 3816 322906 3828
rect 325513 3825 325525 3828
rect 325559 3825 325571 3859
rect 325513 3819 325571 3825
rect 325602 3816 325608 3868
rect 325660 3856 325666 3868
rect 332686 3856 332692 3868
rect 325660 3828 332692 3856
rect 325660 3816 325666 3828
rect 332686 3816 332692 3828
rect 332744 3816 332750 3868
rect 343542 3816 343548 3868
rect 343600 3856 343606 3868
rect 394234 3856 394240 3868
rect 343600 3828 394240 3856
rect 343600 3816 343606 3828
rect 394234 3816 394240 3828
rect 394292 3816 394298 3868
rect 416590 3816 416596 3868
rect 416648 3856 416654 3868
rect 557350 3856 557356 3868
rect 416648 3828 557356 3856
rect 416648 3816 416654 3828
rect 557350 3816 557356 3828
rect 557408 3816 557414 3868
rect 283098 3748 283104 3800
rect 283156 3788 283162 3800
rect 294046 3788 294052 3800
rect 283156 3760 294052 3788
rect 283156 3748 283162 3760
rect 294046 3748 294052 3760
rect 294104 3748 294110 3800
rect 318702 3748 318708 3800
rect 318760 3788 318766 3800
rect 336274 3788 336280 3800
rect 318760 3760 336280 3788
rect 318760 3748 318766 3760
rect 336274 3748 336280 3760
rect 336332 3748 336338 3800
rect 346302 3748 346308 3800
rect 346360 3788 346366 3800
rect 397730 3788 397736 3800
rect 346360 3760 397736 3788
rect 346360 3748 346366 3760
rect 397730 3748 397736 3760
rect 397788 3748 397794 3800
rect 418062 3748 418068 3800
rect 418120 3788 418126 3800
rect 560846 3788 560852 3800
rect 418120 3760 560852 3788
rect 418120 3748 418126 3760
rect 560846 3748 560852 3760
rect 560904 3748 560910 3800
rect 274959 3692 279464 3720
rect 274959 3689 274971 3692
rect 274913 3683 274971 3689
rect 279510 3680 279516 3732
rect 279568 3720 279574 3732
rect 279568 3692 287054 3720
rect 279568 3680 279574 3692
rect 29638 3652 29644 3664
rect 26206 3624 29644 3652
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 26206 3584 26234 3624
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 184934 3652 184940 3664
rect 39632 3624 184940 3652
rect 39632 3612 39638 3624
rect 184934 3612 184940 3624
rect 184992 3612 184998 3664
rect 238110 3612 238116 3664
rect 238168 3652 238174 3664
rect 272429 3655 272487 3661
rect 238168 3624 270816 3652
rect 238168 3612 238174 3624
rect 19484 3556 26234 3584
rect 19484 3544 19490 3556
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 35158 3584 35164 3596
rect 28960 3556 35164 3584
rect 28960 3544 28966 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 183554 3584 183560 3596
rect 36044 3556 183560 3584
rect 36044 3544 36050 3556
rect 183554 3544 183560 3556
rect 183612 3544 183618 3596
rect 227530 3544 227536 3596
rect 227588 3584 227594 3596
rect 227588 3556 229094 3584
rect 227588 3544 227594 3556
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 22738 3516 22744 3528
rect 18288 3488 22744 3516
rect 18288 3476 18294 3488
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 23014 3476 23020 3528
rect 23072 3516 23078 3528
rect 25590 3516 25596 3528
rect 23072 3488 25596 3516
rect 23072 3476 23078 3488
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 32456 3488 171916 3516
rect 32456 3476 32462 3488
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 21358 3448 21364 3460
rect 13596 3420 21364 3448
rect 13596 3408 13602 3420
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 171781 3451 171839 3457
rect 171781 3448 171793 3451
rect 25372 3420 171793 3448
rect 25372 3408 25378 3420
rect 171781 3417 171793 3420
rect 171827 3417 171839 3451
rect 171888 3448 171916 3488
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 172422 3516 172428 3528
rect 172020 3488 172428 3516
rect 172020 3476 172026 3488
rect 172422 3476 172428 3488
rect 172480 3476 172486 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177942 3516 177948 3528
rect 176712 3488 177948 3516
rect 176712 3476 176718 3488
rect 177942 3476 177948 3488
rect 178000 3476 178006 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 181438 3476 181444 3528
rect 181496 3516 181502 3528
rect 182082 3516 182088 3528
rect 181496 3488 182088 3516
rect 181496 3476 181502 3488
rect 182082 3476 182088 3488
rect 182140 3476 182146 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 188522 3476 188528 3528
rect 188580 3516 188586 3528
rect 188982 3516 188988 3528
rect 188580 3488 188988 3516
rect 188580 3476 188586 3488
rect 188982 3476 188988 3488
rect 189040 3476 189046 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 193122 3516 193128 3528
rect 192076 3488 193128 3516
rect 192076 3476 192082 3488
rect 193122 3476 193128 3488
rect 193180 3476 193186 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 200022 3516 200028 3528
rect 199160 3488 200028 3516
rect 199160 3476 199166 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 209682 3516 209688 3528
rect 208636 3488 209688 3516
rect 208636 3476 208642 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 216582 3516 216588 3528
rect 215720 3488 216588 3516
rect 215720 3476 215726 3488
rect 216582 3476 216588 3488
rect 216640 3476 216646 3528
rect 216858 3476 216864 3528
rect 216916 3516 216922 3528
rect 217962 3516 217968 3528
rect 216916 3488 217968 3516
rect 216916 3476 216922 3488
rect 217962 3476 217968 3488
rect 218020 3476 218026 3528
rect 222746 3476 222752 3528
rect 222804 3516 222810 3528
rect 223482 3516 223488 3528
rect 222804 3488 223488 3516
rect 222804 3476 222810 3488
rect 223482 3476 223488 3488
rect 223540 3476 223546 3528
rect 226334 3476 226340 3528
rect 226392 3516 226398 3528
rect 227622 3516 227628 3528
rect 226392 3488 227628 3516
rect 226392 3476 226398 3488
rect 227622 3476 227628 3488
rect 227680 3476 227686 3528
rect 229066 3516 229094 3556
rect 229830 3544 229836 3596
rect 229888 3584 229894 3596
rect 230382 3584 230388 3596
rect 229888 3556 230388 3584
rect 229888 3544 229894 3556
rect 230382 3544 230388 3556
rect 230440 3544 230446 3596
rect 231026 3544 231032 3596
rect 231084 3584 231090 3596
rect 231762 3584 231768 3596
rect 231084 3556 231768 3584
rect 231084 3544 231090 3556
rect 231762 3544 231768 3556
rect 231820 3544 231826 3596
rect 232222 3544 232228 3596
rect 232280 3584 232286 3596
rect 233142 3584 233148 3596
rect 232280 3556 233148 3584
rect 232280 3544 232286 3556
rect 233142 3544 233148 3556
rect 233200 3544 233206 3596
rect 233418 3544 233424 3596
rect 233476 3584 233482 3596
rect 270678 3584 270684 3596
rect 233476 3556 270684 3584
rect 233476 3544 233482 3556
rect 270678 3544 270684 3556
rect 270736 3544 270742 3596
rect 270788 3584 270816 3624
rect 272429 3621 272441 3655
rect 272475 3652 272487 3655
rect 277486 3652 277492 3664
rect 272475 3624 277492 3652
rect 272475 3621 272487 3624
rect 272429 3615 272487 3621
rect 277486 3612 277492 3624
rect 277544 3612 277550 3664
rect 278041 3655 278099 3661
rect 278041 3621 278053 3655
rect 278087 3652 278099 3655
rect 280246 3652 280252 3664
rect 278087 3624 280252 3652
rect 278087 3621 278099 3624
rect 278041 3615 278099 3621
rect 280246 3612 280252 3624
rect 280304 3612 280310 3664
rect 284294 3612 284300 3664
rect 284352 3652 284358 3664
rect 285490 3652 285496 3664
rect 284352 3624 285496 3652
rect 284352 3612 284358 3624
rect 285490 3612 285496 3624
rect 285548 3612 285554 3664
rect 287026 3652 287054 3692
rect 321462 3680 321468 3732
rect 321520 3720 321526 3732
rect 325605 3723 325663 3729
rect 321520 3692 325556 3720
rect 321520 3680 321526 3692
rect 291286 3652 291292 3664
rect 287026 3624 291292 3652
rect 291286 3612 291292 3624
rect 291344 3612 291350 3664
rect 313918 3612 313924 3664
rect 313976 3652 313982 3664
rect 319714 3652 319720 3664
rect 313976 3624 319720 3652
rect 313976 3612 313982 3624
rect 319714 3612 319720 3624
rect 319772 3612 319778 3664
rect 325528 3652 325556 3692
rect 325605 3689 325617 3723
rect 325651 3720 325663 3723
rect 337470 3720 337476 3732
rect 325651 3692 337476 3720
rect 325651 3689 325663 3692
rect 325605 3683 325663 3689
rect 337470 3680 337476 3692
rect 337528 3680 337534 3732
rect 347682 3680 347688 3732
rect 347740 3720 347746 3732
rect 401318 3720 401324 3732
rect 347740 3692 401324 3720
rect 347740 3680 347746 3692
rect 401318 3680 401324 3692
rect 401376 3680 401382 3732
rect 419442 3680 419448 3732
rect 419500 3720 419506 3732
rect 564434 3720 564440 3732
rect 419500 3692 564440 3720
rect 419500 3680 419506 3692
rect 564434 3680 564440 3692
rect 564492 3680 564498 3732
rect 344554 3652 344560 3664
rect 325528 3624 344560 3652
rect 344554 3612 344560 3624
rect 344612 3612 344618 3664
rect 349062 3612 349068 3664
rect 349120 3652 349126 3664
rect 404814 3652 404820 3664
rect 349120 3624 404820 3652
rect 349120 3612 349126 3624
rect 404814 3612 404820 3624
rect 404872 3612 404878 3664
rect 420822 3612 420828 3664
rect 420880 3652 420886 3664
rect 568022 3652 568028 3664
rect 420880 3624 568028 3652
rect 420880 3612 420886 3624
rect 568022 3612 568028 3624
rect 568080 3612 568086 3664
rect 273346 3584 273352 3596
rect 270788 3556 273352 3584
rect 273346 3544 273352 3556
rect 273404 3544 273410 3596
rect 274913 3587 274971 3593
rect 274913 3584 274925 3587
rect 273456 3556 274925 3584
rect 258169 3519 258227 3525
rect 258169 3516 258181 3519
rect 229066 3488 258181 3516
rect 258169 3485 258181 3488
rect 258215 3485 258227 3519
rect 258169 3479 258227 3485
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 267734 3476 267740 3528
rect 267792 3516 267798 3528
rect 269022 3516 269028 3528
rect 267792 3488 269028 3516
rect 267792 3476 267798 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 271782 3516 271788 3528
rect 271288 3488 271788 3516
rect 271288 3476 271294 3488
rect 271782 3476 271788 3488
rect 271840 3476 271846 3528
rect 271877 3519 271935 3525
rect 271877 3485 271889 3519
rect 271923 3516 271935 3519
rect 272613 3519 272671 3525
rect 272613 3516 272625 3519
rect 271923 3488 272625 3516
rect 271923 3485 271935 3488
rect 271877 3479 271935 3485
rect 272613 3485 272625 3488
rect 272659 3485 272671 3519
rect 272613 3479 272671 3485
rect 272702 3476 272708 3528
rect 272760 3516 272766 3528
rect 273456 3516 273484 3556
rect 274913 3553 274925 3556
rect 274959 3553 274971 3587
rect 274913 3547 274971 3553
rect 275002 3544 275008 3596
rect 275060 3584 275066 3596
rect 275925 3587 275983 3593
rect 275925 3584 275937 3587
rect 275060 3556 275937 3584
rect 275060 3544 275066 3556
rect 275925 3553 275937 3556
rect 275971 3553 275983 3587
rect 275925 3547 275983 3553
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 288526 3584 288532 3596
rect 277228 3556 288532 3584
rect 272760 3488 273484 3516
rect 272760 3476 272766 3488
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 277228 3516 277256 3556
rect 288526 3544 288532 3556
rect 288584 3544 288590 3596
rect 306190 3544 306196 3596
rect 306248 3584 306254 3596
rect 307938 3584 307944 3596
rect 306248 3556 307944 3584
rect 306248 3544 306254 3556
rect 307938 3544 307944 3556
rect 307996 3544 308002 3596
rect 325418 3544 325424 3596
rect 325476 3544 325482 3596
rect 325513 3587 325571 3593
rect 325513 3553 325525 3587
rect 325559 3584 325571 3587
rect 348050 3584 348056 3596
rect 325559 3556 348056 3584
rect 325559 3553 325571 3556
rect 325513 3547 325571 3553
rect 348050 3544 348056 3556
rect 348108 3544 348114 3596
rect 351822 3544 351828 3596
rect 351880 3584 351886 3596
rect 411898 3584 411904 3596
rect 351880 3556 411904 3584
rect 351880 3544 351886 3556
rect 411898 3544 411904 3556
rect 411956 3544 411962 3596
rect 423582 3544 423588 3596
rect 423640 3584 423646 3596
rect 571518 3584 571524 3596
rect 423640 3556 571524 3584
rect 423640 3544 423646 3556
rect 571518 3544 571524 3556
rect 571576 3544 571582 3596
rect 273680 3488 277256 3516
rect 277305 3519 277363 3525
rect 273680 3476 273686 3488
rect 277305 3485 277317 3519
rect 277351 3516 277363 3519
rect 287330 3516 287336 3528
rect 277351 3488 287336 3516
rect 277351 3485 277363 3488
rect 277305 3479 277363 3485
rect 287330 3476 287336 3488
rect 287388 3476 287394 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 292482 3516 292488 3528
rect 291436 3488 292488 3516
rect 291436 3476 291442 3488
rect 292482 3476 292488 3488
rect 292540 3476 292546 3528
rect 293678 3476 293684 3528
rect 293736 3516 293742 3528
rect 294598 3516 294604 3528
rect 293736 3488 294604 3516
rect 293736 3476 293742 3488
rect 294598 3476 294604 3488
rect 294656 3476 294662 3528
rect 296070 3476 296076 3528
rect 296128 3516 296134 3528
rect 296622 3516 296628 3528
rect 296128 3488 296628 3516
rect 296128 3476 296134 3488
rect 296622 3476 296628 3488
rect 296680 3476 296686 3528
rect 298462 3476 298468 3528
rect 298520 3516 298526 3528
rect 299382 3516 299388 3528
rect 298520 3488 299388 3516
rect 298520 3476 298526 3488
rect 299382 3476 299388 3488
rect 299440 3476 299446 3528
rect 302326 3476 302332 3528
rect 302384 3516 302390 3528
rect 303154 3516 303160 3528
rect 302384 3488 303160 3516
rect 302384 3476 302390 3488
rect 303154 3476 303160 3488
rect 303212 3476 303218 3528
rect 304902 3476 304908 3528
rect 304960 3516 304966 3528
rect 305546 3516 305552 3528
rect 304960 3488 305552 3516
rect 304960 3476 304966 3488
rect 305546 3476 305552 3488
rect 305604 3476 305610 3528
rect 313182 3476 313188 3528
rect 313240 3516 313246 3528
rect 324406 3516 324412 3528
rect 313240 3488 324412 3516
rect 313240 3476 313246 3488
rect 324406 3476 324412 3488
rect 324464 3476 324470 3528
rect 325436 3516 325464 3544
rect 351638 3516 351644 3528
rect 325436 3488 351644 3516
rect 351638 3476 351644 3488
rect 351696 3476 351702 3528
rect 354582 3476 354588 3528
rect 354640 3516 354646 3528
rect 418982 3516 418988 3528
rect 354640 3488 418988 3516
rect 354640 3476 354646 3488
rect 418982 3476 418988 3488
rect 419040 3476 419046 3528
rect 424686 3476 424692 3528
rect 424744 3516 424750 3528
rect 575106 3516 575112 3528
rect 424744 3488 575112 3516
rect 424744 3476 424750 3488
rect 575106 3476 575112 3488
rect 575164 3476 575170 3528
rect 182358 3448 182364 3460
rect 171888 3420 182364 3448
rect 171781 3411 171839 3417
rect 182358 3408 182364 3420
rect 182416 3408 182422 3460
rect 206186 3408 206192 3460
rect 206244 3448 206250 3460
rect 206922 3448 206928 3460
rect 206244 3420 206928 3448
rect 206244 3408 206250 3420
rect 206922 3408 206928 3420
rect 206980 3408 206986 3460
rect 209774 3408 209780 3460
rect 209832 3448 209838 3460
rect 260834 3448 260840 3460
rect 209832 3420 260840 3448
rect 209832 3408 209838 3420
rect 260834 3408 260840 3420
rect 260892 3408 260898 3460
rect 261754 3408 261760 3460
rect 261812 3448 261818 3460
rect 261812 3420 280568 3448
rect 261812 3408 261818 3420
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 50982 3380 50988 3392
rect 50212 3352 50988 3380
rect 50212 3340 50218 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 57882 3380 57888 3392
rect 57296 3352 57888 3380
rect 57296 3340 57302 3352
rect 57882 3340 57888 3352
rect 57940 3340 57946 3392
rect 60826 3340 60832 3392
rect 60884 3380 60890 3392
rect 61930 3380 61936 3392
rect 60884 3352 61936 3380
rect 60884 3340 60890 3352
rect 61930 3340 61936 3352
rect 61988 3340 61994 3392
rect 64322 3340 64328 3392
rect 64380 3380 64386 3392
rect 64782 3380 64788 3392
rect 64380 3352 64788 3380
rect 64380 3340 64386 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 68922 3380 68928 3392
rect 67968 3352 68928 3380
rect 67968 3340 67974 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 85482 3380 85488 3392
rect 84528 3352 85488 3380
rect 84528 3340 84534 3352
rect 85482 3340 85488 3352
rect 85540 3340 85546 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 92382 3380 92388 3392
rect 91612 3352 92388 3380
rect 91612 3340 91618 3352
rect 92382 3340 92388 3352
rect 92440 3340 92446 3392
rect 207290 3380 207296 3392
rect 92492 3352 207296 3380
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 92492 3312 92520 3352
rect 207290 3340 207296 3352
rect 207348 3340 207354 3392
rect 241698 3340 241704 3392
rect 241756 3380 241762 3392
rect 242802 3380 242808 3392
rect 241756 3352 242808 3380
rect 241756 3340 241762 3352
rect 242802 3340 242808 3352
rect 242860 3340 242866 3392
rect 249978 3340 249984 3392
rect 250036 3380 250042 3392
rect 251082 3380 251088 3392
rect 250036 3352 251088 3380
rect 250036 3340 250042 3352
rect 251082 3340 251088 3352
rect 251140 3340 251146 3392
rect 251174 3340 251180 3392
rect 251232 3380 251238 3392
rect 272521 3383 272579 3389
rect 272521 3380 272533 3383
rect 251232 3352 272533 3380
rect 251232 3340 251238 3352
rect 272521 3349 272533 3352
rect 272567 3349 272579 3383
rect 272521 3343 272579 3349
rect 272613 3383 272671 3389
rect 272613 3349 272625 3383
rect 272659 3380 272671 3383
rect 277213 3383 277271 3389
rect 277213 3380 277225 3383
rect 272659 3352 277225 3380
rect 272659 3349 272671 3352
rect 272613 3343 272671 3349
rect 277213 3349 277225 3352
rect 277259 3349 277271 3383
rect 277213 3343 277271 3349
rect 277302 3340 277308 3392
rect 277360 3380 277366 3392
rect 277578 3380 277584 3392
rect 277360 3352 277584 3380
rect 277360 3340 277366 3352
rect 277578 3340 277584 3352
rect 277636 3340 277642 3392
rect 89220 3284 92520 3312
rect 89220 3272 89226 3284
rect 92750 3272 92756 3324
rect 92808 3312 92814 3324
rect 208670 3312 208676 3324
rect 92808 3284 208676 3312
rect 92808 3272 92814 3284
rect 208670 3272 208676 3284
rect 208728 3272 208734 3324
rect 254670 3272 254676 3324
rect 254728 3312 254734 3324
rect 278041 3315 278099 3321
rect 278041 3312 278053 3315
rect 254728 3284 278053 3312
rect 254728 3272 254734 3284
rect 278041 3281 278053 3284
rect 278087 3281 278099 3315
rect 280540 3312 280568 3420
rect 280706 3408 280712 3460
rect 280764 3448 280770 3460
rect 281442 3448 281448 3460
rect 280764 3420 281448 3448
rect 280764 3408 280770 3420
rect 281442 3408 281448 3420
rect 281500 3408 281506 3460
rect 281902 3408 281908 3460
rect 281960 3448 281966 3460
rect 282822 3448 282828 3460
rect 281960 3420 282828 3448
rect 281960 3408 281966 3420
rect 282822 3408 282828 3420
rect 282880 3408 282886 3460
rect 290182 3408 290188 3460
rect 290240 3448 290246 3460
rect 291838 3448 291844 3460
rect 290240 3420 291844 3448
rect 290240 3408 290246 3420
rect 291838 3408 291844 3420
rect 291896 3408 291902 3460
rect 314562 3408 314568 3460
rect 314620 3448 314626 3460
rect 327994 3448 328000 3460
rect 314620 3420 328000 3448
rect 314620 3408 314626 3420
rect 327994 3408 328000 3420
rect 328052 3408 328058 3460
rect 328178 3408 328184 3460
rect 328236 3448 328242 3460
rect 358722 3448 358728 3460
rect 328236 3420 358728 3448
rect 328236 3408 328242 3420
rect 358722 3408 358728 3420
rect 358780 3408 358786 3460
rect 358814 3408 358820 3460
rect 358872 3448 358878 3460
rect 426158 3448 426164 3460
rect 358872 3420 426164 3448
rect 358872 3408 358878 3420
rect 426158 3408 426164 3420
rect 426216 3408 426222 3460
rect 426250 3408 426256 3460
rect 426308 3448 426314 3460
rect 578602 3448 578608 3460
rect 426308 3420 578608 3448
rect 426308 3408 426314 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 287790 3340 287796 3392
rect 287848 3380 287854 3392
rect 295426 3380 295432 3392
rect 287848 3352 295432 3380
rect 287848 3340 287854 3352
rect 295426 3340 295432 3352
rect 295484 3340 295490 3392
rect 310422 3340 310428 3392
rect 310480 3380 310486 3392
rect 317322 3380 317328 3392
rect 310480 3352 317328 3380
rect 310480 3340 310486 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 327718 3340 327724 3392
rect 327776 3380 327782 3392
rect 329190 3380 329196 3392
rect 327776 3352 329196 3380
rect 327776 3340 327782 3352
rect 329190 3340 329196 3352
rect 329248 3340 329254 3392
rect 336642 3340 336648 3392
rect 336700 3380 336706 3392
rect 376478 3380 376484 3392
rect 336700 3352 376484 3380
rect 336700 3340 336706 3352
rect 376478 3340 376484 3352
rect 376536 3340 376542 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 408494 3340 408500 3392
rect 408552 3380 408558 3392
rect 539594 3380 539600 3392
rect 408552 3352 539600 3380
rect 408552 3340 408558 3352
rect 539594 3340 539600 3352
rect 539652 3340 539658 3392
rect 284570 3312 284576 3324
rect 280540 3284 284576 3312
rect 278041 3275 278099 3281
rect 284570 3272 284576 3284
rect 284628 3272 284634 3324
rect 311158 3272 311164 3324
rect 311216 3312 311222 3324
rect 315022 3312 315028 3324
rect 311216 3284 315028 3312
rect 311216 3272 311222 3284
rect 315022 3272 315028 3284
rect 315080 3272 315086 3324
rect 335262 3272 335268 3324
rect 335320 3312 335326 3324
rect 372890 3312 372896 3324
rect 335320 3284 372896 3312
rect 335320 3272 335326 3284
rect 372890 3272 372896 3284
rect 372948 3272 372954 3324
rect 373994 3272 374000 3324
rect 374052 3312 374058 3324
rect 375282 3312 375288 3324
rect 374052 3284 375288 3312
rect 374052 3272 374058 3284
rect 375282 3272 375288 3284
rect 375340 3272 375346 3324
rect 380802 3272 380808 3324
rect 380860 3312 380866 3324
rect 380860 3284 470594 3312
rect 380860 3272 380866 3284
rect 31294 3204 31300 3256
rect 31352 3244 31358 3256
rect 36538 3244 36544 3256
rect 31352 3216 36544 3244
rect 31352 3204 31358 3216
rect 36538 3204 36544 3216
rect 36596 3204 36602 3256
rect 98638 3204 98644 3256
rect 98696 3244 98702 3256
rect 99282 3244 99288 3256
rect 98696 3216 99288 3244
rect 98696 3204 98702 3216
rect 99282 3204 99288 3216
rect 99340 3204 99346 3256
rect 209958 3244 209964 3256
rect 99392 3216 209964 3244
rect 41874 3136 41880 3188
rect 41932 3176 41938 3188
rect 43438 3176 43444 3188
rect 41932 3148 43444 3176
rect 41932 3136 41938 3148
rect 43438 3136 43444 3148
rect 43496 3136 43502 3188
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 99392 3176 99420 3216
rect 209958 3204 209964 3216
rect 210016 3204 210022 3256
rect 255866 3204 255872 3256
rect 255924 3244 255930 3256
rect 278133 3247 278191 3253
rect 278133 3244 278145 3247
rect 255924 3216 278145 3244
rect 255924 3204 255930 3216
rect 278133 3213 278145 3216
rect 278179 3213 278191 3247
rect 281626 3244 281632 3256
rect 278133 3207 278191 3213
rect 278240 3216 281632 3244
rect 96304 3148 99420 3176
rect 96304 3136 96310 3148
rect 102226 3136 102232 3188
rect 102284 3176 102290 3188
rect 103422 3176 103428 3188
rect 102284 3148 103428 3176
rect 102284 3136 102290 3148
rect 103422 3136 103428 3148
rect 103480 3136 103486 3188
rect 105722 3136 105728 3188
rect 105780 3176 105786 3188
rect 106182 3176 106188 3188
rect 105780 3148 106188 3176
rect 105780 3136 105786 3148
rect 106182 3136 106188 3148
rect 106240 3136 106246 3188
rect 109310 3136 109316 3188
rect 109368 3176 109374 3188
rect 110322 3176 110328 3188
rect 109368 3148 110328 3176
rect 109368 3136 109374 3148
rect 110322 3136 110328 3148
rect 110380 3136 110386 3188
rect 110417 3179 110475 3185
rect 110417 3145 110429 3179
rect 110463 3176 110475 3179
rect 211338 3176 211344 3188
rect 110463 3148 211344 3176
rect 110463 3145 110475 3148
rect 110417 3139 110475 3145
rect 211338 3136 211344 3148
rect 211396 3136 211402 3188
rect 257062 3136 257068 3188
rect 257120 3176 257126 3188
rect 278240 3176 278268 3216
rect 281626 3204 281632 3216
rect 281684 3204 281690 3256
rect 299658 3204 299664 3256
rect 299716 3244 299722 3256
rect 300946 3244 300952 3256
rect 299716 3216 300952 3244
rect 299716 3204 299722 3216
rect 300946 3204 300952 3216
rect 301004 3204 301010 3256
rect 307662 3204 307668 3256
rect 307720 3244 307726 3256
rect 311434 3244 311440 3256
rect 307720 3216 311440 3244
rect 307720 3204 307726 3216
rect 311434 3204 311440 3216
rect 311492 3204 311498 3256
rect 332502 3204 332508 3256
rect 332560 3244 332566 3256
rect 369394 3244 369400 3256
rect 332560 3216 369400 3244
rect 332560 3204 332566 3216
rect 369394 3204 369400 3216
rect 369452 3204 369458 3256
rect 376662 3204 376668 3256
rect 376720 3244 376726 3256
rect 468662 3244 468668 3256
rect 376720 3216 468668 3244
rect 376720 3204 376726 3216
rect 468662 3204 468668 3216
rect 468720 3204 468726 3256
rect 470566 3244 470594 3284
rect 473354 3272 473360 3324
rect 473412 3312 473418 3324
rect 474550 3312 474556 3324
rect 473412 3284 474556 3312
rect 473412 3272 473418 3284
rect 474550 3272 474556 3284
rect 474608 3272 474614 3324
rect 481634 3272 481640 3324
rect 481692 3312 481698 3324
rect 482830 3312 482836 3324
rect 481692 3284 482836 3312
rect 481692 3272 481698 3284
rect 482830 3272 482836 3284
rect 482888 3272 482894 3324
rect 489914 3272 489920 3324
rect 489972 3312 489978 3324
rect 491110 3312 491116 3324
rect 489972 3284 491116 3312
rect 489972 3272 489978 3284
rect 491110 3272 491116 3284
rect 491168 3272 491174 3324
rect 506474 3272 506480 3324
rect 506532 3312 506538 3324
rect 507670 3312 507676 3324
rect 506532 3284 507676 3312
rect 506532 3272 506538 3284
rect 507670 3272 507676 3284
rect 507728 3272 507734 3324
rect 531314 3272 531320 3324
rect 531372 3312 531378 3324
rect 532510 3312 532516 3324
rect 531372 3284 532516 3312
rect 531372 3272 531378 3284
rect 532510 3272 532516 3284
rect 532568 3272 532574 3324
rect 475746 3244 475752 3256
rect 470566 3216 475752 3244
rect 475746 3204 475752 3216
rect 475804 3204 475810 3256
rect 257120 3148 278268 3176
rect 257120 3136 257126 3148
rect 278314 3136 278320 3188
rect 278372 3176 278378 3188
rect 280798 3176 280804 3188
rect 278372 3148 280804 3176
rect 278372 3136 278378 3148
rect 280798 3136 280804 3148
rect 280856 3136 280862 3188
rect 297266 3136 297272 3188
rect 297324 3176 297330 3188
rect 299750 3176 299756 3188
rect 297324 3148 299756 3176
rect 297324 3136 297330 3148
rect 299750 3136 299756 3148
rect 299808 3136 299814 3188
rect 331122 3136 331128 3188
rect 331180 3176 331186 3188
rect 365806 3176 365812 3188
rect 331180 3148 365812 3176
rect 331180 3136 331186 3148
rect 365806 3136 365812 3148
rect 365864 3136 365870 3188
rect 373718 3136 373724 3188
rect 373776 3176 373782 3188
rect 461578 3176 461584 3188
rect 373776 3148 461584 3176
rect 373776 3136 373782 3148
rect 461578 3136 461584 3148
rect 461636 3136 461642 3188
rect 38378 3068 38384 3120
rect 38436 3108 38442 3120
rect 40678 3108 40684 3120
rect 38436 3080 40684 3108
rect 38436 3068 38442 3080
rect 40678 3068 40684 3080
rect 40736 3068 40742 3120
rect 103330 3068 103336 3120
rect 103388 3108 103394 3120
rect 214190 3108 214196 3120
rect 103388 3080 214196 3108
rect 103388 3068 103394 3080
rect 214190 3068 214196 3080
rect 214248 3068 214254 3120
rect 259454 3068 259460 3120
rect 259512 3108 259518 3120
rect 283006 3108 283012 3120
rect 259512 3080 283012 3108
rect 259512 3068 259518 3080
rect 283006 3068 283012 3080
rect 283064 3068 283070 3120
rect 329742 3068 329748 3120
rect 329800 3108 329806 3120
rect 362310 3108 362316 3120
rect 329800 3080 362316 3108
rect 329800 3068 329806 3080
rect 362310 3068 362316 3080
rect 362368 3068 362374 3120
rect 371142 3068 371148 3120
rect 371200 3108 371206 3120
rect 454494 3108 454500 3120
rect 371200 3080 454500 3108
rect 371200 3068 371206 3080
rect 454494 3068 454500 3080
rect 454552 3068 454558 3120
rect 456794 3068 456800 3120
rect 456852 3108 456858 3120
rect 458082 3108 458088 3120
rect 456852 3080 458088 3108
rect 456852 3068 456858 3080
rect 458082 3068 458088 3080
rect 458140 3068 458146 3120
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 18598 3040 18604 3052
rect 11204 3012 18604 3040
rect 11204 3000 11210 3012
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 33778 3040 33784 3052
rect 27764 3012 33784 3040
rect 27764 3000 27770 3012
rect 33778 3000 33784 3012
rect 33836 3000 33842 3052
rect 99834 3000 99840 3052
rect 99892 3040 99898 3052
rect 110417 3043 110475 3049
rect 110417 3040 110429 3043
rect 99892 3012 110429 3040
rect 99892 3000 99898 3012
rect 110417 3009 110429 3012
rect 110463 3009 110475 3043
rect 110417 3003 110475 3009
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 114462 3040 114468 3052
rect 114060 3012 114468 3040
rect 114060 3000 114066 3012
rect 114462 3000 114468 3012
rect 114520 3000 114526 3052
rect 116394 3000 116400 3052
rect 116452 3040 116458 3052
rect 117222 3040 117228 3052
rect 116452 3012 117228 3040
rect 116452 3000 116458 3012
rect 117222 3000 117228 3012
rect 117280 3000 117286 3052
rect 117961 3043 118019 3049
rect 117961 3009 117973 3043
rect 118007 3040 118019 3043
rect 215478 3040 215484 3052
rect 118007 3012 215484 3040
rect 118007 3009 118019 3012
rect 117961 3003 118019 3009
rect 215478 3000 215484 3012
rect 215536 3000 215542 3052
rect 262950 3000 262956 3052
rect 263008 3040 263014 3052
rect 284478 3040 284484 3052
rect 263008 3012 284484 3040
rect 263008 3000 263014 3012
rect 284478 3000 284484 3012
rect 284536 3000 284542 3052
rect 292574 3000 292580 3052
rect 292632 3040 292638 3052
rect 298186 3040 298192 3052
rect 292632 3012 298192 3040
rect 292632 3000 292638 3012
rect 298186 3000 298192 3012
rect 298244 3000 298250 3052
rect 310330 3000 310336 3052
rect 310388 3040 310394 3052
rect 316218 3040 316224 3052
rect 310388 3012 316224 3040
rect 310388 3000 310394 3012
rect 316218 3000 316224 3012
rect 316276 3000 316282 3052
rect 326982 3000 326988 3052
rect 327040 3040 327046 3052
rect 355226 3040 355232 3052
rect 327040 3012 355232 3040
rect 327040 3000 327046 3012
rect 355226 3000 355232 3012
rect 355284 3000 355290 3052
rect 368382 3000 368388 3052
rect 368440 3040 368446 3052
rect 447410 3040 447416 3052
rect 368440 3012 447416 3040
rect 368440 3000 368446 3012
rect 447410 3000 447416 3012
rect 447468 3000 447474 3052
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 11698 2972 11704 2984
rect 10008 2944 11704 2972
rect 10008 2932 10014 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 216766 2972 216772 2984
rect 110564 2944 216772 2972
rect 110564 2932 110570 2944
rect 216766 2932 216772 2944
rect 216824 2932 216830 2984
rect 223942 2932 223948 2984
rect 224000 2972 224006 2984
rect 224862 2972 224868 2984
rect 224000 2944 224868 2972
rect 224000 2932 224006 2944
rect 224862 2932 224868 2944
rect 224920 2932 224926 2984
rect 265342 2932 265348 2984
rect 265400 2972 265406 2984
rect 285766 2972 285772 2984
rect 265400 2944 285772 2972
rect 265400 2932 265406 2944
rect 285766 2932 285772 2944
rect 285824 2932 285830 2984
rect 364242 2932 364248 2984
rect 364300 2972 364306 2984
rect 440234 2972 440240 2984
rect 364300 2944 440240 2972
rect 364300 2932 364306 2944
rect 440234 2932 440240 2944
rect 440292 2932 440298 2984
rect 440326 2932 440332 2984
rect 440384 2972 440390 2984
rect 441522 2972 441528 2984
rect 440384 2944 441528 2972
rect 440384 2932 440390 2944
rect 441522 2932 441528 2944
rect 441580 2932 441586 2984
rect 106918 2864 106924 2916
rect 106976 2904 106982 2916
rect 117961 2907 118019 2913
rect 117961 2904 117973 2907
rect 106976 2876 117973 2904
rect 106976 2864 106982 2876
rect 117961 2873 117973 2876
rect 118007 2873 118019 2907
rect 219618 2904 219624 2916
rect 117961 2867 118019 2873
rect 118068 2876 219624 2904
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 118068 2836 118096 2876
rect 219618 2864 219624 2876
rect 219676 2864 219682 2916
rect 258169 2907 258227 2913
rect 258169 2873 258181 2907
rect 258215 2904 258227 2907
rect 268746 2904 268752 2916
rect 258215 2876 268752 2904
rect 258215 2873 258227 2876
rect 258169 2867 258227 2873
rect 268746 2864 268752 2876
rect 268804 2864 268810 2916
rect 268838 2864 268844 2916
rect 268896 2904 268902 2916
rect 287146 2904 287152 2916
rect 268896 2876 287152 2904
rect 268896 2864 268902 2876
rect 287146 2864 287152 2876
rect 287204 2864 287210 2916
rect 361482 2864 361488 2916
rect 361540 2904 361546 2916
rect 433242 2904 433248 2916
rect 361540 2876 433248 2904
rect 361540 2864 361546 2876
rect 433242 2864 433248 2876
rect 433300 2864 433306 2916
rect 117648 2808 118096 2836
rect 117648 2796 117654 2808
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 221090 2836 221096 2848
rect 121144 2808 221096 2836
rect 121144 2796 121150 2808
rect 221090 2796 221096 2808
rect 221148 2796 221154 2848
rect 266538 2796 266544 2848
rect 266596 2836 266602 2848
rect 285858 2836 285864 2848
rect 266596 2808 285864 2836
rect 266596 2796 266602 2808
rect 285858 2796 285864 2808
rect 285916 2796 285922 2848
rect 360102 2796 360108 2848
rect 360160 2836 360166 2848
rect 429654 2836 429660 2848
rect 360160 2808 429660 2836
rect 360160 2796 360166 2808
rect 429654 2796 429660 2808
rect 429712 2796 429718 2848
<< via1 >>
rect 360108 700884 360160 700936
rect 429844 700884 429896 700936
rect 367008 700816 367060 700868
rect 446128 700816 446180 700868
rect 373908 700748 373960 700800
rect 462320 700748 462372 700800
rect 382188 700680 382240 700732
rect 478512 700680 478564 700732
rect 389088 700612 389140 700664
rect 494796 700612 494848 700664
rect 395988 700544 396040 700596
rect 510988 700544 511040 700596
rect 331128 700476 331180 700528
rect 364984 700476 365036 700528
rect 402888 700476 402940 700528
rect 527180 700476 527232 700528
rect 338028 700408 338080 700460
rect 381176 700408 381228 700460
rect 411168 700408 411220 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 235172 700340 235224 700392
rect 235908 700340 235960 700392
rect 317328 700340 317380 700392
rect 332508 700340 332560 700392
rect 344928 700340 344980 700392
rect 397460 700340 397512 700392
rect 418068 700340 418120 700392
rect 559656 700340 559708 700392
rect 324228 700272 324280 700324
rect 348792 700272 348844 700324
rect 353208 700272 353260 700324
rect 413652 700272 413704 700324
rect 424968 700272 425020 700324
rect 575848 700272 575900 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 56784 700136 56836 700188
rect 57888 700136 57940 700188
rect 186504 700136 186556 700188
rect 187608 700136 187660 700188
rect 251456 700068 251508 700120
rect 252468 700068 252520 700120
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 121644 699660 121696 699712
rect 122748 699660 122800 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 309784 699660 309836 699712
rect 316316 699660 316368 699712
rect 429844 696940 429896 696992
rect 580172 696940 580224 696992
rect 429936 683136 429988 683188
rect 580172 683136 580224 683188
rect 430028 670692 430080 670744
rect 580172 670692 580224 670744
rect 430120 643084 430172 643136
rect 580172 643084 580224 643136
rect 430212 630640 430264 630692
rect 579988 630640 580040 630692
rect 430304 616836 430356 616888
rect 580172 616836 580224 616888
rect 430396 590656 430448 590708
rect 579620 590656 579672 590708
rect 430488 576852 430540 576904
rect 579620 576852 579672 576904
rect 429752 563048 429804 563100
rect 579896 563048 579948 563100
rect 429660 536800 429712 536852
rect 580172 536800 580224 536852
rect 429568 524424 429620 524476
rect 580172 524424 580224 524476
rect 171048 500896 171100 500948
rect 243820 500896 243872 500948
rect 300768 500896 300820 500948
rect 301596 500896 301648 500948
rect 308772 500896 308824 500948
rect 309784 500896 309836 500948
rect 359372 500896 359424 500948
rect 360108 500896 360160 500948
rect 380992 500896 381044 500948
rect 382188 500896 382240 500948
rect 388260 500896 388312 500948
rect 389088 500896 389140 500948
rect 417148 500896 417200 500948
rect 418068 500896 418120 500948
rect 154488 500828 154540 500880
rect 236552 500828 236604 500880
rect 137928 500760 137980 500812
rect 229376 500760 229428 500812
rect 122748 500692 122800 500744
rect 222108 500692 222160 500744
rect 106188 500624 106240 500676
rect 214932 500624 214984 500676
rect 89628 500556 89680 500608
rect 207664 500556 207716 500608
rect 316040 500556 316092 500608
rect 317328 500556 317380 500608
rect 409880 500556 409932 500608
rect 411168 500556 411220 500608
rect 73068 500488 73120 500540
rect 200488 500488 200540 500540
rect 323216 500488 323268 500540
rect 324228 500488 324280 500540
rect 57888 500420 57940 500472
rect 193220 500420 193272 500472
rect 235908 500420 235960 500472
rect 272708 500420 272760 500472
rect 352104 500420 352156 500472
rect 353208 500420 353260 500472
rect 41328 500352 41380 500404
rect 186044 500352 186096 500404
rect 219348 500352 219400 500404
rect 265440 500352 265492 500404
rect 24768 500284 24820 500336
rect 178776 500284 178828 500336
rect 202788 500284 202840 500336
rect 258264 500284 258316 500336
rect 267648 500284 267700 500336
rect 287152 500284 287204 500336
rect 8208 500216 8260 500268
rect 171600 500216 171652 500268
rect 187608 500216 187660 500268
rect 250996 500216 251048 500268
rect 252468 500216 252520 500268
rect 279884 500216 279936 500268
rect 284208 500216 284260 500268
rect 294328 500216 294380 500268
rect 3424 493960 3476 494012
rect 165620 493960 165672 494012
rect 3516 491240 3568 491292
rect 165620 491240 165672 491292
rect 3608 488452 3660 488504
rect 165620 488452 165672 488504
rect 429384 488452 429436 488504
rect 580264 488452 580316 488504
rect 3700 485732 3752 485784
rect 165620 485732 165672 485784
rect 429844 484372 429896 484424
rect 579620 484372 579672 484424
rect 3792 481584 3844 481636
rect 165620 481584 165672 481636
rect 3884 478796 3936 478848
rect 165620 478796 165672 478848
rect 3976 476008 4028 476060
rect 165620 476008 165672 476060
rect 429476 476008 429528 476060
rect 580356 476008 580408 476060
rect 4068 473288 4120 473340
rect 165620 473288 165672 473340
rect 429936 470568 429988 470620
rect 579620 470568 579672 470620
rect 3332 470500 3384 470552
rect 165620 470500 165672 470552
rect 3240 467780 3292 467832
rect 165620 467780 165672 467832
rect 3148 464992 3200 465044
rect 165620 464992 165672 465044
rect 429200 463632 429252 463684
rect 580448 463632 580500 463684
rect 3056 460844 3108 460896
rect 165620 460844 165672 460896
rect 2964 458124 3016 458176
rect 165620 458124 165672 458176
rect 430028 456764 430080 456816
rect 580172 456764 580224 456816
rect 2872 455336 2924 455388
rect 165620 455336 165672 455388
rect 429200 455336 429252 455388
rect 580540 455336 580592 455388
rect 2780 452548 2832 452600
rect 165620 452548 165672 452600
rect 429568 451188 429620 451240
rect 580632 451188 580684 451240
rect 3424 449828 3476 449880
rect 165620 449828 165672 449880
rect 3516 447040 3568 447092
rect 165620 447040 165672 447092
rect 429844 444388 429896 444440
rect 580172 444388 580224 444440
rect 3608 444320 3660 444372
rect 165620 444320 165672 444372
rect 3700 440172 3752 440224
rect 165620 440172 165672 440224
rect 3424 436704 3476 436756
rect 165620 436704 165672 436756
rect 3424 433304 3476 433356
rect 165620 433304 165672 433356
rect 429936 431876 429988 431928
rect 579804 431876 579856 431928
rect 3792 430584 3844 430636
rect 165620 430584 165672 430636
rect 3700 427796 3752 427848
rect 165620 427796 165672 427848
rect 3608 420928 3660 420980
rect 165620 420928 165672 420980
rect 429844 419432 429896 419484
rect 580172 419432 580224 419484
rect 3516 418140 3568 418192
rect 165620 418140 165672 418192
rect 3424 415420 3476 415472
rect 165620 415420 165672 415472
rect 429568 414808 429620 414860
rect 433984 414808 434036 414860
rect 429568 411272 429620 411324
rect 435364 411272 435416 411324
rect 429476 408484 429528 408536
rect 461584 408484 461636 408536
rect 3148 407124 3200 407176
rect 165620 407124 165672 407176
rect 430212 405628 430264 405680
rect 580172 405628 580224 405680
rect 3240 404336 3292 404388
rect 165620 404336 165672 404388
rect 429568 402704 429620 402756
rect 432604 402704 432656 402756
rect 22744 394680 22796 394732
rect 165620 394680 165672 394732
rect 7564 391960 7616 392012
rect 165620 391960 165672 392012
rect 430120 391892 430172 391944
rect 580172 391892 580224 391944
rect 429568 390736 429620 390788
rect 431224 390736 431276 390788
rect 429568 387812 429620 387864
rect 454684 387812 454736 387864
rect 3332 384956 3384 385008
rect 166264 384956 166316 385008
rect 3332 383664 3384 383716
rect 165620 383664 165672 383716
rect 14464 379516 14516 379568
rect 165620 379516 165672 379568
rect 430028 379448 430080 379500
rect 580172 379448 580224 379500
rect 4068 374008 4120 374060
rect 165620 374008 165672 374060
rect 25504 371220 25556 371272
rect 165620 371220 165672 371272
rect 3976 368500 4028 368552
rect 165620 368500 165672 368552
rect 429936 368500 429988 368552
rect 447784 368500 447836 368552
rect 430028 365644 430080 365696
rect 580172 365644 580224 365696
rect 3884 362924 3936 362976
rect 165620 362924 165672 362976
rect 3792 358776 3844 358828
rect 165620 358776 165672 358828
rect 15844 356056 15896 356108
rect 165620 356056 165672 356108
rect 3700 353268 3752 353320
rect 165620 353268 165672 353320
rect 429936 353200 429988 353252
rect 580172 353200 580224 353252
rect 32404 350548 32456 350600
rect 165620 350548 165672 350600
rect 429844 350548 429896 350600
rect 442264 350548 442316 350600
rect 3608 347760 3660 347812
rect 165620 347760 165672 347812
rect 429844 347760 429896 347812
rect 439504 347760 439556 347812
rect 3516 345040 3568 345092
rect 165620 345040 165672 345092
rect 3424 342252 3476 342304
rect 165620 342252 165672 342304
rect 429108 339464 429160 339516
rect 489184 339464 489236 339516
rect 433984 339396 434036 339448
rect 579988 339396 580040 339448
rect 17224 338104 17276 338156
rect 165620 338104 165672 338156
rect 178040 336676 178092 336728
rect 178316 336676 178368 336728
rect 188344 336676 188396 336728
rect 190276 336676 190328 336728
rect 191840 336676 191892 336728
rect 192116 336676 192168 336728
rect 236000 336676 236052 336728
rect 236276 336676 236328 336728
rect 231768 336608 231820 336660
rect 270500 336676 270552 336728
rect 270684 336676 270736 336728
rect 271420 336676 271472 336728
rect 286968 336676 287020 336728
rect 295524 336676 295576 336728
rect 303896 336676 303948 336728
rect 304908 336676 304960 336728
rect 306564 336676 306616 336728
rect 307668 336676 307720 336728
rect 308680 336676 308732 336728
rect 309784 336676 309836 336728
rect 312912 336676 312964 336728
rect 270224 336608 270276 336660
rect 285588 336608 285640 336660
rect 294972 336608 295024 336660
rect 308128 336608 308180 336660
rect 311164 336608 311216 336660
rect 312360 336608 312412 336660
rect 313188 336608 313240 336660
rect 316592 336676 316644 336728
rect 317328 336676 317380 336728
rect 318708 336676 318760 336728
rect 319444 336676 319496 336728
rect 320272 336676 320324 336728
rect 321376 336676 321428 336728
rect 321836 336676 321888 336728
rect 322664 336676 322716 336728
rect 326068 336676 326120 336728
rect 326988 336676 327040 336728
rect 327080 336676 327132 336728
rect 328276 336676 328328 336728
rect 332876 336676 332928 336728
rect 333888 336676 333940 336728
rect 334440 336676 334492 336728
rect 335176 336676 335228 336728
rect 335544 336676 335596 336728
rect 336648 336676 336700 336728
rect 337108 336676 337160 336728
rect 338028 336676 338080 336728
rect 338120 336676 338172 336728
rect 339224 336676 339276 336728
rect 339684 336676 339736 336728
rect 340604 336676 340656 336728
rect 341340 336676 341392 336728
rect 342076 336676 342128 336728
rect 342352 336676 342404 336728
rect 343456 336676 343508 336728
rect 343916 336676 343968 336728
rect 344928 336676 344980 336728
rect 345480 336676 345532 336728
rect 346216 336676 346268 336728
rect 347136 336676 347188 336728
rect 347596 336676 347648 336728
rect 348148 336676 348200 336728
rect 349068 336676 349120 336728
rect 352380 336676 352432 336728
rect 353208 336676 353260 336728
rect 353392 336676 353444 336728
rect 354496 336676 354548 336728
rect 320456 336608 320508 336660
rect 333980 336608 334032 336660
rect 335268 336608 335320 336660
rect 338672 336608 338724 336660
rect 339408 336608 339460 336660
rect 349712 336608 349764 336660
rect 224868 336540 224920 336592
rect 267648 336540 267700 336592
rect 282828 336540 282880 336592
rect 293408 336540 293460 336592
rect 310796 336540 310848 336592
rect 316040 336540 316092 336592
rect 317236 336540 317288 336592
rect 317604 336540 317656 336592
rect 318708 336540 318760 336592
rect 329196 336540 329248 336592
rect 329748 336540 329800 336592
rect 336004 336540 336056 336592
rect 336556 336540 336608 336592
rect 351276 336540 351328 336592
rect 351828 336540 351880 336592
rect 352840 336608 352892 336660
rect 354956 336676 355008 336728
rect 355968 336676 356020 336728
rect 356520 336676 356572 336728
rect 357348 336676 357400 336728
rect 357624 336676 357676 336728
rect 358728 336676 358780 336728
rect 359188 336676 359240 336728
rect 360108 336676 360160 336728
rect 360752 336676 360804 336728
rect 361488 336676 361540 336728
rect 361856 336676 361908 336728
rect 362868 336676 362920 336728
rect 363420 336676 363472 336728
rect 364156 336676 364208 336728
rect 364432 336676 364484 336728
rect 365628 336676 365680 336728
rect 365996 336676 366048 336728
rect 367008 336676 367060 336728
rect 367100 336676 367152 336728
rect 368388 336676 368440 336728
rect 370228 336676 370280 336728
rect 371148 336676 371200 336728
rect 371332 336676 371384 336728
rect 372436 336676 372488 336728
rect 374460 336676 374512 336728
rect 375288 336676 375340 336728
rect 375472 336676 375524 336728
rect 376576 336676 376628 336728
rect 377128 336676 377180 336728
rect 378048 336676 378100 336728
rect 378692 336676 378744 336728
rect 379428 336676 379480 336728
rect 380624 336676 380676 336728
rect 380808 336676 380860 336728
rect 382372 336676 382424 336728
rect 383568 336676 383620 336728
rect 384948 336676 385000 336728
rect 385684 336676 385736 336728
rect 388168 336676 388220 336728
rect 388996 336676 389048 336728
rect 390744 336676 390796 336728
rect 391756 336676 391808 336728
rect 392308 336676 392360 336728
rect 393136 336676 393188 336728
rect 394976 336676 395028 336728
rect 395988 336676 396040 336728
rect 396540 336676 396592 336728
rect 397276 336676 397328 336728
rect 398104 336676 398156 336728
rect 398656 336676 398708 336728
rect 399208 336676 399260 336728
rect 400128 336676 400180 336728
rect 400220 336676 400272 336728
rect 401324 336676 401376 336728
rect 402336 336676 402388 336728
rect 402888 336676 402940 336728
rect 404452 336676 404504 336728
rect 405556 336676 405608 336728
rect 406016 336676 406068 336728
rect 407028 336676 407080 336728
rect 407120 336676 407172 336728
rect 408316 336676 408368 336728
rect 408684 336676 408736 336728
rect 409696 336676 409748 336728
rect 410248 336676 410300 336728
rect 411168 336676 411220 336728
rect 411812 336676 411864 336728
rect 412456 336676 412508 336728
rect 413376 336676 413428 336728
rect 413836 336676 413888 336728
rect 414480 336676 414532 336728
rect 415308 336676 415360 336728
rect 415492 336676 415544 336728
rect 416504 336676 416556 336728
rect 418160 336676 418212 336728
rect 419356 336676 419408 336728
rect 419724 336676 419776 336728
rect 420736 336676 420788 336728
rect 422852 336676 422904 336728
rect 423496 336676 423548 336728
rect 424416 336676 424468 336728
rect 424876 336676 424928 336728
rect 159364 336472 159416 336524
rect 203984 336472 204036 336524
rect 227628 336472 227680 336524
rect 268660 336472 268712 336524
rect 280896 336472 280948 336524
rect 291476 336472 291528 336524
rect 311808 336472 311860 336524
rect 323124 336472 323176 336524
rect 407396 336608 407448 336660
rect 416044 336608 416096 336660
rect 416688 336608 416740 336660
rect 417056 336608 417108 336660
rect 417976 336608 418028 336660
rect 421288 336608 421340 336660
rect 422208 336608 422260 336660
rect 422392 336608 422444 336660
rect 423588 336608 423640 336660
rect 415676 336540 415728 336592
rect 426532 336540 426584 336592
rect 427544 336540 427596 336592
rect 125508 336404 125560 336456
rect 223396 336404 223448 336456
rect 223488 336404 223540 336456
rect 267096 336404 267148 336456
rect 278044 336404 278096 336456
rect 290280 336404 290332 336456
rect 313372 336404 313424 336456
rect 318064 336404 318116 336456
rect 319168 336404 319220 336456
rect 320088 336404 320140 336456
rect 356060 336404 356112 336456
rect 422576 336472 422628 336524
rect 362316 336404 362368 336456
rect 436100 336404 436152 336456
rect 114468 336336 114520 336388
rect 218704 336336 218756 336388
rect 220728 336336 220780 336388
rect 266084 336336 266136 336388
rect 281448 336336 281500 336388
rect 292856 336336 292908 336388
rect 294604 336336 294656 336388
rect 298652 336336 298704 336388
rect 306012 336336 306064 336388
rect 309324 336336 309376 336388
rect 310244 336336 310296 336388
rect 313924 336336 313976 336388
rect 324412 336336 324464 336388
rect 369216 336336 369268 336388
rect 370504 336336 370556 336388
rect 35164 336268 35216 336320
rect 180800 336268 180852 336320
rect 217968 336268 218020 336320
rect 264428 336268 264480 336320
rect 277216 336268 277268 336320
rect 290740 336268 290792 336320
rect 311348 336268 311400 336320
rect 321836 336268 321888 336320
rect 330208 336268 330260 336320
rect 352564 336268 352616 336320
rect 29644 336200 29696 336252
rect 176568 336200 176620 336252
rect 219256 336200 219308 336252
rect 265532 336200 265584 336252
rect 277308 336200 277360 336252
rect 291292 336200 291344 336252
rect 307576 336200 307628 336252
rect 313372 336200 313424 336252
rect 314476 336200 314528 336252
rect 327724 336200 327776 336252
rect 328644 336200 328696 336252
rect 349804 336200 349856 336252
rect 365536 336200 365588 336252
rect 443000 336336 443052 336388
rect 28264 336132 28316 336184
rect 177120 336132 177172 336184
rect 213828 336132 213880 336184
rect 262864 336132 262916 336184
rect 271788 336132 271840 336184
rect 288716 336132 288768 336184
rect 292488 336132 292540 336184
rect 297640 336132 297692 336184
rect 305000 336132 305052 336184
rect 306196 336132 306248 336184
rect 319720 336132 319772 336184
rect 341064 336132 341116 336184
rect 344468 336132 344520 336184
rect 358084 336132 358136 336184
rect 368664 336132 368716 336184
rect 449900 336268 449952 336320
rect 371792 336200 371844 336252
rect 456800 336200 456852 336252
rect 379704 336132 379756 336184
rect 380808 336132 380860 336184
rect 465080 336132 465132 336184
rect 18604 336064 18656 336116
rect 172888 336064 172940 336116
rect 191104 336064 191156 336116
rect 216220 336064 216272 336116
rect 216588 336064 216640 336116
rect 263968 336064 264020 336116
rect 269028 336064 269080 336116
rect 287060 336064 287112 336116
rect 289728 336064 289780 336116
rect 296536 336064 296588 336116
rect 296628 336064 296680 336116
rect 299756 336064 299808 336116
rect 315028 336064 315080 336116
rect 330024 336064 330076 336116
rect 349160 336064 349212 336116
rect 350356 336064 350408 336116
rect 378140 336064 378192 336116
rect 471980 336064 472032 336116
rect 10324 335996 10376 336048
rect 170220 335996 170272 336048
rect 212448 335996 212500 336048
rect 262312 335996 262364 336048
rect 264888 335996 264940 336048
rect 285220 335996 285272 336048
rect 285496 335996 285548 336048
rect 294420 335996 294472 336048
rect 326528 335996 326580 336048
rect 230388 335928 230440 335980
rect 242808 335928 242860 335980
rect 275560 335928 275612 335980
rect 309692 335928 309744 335980
rect 317512 335928 317564 335980
rect 324504 335928 324556 335980
rect 325424 335928 325476 335980
rect 358176 335996 358228 336048
rect 374644 335996 374696 336048
rect 375012 335996 375064 336048
rect 381268 335996 381320 336048
rect 478880 335996 478932 336048
rect 356152 335928 356204 335980
rect 385500 335928 385552 335980
rect 386328 335928 386380 335980
rect 389180 335928 389232 335980
rect 390284 335928 390336 335980
rect 393412 335928 393464 335980
rect 394424 335928 394476 335980
rect 396080 335928 396132 335980
rect 397368 335928 397420 335980
rect 397644 335928 397696 335980
rect 398748 335928 398800 335980
rect 400772 335928 400824 335980
rect 401508 335928 401560 335980
rect 240784 335860 240836 335912
rect 243452 335860 243504 335912
rect 251088 335860 251140 335912
rect 279240 335860 279292 335912
rect 345020 335860 345072 335912
rect 346308 335860 346360 335912
rect 253848 335792 253900 335844
rect 280804 335792 280856 335844
rect 259368 335724 259420 335776
rect 282920 335724 282972 335776
rect 331312 335724 331364 335776
rect 332416 335724 332468 335776
rect 210516 335656 210568 335708
rect 211804 335656 211856 335708
rect 304448 335656 304500 335708
rect 306656 335656 306708 335708
rect 340236 335656 340288 335708
rect 340788 335656 340840 335708
rect 260748 335588 260800 335640
rect 283932 335588 283984 335640
rect 291844 335588 291896 335640
rect 297088 335588 297140 335640
rect 299388 335588 299440 335640
rect 300768 335588 300820 335640
rect 360292 335588 360344 335640
rect 361396 335588 361448 335640
rect 309232 335520 309284 335572
rect 310428 335520 310480 335572
rect 346584 335520 346636 335572
rect 347688 335520 347740 335572
rect 411260 335520 411312 335572
rect 412548 335520 412600 335572
rect 307116 335452 307168 335504
rect 312084 335452 312136 335504
rect 283564 335316 283616 335368
rect 289176 335316 289228 335368
rect 383936 335316 383988 335368
rect 412916 335316 412968 335368
rect 384948 335180 385000 335232
rect 423956 335316 424008 335368
rect 413928 335180 413980 335232
rect 424968 335180 425020 335232
rect 126888 334636 126940 334688
rect 223948 334636 224000 334688
rect 386604 334636 386656 334688
rect 489920 334636 489972 334688
rect 39304 334568 39356 334620
rect 183376 334568 183428 334620
rect 202788 334568 202840 334620
rect 258172 334568 258224 334620
rect 324964 334568 325016 334620
rect 351920 334568 351972 334620
rect 405004 334568 405056 334620
rect 531320 334568 531372 334620
rect 206928 333344 206980 333396
rect 259736 333344 259788 333396
rect 161388 333276 161440 333328
rect 95148 333208 95200 333260
rect 210240 333140 210292 333192
rect 372896 333276 372948 333328
rect 459560 333276 459612 333328
rect 328184 333208 328236 333260
rect 358820 333208 358872 333260
rect 394608 333208 394660 333260
rect 507860 333208 507912 333260
rect 239772 333140 239824 333192
rect 3056 332528 3108 332580
rect 166908 332528 166960 332580
rect 195888 331916 195940 331968
rect 254952 331916 255004 331968
rect 383384 331916 383436 331968
rect 483020 331916 483072 331968
rect 140688 331848 140740 331900
rect 230296 331848 230348 331900
rect 401784 331848 401836 331900
rect 524420 331848 524472 331900
rect 193404 331168 193456 331220
rect 193588 331168 193640 331220
rect 214196 331168 214248 331220
rect 214380 331168 214432 331220
rect 232044 331168 232096 331220
rect 232228 331168 232280 331220
rect 276204 330760 276256 330812
rect 165528 330556 165580 330608
rect 241336 330556 241388 330608
rect 276204 330556 276256 330608
rect 350816 330556 350868 330608
rect 409880 330556 409932 330608
rect 21364 330488 21416 330540
rect 173900 330488 173952 330540
rect 175372 330488 175424 330540
rect 175648 330488 175700 330540
rect 197360 330488 197412 330540
rect 198372 330488 198424 330540
rect 200120 330488 200172 330540
rect 200948 330488 201000 330540
rect 202972 330488 203024 330540
rect 203156 330488 203208 330540
rect 269212 330488 269264 330540
rect 269396 330488 269448 330540
rect 270592 330488 270644 330540
rect 271052 330488 271104 330540
rect 276112 330488 276164 330540
rect 276756 330488 276808 330540
rect 277400 330488 277452 330540
rect 278412 330488 278464 330540
rect 280252 330488 280304 330540
rect 280988 330488 281040 330540
rect 281632 330488 281684 330540
rect 282092 330488 282144 330540
rect 284484 330488 284536 330540
rect 284668 330488 284720 330540
rect 300860 330488 300912 330540
rect 301596 330488 301648 330540
rect 391296 330488 391348 330540
rect 500960 330488 501012 330540
rect 168380 330420 168432 330472
rect 168932 330420 168984 330472
rect 195980 329536 196032 329588
rect 196716 329536 196768 329588
rect 129648 329128 129700 329180
rect 225512 329128 225564 329180
rect 362776 329128 362828 329180
rect 437480 329128 437532 329180
rect 119988 329060 120040 329112
rect 221280 329060 221332 329112
rect 235908 329060 235960 329112
rect 272892 329060 272944 329112
rect 380624 329060 380676 329112
rect 477500 329060 477552 329112
rect 198740 328040 198792 328092
rect 199476 328040 199528 328092
rect 131028 327768 131080 327820
rect 225696 327768 225748 327820
rect 368020 327768 368072 327820
rect 448520 327768 448572 327820
rect 11704 327700 11756 327752
rect 172060 327700 172112 327752
rect 176568 327700 176620 327752
rect 245752 327700 245804 327752
rect 398564 327700 398616 327752
rect 517520 327700 517572 327752
rect 248604 326816 248656 326868
rect 248604 326612 248656 326664
rect 169668 326408 169720 326460
rect 242992 326408 243044 326460
rect 247132 326408 247184 326460
rect 362868 326408 362920 326460
rect 434720 326408 434772 326460
rect 88248 326340 88300 326392
rect 186320 326272 186372 326324
rect 186780 326272 186832 326324
rect 187700 326272 187752 326324
rect 188436 326272 188488 326324
rect 189172 326272 189224 326324
rect 189356 326272 189408 326324
rect 193312 326272 193364 326324
rect 194140 326272 194192 326324
rect 194600 326272 194652 326324
rect 195244 326272 195296 326324
rect 207112 326340 207164 326392
rect 207756 326340 207808 326392
rect 208492 326340 208544 326392
rect 209412 326340 209464 326392
rect 214104 326340 214156 326392
rect 214748 326340 214800 326392
rect 216772 326340 216824 326392
rect 217324 326340 217376 326392
rect 222292 326340 222344 326392
rect 222476 326340 222528 326392
rect 230480 326340 230532 326392
rect 230940 326340 230992 326392
rect 231952 326340 232004 326392
rect 232596 326340 232648 326392
rect 237380 326340 237432 326392
rect 237656 326340 237708 326392
rect 241520 326340 241572 326392
rect 241980 326340 242032 326392
rect 244280 326340 244332 326392
rect 245108 326340 245160 326392
rect 207204 326272 207256 326324
rect 248512 326340 248564 326392
rect 249340 326340 249392 326392
rect 258172 326340 258224 326392
rect 258908 326340 258960 326392
rect 259552 326340 259604 326392
rect 260380 326340 260432 326392
rect 333796 326340 333848 326392
rect 371240 326340 371292 326392
rect 387616 326340 387668 326392
rect 492680 326340 492732 326392
rect 237472 326204 237524 326256
rect 238300 326204 238352 326256
rect 247132 326204 247184 326256
rect 435364 325592 435416 325644
rect 580172 325592 580224 325644
rect 133788 324980 133840 325032
rect 226616 324980 226668 325032
rect 40684 324912 40736 324964
rect 185124 324912 185176 324964
rect 347504 324912 347556 324964
rect 402980 324912 403032 324964
rect 186412 324572 186464 324624
rect 187332 324572 187384 324624
rect 178132 324368 178184 324420
rect 178868 324368 178920 324420
rect 180892 324368 180944 324420
rect 181444 324368 181496 324420
rect 236092 324368 236144 324420
rect 236828 324368 236880 324420
rect 136548 323620 136600 323672
rect 228272 323620 228324 323672
rect 355876 323620 355928 323672
rect 420920 323620 420972 323672
rect 53748 323552 53800 323604
rect 192024 323552 192076 323604
rect 248420 323552 248472 323604
rect 248696 323552 248748 323604
rect 391756 323552 391808 323604
rect 499580 323552 499632 323604
rect 182272 323484 182324 323536
rect 182456 323484 182508 323536
rect 251180 323416 251232 323468
rect 252100 323416 252152 323468
rect 147588 322192 147640 322244
rect 233424 322192 233476 322244
rect 366916 322192 366968 322244
rect 445760 322192 445812 322244
rect 247040 321648 247092 321700
rect 247224 321648 247276 321700
rect 215392 321308 215444 321360
rect 215576 321308 215628 321360
rect 144828 320832 144880 320884
rect 232228 320832 232280 320884
rect 369768 320832 369820 320884
rect 452660 320832 452712 320884
rect 3056 320084 3108 320136
rect 166816 320084 166868 320136
rect 254032 319472 254084 319524
rect 254216 319472 254268 319524
rect 375288 319404 375340 319456
rect 463700 319404 463752 319456
rect 180708 318112 180760 318164
rect 247776 318112 247828 318164
rect 113088 318044 113140 318096
rect 218152 318044 218204 318096
rect 377956 318044 378008 318096
rect 470600 318044 470652 318096
rect 137928 316684 137980 316736
rect 229192 316684 229244 316736
rect 376484 316684 376536 316736
rect 466460 316684 466512 316736
rect 162768 315256 162820 315308
rect 240232 315256 240284 315308
rect 383476 315256 383528 315308
rect 481640 315256 481692 315308
rect 142068 313896 142120 313948
rect 230572 313896 230624 313948
rect 390284 313896 390336 313948
rect 496820 313896 496872 313948
rect 461584 313216 461636 313268
rect 580172 313216 580224 313268
rect 143448 312536 143500 312588
rect 230480 312536 230532 312588
rect 99288 311108 99340 311160
rect 210424 311108 210476 311160
rect 384856 311108 384908 311160
rect 485780 311108 485832 311160
rect 33784 309748 33836 309800
rect 179512 309748 179564 309800
rect 393136 309748 393188 309800
rect 503720 309748 503772 309800
rect 124128 308388 124180 308440
rect 222292 308388 222344 308440
rect 395896 308388 395948 308440
rect 510620 308388 510672 308440
rect 106188 307028 106240 307080
rect 214104 307028 214156 307080
rect 394516 307028 394568 307080
rect 506480 307028 506532 307080
rect 43444 305600 43496 305652
rect 186504 305600 186556 305652
rect 397184 305600 397236 305652
rect 514760 305600 514812 305652
rect 36544 304240 36596 304292
rect 180892 304240 180944 304292
rect 406936 304240 406988 304292
rect 535460 304240 535512 304292
rect 57888 302880 57940 302932
rect 193404 302880 193456 302932
rect 401324 302880 401376 302932
rect 521660 302880 521712 302932
rect 50988 301452 51040 301504
rect 188344 301452 188396 301504
rect 404176 301452 404228 301504
rect 528560 301452 528612 301504
rect 46204 300092 46256 300144
rect 187792 300092 187844 300144
rect 429200 299412 429252 299464
rect 580172 299412 580224 299464
rect 61936 298732 61988 298784
rect 194692 298732 194744 298784
rect 64788 297372 64840 297424
rect 196164 297372 196216 297424
rect 68928 294584 68980 294636
rect 197544 294584 197596 294636
rect 177948 290436 178000 290488
rect 245660 290436 245712 290488
rect 173808 286288 173860 286340
rect 244464 286288 244516 286340
rect 432604 285608 432656 285660
rect 580172 285608 580224 285660
rect 3240 280100 3292 280152
rect 166724 280100 166776 280152
rect 429292 273164 429344 273216
rect 580172 273164 580224 273216
rect 135168 268336 135220 268388
rect 226432 268336 226484 268388
rect 3056 267656 3108 267708
rect 166632 267656 166684 267708
rect 429384 259360 429436 259412
rect 580172 259360 580224 259412
rect 117228 255960 117280 256012
rect 219532 255960 219584 256012
rect 3240 255212 3292 255264
rect 22744 255212 22796 255264
rect 22744 253172 22796 253224
rect 175372 253172 175424 253224
rect 386236 251812 386288 251864
rect 490012 251812 490064 251864
rect 429476 245556 429528 245608
rect 580172 245556 580224 245608
rect 3240 241204 3292 241256
rect 7564 241204 7616 241256
rect 431224 233180 431276 233232
rect 579988 233180 580040 233232
rect 360016 232500 360068 232552
rect 430580 232500 430632 232552
rect 3240 229032 3292 229084
rect 166540 229032 166592 229084
rect 454684 219376 454736 219428
rect 580172 219376 580224 219428
rect 3240 215228 3292 215280
rect 166448 215228 166500 215280
rect 429568 206932 429620 206984
rect 579804 206932 579856 206984
rect 429660 193128 429712 193180
rect 580172 193128 580224 193180
rect 3332 188980 3384 189032
rect 14464 188980 14516 189032
rect 429752 179324 429804 179376
rect 580172 179324 580224 179376
rect 25596 177284 25648 177336
rect 178224 177284 178276 177336
rect 3332 176604 3384 176656
rect 166356 176604 166408 176656
rect 372436 175924 372488 175976
rect 456892 175924 456944 175976
rect 166908 174496 166960 174548
rect 241612 174496 241664 174548
rect 365536 174496 365588 174548
rect 441620 174496 441672 174548
rect 430488 166948 430540 167000
rect 580172 166948 580224 167000
rect 430396 153144 430448 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 25504 150356 25556 150408
rect 447784 139340 447836 139392
rect 580172 139340 580224 139392
rect 430304 126896 430356 126948
rect 580172 126896 580224 126948
rect 3148 124108 3200 124160
rect 166264 124108 166316 124160
rect 430212 113092 430264 113144
rect 579804 113092 579856 113144
rect 430120 100648 430172 100700
rect 580172 100648 580224 100700
rect 430028 86912 430080 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 15844 85484 15896 85536
rect 429936 73108 429988 73160
rect 580172 73108 580224 73160
rect 442264 60664 442316 60716
rect 580172 60664 580224 60716
rect 2872 59304 2924 59356
rect 32404 59304 32456 59356
rect 439504 46860 439556 46912
rect 580172 46860 580224 46912
rect 364156 44820 364208 44872
rect 438860 44820 438912 44872
rect 136456 35164 136508 35216
rect 227720 35164 227772 35216
rect 368296 35164 368348 35216
rect 448612 35164 448664 35216
rect 429844 33056 429896 33108
rect 580172 33056 580224 33108
rect 209688 31016 209740 31068
rect 259552 31016 259604 31068
rect 354404 31016 354456 31068
rect 416780 31016 416832 31068
rect 346124 29588 346176 29640
rect 398840 29588 398892 29640
rect 92388 28228 92440 28280
rect 208584 28228 208636 28280
rect 353208 28228 353260 28280
rect 414020 28228 414072 28280
rect 146208 26868 146260 26920
rect 231952 26868 232004 26920
rect 358084 26868 358136 26920
rect 396080 26868 396132 26920
rect 343364 25576 343416 25628
rect 391940 25576 391992 25628
rect 139308 25508 139360 25560
rect 229284 25508 229336 25560
rect 379336 25508 379388 25560
rect 473360 25508 473412 25560
rect 200028 24080 200080 24132
rect 255504 24080 255556 24132
rect 372528 24080 372580 24132
rect 458180 24080 458232 24132
rect 177856 22720 177908 22772
rect 247132 22720 247184 22772
rect 371056 22720 371108 22772
rect 455420 22720 455472 22772
rect 188988 21360 189040 21412
rect 251364 21360 251416 21412
rect 370504 21360 370556 21412
rect 451280 21360 451332 21412
rect 336464 20000 336516 20052
rect 378140 20000 378192 20052
rect 182088 19932 182140 19984
rect 248604 19932 248656 19984
rect 357256 19932 357308 19984
rect 423680 19932 423732 19984
rect 187608 18640 187660 18692
rect 251272 18640 251324 18692
rect 332324 18640 332376 18692
rect 367100 18640 367152 18692
rect 103428 18572 103480 18624
rect 212632 18572 212684 18624
rect 367008 18572 367060 18624
rect 444380 18572 444432 18624
rect 184848 17280 184900 17332
rect 248512 17280 248564 17332
rect 85488 17212 85540 17264
rect 204444 17212 204496 17264
rect 328276 17212 328328 17264
rect 357532 17212 357584 17264
rect 365628 17212 365680 17264
rect 440332 17212 440384 17264
rect 169576 15852 169628 15904
rect 240784 15852 240836 15904
rect 324136 15852 324188 15904
rect 349252 15852 349304 15904
rect 349804 15852 349856 15904
rect 361120 15852 361172 15904
rect 361304 15852 361356 15904
rect 434444 15852 434496 15904
rect 128268 14424 128320 14476
rect 223672 14424 223724 14476
rect 233148 14424 233200 14476
rect 270592 14424 270644 14476
rect 320088 14424 320140 14476
rect 339868 14424 339920 14476
rect 340604 14424 340656 14476
rect 385960 14424 386012 14476
rect 390376 14424 390428 14476
rect 498200 14424 498252 14476
rect 183468 13132 183520 13184
rect 248420 13132 248472 13184
rect 342076 13132 342128 13184
rect 389456 13132 389508 13184
rect 131764 13064 131816 13116
rect 226340 13064 226392 13116
rect 321284 13064 321336 13116
rect 343364 13064 343416 13116
rect 388996 13064 389048 13116
rect 494704 13064 494756 13116
rect 179052 11772 179104 11824
rect 247040 11772 247092 11824
rect 322664 11772 322716 11824
rect 345756 11772 345808 11824
rect 489184 11772 489236 11824
rect 580264 11772 580316 11824
rect 110328 11704 110380 11756
rect 191104 11704 191156 11756
rect 193128 11704 193180 11756
rect 252652 11704 252704 11756
rect 339224 11704 339276 11756
rect 382372 11704 382424 11756
rect 393228 11704 393280 11756
rect 505376 11704 505428 11756
rect 186136 10344 186188 10396
rect 249892 10344 249944 10396
rect 319444 10344 319496 10396
rect 338672 10344 338724 10396
rect 350356 10344 350408 10396
rect 407212 10344 407264 10396
rect 81348 10276 81400 10328
rect 159364 10276 159416 10328
rect 172428 10276 172480 10328
rect 244372 10276 244424 10328
rect 335084 10276 335136 10328
rect 374000 10276 374052 10328
rect 385684 10276 385736 10328
rect 487620 10276 487672 10328
rect 185124 9188 185176 9240
rect 249800 9188 249852 9240
rect 77392 9120 77444 9172
rect 201592 9120 201644 9172
rect 73804 9052 73856 9104
rect 200304 9052 200356 9104
rect 70308 8984 70360 9036
rect 198832 8984 198884 9036
rect 321376 8984 321428 9036
rect 342168 8984 342220 9036
rect 374644 8984 374696 9036
rect 427268 8984 427320 9036
rect 66720 8916 66772 8968
rect 197452 8916 197504 8968
rect 228732 8916 228784 8968
rect 269212 8916 269264 8968
rect 325516 8916 325568 8968
rect 354036 8916 354088 8968
rect 382188 8916 382240 8968
rect 480536 8916 480588 8968
rect 424692 8304 424744 8356
rect 424968 8304 425020 8356
rect 108120 8236 108172 8288
rect 215392 8236 215444 8288
rect 409604 8236 409656 8288
rect 541992 8236 542044 8288
rect 104532 8168 104584 8220
rect 214012 8168 214064 8220
rect 411076 8168 411128 8220
rect 545488 8168 545540 8220
rect 101036 8100 101088 8152
rect 212540 8100 212592 8152
rect 412364 8100 412416 8152
rect 549076 8100 549128 8152
rect 97448 8032 97500 8084
rect 211252 8032 211304 8084
rect 413744 8032 413796 8084
rect 552664 8032 552716 8084
rect 93952 7964 94004 8016
rect 208492 7964 208544 8016
rect 416504 7964 416556 8016
rect 556160 7964 556212 8016
rect 90364 7896 90416 7948
rect 207112 7896 207164 7948
rect 417976 7896 418028 7948
rect 559748 7896 559800 7948
rect 86868 7828 86920 7880
rect 205732 7828 205784 7880
rect 420644 7828 420696 7880
rect 63224 7760 63276 7812
rect 196072 7760 196124 7812
rect 422116 7760 422168 7812
rect 563244 7828 563296 7880
rect 59636 7692 59688 7744
rect 193312 7692 193364 7744
rect 423404 7692 423456 7744
rect 566832 7760 566884 7812
rect 56048 7624 56100 7676
rect 191932 7624 191984 7676
rect 317144 7624 317196 7676
rect 335084 7624 335136 7676
rect 424784 7624 424836 7676
rect 570328 7692 570380 7744
rect 52552 7556 52604 7608
rect 190552 7556 190604 7608
rect 239312 7556 239364 7608
rect 273444 7556 273496 7608
rect 324228 7556 324280 7608
rect 350356 7556 350408 7608
rect 423680 7556 423732 7608
rect 424968 7556 425020 7608
rect 573916 7624 573968 7676
rect 577412 7556 577464 7608
rect 111616 7488 111668 7540
rect 216772 7488 216824 7540
rect 408224 7488 408276 7540
rect 538404 7488 538456 7540
rect 115204 7420 115256 7472
rect 218244 7420 218296 7472
rect 407028 7420 407080 7472
rect 534908 7420 534960 7472
rect 118792 7352 118844 7404
rect 220912 7352 220964 7404
rect 405556 7352 405608 7404
rect 531412 7352 531464 7404
rect 122288 7284 122340 7336
rect 222384 7284 222436 7336
rect 402796 7284 402848 7336
rect 527824 7284 527876 7336
rect 153016 7216 153068 7268
rect 236184 7216 236236 7268
rect 361396 7216 361448 7268
rect 432052 7216 432104 7268
rect 149520 7148 149572 7200
rect 233332 7148 233384 7200
rect 358636 7148 358688 7200
rect 428464 7148 428516 7200
rect 156604 7080 156656 7132
rect 237564 7080 237616 7132
rect 419264 7080 419316 7132
rect 160100 7012 160152 7064
rect 238760 7012 238812 7064
rect 3424 6808 3476 6860
rect 17224 6808 17276 6860
rect 83280 6808 83332 6860
rect 204352 6808 204404 6860
rect 386328 6808 386380 6860
rect 488816 6808 488868 6860
rect 48964 6740 49016 6792
rect 189172 6740 189224 6792
rect 387524 6740 387576 6792
rect 492312 6740 492364 6792
rect 44272 6672 44324 6724
rect 186412 6672 186464 6724
rect 389088 6672 389140 6724
rect 495900 6672 495952 6724
rect 40776 6604 40828 6656
rect 185032 6604 185084 6656
rect 390468 6604 390520 6656
rect 499396 6604 499448 6656
rect 37188 6536 37240 6588
rect 183652 6536 183704 6588
rect 205088 6536 205140 6588
rect 258172 6536 258224 6588
rect 391848 6536 391900 6588
rect 502984 6536 503036 6588
rect 33600 6468 33652 6520
rect 182272 6468 182324 6520
rect 201592 6468 201644 6520
rect 256792 6468 256844 6520
rect 394424 6468 394476 6520
rect 506572 6468 506624 6520
rect 30104 6400 30156 6452
rect 180984 6400 181036 6452
rect 197912 6400 197964 6452
rect 255412 6400 255464 6452
rect 395988 6400 396040 6452
rect 510068 6400 510120 6452
rect 26516 6332 26568 6384
rect 179420 6332 179472 6384
rect 194416 6332 194468 6384
rect 254032 6332 254084 6384
rect 397276 6332 397328 6384
rect 513564 6332 513616 6384
rect 21824 6264 21876 6316
rect 176752 6264 176804 6316
rect 190828 6264 190880 6316
rect 252560 6264 252612 6316
rect 398656 6264 398708 6316
rect 517152 6264 517204 6316
rect 8760 6196 8812 6248
rect 171232 6196 171284 6248
rect 174268 6196 174320 6248
rect 244280 6196 244332 6248
rect 315948 6196 316000 6248
rect 331588 6196 331640 6248
rect 400036 6196 400088 6248
rect 520740 6196 520792 6248
rect 4068 6128 4120 6180
rect 169852 6128 169904 6180
rect 170772 6128 170824 6180
rect 243084 6128 243136 6180
rect 322756 6128 322808 6180
rect 346952 6128 347004 6180
rect 352564 6128 352616 6180
rect 364616 6128 364668 6180
rect 401416 6128 401468 6180
rect 524236 6128 524288 6180
rect 128176 6060 128228 6112
rect 224960 6060 225012 6112
rect 384948 6060 385000 6112
rect 485228 6060 485280 6112
rect 144736 5992 144788 6044
rect 231860 5992 231912 6044
rect 383568 5992 383620 6044
rect 481732 5992 481784 6044
rect 148324 5924 148376 5976
rect 233240 5924 233292 5976
rect 380716 5924 380768 5976
rect 476948 5924 477000 5976
rect 151820 5856 151872 5908
rect 234712 5856 234764 5908
rect 379428 5856 379480 5908
rect 473452 5856 473504 5908
rect 155408 5788 155460 5840
rect 236092 5788 236144 5840
rect 378048 5788 378100 5840
rect 469864 5788 469916 5840
rect 158904 5720 158956 5772
rect 237472 5720 237524 5772
rect 376576 5720 376628 5772
rect 466276 5720 466328 5772
rect 163688 5652 163740 5704
rect 240324 5652 240376 5704
rect 373816 5652 373868 5704
rect 462780 5652 462832 5704
rect 167184 5584 167236 5636
rect 241520 5584 241572 5636
rect 62028 5448 62080 5500
rect 194600 5448 194652 5500
rect 225144 5448 225196 5500
rect 267832 5448 267884 5500
rect 343456 5448 343508 5500
rect 391848 5448 391900 5500
rect 409696 5448 409748 5500
rect 540796 5448 540848 5500
rect 58440 5380 58492 5432
rect 193220 5380 193272 5432
rect 221556 5380 221608 5432
rect 266452 5380 266504 5432
rect 340696 5380 340748 5432
rect 388260 5380 388312 5432
rect 411168 5380 411220 5432
rect 544384 5380 544436 5432
rect 54944 5312 54996 5364
rect 191840 5312 191892 5364
rect 218060 5312 218112 5364
rect 265072 5312 265124 5364
rect 344928 5312 344980 5364
rect 395344 5312 395396 5364
rect 412456 5312 412508 5364
rect 547880 5312 547932 5364
rect 51356 5244 51408 5296
rect 190460 5244 190512 5296
rect 214472 5244 214524 5296
rect 262312 5244 262364 5296
rect 346216 5244 346268 5296
rect 398932 5244 398984 5296
rect 413836 5244 413888 5296
rect 551468 5244 551520 5296
rect 47860 5176 47912 5228
rect 189264 5176 189316 5228
rect 210976 5176 211028 5228
rect 260932 5176 260984 5228
rect 347596 5176 347648 5228
rect 402520 5176 402572 5228
rect 415216 5176 415268 5228
rect 554964 5176 555016 5228
rect 17040 5108 17092 5160
rect 175464 5108 175516 5160
rect 207388 5108 207440 5160
rect 259644 5108 259696 5160
rect 348976 5108 349028 5160
rect 406016 5108 406068 5160
rect 416596 5108 416648 5160
rect 558552 5108 558604 5160
rect 12348 5040 12400 5092
rect 162768 5040 162820 5092
rect 7656 4972 7708 5024
rect 171140 5040 171192 5092
rect 203892 5040 203944 5092
rect 258264 5040 258316 5092
rect 350448 5040 350500 5092
rect 409604 5040 409656 5092
rect 419356 5040 419408 5092
rect 562048 5040 562100 5092
rect 168472 4972 168524 5024
rect 2872 4904 2924 4956
rect 162768 4904 162820 4956
rect 172612 4972 172664 5024
rect 200304 4972 200356 5024
rect 256700 4972 256752 5024
rect 351736 4972 351788 5024
rect 413100 4972 413152 5024
rect 420736 4972 420788 5024
rect 565636 4972 565688 5024
rect 196808 4904 196860 4956
rect 255320 4904 255372 4956
rect 354496 4904 354548 4956
rect 416504 4904 416556 4956
rect 422208 4904 422260 4956
rect 569132 4904 569184 4956
rect 572 4836 624 4888
rect 167000 4836 167052 4888
rect 193220 4836 193272 4888
rect 254124 4836 254176 4888
rect 355968 4836 356020 4888
rect 420184 4836 420236 4888
rect 423496 4836 423548 4888
rect 572720 4836 572772 4888
rect 1676 4768 1728 4820
rect 168380 4768 168432 4820
rect 189724 4768 189776 4820
rect 251180 4768 251232 4820
rect 357348 4768 357400 4820
rect 423772 4768 423824 4820
rect 424876 4768 424928 4820
rect 576308 4768 576360 4820
rect 65524 4700 65576 4752
rect 195980 4700 196032 4752
rect 339316 4700 339368 4752
rect 384764 4700 384816 4752
rect 408316 4700 408368 4752
rect 537208 4700 537260 4752
rect 72608 4632 72660 4684
rect 200212 4632 200264 4684
rect 337936 4632 337988 4684
rect 381176 4632 381228 4684
rect 405464 4632 405516 4684
rect 533712 4632 533764 4684
rect 69112 4564 69164 4616
rect 197360 4564 197412 4616
rect 336556 4564 336608 4616
rect 377680 4564 377732 4616
rect 404268 4564 404320 4616
rect 530124 4564 530176 4616
rect 76196 4496 76248 4548
rect 201500 4496 201552 4548
rect 335176 4496 335228 4548
rect 79692 4428 79744 4480
rect 202972 4428 203024 4480
rect 333888 4428 333940 4480
rect 402888 4496 402940 4548
rect 526628 4496 526680 4548
rect 150624 4360 150676 4412
rect 234620 4360 234672 4412
rect 332416 4360 332468 4412
rect 367008 4360 367060 4412
rect 374092 4428 374144 4480
rect 401508 4428 401560 4480
rect 523040 4428 523092 4480
rect 370596 4360 370648 4412
rect 400128 4360 400180 4412
rect 519544 4360 519596 4412
rect 154212 4292 154264 4344
rect 236000 4292 236052 4344
rect 329656 4292 329708 4344
rect 363512 4292 363564 4344
rect 398748 4292 398800 4344
rect 515956 4292 516008 4344
rect 157800 4224 157852 4276
rect 237380 4224 237432 4276
rect 397368 4224 397420 4276
rect 512460 4224 512512 4276
rect 126980 4156 127032 4208
rect 128268 4156 128320 4208
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 143540 4156 143592 4208
rect 144828 4156 144880 4208
rect 168380 4156 168432 4208
rect 169668 4156 169720 4208
rect 178132 4156 178184 4208
rect 20628 4088 20680 4140
rect 28264 4088 28316 4140
rect 45468 4088 45520 4140
rect 46204 4088 46256 4140
rect 85672 4088 85724 4140
rect 205640 4088 205692 4140
rect 252376 4088 252428 4140
rect 448612 4156 448664 4208
rect 449808 4156 449860 4208
rect 82084 4020 82136 4072
rect 204260 4020 204312 4072
rect 248788 4020 248840 4072
rect 280344 4088 280396 4140
rect 306288 4088 306340 4140
rect 309048 4088 309100 4140
rect 309784 4088 309836 4140
rect 310336 4088 310388 4140
rect 318616 4088 318668 4140
rect 338028 4088 338080 4140
rect 379980 4088 380032 4140
rect 409788 4088 409840 4140
rect 543188 4088 543240 4140
rect 277216 4020 277268 4072
rect 294880 4020 294932 4072
rect 298284 4020 298336 4072
rect 317236 4020 317288 4072
rect 325516 4020 325568 4072
rect 339408 4020 339460 4072
rect 383568 4020 383620 4072
rect 412548 4020 412600 4072
rect 546684 4020 546736 4072
rect 78588 3952 78640 4004
rect 203064 3952 203116 4004
rect 247592 3952 247644 4004
rect 276204 3952 276256 4004
rect 278044 3952 278096 4004
rect 317328 3952 317380 4004
rect 333888 3952 333940 4004
rect 340788 3952 340840 4004
rect 387156 3952 387208 4004
rect 413928 3952 413980 4004
rect 550272 3952 550324 4004
rect 75000 3884 75052 3936
rect 200120 3884 200172 3936
rect 246396 3884 246448 3936
rect 277400 3884 277452 3936
rect 281724 3884 281776 3936
rect 318064 3884 318116 3936
rect 326804 3884 326856 3936
rect 342076 3884 342128 3936
rect 390652 3884 390704 3936
rect 415308 3884 415360 3936
rect 553768 3884 553820 3936
rect 71504 3816 71556 3868
rect 198740 3816 198792 3868
rect 245200 3816 245252 3868
rect 34796 3748 34848 3800
rect 39304 3748 39356 3800
rect 46664 3748 46716 3800
rect 187700 3748 187752 3800
rect 242900 3748 242952 3800
rect 270040 3748 270092 3800
rect 278964 3816 279016 3868
rect 276112 3748 276164 3800
rect 277032 3748 277084 3800
rect 277308 3748 277360 3800
rect 43076 3680 43128 3732
rect 186320 3680 186372 3732
rect 240508 3680 240560 3732
rect 274824 3680 274876 3732
rect 283564 3816 283616 3868
rect 322848 3816 322900 3868
rect 325608 3816 325660 3868
rect 332692 3816 332744 3868
rect 343548 3816 343600 3868
rect 394240 3816 394292 3868
rect 416596 3816 416648 3868
rect 557356 3816 557408 3868
rect 283104 3748 283156 3800
rect 294052 3748 294104 3800
rect 318708 3748 318760 3800
rect 336280 3748 336332 3800
rect 346308 3748 346360 3800
rect 397736 3748 397788 3800
rect 418068 3748 418120 3800
rect 560852 3748 560904 3800
rect 279516 3680 279568 3732
rect 19432 3544 19484 3596
rect 29644 3612 29696 3664
rect 39580 3612 39632 3664
rect 184940 3612 184992 3664
rect 238116 3612 238168 3664
rect 28908 3544 28960 3596
rect 35164 3544 35216 3596
rect 35992 3544 36044 3596
rect 183560 3544 183612 3596
rect 227536 3544 227588 3596
rect 18236 3476 18288 3528
rect 22744 3476 22796 3528
rect 23020 3476 23072 3528
rect 25596 3476 25648 3528
rect 32404 3476 32456 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 13544 3408 13596 3460
rect 21364 3408 21416 3460
rect 25320 3408 25372 3460
rect 171968 3476 172020 3528
rect 172428 3476 172480 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 176660 3476 176712 3528
rect 177948 3476 178000 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 181444 3476 181496 3528
rect 182088 3476 182140 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 188528 3476 188580 3528
rect 188988 3476 189040 3528
rect 192024 3476 192076 3528
rect 193128 3476 193180 3528
rect 199108 3476 199160 3528
rect 200028 3476 200080 3528
rect 208584 3476 208636 3528
rect 209688 3476 209740 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 215668 3476 215720 3528
rect 216588 3476 216640 3528
rect 216864 3476 216916 3528
rect 217968 3476 218020 3528
rect 222752 3476 222804 3528
rect 223488 3476 223540 3528
rect 226340 3476 226392 3528
rect 227628 3476 227680 3528
rect 229836 3544 229888 3596
rect 230388 3544 230440 3596
rect 231032 3544 231084 3596
rect 231768 3544 231820 3596
rect 232228 3544 232280 3596
rect 233148 3544 233200 3596
rect 233424 3544 233476 3596
rect 270684 3544 270736 3596
rect 277492 3612 277544 3664
rect 280252 3612 280304 3664
rect 284300 3612 284352 3664
rect 285496 3612 285548 3664
rect 321468 3680 321520 3732
rect 291292 3612 291344 3664
rect 313924 3612 313976 3664
rect 319720 3612 319772 3664
rect 337476 3680 337528 3732
rect 347688 3680 347740 3732
rect 401324 3680 401376 3732
rect 419448 3680 419500 3732
rect 564440 3680 564492 3732
rect 344560 3612 344612 3664
rect 349068 3612 349120 3664
rect 404820 3612 404872 3664
rect 420828 3612 420880 3664
rect 568028 3612 568080 3664
rect 273352 3544 273404 3596
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 267740 3476 267792 3528
rect 269028 3476 269080 3528
rect 271236 3476 271288 3528
rect 271788 3476 271840 3528
rect 272708 3476 272760 3528
rect 275008 3544 275060 3596
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 273628 3476 273680 3528
rect 288532 3544 288584 3596
rect 306196 3544 306248 3596
rect 307944 3544 307996 3596
rect 325424 3544 325476 3596
rect 348056 3544 348108 3596
rect 351828 3544 351880 3596
rect 411904 3544 411956 3596
rect 423588 3544 423640 3596
rect 571524 3544 571576 3596
rect 287336 3476 287388 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 291384 3476 291436 3528
rect 292488 3476 292540 3528
rect 293684 3476 293736 3528
rect 294604 3476 294656 3528
rect 296076 3476 296128 3528
rect 296628 3476 296680 3528
rect 298468 3476 298520 3528
rect 299388 3476 299440 3528
rect 302332 3476 302384 3528
rect 303160 3476 303212 3528
rect 304908 3476 304960 3528
rect 305552 3476 305604 3528
rect 313188 3476 313240 3528
rect 324412 3476 324464 3528
rect 351644 3476 351696 3528
rect 354588 3476 354640 3528
rect 418988 3476 419040 3528
rect 424692 3476 424744 3528
rect 575112 3476 575164 3528
rect 182364 3408 182416 3460
rect 206192 3408 206244 3460
rect 206928 3408 206980 3460
rect 209780 3408 209832 3460
rect 260840 3408 260892 3460
rect 261760 3408 261812 3460
rect 50160 3340 50212 3392
rect 50988 3340 51040 3392
rect 57244 3340 57296 3392
rect 57888 3340 57940 3392
rect 60832 3340 60884 3392
rect 61936 3340 61988 3392
rect 64328 3340 64380 3392
rect 64788 3340 64840 3392
rect 67916 3340 67968 3392
rect 68928 3340 68980 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 84476 3340 84528 3392
rect 85488 3340 85540 3392
rect 91560 3340 91612 3392
rect 92388 3340 92440 3392
rect 89168 3272 89220 3324
rect 207296 3340 207348 3392
rect 241704 3340 241756 3392
rect 242808 3340 242860 3392
rect 249984 3340 250036 3392
rect 251088 3340 251140 3392
rect 251180 3340 251232 3392
rect 277308 3340 277360 3392
rect 277584 3340 277636 3392
rect 92756 3272 92808 3324
rect 208676 3272 208728 3324
rect 254676 3272 254728 3324
rect 280712 3408 280764 3460
rect 281448 3408 281500 3460
rect 281908 3408 281960 3460
rect 282828 3408 282880 3460
rect 290188 3408 290240 3460
rect 291844 3408 291896 3460
rect 314568 3408 314620 3460
rect 328000 3408 328052 3460
rect 328184 3408 328236 3460
rect 358728 3408 358780 3460
rect 358820 3408 358872 3460
rect 426164 3408 426216 3460
rect 426256 3408 426308 3460
rect 578608 3408 578660 3460
rect 287796 3340 287848 3392
rect 295432 3340 295484 3392
rect 310428 3340 310480 3392
rect 317328 3340 317380 3392
rect 327724 3340 327776 3392
rect 329196 3340 329248 3392
rect 336648 3340 336700 3392
rect 376484 3340 376536 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 408500 3340 408552 3392
rect 539600 3340 539652 3392
rect 284576 3272 284628 3324
rect 311164 3272 311216 3324
rect 315028 3272 315080 3324
rect 335268 3272 335320 3324
rect 372896 3272 372948 3324
rect 374000 3272 374052 3324
rect 375288 3272 375340 3324
rect 380808 3272 380860 3324
rect 31300 3204 31352 3256
rect 36544 3204 36596 3256
rect 98644 3204 98696 3256
rect 99288 3204 99340 3256
rect 41880 3136 41932 3188
rect 43444 3136 43496 3188
rect 96252 3136 96304 3188
rect 209964 3204 210016 3256
rect 255872 3204 255924 3256
rect 102232 3136 102284 3188
rect 103428 3136 103480 3188
rect 105728 3136 105780 3188
rect 106188 3136 106240 3188
rect 109316 3136 109368 3188
rect 110328 3136 110380 3188
rect 211344 3136 211396 3188
rect 257068 3136 257120 3188
rect 281632 3204 281684 3256
rect 299664 3204 299716 3256
rect 300952 3204 301004 3256
rect 307668 3204 307720 3256
rect 311440 3204 311492 3256
rect 332508 3204 332560 3256
rect 369400 3204 369452 3256
rect 376668 3204 376720 3256
rect 468668 3204 468720 3256
rect 473360 3272 473412 3324
rect 474556 3272 474608 3324
rect 481640 3272 481692 3324
rect 482836 3272 482888 3324
rect 489920 3272 489972 3324
rect 491116 3272 491168 3324
rect 506480 3272 506532 3324
rect 507676 3272 507728 3324
rect 531320 3272 531372 3324
rect 532516 3272 532568 3324
rect 475752 3204 475804 3256
rect 278320 3136 278372 3188
rect 280804 3136 280856 3188
rect 297272 3136 297324 3188
rect 299756 3136 299808 3188
rect 331128 3136 331180 3188
rect 365812 3136 365864 3188
rect 373724 3136 373776 3188
rect 461584 3136 461636 3188
rect 38384 3068 38436 3120
rect 40684 3068 40736 3120
rect 103336 3068 103388 3120
rect 214196 3068 214248 3120
rect 259460 3068 259512 3120
rect 283012 3068 283064 3120
rect 329748 3068 329800 3120
rect 362316 3068 362368 3120
rect 371148 3068 371200 3120
rect 454500 3068 454552 3120
rect 456800 3068 456852 3120
rect 458088 3068 458140 3120
rect 11152 3000 11204 3052
rect 18604 3000 18656 3052
rect 27712 3000 27764 3052
rect 33784 3000 33836 3052
rect 99840 3000 99892 3052
rect 114008 3000 114060 3052
rect 114468 3000 114520 3052
rect 116400 3000 116452 3052
rect 117228 3000 117280 3052
rect 215484 3000 215536 3052
rect 262956 3000 263008 3052
rect 284484 3000 284536 3052
rect 292580 3000 292632 3052
rect 298192 3000 298244 3052
rect 310336 3000 310388 3052
rect 316224 3000 316276 3052
rect 326988 3000 327040 3052
rect 355232 3000 355284 3052
rect 368388 3000 368440 3052
rect 447416 3000 447468 3052
rect 9956 2932 10008 2984
rect 11704 2932 11756 2984
rect 110512 2932 110564 2984
rect 216772 2932 216824 2984
rect 223948 2932 224000 2984
rect 224868 2932 224920 2984
rect 265348 2932 265400 2984
rect 285772 2932 285824 2984
rect 364248 2932 364300 2984
rect 440240 2932 440292 2984
rect 440332 2932 440384 2984
rect 441528 2932 441580 2984
rect 106924 2864 106976 2916
rect 117596 2796 117648 2848
rect 219624 2864 219676 2916
rect 268752 2864 268804 2916
rect 268844 2864 268896 2916
rect 287152 2864 287204 2916
rect 361488 2864 361540 2916
rect 433248 2864 433300 2916
rect 121092 2796 121144 2848
rect 221096 2796 221148 2848
rect 266544 2796 266596 2848
rect 285864 2796 285916 2848
rect 360108 2796 360160 2848
rect 429660 2796 429712 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3054 540832 3110 540841
rect 3054 540767 3110 540776
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2870 514856 2926 514865
rect 2870 514791 2926 514800
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2792 452606 2820 501735
rect 2884 455394 2912 514791
rect 2976 458182 3004 527847
rect 3068 460902 3096 540767
rect 3160 465050 3188 553823
rect 3252 467838 3280 566879
rect 3344 470558 3372 579935
rect 3436 494018 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3424 494012 3476 494018
rect 3424 493954 3476 493960
rect 3528 491298 3556 671191
rect 3606 658200 3662 658209
rect 3606 658135 3662 658144
rect 3516 491292 3568 491298
rect 3516 491234 3568 491240
rect 3422 488744 3478 488753
rect 3422 488679 3478 488688
rect 3332 470552 3384 470558
rect 3332 470494 3384 470500
rect 3240 467832 3292 467838
rect 3240 467774 3292 467780
rect 3148 465044 3200 465050
rect 3148 464986 3200 464992
rect 3056 460896 3108 460902
rect 3056 460838 3108 460844
rect 2964 458176 3016 458182
rect 2964 458118 3016 458124
rect 2872 455388 2924 455394
rect 2872 455330 2924 455336
rect 2780 452600 2832 452606
rect 2780 452542 2832 452548
rect 3436 449886 3464 488679
rect 3620 488510 3648 658135
rect 3698 645144 3754 645153
rect 3698 645079 3754 645088
rect 3608 488504 3660 488510
rect 3608 488446 3660 488452
rect 3712 485790 3740 645079
rect 3790 632088 3846 632097
rect 3790 632023 3846 632032
rect 3700 485784 3752 485790
rect 3700 485726 3752 485732
rect 3804 481642 3832 632023
rect 3882 619168 3938 619177
rect 3882 619103 3938 619112
rect 3792 481636 3844 481642
rect 3792 481578 3844 481584
rect 3896 478854 3924 619103
rect 3974 606112 4030 606121
rect 3974 606047 4030 606056
rect 3884 478848 3936 478854
rect 3884 478790 3936 478796
rect 3988 476066 4016 606047
rect 4066 593056 4122 593065
rect 4066 592991 4122 593000
rect 3976 476060 4028 476066
rect 3976 476002 4028 476008
rect 3514 475688 3570 475697
rect 3514 475623 3570 475632
rect 3424 449880 3476 449886
rect 3424 449822 3476 449828
rect 3528 447098 3556 475623
rect 4080 473346 4108 592991
rect 8220 500274 8248 702406
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 24780 500342 24808 699654
rect 41340 500410 41368 700334
rect 56796 700194 56824 703520
rect 72988 702434 73016 703520
rect 72988 702406 73108 702434
rect 56784 700188 56836 700194
rect 56784 700130 56836 700136
rect 57888 700188 57940 700194
rect 57888 700130 57940 700136
rect 57900 500478 57928 700130
rect 73080 500546 73108 702406
rect 89180 699718 89208 703520
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 89640 500614 89668 699654
rect 106200 500682 106228 700334
rect 121656 699718 121684 703520
rect 137848 702434 137876 703520
rect 154132 702434 154160 703520
rect 137848 702406 137968 702434
rect 154132 702406 154528 702434
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 122748 699712 122800 699718
rect 122748 699654 122800 699660
rect 122760 500750 122788 699654
rect 137940 500818 137968 702406
rect 154500 500886 154528 702406
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 171060 500954 171088 700198
rect 186516 700194 186544 703520
rect 186504 700188 186556 700194
rect 186504 700130 186556 700136
rect 187608 700188 187660 700194
rect 187608 700130 187660 700136
rect 171048 500948 171100 500954
rect 171048 500890 171100 500896
rect 154488 500880 154540 500886
rect 154488 500822 154540 500828
rect 137928 500812 137980 500818
rect 137928 500754 137980 500760
rect 122748 500744 122800 500750
rect 122748 500686 122800 500692
rect 106188 500676 106240 500682
rect 106188 500618 106240 500624
rect 89628 500608 89680 500614
rect 89628 500550 89680 500556
rect 73068 500540 73120 500546
rect 73068 500482 73120 500488
rect 57888 500472 57940 500478
rect 57888 500414 57940 500420
rect 41328 500404 41380 500410
rect 41328 500346 41380 500352
rect 186044 500404 186096 500410
rect 186044 500346 186096 500352
rect 24768 500336 24820 500342
rect 24768 500278 24820 500284
rect 178776 500336 178828 500342
rect 178776 500278 178828 500284
rect 8208 500268 8260 500274
rect 8208 500210 8260 500216
rect 171600 500268 171652 500274
rect 171600 500210 171652 500216
rect 171612 497964 171640 500210
rect 178788 497964 178816 500278
rect 186056 497964 186084 500346
rect 187620 500274 187648 700130
rect 200488 500540 200540 500546
rect 200488 500482 200540 500488
rect 193220 500472 193272 500478
rect 193220 500414 193272 500420
rect 187608 500268 187660 500274
rect 187608 500210 187660 500216
rect 193232 497964 193260 500414
rect 200500 497964 200528 500482
rect 202800 500342 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 214932 500676 214984 500682
rect 214932 500618 214984 500624
rect 207664 500608 207716 500614
rect 207664 500550 207716 500556
rect 202788 500336 202840 500342
rect 202788 500278 202840 500284
rect 207676 497964 207704 500550
rect 214944 497964 214972 500618
rect 219360 500410 219388 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 235908 700392 235960 700398
rect 235908 700334 235960 700340
rect 229376 500812 229428 500818
rect 229376 500754 229428 500760
rect 222108 500744 222160 500750
rect 222108 500686 222160 500692
rect 219348 500404 219400 500410
rect 219348 500346 219400 500352
rect 222120 497964 222148 500686
rect 229388 497964 229416 500754
rect 235920 500478 235948 700334
rect 251468 700126 251496 703520
rect 251456 700120 251508 700126
rect 251456 700062 251508 700068
rect 252468 700120 252520 700126
rect 252468 700062 252520 700068
rect 243820 500948 243872 500954
rect 243820 500890 243872 500896
rect 236552 500880 236604 500886
rect 236552 500822 236604 500828
rect 235908 500472 235960 500478
rect 235908 500414 235960 500420
rect 236564 497964 236592 500822
rect 243832 497964 243860 500890
rect 252480 500274 252508 700062
rect 265440 500404 265492 500410
rect 265440 500346 265492 500352
rect 258264 500336 258316 500342
rect 258264 500278 258316 500284
rect 250996 500268 251048 500274
rect 250996 500210 251048 500216
rect 252468 500268 252520 500274
rect 252468 500210 252520 500216
rect 251008 497964 251036 500210
rect 258276 497964 258304 500278
rect 265452 497964 265480 500346
rect 267660 500342 267688 703520
rect 283852 702434 283880 703520
rect 283852 702406 284248 702434
rect 272708 500472 272760 500478
rect 272708 500414 272760 500420
rect 267648 500336 267700 500342
rect 267648 500278 267700 500284
rect 272720 497964 272748 500414
rect 284220 500274 284248 702406
rect 300136 699718 300164 703520
rect 316328 699718 316356 703520
rect 331128 700528 331180 700534
rect 331128 700470 331180 700476
rect 317328 700392 317380 700398
rect 317328 700334 317380 700340
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 309784 699712 309836 699718
rect 309784 699654 309836 699660
rect 316316 699712 316368 699718
rect 316316 699654 316368 699660
rect 300780 500954 300808 699654
rect 309796 500954 309824 699654
rect 300768 500948 300820 500954
rect 300768 500890 300820 500896
rect 301596 500948 301648 500954
rect 301596 500890 301648 500896
rect 308772 500948 308824 500954
rect 308772 500890 308824 500896
rect 309784 500948 309836 500954
rect 309784 500890 309836 500896
rect 287152 500336 287204 500342
rect 287152 500278 287204 500284
rect 279884 500268 279936 500274
rect 279884 500210 279936 500216
rect 284208 500268 284260 500274
rect 284208 500210 284260 500216
rect 279896 497964 279924 500210
rect 287164 497964 287192 500278
rect 294328 500268 294380 500274
rect 294328 500210 294380 500216
rect 294340 497964 294368 500210
rect 301608 497964 301636 500890
rect 308784 497964 308812 500890
rect 317340 500614 317368 700334
rect 324228 700324 324280 700330
rect 324228 700266 324280 700272
rect 316040 500608 316092 500614
rect 316040 500550 316092 500556
rect 317328 500608 317380 500614
rect 317328 500550 317380 500556
rect 316052 497964 316080 500550
rect 324240 500546 324268 700266
rect 323216 500540 323268 500546
rect 323216 500482 323268 500488
rect 324228 500540 324280 500546
rect 324228 500482 324280 500488
rect 323228 497964 323256 500482
rect 331140 499574 331168 700470
rect 332520 700398 332548 703520
rect 338028 700460 338080 700466
rect 338028 700402 338080 700408
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 330864 499546 331168 499574
rect 330864 497978 330892 499546
rect 338040 497978 338068 700402
rect 344928 700392 344980 700398
rect 344928 700334 344980 700340
rect 330510 497950 330892 497978
rect 337686 497950 338068 497978
rect 344940 497964 344968 700334
rect 348804 700330 348832 703520
rect 360108 700936 360160 700942
rect 360108 700878 360160 700884
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 353208 700324 353260 700330
rect 353208 700266 353260 700272
rect 353220 500478 353248 700266
rect 360120 500954 360148 700878
rect 364996 700534 365024 703520
rect 367008 700868 367060 700874
rect 367008 700810 367060 700816
rect 364984 700528 365036 700534
rect 364984 700470 365036 700476
rect 359372 500948 359424 500954
rect 359372 500890 359424 500896
rect 360108 500948 360160 500954
rect 360108 500890 360160 500896
rect 352104 500472 352156 500478
rect 352104 500414 352156 500420
rect 353208 500472 353260 500478
rect 353208 500414 353260 500420
rect 352116 497964 352144 500414
rect 359384 497964 359412 500890
rect 367020 499574 367048 700810
rect 373908 700800 373960 700806
rect 373908 700742 373960 700748
rect 366928 499546 367048 499574
rect 366928 497978 366956 499546
rect 373920 497978 373948 700742
rect 381188 700466 381216 703520
rect 382188 700732 382240 700738
rect 382188 700674 382240 700680
rect 381176 700460 381228 700466
rect 381176 700402 381228 700408
rect 382200 500954 382228 700674
rect 389088 700664 389140 700670
rect 389088 700606 389140 700612
rect 389100 500954 389128 700606
rect 395988 700596 396040 700602
rect 395988 700538 396040 700544
rect 380992 500948 381044 500954
rect 380992 500890 381044 500896
rect 382188 500948 382240 500954
rect 382188 500890 382240 500896
rect 388260 500948 388312 500954
rect 388260 500890 388312 500896
rect 389088 500948 389140 500954
rect 389088 500890 389140 500896
rect 366574 497950 366956 497978
rect 373842 497950 373948 497978
rect 381004 497964 381032 500890
rect 388272 497964 388300 500890
rect 396000 499574 396028 700538
rect 397472 700398 397500 703520
rect 402888 700528 402940 700534
rect 402888 700470 402940 700476
rect 397460 700392 397512 700398
rect 397460 700334 397512 700340
rect 395816 499546 396028 499574
rect 395816 497978 395844 499546
rect 402900 497978 402928 700470
rect 411168 700460 411220 700466
rect 411168 700402 411220 700408
rect 411180 500614 411208 700402
rect 413664 700330 413692 703520
rect 429856 700942 429884 703520
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 446140 700874 446168 703520
rect 446128 700868 446180 700874
rect 446128 700810 446180 700816
rect 462332 700806 462360 703520
rect 462320 700800 462372 700806
rect 462320 700742 462372 700748
rect 478524 700738 478552 703520
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 511000 700602 511028 703520
rect 510988 700596 511040 700602
rect 510988 700538 511040 700544
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 418068 700392 418120 700398
rect 418068 700334 418120 700340
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 418080 500954 418108 700334
rect 575860 700330 575888 703520
rect 424968 700324 425020 700330
rect 424968 700266 425020 700272
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 417148 500948 417200 500954
rect 417148 500890 417200 500896
rect 418068 500948 418120 500954
rect 418068 500890 418120 500896
rect 409880 500608 409932 500614
rect 409880 500550 409932 500556
rect 411168 500608 411220 500614
rect 411168 500550 411220 500556
rect 395462 497950 395844 497978
rect 402730 497950 402928 497978
rect 409892 497964 409920 500550
rect 417160 497964 417188 500890
rect 424980 499574 425008 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 429844 696992 429896 696998
rect 429844 696934 429896 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 429752 563100 429804 563106
rect 429752 563042 429804 563048
rect 429660 536852 429712 536858
rect 429660 536794 429712 536800
rect 429568 524476 429620 524482
rect 429568 524418 429620 524424
rect 424704 499546 425008 499574
rect 424704 497978 424732 499546
rect 424350 497950 424732 497978
rect 165620 494012 165672 494018
rect 165620 493954 165672 493960
rect 165632 493377 165660 493954
rect 165618 493368 165674 493377
rect 165618 493303 165674 493312
rect 165620 491292 165672 491298
rect 165620 491234 165672 491240
rect 165632 490385 165660 491234
rect 165618 490376 165674 490385
rect 165618 490311 165674 490320
rect 165620 488504 165672 488510
rect 165620 488446 165672 488452
rect 429384 488504 429436 488510
rect 429384 488446 429436 488452
rect 165632 487393 165660 488446
rect 429396 487393 429424 488446
rect 165618 487384 165674 487393
rect 165618 487319 165674 487328
rect 429382 487384 429438 487393
rect 429382 487319 429438 487328
rect 165620 485784 165672 485790
rect 165620 485726 165672 485732
rect 165632 484537 165660 485726
rect 165618 484528 165674 484537
rect 165618 484463 165674 484472
rect 165620 481636 165672 481642
rect 165620 481578 165672 481584
rect 165632 481545 165660 481578
rect 165618 481536 165674 481545
rect 165618 481471 165674 481480
rect 165620 478848 165672 478854
rect 165620 478790 165672 478796
rect 165632 478553 165660 478790
rect 165618 478544 165674 478553
rect 165618 478479 165674 478488
rect 165620 476060 165672 476066
rect 165620 476002 165672 476008
rect 429476 476060 429528 476066
rect 429476 476002 429528 476008
rect 165632 475561 165660 476002
rect 165618 475552 165674 475561
rect 165618 475487 165674 475496
rect 429488 475289 429516 476002
rect 429474 475280 429530 475289
rect 429474 475215 429530 475224
rect 4068 473340 4120 473346
rect 4068 473282 4120 473288
rect 165620 473340 165672 473346
rect 165620 473282 165672 473288
rect 165632 472705 165660 473282
rect 165618 472696 165674 472705
rect 165618 472631 165674 472640
rect 165620 470552 165672 470558
rect 165620 470494 165672 470500
rect 165632 469713 165660 470494
rect 165618 469704 165674 469713
rect 165618 469639 165674 469648
rect 165620 467832 165672 467838
rect 165620 467774 165672 467780
rect 165632 466721 165660 467774
rect 165618 466712 165674 466721
rect 165618 466647 165674 466656
rect 165620 465044 165672 465050
rect 165620 464986 165672 464992
rect 165632 463729 165660 464986
rect 165618 463720 165674 463729
rect 165618 463655 165674 463664
rect 429200 463684 429252 463690
rect 429200 463626 429252 463632
rect 429212 463185 429240 463626
rect 429198 463176 429254 463185
rect 429198 463111 429254 463120
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3516 447092 3568 447098
rect 3516 447034 3568 447040
rect 3620 444378 3648 462567
rect 165620 460896 165672 460902
rect 165620 460838 165672 460844
rect 165632 460737 165660 460838
rect 165618 460728 165674 460737
rect 165618 460663 165674 460672
rect 165620 458176 165672 458182
rect 165620 458118 165672 458124
rect 165632 457881 165660 458118
rect 165618 457872 165674 457881
rect 165618 457807 165674 457816
rect 429580 457201 429608 524418
rect 429672 460193 429700 536794
rect 429764 466177 429792 563042
rect 429856 496369 429884 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 429936 683188 429988 683194
rect 429936 683130 429988 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 429842 496360 429898 496369
rect 429842 496295 429898 496304
rect 429948 493377 429976 683130
rect 430028 670744 430080 670750
rect 580172 670744 580224 670750
rect 430028 670686 430080 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 429934 493368 429990 493377
rect 429934 493303 429990 493312
rect 430040 490385 430068 670686
rect 580170 670647 580226 670656
rect 580262 657384 580318 657393
rect 580262 657319 580318 657328
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 430120 643136 430172 643142
rect 430120 643078 430172 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 430026 490376 430082 490385
rect 430026 490311 430082 490320
rect 429844 484424 429896 484430
rect 430132 484401 430160 643078
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 430212 630692 430264 630698
rect 430212 630634 430264 630640
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 429844 484366 429896 484372
rect 430118 484392 430174 484401
rect 429750 466168 429806 466177
rect 429750 466103 429806 466112
rect 429658 460184 429714 460193
rect 429658 460119 429714 460128
rect 429566 457192 429622 457201
rect 429566 457127 429622 457136
rect 165620 455388 165672 455394
rect 165620 455330 165672 455336
rect 429200 455388 429252 455394
rect 429200 455330 429252 455336
rect 165632 454889 165660 455330
rect 165618 454880 165674 454889
rect 165618 454815 165674 454824
rect 429212 454209 429240 455330
rect 429198 454200 429254 454209
rect 429198 454135 429254 454144
rect 165620 452600 165672 452606
rect 165620 452542 165672 452548
rect 165632 451897 165660 452542
rect 165618 451888 165674 451897
rect 165618 451823 165674 451832
rect 429568 451240 429620 451246
rect 429568 451182 429620 451188
rect 429580 451081 429608 451182
rect 429566 451072 429622 451081
rect 429566 451007 429622 451016
rect 165620 449880 165672 449886
rect 165620 449822 165672 449828
rect 3698 449576 3754 449585
rect 3698 449511 3754 449520
rect 3608 444372 3660 444378
rect 3608 444314 3660 444320
rect 3712 440230 3740 449511
rect 165632 448905 165660 449822
rect 165618 448896 165674 448905
rect 165618 448831 165674 448840
rect 429856 448089 429884 484366
rect 430118 484327 430174 484336
rect 430224 481273 430252 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 430304 616888 430356 616894
rect 430304 616830 430356 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 430210 481264 430266 481273
rect 430210 481199 430266 481208
rect 430316 478281 430344 616830
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 430396 590708 430448 590714
rect 430396 590650 430448 590656
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 430302 478272 430358 478281
rect 430302 478207 430358 478216
rect 430408 472297 430436 590650
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 430488 576904 430540 576910
rect 430488 576846 430540 576852
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 430394 472288 430450 472297
rect 430394 472223 430450 472232
rect 429936 470620 429988 470626
rect 429936 470562 429988 470568
rect 429842 448080 429898 448089
rect 429842 448015 429898 448024
rect 165620 447092 165672 447098
rect 165620 447034 165672 447040
rect 165632 446049 165660 447034
rect 165618 446040 165674 446049
rect 165618 445975 165674 445984
rect 429948 445097 429976 470562
rect 430500 469305 430528 576846
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580276 488510 580304 657319
rect 580354 604208 580410 604217
rect 580354 604143 580410 604152
rect 580264 488504 580316 488510
rect 580264 488446 580316 488452
rect 579618 484664 579674 484673
rect 579618 484599 579674 484608
rect 579632 484430 579660 484599
rect 579620 484424 579672 484430
rect 579620 484366 579672 484372
rect 580368 476066 580396 604143
rect 580446 551168 580502 551177
rect 580446 551103 580502 551112
rect 580356 476060 580408 476066
rect 580356 476002 580408 476008
rect 579618 471472 579674 471481
rect 579618 471407 579674 471416
rect 579632 470626 579660 471407
rect 579620 470620 579672 470626
rect 579620 470562 579672 470568
rect 430486 469296 430542 469305
rect 430486 469231 430542 469240
rect 580460 463690 580488 551103
rect 580538 511320 580594 511329
rect 580538 511255 580594 511264
rect 580448 463684 580500 463690
rect 580448 463626 580500 463632
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 430028 456816 430080 456822
rect 430028 456758 430080 456764
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 429934 445088 429990 445097
rect 429934 445023 429990 445032
rect 429844 444440 429896 444446
rect 429844 444382 429896 444388
rect 165620 444372 165672 444378
rect 165620 444314 165672 444320
rect 165632 443057 165660 444314
rect 165618 443048 165674 443057
rect 165618 442983 165674 442992
rect 3700 440224 3752 440230
rect 3700 440166 3752 440172
rect 165620 440224 165672 440230
rect 165620 440166 165672 440172
rect 165632 440065 165660 440166
rect 165618 440056 165674 440065
rect 165618 439991 165674 440000
rect 429856 439113 429884 444382
rect 430040 442105 430068 456758
rect 580552 455394 580580 511255
rect 580630 497992 580686 498001
rect 580630 497927 580686 497936
rect 580540 455388 580592 455394
rect 580540 455330 580592 455336
rect 580644 451246 580672 497927
rect 580632 451240 580684 451246
rect 580632 451182 580684 451188
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580184 444446 580212 444751
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 430026 442096 430082 442105
rect 430026 442031 430082 442040
rect 429842 439104 429898 439113
rect 429842 439039 429898 439048
rect 165618 437064 165674 437073
rect 165618 436999 165674 437008
rect 165632 436762 165660 436999
rect 3424 436756 3476 436762
rect 3424 436698 3476 436704
rect 165620 436756 165672 436762
rect 165620 436698 165672 436704
rect 3436 436665 3464 436698
rect 3422 436656 3478 436665
rect 3422 436591 3478 436600
rect 429934 436112 429990 436121
rect 429934 436047 429990 436056
rect 165618 434072 165674 434081
rect 165618 434007 165674 434016
rect 165632 433362 165660 434007
rect 3424 433356 3476 433362
rect 3424 433298 3476 433304
rect 165620 433356 165672 433362
rect 165620 433298 165672 433304
rect 3436 423609 3464 433298
rect 429842 432984 429898 432993
rect 429842 432919 429898 432928
rect 165618 431216 165674 431225
rect 165618 431151 165674 431160
rect 165632 430642 165660 431151
rect 3792 430636 3844 430642
rect 3792 430578 3844 430584
rect 165620 430636 165672 430642
rect 165620 430578 165672 430584
rect 3700 427848 3752 427854
rect 3700 427790 3752 427796
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3608 420980 3660 420986
rect 3608 420922 3660 420928
rect 3516 418192 3568 418198
rect 3516 418134 3568 418140
rect 3424 415472 3476 415478
rect 3424 415414 3476 415420
rect 3148 407176 3200 407182
rect 3148 407118 3200 407124
rect 3056 332580 3108 332586
rect 3056 332522 3108 332528
rect 3068 332353 3096 332522
rect 3054 332344 3110 332353
rect 3054 332279 3110 332288
rect 3056 320136 3108 320142
rect 3056 320078 3108 320084
rect 3068 319297 3096 320078
rect 3054 319288 3110 319297
rect 3054 319223 3110 319232
rect 3160 306241 3188 407118
rect 3240 404388 3292 404394
rect 3240 404330 3292 404336
rect 3146 306232 3202 306241
rect 3146 306167 3202 306176
rect 3252 293185 3280 404330
rect 3332 385008 3384 385014
rect 3332 384950 3384 384956
rect 3344 384441 3372 384950
rect 3330 384432 3386 384441
rect 3330 384367 3386 384376
rect 3332 383716 3384 383722
rect 3332 383658 3384 383664
rect 3238 293176 3294 293185
rect 3238 293111 3294 293120
rect 3240 280152 3292 280158
rect 3238 280120 3240 280129
rect 3292 280120 3294 280129
rect 3238 280055 3294 280064
rect 3056 267708 3108 267714
rect 3056 267650 3108 267656
rect 3068 267209 3096 267650
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3240 255264 3292 255270
rect 3240 255206 3292 255212
rect 3252 254153 3280 255206
rect 3238 254144 3294 254153
rect 3238 254079 3294 254088
rect 3240 241256 3292 241262
rect 3240 241198 3292 241204
rect 3252 241097 3280 241198
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3240 229084 3292 229090
rect 3240 229026 3292 229032
rect 3252 228041 3280 229026
rect 3238 228032 3294 228041
rect 3238 227967 3294 227976
rect 3240 215280 3292 215286
rect 3240 215222 3292 215228
rect 3252 214985 3280 215222
rect 3238 214976 3294 214985
rect 3238 214911 3294 214920
rect 3344 201929 3372 383658
rect 3436 345409 3464 415414
rect 3528 358465 3556 418134
rect 3620 371385 3648 420922
rect 3712 397497 3740 427790
rect 3804 410553 3832 430578
rect 165618 428224 165674 428233
rect 165618 428159 165674 428168
rect 165632 427854 165660 428159
rect 165620 427848 165672 427854
rect 165620 427790 165672 427796
rect 166262 425232 166318 425241
rect 166262 425167 166318 425176
rect 165618 422240 165674 422249
rect 165618 422175 165674 422184
rect 165632 420986 165660 422175
rect 165620 420980 165672 420986
rect 165620 420922 165672 420928
rect 165618 419384 165674 419393
rect 165618 419319 165674 419328
rect 165632 418198 165660 419319
rect 165620 418192 165672 418198
rect 165620 418134 165672 418140
rect 165618 416392 165674 416401
rect 165618 416327 165674 416336
rect 165632 415478 165660 416327
rect 165620 415472 165672 415478
rect 165620 415414 165672 415420
rect 3790 410544 3846 410553
rect 3790 410479 3846 410488
rect 165618 407416 165674 407425
rect 165618 407351 165674 407360
rect 165632 407182 165660 407351
rect 165620 407176 165672 407182
rect 165620 407118 165672 407124
rect 165618 404560 165674 404569
rect 165618 404495 165674 404504
rect 165632 404394 165660 404495
rect 165620 404388 165672 404394
rect 165620 404330 165672 404336
rect 3698 397488 3754 397497
rect 3698 397423 3754 397432
rect 165618 395584 165674 395593
rect 165618 395519 165674 395528
rect 165632 394738 165660 395519
rect 22744 394732 22796 394738
rect 22744 394674 22796 394680
rect 165620 394732 165672 394738
rect 165620 394674 165672 394680
rect 7564 392012 7616 392018
rect 7564 391954 7616 391960
rect 4068 374060 4120 374066
rect 4068 374002 4120 374008
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3976 368552 4028 368558
rect 3976 368494 4028 368500
rect 3884 362976 3936 362982
rect 3884 362918 3936 362924
rect 3792 358828 3844 358834
rect 3792 358770 3844 358776
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3700 353320 3752 353326
rect 3700 353262 3752 353268
rect 3608 347812 3660 347818
rect 3608 347754 3660 347760
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3516 345092 3568 345098
rect 3516 345034 3568 345040
rect 3424 342304 3476 342310
rect 3424 342246 3476 342252
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3332 176656 3384 176662
rect 3332 176598 3384 176604
rect 3344 175953 3372 176598
rect 3330 175944 3386 175953
rect 3330 175879 3386 175888
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3148 124160 3200 124166
rect 3148 124102 3200 124108
rect 3160 123729 3188 124102
rect 3146 123720 3202 123729
rect 3146 123655 3202 123664
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 2872 59356 2924 59362
rect 2872 59298 2924 59304
rect 2884 58585 2912 59298
rect 2870 58576 2926 58585
rect 2870 58511 2926 58520
rect 3436 19417 3464 342246
rect 3528 32473 3556 345034
rect 3620 45529 3648 347754
rect 3712 71641 3740 353262
rect 3804 97617 3832 358770
rect 3896 110673 3924 362918
rect 3988 136785 4016 368494
rect 4080 162897 4108 374002
rect 7576 241262 7604 391954
rect 14464 379568 14516 379574
rect 14464 379510 14516 379516
rect 10324 336048 10376 336054
rect 10324 335990 10376 335996
rect 7564 241256 7616 241262
rect 7564 241198 7616 241204
rect 4066 162888 4122 162897
rect 4066 162823 4122 162832
rect 3974 136776 4030 136785
rect 3974 136711 4030 136720
rect 3882 110664 3938 110673
rect 3882 110599 3938 110608
rect 3790 97608 3846 97617
rect 3790 97543 3846 97552
rect 3698 71632 3754 71641
rect 3698 71567 3754 71576
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8772 480 8800 6190
rect 10336 3466 10364 335990
rect 11704 327752 11756 327758
rect 11704 327694 11756 327700
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 480 9996 2926
rect 11164 480 11192 2994
rect 11716 2990 11744 327694
rect 14476 189038 14504 379510
rect 15844 356108 15896 356114
rect 15844 356050 15896 356056
rect 14464 189032 14516 189038
rect 14464 188974 14516 188980
rect 15856 85542 15884 356050
rect 17224 338156 17276 338162
rect 17224 338098 17276 338104
rect 15844 85536 15896 85542
rect 15844 85478 15896 85484
rect 17236 6866 17264 338098
rect 18604 336116 18656 336122
rect 18604 336058 18656 336064
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 12360 480 12388 5034
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 14738 3496 14794 3505
rect 13544 3460 13596 3466
rect 14738 3431 14794 3440
rect 13544 3402 13596 3408
rect 13556 480 13584 3402
rect 14752 480 14780 3431
rect 15948 480 15976 3567
rect 17052 480 17080 5102
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 480 18276 3470
rect 18616 3058 18644 336058
rect 21364 330540 21416 330546
rect 21364 330482 21416 330488
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 19444 480 19472 3538
rect 20640 480 20668 4082
rect 21376 3466 21404 330482
rect 22756 255270 22784 394674
rect 165618 392728 165674 392737
rect 165618 392663 165674 392672
rect 165632 392018 165660 392663
rect 165620 392012 165672 392018
rect 165620 391954 165672 391960
rect 166276 385014 166304 425167
rect 429856 419490 429884 432919
rect 429948 431934 429976 436047
rect 429936 431928 429988 431934
rect 429936 431870 429988 431876
rect 579804 431928 579856 431934
rect 579804 431870 579856 431876
rect 579816 431633 579844 431870
rect 579802 431624 579858 431633
rect 579802 431559 579858 431568
rect 430210 429992 430266 430001
rect 430210 429927 430266 429936
rect 430118 427000 430174 427009
rect 430118 426935 430174 426944
rect 430026 424008 430082 424017
rect 430026 423943 430082 423952
rect 429934 421016 429990 421025
rect 429934 420951 429990 420960
rect 429844 419484 429896 419490
rect 429844 419426 429896 419432
rect 429842 417888 429898 417897
rect 429842 417823 429898 417832
rect 429566 414896 429622 414905
rect 429566 414831 429568 414840
rect 429620 414831 429622 414840
rect 429568 414802 429620 414808
rect 166906 413400 166962 413409
rect 166906 413335 166962 413344
rect 166814 410408 166870 410417
rect 166814 410343 166870 410352
rect 166722 401568 166778 401577
rect 166722 401503 166778 401512
rect 166630 398576 166686 398585
rect 166630 398511 166686 398520
rect 166538 389736 166594 389745
rect 166538 389671 166594 389680
rect 166446 386744 166502 386753
rect 166446 386679 166502 386688
rect 166264 385008 166316 385014
rect 166264 384950 166316 384956
rect 165618 383752 165674 383761
rect 165618 383687 165620 383696
rect 165672 383687 165674 383696
rect 165620 383658 165672 383664
rect 165618 380760 165674 380769
rect 165618 380695 165674 380704
rect 165632 379574 165660 380695
rect 165620 379568 165672 379574
rect 165620 379510 165672 379516
rect 166354 377904 166410 377913
rect 166354 377839 166410 377848
rect 165618 374912 165674 374921
rect 165618 374847 165674 374856
rect 165632 374066 165660 374847
rect 165620 374060 165672 374066
rect 165620 374002 165672 374008
rect 165618 371920 165674 371929
rect 165618 371855 165674 371864
rect 165632 371278 165660 371855
rect 25504 371272 25556 371278
rect 25504 371214 25556 371220
rect 165620 371272 165672 371278
rect 165620 371214 165672 371220
rect 22744 255264 22796 255270
rect 22744 255206 22796 255212
rect 22744 253224 22796 253230
rect 22744 253166 22796 253172
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21836 480 21864 6258
rect 22756 3534 22784 253166
rect 25516 150414 25544 371214
rect 165618 368928 165674 368937
rect 165618 368863 165674 368872
rect 165632 368558 165660 368863
rect 165620 368552 165672 368558
rect 165620 368494 165672 368500
rect 166262 366072 166318 366081
rect 166262 366007 166318 366016
rect 165618 363080 165674 363089
rect 165618 363015 165674 363024
rect 165632 362982 165660 363015
rect 165620 362976 165672 362982
rect 165620 362918 165672 362924
rect 165618 360088 165674 360097
rect 165618 360023 165674 360032
rect 165632 358834 165660 360023
rect 165620 358828 165672 358834
rect 165620 358770 165672 358776
rect 165618 357096 165674 357105
rect 165618 357031 165674 357040
rect 165632 356114 165660 357031
rect 165620 356108 165672 356114
rect 165620 356050 165672 356056
rect 165618 354104 165674 354113
rect 165618 354039 165674 354048
rect 165632 353326 165660 354039
rect 165620 353320 165672 353326
rect 165620 353262 165672 353268
rect 165618 351248 165674 351257
rect 165618 351183 165674 351192
rect 165632 350606 165660 351183
rect 32404 350600 32456 350606
rect 32404 350542 32456 350548
rect 165620 350600 165672 350606
rect 165620 350542 165672 350548
rect 29644 336252 29696 336258
rect 29644 336194 29696 336200
rect 28264 336184 28316 336190
rect 28264 336126 28316 336132
rect 25596 177336 25648 177342
rect 25596 177278 25648 177284
rect 25504 150408 25556 150414
rect 25504 150350 25556 150356
rect 24214 3768 24270 3777
rect 24214 3703 24270 3712
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23032 480 23060 3470
rect 24228 480 24256 3703
rect 25608 3534 25636 177278
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25332 480 25360 3402
rect 26528 480 26556 6326
rect 28276 4146 28304 336126
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 29656 3670 29684 336194
rect 32416 59362 32444 350542
rect 165618 348256 165674 348265
rect 165618 348191 165674 348200
rect 165632 347818 165660 348191
rect 165620 347812 165672 347818
rect 165620 347754 165672 347760
rect 165618 345264 165674 345273
rect 165618 345199 165674 345208
rect 165632 345098 165660 345199
rect 165620 345092 165672 345098
rect 165620 345034 165672 345040
rect 165620 342304 165672 342310
rect 165618 342272 165620 342281
rect 165672 342272 165674 342281
rect 165618 342207 165674 342216
rect 165618 339416 165674 339425
rect 165618 339351 165674 339360
rect 165632 338162 165660 339351
rect 165620 338156 165672 338162
rect 165620 338098 165672 338104
rect 159364 336524 159416 336530
rect 159364 336466 159416 336472
rect 125508 336456 125560 336462
rect 125508 336398 125560 336404
rect 114468 336388 114520 336394
rect 114468 336330 114520 336336
rect 35164 336320 35216 336326
rect 35164 336262 35216 336268
rect 33784 309800 33836 309806
rect 33784 309742 33836 309748
rect 32404 59356 32456 59362
rect 32404 59298 32456 59304
rect 33600 6520 33652 6526
rect 33600 6462 33652 6468
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28920 480 28948 3538
rect 30116 480 30144 6394
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31300 3256 31352 3262
rect 31300 3198 31352 3204
rect 31312 480 31340 3198
rect 32416 480 32444 3470
rect 33612 480 33640 6462
rect 33796 3058 33824 309742
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 33784 3052 33836 3058
rect 33784 2994 33836 3000
rect 34808 480 34836 3742
rect 35176 3602 35204 336262
rect 39304 334620 39356 334626
rect 39304 334562 39356 334568
rect 36544 304292 36596 304298
rect 36544 304234 36596 304240
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 36004 480 36032 3538
rect 36556 3262 36584 304234
rect 37188 6588 37240 6594
rect 37188 6530 37240 6536
rect 36544 3256 36596 3262
rect 36544 3198 36596 3204
rect 37200 480 37228 6530
rect 39316 3806 39344 334562
rect 95148 333260 95200 333266
rect 95148 333202 95200 333208
rect 88248 326392 88300 326398
rect 88248 326334 88300 326340
rect 40684 324964 40736 324970
rect 40684 324906 40736 324912
rect 39304 3800 39356 3806
rect 39304 3742 39356 3748
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 38384 3120 38436 3126
rect 38384 3062 38436 3068
rect 38396 480 38424 3062
rect 39592 480 39620 3606
rect 40696 3126 40724 324906
rect 53748 323604 53800 323610
rect 53748 323546 53800 323552
rect 43444 305652 43496 305658
rect 43444 305594 43496 305600
rect 40776 6656 40828 6662
rect 40776 6598 40828 6604
rect 40684 3120 40736 3126
rect 40684 3062 40736 3068
rect 40788 2938 40816 6598
rect 43076 3732 43128 3738
rect 43076 3674 43128 3680
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 40696 2910 40816 2938
rect 40696 480 40724 2910
rect 41892 480 41920 3130
rect 43088 480 43116 3674
rect 43456 3194 43484 305594
rect 50988 301504 51040 301510
rect 50988 301446 51040 301452
rect 46204 300144 46256 300150
rect 46204 300086 46256 300092
rect 44272 6724 44324 6730
rect 44272 6666 44324 6672
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 44284 480 44312 6666
rect 46216 4146 46244 300086
rect 48964 6792 49016 6798
rect 48964 6734 49016 6740
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 45480 480 45508 4082
rect 46664 3800 46716 3806
rect 46664 3742 46716 3748
rect 46676 480 46704 3742
rect 47872 480 47900 5170
rect 48976 480 49004 6734
rect 51000 3398 51028 301446
rect 52552 7608 52604 7614
rect 52552 7550 52604 7556
rect 51356 5296 51408 5302
rect 51356 5238 51408 5244
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 50172 480 50200 3334
rect 51368 480 51396 5238
rect 52564 480 52592 7550
rect 53760 480 53788 323546
rect 57888 302932 57940 302938
rect 57888 302874 57940 302880
rect 56048 7676 56100 7682
rect 56048 7618 56100 7624
rect 54944 5364 54996 5370
rect 54944 5306 54996 5312
rect 54956 480 54984 5306
rect 56060 480 56088 7618
rect 57900 3398 57928 302874
rect 61936 298784 61988 298790
rect 61936 298726 61988 298732
rect 59636 7744 59688 7750
rect 59636 7686 59688 7692
rect 58440 5432 58492 5438
rect 58440 5374 58492 5380
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 57256 480 57284 3334
rect 58452 480 58480 5374
rect 59648 480 59676 7686
rect 61948 3398 61976 298726
rect 64788 297424 64840 297430
rect 64788 297366 64840 297372
rect 63224 7812 63276 7818
rect 63224 7754 63276 7760
rect 62028 5500 62080 5506
rect 62028 5442 62080 5448
rect 60832 3392 60884 3398
rect 60832 3334 60884 3340
rect 61936 3392 61988 3398
rect 61936 3334 61988 3340
rect 60844 480 60872 3334
rect 62040 480 62068 5442
rect 63236 480 63264 7754
rect 64800 3398 64828 297366
rect 68928 294636 68980 294642
rect 68928 294578 68980 294584
rect 66720 8968 66772 8974
rect 66720 8910 66772 8916
rect 65524 4752 65576 4758
rect 65524 4694 65576 4700
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64340 480 64368 3334
rect 65536 480 65564 4694
rect 66732 480 66760 8910
rect 68940 3398 68968 294578
rect 85488 17264 85540 17270
rect 85488 17206 85540 17212
rect 81348 10328 81400 10334
rect 81348 10270 81400 10276
rect 77392 9172 77444 9178
rect 77392 9114 77444 9120
rect 73804 9104 73856 9110
rect 73804 9046 73856 9052
rect 70308 9036 70360 9042
rect 70308 8978 70360 8984
rect 69112 4616 69164 4622
rect 69112 4558 69164 4564
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 67928 480 67956 3334
rect 69124 480 69152 4558
rect 70320 480 70348 8978
rect 72608 4684 72660 4690
rect 72608 4626 72660 4632
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 71516 480 71544 3810
rect 72620 480 72648 4626
rect 73816 480 73844 9046
rect 76196 4548 76248 4554
rect 76196 4490 76248 4496
rect 75000 3936 75052 3942
rect 75000 3878 75052 3884
rect 75012 480 75040 3878
rect 76208 480 76236 4490
rect 77404 480 77432 9114
rect 79692 4480 79744 4486
rect 79692 4422 79744 4428
rect 78588 4004 78640 4010
rect 78588 3946 78640 3952
rect 78600 480 78628 3946
rect 79704 480 79732 4422
rect 81360 3398 81388 10270
rect 83280 6860 83332 6866
rect 83280 6802 83332 6808
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82096 480 82124 4014
rect 83292 480 83320 6802
rect 85500 3398 85528 17206
rect 86868 7880 86920 7886
rect 86868 7822 86920 7828
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 85488 3392 85540 3398
rect 85488 3334 85540 3340
rect 84488 480 84516 3334
rect 85684 480 85712 4082
rect 86880 480 86908 7822
rect 88260 6914 88288 326334
rect 92388 28280 92440 28286
rect 92388 28222 92440 28228
rect 90364 7948 90416 7954
rect 90364 7890 90416 7896
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 89180 480 89208 3266
rect 90376 480 90404 7890
rect 92400 3398 92428 28222
rect 93952 8016 94004 8022
rect 93952 7958 94004 7964
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 92388 3392 92440 3398
rect 92388 3334 92440 3340
rect 91572 480 91600 3334
rect 92756 3324 92808 3330
rect 92756 3266 92808 3272
rect 92768 480 92796 3266
rect 93964 480 93992 7958
rect 95160 480 95188 333202
rect 113088 318096 113140 318102
rect 113088 318038 113140 318044
rect 99288 311160 99340 311166
rect 99288 311102 99340 311108
rect 97448 8084 97500 8090
rect 97448 8026 97500 8032
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96264 480 96292 3130
rect 97460 480 97488 8026
rect 99300 3262 99328 311102
rect 106188 307080 106240 307086
rect 106188 307022 106240 307028
rect 103428 18624 103480 18630
rect 103428 18566 103480 18572
rect 101036 8152 101088 8158
rect 101036 8094 101088 8100
rect 98644 3256 98696 3262
rect 98644 3198 98696 3204
rect 99288 3256 99340 3262
rect 99288 3198 99340 3204
rect 98656 480 98684 3198
rect 99840 3052 99892 3058
rect 99840 2994 99892 3000
rect 99852 480 99880 2994
rect 101048 480 101076 8094
rect 103440 3194 103468 18566
rect 104532 8220 104584 8226
rect 104532 8162 104584 8168
rect 102232 3188 102284 3194
rect 102232 3130 102284 3136
rect 103428 3188 103480 3194
rect 103428 3130 103480 3136
rect 102244 480 102272 3130
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 103348 480 103376 3062
rect 104544 480 104572 8162
rect 106200 3194 106228 307022
rect 110328 11756 110380 11762
rect 110328 11698 110380 11704
rect 108120 8288 108172 8294
rect 108120 8230 108172 8236
rect 105728 3188 105780 3194
rect 105728 3130 105780 3136
rect 106188 3188 106240 3194
rect 106188 3130 106240 3136
rect 105740 480 105768 3130
rect 106924 2916 106976 2922
rect 106924 2858 106976 2864
rect 106936 480 106964 2858
rect 108132 480 108160 8230
rect 110340 3194 110368 11698
rect 111616 7540 111668 7546
rect 111616 7482 111668 7488
rect 109316 3188 109368 3194
rect 109316 3130 109368 3136
rect 110328 3188 110380 3194
rect 110328 3130 110380 3136
rect 109328 480 109356 3130
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110524 480 110552 2926
rect 111628 480 111656 7482
rect 113100 6914 113128 318038
rect 112824 6886 113128 6914
rect 112824 480 112852 6886
rect 114480 3058 114508 336330
rect 119988 329112 120040 329118
rect 119988 329054 120040 329060
rect 117228 256012 117280 256018
rect 117228 255954 117280 255960
rect 115204 7472 115256 7478
rect 115204 7414 115256 7420
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 114468 3052 114520 3058
rect 114468 2994 114520 3000
rect 114020 480 114048 2994
rect 115216 480 115244 7414
rect 117240 3058 117268 255954
rect 118792 7404 118844 7410
rect 118792 7346 118844 7352
rect 116400 3052 116452 3058
rect 116400 2994 116452 3000
rect 117228 3052 117280 3058
rect 117228 2994 117280 3000
rect 116412 480 116440 2994
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 117608 480 117636 2790
rect 118804 480 118832 7346
rect 120000 6914 120028 329054
rect 124128 308440 124180 308446
rect 124128 308382 124180 308388
rect 122288 7336 122340 7342
rect 122288 7278 122340 7284
rect 119908 6886 120028 6914
rect 119908 480 119936 6886
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 121104 480 121132 2790
rect 122300 480 122328 7278
rect 124140 6914 124168 308382
rect 125520 6914 125548 336398
rect 126888 334688 126940 334694
rect 126888 334630 126940 334636
rect 126900 6914 126928 334630
rect 140688 331900 140740 331906
rect 140688 331842 140740 331848
rect 129648 329180 129700 329186
rect 129648 329122 129700 329128
rect 128268 14476 128320 14482
rect 128268 14418 128320 14424
rect 123496 6886 124168 6914
rect 124692 6886 125548 6914
rect 125888 6886 126928 6914
rect 123496 480 123524 6886
rect 124692 480 124720 6886
rect 125888 480 125916 6886
rect 128176 6112 128228 6118
rect 128176 6054 128228 6060
rect 126980 4208 127032 4214
rect 126980 4150 127032 4156
rect 126992 480 127020 4150
rect 128188 480 128216 6054
rect 128280 4214 128308 14418
rect 129660 6914 129688 329122
rect 131028 327820 131080 327826
rect 131028 327762 131080 327768
rect 131040 6914 131068 327762
rect 133788 325032 133840 325038
rect 133788 324974 133840 324980
rect 131764 13116 131816 13122
rect 131764 13058 131816 13064
rect 129384 6886 129688 6914
rect 130580 6886 131068 6914
rect 128268 4208 128320 4214
rect 128268 4150 128320 4156
rect 129384 480 129412 6886
rect 130580 480 130608 6886
rect 131776 480 131804 13058
rect 133800 6914 133828 324974
rect 136548 323672 136600 323678
rect 136548 323614 136600 323620
rect 135168 268388 135220 268394
rect 135168 268330 135220 268336
rect 135180 6914 135208 268330
rect 136456 35216 136508 35222
rect 136456 35158 136508 35164
rect 132972 6886 133828 6914
rect 134168 6886 135208 6914
rect 132972 480 133000 6886
rect 134168 480 134196 6886
rect 136468 4214 136496 35158
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 480 135300 4150
rect 136560 1442 136588 323614
rect 137928 316736 137980 316742
rect 137928 316678 137980 316684
rect 137940 6914 137968 316678
rect 139308 25560 139360 25566
rect 139308 25502 139360 25508
rect 139320 6914 139348 25502
rect 140700 6914 140728 331842
rect 147588 322244 147640 322250
rect 147588 322186 147640 322192
rect 144828 320884 144880 320890
rect 144828 320826 144880 320832
rect 142068 313948 142120 313954
rect 142068 313890 142120 313896
rect 142080 6914 142108 313890
rect 143448 312588 143500 312594
rect 143448 312530 143500 312536
rect 143460 6914 143488 312530
rect 136468 1414 136588 1442
rect 137664 6886 137968 6914
rect 138860 6886 139348 6914
rect 140056 6886 140728 6914
rect 141252 6886 142108 6914
rect 142448 6886 143488 6914
rect 136468 480 136496 1414
rect 137664 480 137692 6886
rect 138860 480 138888 6886
rect 140056 480 140084 6886
rect 141252 480 141280 6886
rect 142448 480 142476 6886
rect 144736 6044 144788 6050
rect 144736 5986 144788 5992
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 144748 480 144776 5986
rect 144840 4214 144868 320826
rect 146208 26920 146260 26926
rect 146208 26862 146260 26868
rect 146220 6914 146248 26862
rect 147600 6914 147628 322186
rect 159376 10334 159404 336466
rect 161388 333328 161440 333334
rect 161388 333270 161440 333276
rect 159364 10328 159416 10334
rect 159364 10270 159416 10276
rect 153016 7268 153068 7274
rect 153016 7210 153068 7216
rect 149520 7200 149572 7206
rect 149520 7142 149572 7148
rect 145944 6886 146248 6914
rect 147140 6886 147628 6914
rect 144828 4208 144880 4214
rect 144828 4150 144880 4156
rect 145944 480 145972 6886
rect 147140 480 147168 6886
rect 148324 5976 148376 5982
rect 148324 5918 148376 5924
rect 148336 480 148364 5918
rect 149532 480 149560 7142
rect 151820 5908 151872 5914
rect 151820 5850 151872 5856
rect 150624 4412 150676 4418
rect 150624 4354 150676 4360
rect 150636 480 150664 4354
rect 151832 480 151860 5850
rect 153028 480 153056 7210
rect 156604 7132 156656 7138
rect 156604 7074 156656 7080
rect 155408 5840 155460 5846
rect 155408 5782 155460 5788
rect 154212 4344 154264 4350
rect 154212 4286 154264 4292
rect 154224 480 154252 4286
rect 155420 480 155448 5782
rect 156616 480 156644 7074
rect 160100 7064 160152 7070
rect 160100 7006 160152 7012
rect 158904 5772 158956 5778
rect 158904 5714 158956 5720
rect 157800 4276 157852 4282
rect 157800 4218 157852 4224
rect 157812 480 157840 4218
rect 158916 480 158944 5714
rect 160112 480 160140 7006
rect 161400 6914 161428 333270
rect 165528 330608 165580 330614
rect 165528 330550 165580 330556
rect 162768 315308 162820 315314
rect 162768 315250 162820 315256
rect 162780 6914 162808 315250
rect 165540 6914 165568 330550
rect 166276 124166 166304 366007
rect 166368 176662 166396 377839
rect 166460 215286 166488 386679
rect 166552 229090 166580 389671
rect 166644 267714 166672 398511
rect 166736 280158 166764 401503
rect 166828 320142 166856 410343
rect 166920 332586 166948 413335
rect 429566 411904 429622 411913
rect 429566 411839 429622 411848
rect 429580 411330 429608 411839
rect 429568 411324 429620 411330
rect 429568 411266 429620 411272
rect 429474 408912 429530 408921
rect 429474 408847 429530 408856
rect 429488 408542 429516 408847
rect 429476 408536 429528 408542
rect 429476 408478 429528 408484
rect 429198 405920 429254 405929
rect 429198 405855 429254 405864
rect 429106 339552 429162 339561
rect 429106 339487 429108 339496
rect 429160 339487 429162 339496
rect 429108 339458 429160 339464
rect 167748 338014 168222 338042
rect 168484 338014 168682 338042
rect 168944 338014 169234 338042
rect 169786 338014 169892 338042
rect 166908 332580 166960 332586
rect 166908 332522 166960 332528
rect 166816 320136 166868 320142
rect 166816 320078 166868 320084
rect 167748 316034 167776 338014
rect 168380 330472 168432 330478
rect 168380 330414 168432 330420
rect 167012 316006 167776 316034
rect 166724 280152 166776 280158
rect 166724 280094 166776 280100
rect 166632 267708 166684 267714
rect 166632 267650 166684 267656
rect 166540 229084 166592 229090
rect 166540 229026 166592 229032
rect 166448 215280 166500 215286
rect 166448 215222 166500 215228
rect 166356 176656 166408 176662
rect 166356 176598 166408 176604
rect 166908 174548 166960 174554
rect 166908 174490 166960 174496
rect 166264 124160 166316 124166
rect 166264 124102 166316 124108
rect 166920 6914 166948 174490
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 164896 6886 165568 6914
rect 166092 6886 166948 6914
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 163688 5704 163740 5710
rect 163688 5646 163740 5652
rect 162768 5092 162820 5098
rect 162768 5034 162820 5040
rect 162780 4962 162808 5034
rect 162768 4956 162820 4962
rect 162768 4898 162820 4904
rect 163700 480 163728 5646
rect 164896 480 164924 6886
rect 166092 480 166120 6886
rect 167012 4894 167040 316006
rect 167184 5636 167236 5642
rect 167184 5578 167236 5584
rect 167000 4888 167052 4894
rect 167000 4830 167052 4836
rect 167196 480 167224 5578
rect 168392 4826 168420 330414
rect 168484 5030 168512 338014
rect 168944 330478 168972 338014
rect 168932 330472 168984 330478
rect 168932 330414 168984 330420
rect 169668 326460 169720 326466
rect 169668 326402 169720 326408
rect 169576 15904 169628 15910
rect 169576 15846 169628 15852
rect 168472 5024 168524 5030
rect 168472 4966 168524 4972
rect 168380 4820 168432 4826
rect 168380 4762 168432 4768
rect 168380 4208 168432 4214
rect 168380 4150 168432 4156
rect 168392 480 168420 4150
rect 169588 480 169616 15846
rect 169680 4214 169708 326402
rect 169864 6186 169892 338014
rect 170232 336054 170260 338028
rect 170324 338014 170798 338042
rect 171152 338014 171350 338042
rect 171428 338014 171902 338042
rect 172072 338014 172362 338042
rect 170220 336048 170272 336054
rect 170220 335990 170272 335996
rect 170324 316034 170352 338014
rect 169956 316006 170352 316034
rect 169852 6180 169904 6186
rect 169852 6122 169904 6128
rect 169668 4208 169720 4214
rect 169668 4150 169720 4156
rect 169956 3369 169984 316006
rect 170772 6180 170824 6186
rect 170772 6122 170824 6128
rect 169942 3360 169998 3369
rect 169942 3295 169998 3304
rect 170784 480 170812 6122
rect 171152 5098 171180 338014
rect 171428 335354 171456 338014
rect 171244 335326 171456 335354
rect 171244 6254 171272 335326
rect 172072 327758 172100 338014
rect 172900 336122 172928 338028
rect 173084 338014 173466 338042
rect 172888 336116 172940 336122
rect 172888 336058 172940 336064
rect 172060 327752 172112 327758
rect 172060 327694 172112 327700
rect 173084 316034 173112 338014
rect 173912 330546 173940 338028
rect 174004 338014 174478 338042
rect 174556 338014 175030 338042
rect 175476 338014 175582 338042
rect 175660 338014 176042 338042
rect 173900 330540 173952 330546
rect 173900 330482 173952 330488
rect 172624 316006 173112 316034
rect 172428 10328 172480 10334
rect 172428 10270 172480 10276
rect 171232 6248 171284 6254
rect 171232 6190 171284 6196
rect 171140 5092 171192 5098
rect 171140 5034 171192 5040
rect 172440 3534 172468 10270
rect 172624 5030 172652 316006
rect 173808 286340 173860 286346
rect 173808 286282 173860 286288
rect 172612 5024 172664 5030
rect 172612 4966 172664 4972
rect 173820 3534 173848 286282
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 172428 3528 172480 3534
rect 172428 3470 172480 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 174004 3505 174032 338014
rect 174556 316034 174584 338014
rect 175372 330540 175424 330546
rect 175372 330482 175424 330488
rect 174096 316006 174584 316034
rect 174096 3641 174124 316006
rect 175384 253230 175412 330482
rect 175372 253224 175424 253230
rect 175372 253166 175424 253172
rect 174268 6248 174320 6254
rect 174268 6190 174320 6196
rect 174082 3632 174138 3641
rect 174082 3567 174138 3576
rect 173808 3470 173860 3476
rect 173990 3496 174046 3505
rect 171980 480 172008 3470
rect 173176 480 173204 3470
rect 173990 3431 174046 3440
rect 174280 480 174308 6190
rect 175476 5166 175504 338014
rect 175660 330546 175688 338014
rect 176580 336258 176608 338028
rect 176568 336252 176620 336258
rect 176568 336194 176620 336200
rect 177132 336190 177160 338028
rect 177224 338014 177606 338042
rect 178158 338014 178264 338042
rect 177120 336184 177172 336190
rect 177120 336126 177172 336132
rect 175648 330540 175700 330546
rect 175648 330482 175700 330488
rect 176568 327752 176620 327758
rect 176568 327694 176620 327700
rect 175464 5160 175516 5166
rect 175464 5102 175516 5108
rect 176580 3534 176608 327694
rect 177224 316034 177252 338014
rect 178040 336728 178092 336734
rect 178040 336670 178092 336676
rect 176764 316006 177252 316034
rect 176764 6322 176792 316006
rect 177948 290488 178000 290494
rect 177948 290430 178000 290436
rect 177856 22772 177908 22778
rect 177856 22714 177908 22720
rect 176752 6316 176804 6322
rect 176752 6258 176804 6264
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 175476 480 175504 3470
rect 176672 480 176700 3470
rect 177868 480 177896 22714
rect 177960 3534 177988 290430
rect 178052 3777 178080 336670
rect 178132 324420 178184 324426
rect 178132 324362 178184 324368
rect 178144 4214 178172 324362
rect 178236 177342 178264 338014
rect 178328 338014 178710 338042
rect 178880 338014 179262 338042
rect 179432 338014 179722 338042
rect 179892 338014 180274 338042
rect 178328 336734 178356 338014
rect 178316 336728 178368 336734
rect 178316 336670 178368 336676
rect 178880 324426 178908 338014
rect 178868 324420 178920 324426
rect 178868 324362 178920 324368
rect 178224 177336 178276 177342
rect 178224 177278 178276 177284
rect 179052 11824 179104 11830
rect 179052 11766 179104 11772
rect 178132 4208 178184 4214
rect 178132 4150 178184 4156
rect 178038 3768 178094 3777
rect 178038 3703 178094 3712
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179064 480 179092 11766
rect 179432 6390 179460 338014
rect 179892 316034 179920 338014
rect 180812 336326 180840 338028
rect 180996 338014 181378 338042
rect 181456 338014 181838 338042
rect 180800 336320 180852 336326
rect 180800 336262 180852 336268
rect 180892 324420 180944 324426
rect 180892 324362 180944 324368
rect 180708 318164 180760 318170
rect 180708 318106 180760 318112
rect 179524 316006 179920 316034
rect 179524 309806 179552 316006
rect 179512 309800 179564 309806
rect 179512 309742 179564 309748
rect 179420 6384 179472 6390
rect 179420 6326 179472 6332
rect 180720 3534 180748 318106
rect 180904 304298 180932 324362
rect 180892 304292 180944 304298
rect 180892 304234 180944 304240
rect 180996 6458 181024 338014
rect 181456 324426 181484 338014
rect 182376 328454 182404 338028
rect 182284 328426 182404 328454
rect 182468 338014 182942 338042
rect 181444 324420 181496 324426
rect 181444 324362 181496 324368
rect 182284 323626 182312 328426
rect 182284 323598 182404 323626
rect 182272 323536 182324 323542
rect 182272 323478 182324 323484
rect 182088 19984 182140 19990
rect 182088 19926 182140 19932
rect 180984 6452 181036 6458
rect 180984 6394 181036 6400
rect 182100 3534 182128 19926
rect 182284 6526 182312 323478
rect 182272 6520 182324 6526
rect 182272 6462 182324 6468
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 181444 3528 181496 3534
rect 181444 3470 181496 3476
rect 182088 3528 182140 3534
rect 182088 3470 182140 3476
rect 180260 480 180288 3470
rect 181456 480 181484 3470
rect 182376 3466 182404 323598
rect 182468 323542 182496 338014
rect 183388 334626 183416 338028
rect 183572 338014 183954 338042
rect 184124 338014 184506 338042
rect 185058 338014 185164 338042
rect 183376 334620 183428 334626
rect 183376 334562 183428 334568
rect 182456 323536 182508 323542
rect 182456 323478 182508 323484
rect 183468 13184 183520 13190
rect 183468 13126 183520 13132
rect 183480 3534 183508 13126
rect 183572 3602 183600 338014
rect 184124 316034 184152 338014
rect 185136 324970 185164 338014
rect 185228 338014 185518 338042
rect 185688 338014 186070 338042
rect 186516 338014 186622 338042
rect 186792 338014 187082 338042
rect 187344 338014 187634 338042
rect 187804 338014 188186 338042
rect 188448 338014 188738 338042
rect 189198 338014 189304 338042
rect 185124 324964 185176 324970
rect 185124 324906 185176 324912
rect 185228 324850 185256 338014
rect 183664 316006 184152 316034
rect 184952 324822 185256 324850
rect 183664 6594 183692 316006
rect 184848 17332 184900 17338
rect 184848 17274 184900 17280
rect 183652 6588 183704 6594
rect 183652 6530 183704 6536
rect 183560 3596 183612 3602
rect 183560 3538 183612 3544
rect 184860 3534 184888 17274
rect 184952 3670 184980 324822
rect 185688 321554 185716 338014
rect 186320 326324 186372 326330
rect 186320 326266 186372 326272
rect 185044 321526 185716 321554
rect 185044 6662 185072 321526
rect 186136 10396 186188 10402
rect 186136 10338 186188 10344
rect 185124 9240 185176 9246
rect 185124 9182 185176 9188
rect 185032 6656 185084 6662
rect 185032 6598 185084 6604
rect 184940 3664 184992 3670
rect 184940 3606 184992 3612
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 184848 3528 184900 3534
rect 185136 3482 185164 9182
rect 184848 3470 184900 3476
rect 182364 3460 182416 3466
rect 182364 3402 182416 3408
rect 182560 480 182588 3470
rect 183756 480 183784 3470
rect 184952 3454 185164 3482
rect 184952 480 184980 3454
rect 186148 480 186176 10338
rect 186332 3738 186360 326266
rect 186412 324624 186464 324630
rect 186412 324566 186464 324572
rect 186424 6730 186452 324566
rect 186516 305658 186544 338014
rect 186792 326330 186820 338014
rect 186780 326324 186832 326330
rect 186780 326266 186832 326272
rect 187344 324630 187372 338014
rect 187700 326324 187752 326330
rect 187700 326266 187752 326272
rect 187332 324624 187384 324630
rect 187332 324566 187384 324572
rect 186504 305652 186556 305658
rect 186504 305594 186556 305600
rect 187608 18692 187660 18698
rect 187608 18634 187660 18640
rect 187620 6914 187648 18634
rect 187344 6886 187648 6914
rect 186412 6724 186464 6730
rect 186412 6666 186464 6672
rect 186320 3732 186372 3738
rect 186320 3674 186372 3680
rect 187344 480 187372 6886
rect 187712 3806 187740 326266
rect 187804 300150 187832 338014
rect 188344 336728 188396 336734
rect 188344 336670 188396 336676
rect 188356 301510 188384 336670
rect 188448 326330 188476 338014
rect 188436 326324 188488 326330
rect 188436 326266 188488 326272
rect 189172 326324 189224 326330
rect 189172 326266 189224 326272
rect 188344 301504 188396 301510
rect 188344 301446 188396 301452
rect 187792 300144 187844 300150
rect 187792 300086 187844 300092
rect 188988 21412 189040 21418
rect 188988 21354 189040 21360
rect 187700 3800 187752 3806
rect 187700 3742 187752 3748
rect 189000 3534 189028 21354
rect 189184 6798 189212 326266
rect 189172 6792 189224 6798
rect 189172 6734 189224 6740
rect 189276 5234 189304 338014
rect 189368 338014 189750 338042
rect 189368 326330 189396 338014
rect 190288 336734 190316 338028
rect 190472 338014 190762 338042
rect 190932 338014 191314 338042
rect 191866 338014 192064 338042
rect 190276 336728 190328 336734
rect 190276 336670 190328 336676
rect 189356 326324 189408 326330
rect 189356 326266 189408 326272
rect 190472 5302 190500 338014
rect 190932 316034 190960 338014
rect 191840 336728 191892 336734
rect 191840 336670 191892 336676
rect 191104 336116 191156 336122
rect 191104 336058 191156 336064
rect 190564 316006 190960 316034
rect 190564 7614 190592 316006
rect 191116 11762 191144 336058
rect 191104 11756 191156 11762
rect 191104 11698 191156 11704
rect 190552 7608 190604 7614
rect 190552 7550 190604 7556
rect 190828 6316 190880 6322
rect 190828 6258 190880 6264
rect 190460 5296 190512 5302
rect 190460 5238 190512 5244
rect 189264 5228 189316 5234
rect 189264 5170 189316 5176
rect 189724 4820 189776 4826
rect 189724 4762 189776 4768
rect 188528 3528 188580 3534
rect 188528 3470 188580 3476
rect 188988 3528 189040 3534
rect 188988 3470 189040 3476
rect 188540 480 188568 3470
rect 189736 480 189764 4762
rect 190840 480 190868 6258
rect 191852 5370 191880 336670
rect 192036 323610 192064 338014
rect 192128 338014 192418 338042
rect 192496 338014 192878 338042
rect 192128 336734 192156 338014
rect 192116 336728 192168 336734
rect 192116 336670 192168 336676
rect 192024 323604 192076 323610
rect 192024 323546 192076 323552
rect 192496 321554 192524 338014
rect 193416 331226 193444 338028
rect 193508 338014 193982 338042
rect 194152 338014 194534 338042
rect 194704 338014 194994 338042
rect 195256 338014 195546 338042
rect 193404 331220 193456 331226
rect 193404 331162 193456 331168
rect 193508 326618 193536 338014
rect 193588 331220 193640 331226
rect 193588 331162 193640 331168
rect 191944 321526 192524 321554
rect 193232 326590 193536 326618
rect 191944 7682 191972 321526
rect 193128 11756 193180 11762
rect 193128 11698 193180 11704
rect 191932 7676 191984 7682
rect 191932 7618 191984 7624
rect 191840 5364 191892 5370
rect 191840 5306 191892 5312
rect 193140 3534 193168 11698
rect 193232 5438 193260 326590
rect 193312 326324 193364 326330
rect 193312 326266 193364 326272
rect 193324 7750 193352 326266
rect 193600 316034 193628 331162
rect 194152 326330 194180 338014
rect 194140 326324 194192 326330
rect 194140 326266 194192 326272
rect 194600 326324 194652 326330
rect 194600 326266 194652 326272
rect 193416 316006 193628 316034
rect 193416 302938 193444 316006
rect 193404 302932 193456 302938
rect 193404 302874 193456 302880
rect 193312 7744 193364 7750
rect 193312 7686 193364 7692
rect 194416 6384 194468 6390
rect 194416 6326 194468 6332
rect 193220 5432 193272 5438
rect 193220 5374 193272 5380
rect 193220 4888 193272 4894
rect 193220 4830 193272 4836
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 193128 3528 193180 3534
rect 193128 3470 193180 3476
rect 192036 480 192064 3470
rect 193232 480 193260 4830
rect 194428 480 194456 6326
rect 194612 5506 194640 326266
rect 194704 298790 194732 338014
rect 195256 326330 195284 338014
rect 195888 331968 195940 331974
rect 195888 331910 195940 331916
rect 195244 326324 195296 326330
rect 195244 326266 195296 326272
rect 194692 298784 194744 298790
rect 194692 298726 194744 298732
rect 195900 6914 195928 331910
rect 195980 329588 196032 329594
rect 195980 329530 196032 329536
rect 195624 6886 195928 6914
rect 194600 5500 194652 5506
rect 194600 5442 194652 5448
rect 195624 480 195652 6886
rect 195992 4758 196020 329530
rect 196084 7818 196112 338028
rect 196176 338014 196558 338042
rect 196728 338014 197110 338042
rect 197464 338014 197662 338042
rect 197740 338014 198214 338042
rect 198384 338014 198674 338042
rect 198844 338014 199226 338042
rect 199488 338014 199778 338042
rect 196176 297430 196204 338014
rect 196728 329594 196756 338014
rect 197360 330540 197412 330546
rect 197360 330482 197412 330488
rect 196716 329588 196768 329594
rect 196716 329530 196768 329536
rect 196164 297424 196216 297430
rect 196164 297366 196216 297372
rect 196072 7812 196124 7818
rect 196072 7754 196124 7760
rect 196808 4956 196860 4962
rect 196808 4898 196860 4904
rect 195980 4752 196032 4758
rect 195980 4694 196032 4700
rect 196820 480 196848 4898
rect 197372 4622 197400 330482
rect 197464 8974 197492 338014
rect 197740 316034 197768 338014
rect 198384 330546 198412 338014
rect 198372 330540 198424 330546
rect 198372 330482 198424 330488
rect 198740 328092 198792 328098
rect 198740 328034 198792 328040
rect 197556 316006 197768 316034
rect 197556 294642 197584 316006
rect 197544 294636 197596 294642
rect 197544 294578 197596 294584
rect 197452 8968 197504 8974
rect 197452 8910 197504 8916
rect 197912 6452 197964 6458
rect 197912 6394 197964 6400
rect 197360 4616 197412 4622
rect 197360 4558 197412 4564
rect 197924 480 197952 6394
rect 198752 3874 198780 328034
rect 198844 9042 198872 338014
rect 199488 328098 199516 338014
rect 200120 330540 200172 330546
rect 200120 330482 200172 330488
rect 199476 328092 199528 328098
rect 199476 328034 199528 328040
rect 200028 24132 200080 24138
rect 200028 24074 200080 24080
rect 198832 9036 198884 9042
rect 198832 8978 198884 8984
rect 198740 3868 198792 3874
rect 198740 3810 198792 3816
rect 200040 3534 200068 24074
rect 200132 3942 200160 330482
rect 200224 4690 200252 338028
rect 200316 338014 200790 338042
rect 200960 338014 201342 338042
rect 201512 338014 201894 338042
rect 201972 338014 202354 338042
rect 202906 338014 203104 338042
rect 200316 9110 200344 338014
rect 200960 330546 200988 338014
rect 200948 330540 201000 330546
rect 200948 330482 201000 330488
rect 200304 9104 200356 9110
rect 200304 9046 200356 9052
rect 200304 5024 200356 5030
rect 200304 4966 200356 4972
rect 200212 4684 200264 4690
rect 200212 4626 200264 4632
rect 200120 3936 200172 3942
rect 200120 3878 200172 3884
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 199120 480 199148 3470
rect 200316 480 200344 4966
rect 201512 4554 201540 338014
rect 201972 316034 202000 338014
rect 202788 334620 202840 334626
rect 202788 334562 202840 334568
rect 201604 316006 202000 316034
rect 201604 9178 201632 316006
rect 201592 9172 201644 9178
rect 201592 9114 201644 9120
rect 202800 6914 202828 334562
rect 202972 330540 203024 330546
rect 202972 330482 203024 330488
rect 202708 6886 202828 6914
rect 201592 6520 201644 6526
rect 201592 6462 201644 6468
rect 201500 4548 201552 4554
rect 201500 4490 201552 4496
rect 201604 3244 201632 6462
rect 201512 3216 201632 3244
rect 201512 480 201540 3216
rect 202708 480 202736 6886
rect 202984 4486 203012 330482
rect 202972 4480 203024 4486
rect 202972 4422 203024 4428
rect 203076 4010 203104 338014
rect 203168 338014 203458 338042
rect 203168 330546 203196 338014
rect 203996 336530 204024 338028
rect 204272 338014 204470 338042
rect 204548 338014 205022 338042
rect 205192 338014 205574 338042
rect 205652 338014 206034 338042
rect 206204 338014 206586 338042
rect 207138 338014 207244 338042
rect 203984 336524 204036 336530
rect 203984 336466 204036 336472
rect 203156 330540 203208 330546
rect 203156 330482 203208 330488
rect 203892 5092 203944 5098
rect 203892 5034 203944 5040
rect 203064 4004 203116 4010
rect 203064 3946 203116 3952
rect 203904 480 203932 5034
rect 204272 4078 204300 338014
rect 204548 335354 204576 338014
rect 204364 335326 204576 335354
rect 204364 6866 204392 335326
rect 205192 316034 205220 338014
rect 204456 316006 205220 316034
rect 204456 17270 204484 316006
rect 204444 17264 204496 17270
rect 204444 17206 204496 17212
rect 204352 6860 204404 6866
rect 204352 6802 204404 6808
rect 205088 6588 205140 6594
rect 205088 6530 205140 6536
rect 204260 4072 204312 4078
rect 204260 4014 204312 4020
rect 205100 480 205128 6530
rect 205652 4146 205680 338014
rect 206204 316034 206232 338014
rect 206928 333396 206980 333402
rect 206928 333338 206980 333344
rect 205744 316006 206232 316034
rect 205744 7886 205772 316006
rect 205732 7880 205784 7886
rect 205732 7822 205784 7828
rect 205640 4140 205692 4146
rect 205640 4082 205692 4088
rect 206940 3466 206968 333338
rect 207112 326392 207164 326398
rect 207112 326334 207164 326340
rect 207124 7954 207152 326334
rect 207216 326330 207244 338014
rect 207308 338014 207690 338042
rect 207768 338014 208150 338042
rect 208596 338014 208702 338042
rect 208780 338014 209254 338042
rect 209424 338014 209714 338042
rect 207204 326324 207256 326330
rect 207204 326266 207256 326272
rect 207112 7948 207164 7954
rect 207112 7890 207164 7896
rect 206192 3460 206244 3466
rect 206192 3402 206244 3408
rect 206928 3460 206980 3466
rect 206928 3402 206980 3408
rect 206204 480 206232 3402
rect 207308 3398 207336 338014
rect 207768 326398 207796 338014
rect 207756 326392 207808 326398
rect 207756 326334 207808 326340
rect 208492 326392 208544 326398
rect 208492 326334 208544 326340
rect 208504 8022 208532 326334
rect 208596 28286 208624 338014
rect 208780 316034 208808 338014
rect 209424 326398 209452 338014
rect 210252 333198 210280 338028
rect 210344 338014 210818 338042
rect 211264 338014 211370 338042
rect 210240 333192 210292 333198
rect 210240 333134 210292 333140
rect 209412 326392 209464 326398
rect 209412 326334 209464 326340
rect 210344 316034 210372 338014
rect 210516 335708 210568 335714
rect 210516 335650 210568 335656
rect 210528 316034 210556 335650
rect 208688 316006 208808 316034
rect 209976 316006 210372 316034
rect 210436 316006 210556 316034
rect 208584 28280 208636 28286
rect 208584 28222 208636 28228
rect 208492 8016 208544 8022
rect 208492 7958 208544 7964
rect 207388 5160 207440 5166
rect 207388 5102 207440 5108
rect 207296 3392 207348 3398
rect 207296 3334 207348 3340
rect 207400 480 207428 5102
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 208596 480 208624 3470
rect 208688 3330 208716 316006
rect 209688 31068 209740 31074
rect 209688 31010 209740 31016
rect 209700 3534 209728 31010
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 209780 3460 209832 3466
rect 209780 3402 209832 3408
rect 208676 3324 208728 3330
rect 208676 3266 208728 3272
rect 209792 480 209820 3402
rect 209976 3262 210004 316006
rect 210436 311166 210464 316006
rect 210424 311160 210476 311166
rect 210424 311102 210476 311108
rect 211264 8090 211292 338014
rect 211816 335714 211844 338028
rect 211908 338014 212382 338042
rect 212552 338014 212934 338042
rect 213012 338014 213394 338042
rect 213946 338014 214236 338042
rect 211804 335708 211856 335714
rect 211804 335650 211856 335656
rect 211908 316034 211936 338014
rect 212448 336048 212500 336054
rect 212448 335990 212500 335996
rect 211356 316006 211936 316034
rect 211252 8084 211304 8090
rect 211252 8026 211304 8032
rect 210976 5228 211028 5234
rect 210976 5170 211028 5176
rect 209964 3256 210016 3262
rect 209964 3198 210016 3204
rect 210988 480 211016 5170
rect 211356 3194 211384 316006
rect 212460 6914 212488 335990
rect 212552 8158 212580 338014
rect 213012 316034 213040 338014
rect 213828 336184 213880 336190
rect 213828 336126 213880 336132
rect 212644 316006 213040 316034
rect 212644 18630 212672 316006
rect 212632 18624 212684 18630
rect 212632 18566 212684 18572
rect 212540 8152 212592 8158
rect 212540 8094 212592 8100
rect 212184 6886 212488 6914
rect 211344 3188 211396 3194
rect 211344 3130 211396 3136
rect 212184 480 212212 6886
rect 213840 3534 213868 336126
rect 214208 331226 214236 338014
rect 214300 338014 214498 338042
rect 214760 338014 215050 338042
rect 214196 331220 214248 331226
rect 214196 331162 214248 331168
rect 214300 326618 214328 338014
rect 214380 331220 214432 331226
rect 214380 331162 214432 331168
rect 214024 326590 214328 326618
rect 214024 8226 214052 326590
rect 214104 326392 214156 326398
rect 214104 326334 214156 326340
rect 214116 307086 214144 326334
rect 214392 316034 214420 331162
rect 214760 326398 214788 338014
rect 215496 328454 215524 338028
rect 215404 328426 215524 328454
rect 215588 338014 216062 338042
rect 216232 338014 216614 338042
rect 216876 338014 217166 338042
rect 217336 338014 217626 338042
rect 214748 326392 214800 326398
rect 214748 326334 214800 326340
rect 215404 323626 215432 328426
rect 215404 323598 215524 323626
rect 215392 321360 215444 321366
rect 215392 321302 215444 321308
rect 214208 316006 214420 316034
rect 214104 307080 214156 307086
rect 214104 307022 214156 307028
rect 214012 8220 214064 8226
rect 214012 8162 214064 8168
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 213380 480 213408 3470
rect 214208 3126 214236 316006
rect 215404 8294 215432 321302
rect 215392 8288 215444 8294
rect 215392 8230 215444 8236
rect 214472 5296 214524 5302
rect 214472 5238 214524 5244
rect 214196 3120 214248 3126
rect 214196 3062 214248 3068
rect 214484 480 214512 5238
rect 215496 3058 215524 323598
rect 215588 321366 215616 338014
rect 216232 336122 216260 338014
rect 216220 336116 216272 336122
rect 216220 336058 216272 336064
rect 216588 336116 216640 336122
rect 216588 336058 216640 336064
rect 215576 321360 215628 321366
rect 215576 321302 215628 321308
rect 216600 3534 216628 336058
rect 216772 326392 216824 326398
rect 216772 326334 216824 326340
rect 216784 7546 216812 326334
rect 216772 7540 216824 7546
rect 216772 7482 216824 7488
rect 216876 6914 216904 338014
rect 217336 326398 217364 338014
rect 217968 336320 218020 336326
rect 217968 336262 218020 336268
rect 217324 326392 217376 326398
rect 217324 326334 217376 326340
rect 216784 6886 216904 6914
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 216588 3528 216640 3534
rect 216588 3470 216640 3476
rect 215484 3052 215536 3058
rect 215484 2994 215536 3000
rect 215680 480 215708 3470
rect 216784 2990 216812 6886
rect 217980 3534 218008 336262
rect 218164 318102 218192 338028
rect 218716 336394 218744 338028
rect 218808 338014 219190 338042
rect 219544 338014 219742 338042
rect 219820 338014 220294 338042
rect 220846 338014 220952 338042
rect 218704 336388 218756 336394
rect 218704 336330 218756 336336
rect 218152 318096 218204 318102
rect 218152 318038 218204 318044
rect 218808 316034 218836 338014
rect 219256 336252 219308 336258
rect 219256 336194 219308 336200
rect 218256 316006 218836 316034
rect 218256 7478 218284 316006
rect 218244 7472 218296 7478
rect 218244 7414 218296 7420
rect 218060 5364 218112 5370
rect 218060 5306 218112 5312
rect 216864 3528 216916 3534
rect 216864 3470 216916 3476
rect 217968 3528 218020 3534
rect 217968 3470 218020 3476
rect 216772 2984 216824 2990
rect 216772 2926 216824 2932
rect 216876 480 216904 3470
rect 218072 480 218100 5306
rect 219268 480 219296 336194
rect 219544 256018 219572 338014
rect 219820 316034 219848 338014
rect 220728 336388 220780 336394
rect 220728 336330 220780 336336
rect 219636 316006 219848 316034
rect 219532 256012 219584 256018
rect 219532 255954 219584 255960
rect 219636 2922 219664 316006
rect 220740 6914 220768 336330
rect 220924 7410 220952 338014
rect 221292 329118 221320 338028
rect 221476 338014 221858 338042
rect 221280 329112 221332 329118
rect 221280 329054 221332 329060
rect 221476 316034 221504 338014
rect 222292 326392 222344 326398
rect 222292 326334 222344 326340
rect 221108 316006 221504 316034
rect 220912 7404 220964 7410
rect 220912 7346 220964 7352
rect 220464 6886 220768 6914
rect 219624 2916 219676 2922
rect 219624 2858 219676 2864
rect 220464 480 220492 6886
rect 221108 2854 221136 316006
rect 222304 308446 222332 326334
rect 222292 308440 222344 308446
rect 222292 308382 222344 308388
rect 222396 7342 222424 338028
rect 222488 338014 222870 338042
rect 222488 326398 222516 338014
rect 223408 336462 223436 338028
rect 223396 336456 223448 336462
rect 223396 336398 223448 336404
rect 223488 336456 223540 336462
rect 223488 336398 223540 336404
rect 222476 326392 222528 326398
rect 222476 326334 222528 326340
rect 222384 7336 222436 7342
rect 222384 7278 222436 7284
rect 221556 5432 221608 5438
rect 221556 5374 221608 5380
rect 221096 2848 221148 2854
rect 221096 2790 221148 2796
rect 221568 480 221596 5374
rect 223500 3534 223528 336398
rect 223960 334694 223988 338028
rect 224052 338014 224526 338042
rect 223948 334688 224000 334694
rect 223948 334630 224000 334636
rect 224052 316034 224080 338014
rect 224868 336592 224920 336598
rect 224868 336534 224920 336540
rect 223684 316006 224080 316034
rect 223684 14482 223712 316006
rect 223672 14476 223724 14482
rect 223672 14418 223724 14424
rect 222752 3528 222804 3534
rect 222752 3470 222804 3476
rect 223488 3528 223540 3534
rect 223488 3470 223540 3476
rect 222764 480 222792 3470
rect 224880 2990 224908 336534
rect 224972 6118 225000 338028
rect 225524 329186 225552 338028
rect 225708 338014 226090 338042
rect 226352 338014 226550 338042
rect 226628 338014 227102 338042
rect 227272 338014 227654 338042
rect 227732 338014 228206 338042
rect 228284 338014 228666 338042
rect 225512 329180 225564 329186
rect 225512 329122 225564 329128
rect 225708 327826 225736 338014
rect 225696 327820 225748 327826
rect 225696 327762 225748 327768
rect 226352 13122 226380 338014
rect 226628 325038 226656 338014
rect 226616 325032 226668 325038
rect 226616 324974 226668 324980
rect 227272 321554 227300 338014
rect 227628 336524 227680 336530
rect 227628 336466 227680 336472
rect 226444 321526 227300 321554
rect 226444 268394 226472 321526
rect 226432 268388 226484 268394
rect 226432 268330 226484 268336
rect 226340 13116 226392 13122
rect 226340 13058 226392 13064
rect 224960 6112 225012 6118
rect 224960 6054 225012 6060
rect 225144 5500 225196 5506
rect 225144 5442 225196 5448
rect 223948 2984 224000 2990
rect 223948 2926 224000 2932
rect 224868 2984 224920 2990
rect 224868 2926 224920 2932
rect 223960 480 223988 2926
rect 225156 480 225184 5442
rect 227536 3596 227588 3602
rect 227536 3538 227588 3544
rect 226340 3528 226392 3534
rect 226340 3470 226392 3476
rect 226352 480 226380 3470
rect 227548 480 227576 3538
rect 227640 3534 227668 336466
rect 227732 35222 227760 338014
rect 228284 323678 228312 338014
rect 228272 323672 228324 323678
rect 228272 323614 228324 323620
rect 229204 316742 229232 338028
rect 229388 338014 229770 338042
rect 229192 316736 229244 316742
rect 229192 316678 229244 316684
rect 229388 316034 229416 338014
rect 230308 331906 230336 338028
rect 230584 338014 230782 338042
rect 230952 338014 231334 338042
rect 231886 338014 232084 338042
rect 230388 335980 230440 335986
rect 230388 335922 230440 335928
rect 230296 331900 230348 331906
rect 230296 331842 230348 331848
rect 229296 316006 229416 316034
rect 227720 35216 227772 35222
rect 227720 35158 227772 35164
rect 229296 25566 229324 316006
rect 229284 25560 229336 25566
rect 229284 25502 229336 25508
rect 228732 8968 228784 8974
rect 228732 8910 228784 8916
rect 227628 3528 227680 3534
rect 227628 3470 227680 3476
rect 228744 480 228772 8910
rect 230400 3602 230428 335922
rect 230480 326392 230532 326398
rect 230480 326334 230532 326340
rect 230492 312594 230520 326334
rect 230584 313954 230612 338014
rect 230952 326398 230980 338014
rect 231768 336660 231820 336666
rect 231768 336602 231820 336608
rect 230940 326392 230992 326398
rect 230940 326334 230992 326340
rect 230572 313948 230624 313954
rect 230572 313890 230624 313896
rect 230480 312588 230532 312594
rect 230480 312530 230532 312536
rect 231780 3602 231808 336602
rect 232056 331226 232084 338014
rect 232148 338014 232346 338042
rect 232608 338014 232898 338042
rect 232044 331220 232096 331226
rect 232044 331162 232096 331168
rect 232148 326618 232176 338014
rect 232228 331220 232280 331226
rect 232228 331162 232280 331168
rect 231872 326590 232176 326618
rect 231872 6050 231900 326590
rect 231952 326392 232004 326398
rect 231952 326334 232004 326340
rect 231964 26926 231992 326334
rect 232240 320890 232268 331162
rect 232608 326398 232636 338014
rect 232596 326392 232648 326398
rect 232596 326334 232648 326340
rect 233436 322250 233464 338028
rect 233712 338014 234002 338042
rect 234080 338014 234462 338042
rect 234632 338014 235014 338042
rect 235092 338014 235566 338042
rect 236026 338014 236224 338042
rect 233712 331214 233740 338014
rect 233528 331186 233740 331214
rect 233424 322244 233476 322250
rect 233424 322186 233476 322192
rect 233528 322130 233556 331186
rect 233252 322102 233556 322130
rect 232228 320884 232280 320890
rect 232228 320826 232280 320832
rect 231952 26920 232004 26926
rect 231952 26862 232004 26868
rect 233148 14476 233200 14482
rect 233148 14418 233200 14424
rect 231860 6044 231912 6050
rect 231860 5986 231912 5992
rect 233160 3602 233188 14418
rect 233252 5982 233280 322102
rect 234080 321554 234108 338014
rect 233344 321526 234108 321554
rect 233344 7206 233372 321526
rect 233332 7200 233384 7206
rect 233332 7142 233384 7148
rect 233240 5976 233292 5982
rect 233240 5918 233292 5924
rect 234632 4418 234660 338014
rect 235092 316034 235120 338014
rect 236000 336728 236052 336734
rect 236000 336670 236052 336676
rect 235908 329112 235960 329118
rect 235908 329054 235960 329060
rect 234724 316006 235120 316034
rect 234724 5914 234752 316006
rect 235920 6914 235948 329054
rect 235828 6886 235948 6914
rect 234712 5908 234764 5914
rect 234712 5850 234764 5856
rect 234620 4412 234672 4418
rect 234620 4354 234672 4360
rect 229836 3596 229888 3602
rect 229836 3538 229888 3544
rect 230388 3596 230440 3602
rect 230388 3538 230440 3544
rect 231032 3596 231084 3602
rect 231032 3538 231084 3544
rect 231768 3596 231820 3602
rect 231768 3538 231820 3544
rect 232228 3596 232280 3602
rect 232228 3538 232280 3544
rect 233148 3596 233200 3602
rect 233148 3538 233200 3544
rect 233424 3596 233476 3602
rect 233424 3538 233476 3544
rect 229848 480 229876 3538
rect 231044 480 231072 3538
rect 232240 480 232268 3538
rect 233436 480 233464 3538
rect 234618 3360 234674 3369
rect 234618 3295 234674 3304
rect 234632 480 234660 3295
rect 235828 480 235856 6886
rect 236012 4350 236040 336670
rect 236092 324420 236144 324426
rect 236092 324362 236144 324368
rect 236104 5846 236132 324362
rect 236196 7274 236224 338014
rect 236288 338014 236578 338042
rect 236840 338014 237130 338042
rect 237484 338014 237682 338042
rect 237760 338014 238142 338042
rect 238312 338014 238694 338042
rect 238772 338014 239246 338042
rect 236288 336734 236316 338014
rect 236276 336728 236328 336734
rect 236276 336670 236328 336676
rect 236840 324426 236868 338014
rect 237380 326392 237432 326398
rect 237380 326334 237432 326340
rect 237484 326346 237512 338014
rect 237760 335354 237788 338014
rect 237668 335326 237788 335354
rect 237668 326398 237696 335326
rect 237656 326392 237708 326398
rect 236828 324420 236880 324426
rect 236828 324362 236880 324368
rect 236184 7268 236236 7274
rect 236184 7210 236236 7216
rect 236092 5840 236144 5846
rect 236092 5782 236144 5788
rect 236000 4344 236052 4350
rect 236000 4286 236052 4292
rect 237392 4282 237420 326334
rect 237484 326318 237604 326346
rect 237656 326334 237708 326340
rect 237472 326256 237524 326262
rect 237472 326198 237524 326204
rect 237484 5778 237512 326198
rect 237576 7138 237604 326318
rect 238312 326262 238340 338014
rect 238300 326256 238352 326262
rect 238300 326198 238352 326204
rect 237564 7132 237616 7138
rect 237564 7074 237616 7080
rect 238772 7070 238800 338014
rect 239784 333198 239812 338028
rect 239772 333192 239824 333198
rect 239772 333134 239824 333140
rect 240244 315314 240272 338028
rect 240428 338014 240810 338042
rect 240428 316034 240456 338014
rect 240784 335912 240836 335918
rect 240784 335854 240836 335860
rect 240336 316006 240456 316034
rect 240232 315308 240284 315314
rect 240232 315250 240284 315256
rect 239312 7608 239364 7614
rect 239312 7550 239364 7556
rect 238760 7064 238812 7070
rect 238760 7006 238812 7012
rect 237472 5772 237524 5778
rect 237472 5714 237524 5720
rect 237380 4276 237432 4282
rect 237380 4218 237432 4224
rect 238116 3664 238168 3670
rect 238116 3606 238168 3612
rect 237010 3496 237066 3505
rect 237010 3431 237066 3440
rect 237024 480 237052 3431
rect 238128 480 238156 3606
rect 239324 480 239352 7550
rect 240336 5710 240364 316006
rect 240796 15910 240824 335854
rect 241348 330614 241376 338028
rect 241624 338014 241822 338042
rect 241992 338014 242374 338042
rect 242926 338014 243032 338042
rect 241336 330608 241388 330614
rect 241336 330550 241388 330556
rect 241520 326392 241572 326398
rect 241520 326334 241572 326340
rect 240784 15904 240836 15910
rect 240784 15846 240836 15852
rect 240324 5704 240376 5710
rect 240324 5646 240376 5652
rect 241532 5642 241560 326334
rect 241624 174554 241652 338014
rect 241992 326398 242020 338014
rect 242808 335980 242860 335986
rect 242808 335922 242860 335928
rect 241980 326392 242032 326398
rect 241980 326334 242032 326340
rect 241612 174548 241664 174554
rect 241612 174490 241664 174496
rect 241520 5636 241572 5642
rect 241520 5578 241572 5584
rect 240508 3732 240560 3738
rect 240508 3674 240560 3680
rect 240520 480 240548 3674
rect 242820 3398 242848 335922
rect 243004 326466 243032 338014
rect 243464 335918 243492 338028
rect 243556 338014 243938 338042
rect 244384 338014 244490 338042
rect 244660 338014 245042 338042
rect 245120 338014 245502 338042
rect 245764 338014 246054 338042
rect 246224 338014 246606 338042
rect 243452 335912 243504 335918
rect 243452 335854 243504 335860
rect 242992 326460 243044 326466
rect 242992 326402 243044 326408
rect 243556 316034 243584 338014
rect 244280 326392 244332 326398
rect 244280 326334 244332 326340
rect 243096 316006 243584 316034
rect 243096 6186 243124 316006
rect 244292 6254 244320 326334
rect 244384 10334 244412 338014
rect 244660 316034 244688 338014
rect 245120 326398 245148 338014
rect 245764 327758 245792 338014
rect 245752 327752 245804 327758
rect 245752 327694 245804 327700
rect 245108 326392 245160 326398
rect 245108 326334 245160 326340
rect 246224 316034 246252 338014
rect 247144 326466 247172 338028
rect 247236 338014 247618 338042
rect 247788 338014 248170 338042
rect 248616 338014 248722 338042
rect 248800 338014 249182 338042
rect 249352 338014 249734 338042
rect 249812 338014 250286 338042
rect 250364 338014 250838 338042
rect 247132 326460 247184 326466
rect 247132 326402 247184 326408
rect 247132 326256 247184 326262
rect 247132 326198 247184 326204
rect 247040 321700 247092 321706
rect 247040 321642 247092 321648
rect 244476 316006 244688 316034
rect 245672 316006 246252 316034
rect 244476 286346 244504 316006
rect 245672 290494 245700 316006
rect 245660 290488 245712 290494
rect 245660 290430 245712 290436
rect 244464 286340 244516 286346
rect 244464 286282 244516 286288
rect 247052 11830 247080 321642
rect 247144 22778 247172 326198
rect 247236 321706 247264 338014
rect 247224 321700 247276 321706
rect 247224 321642 247276 321648
rect 247788 318170 247816 338014
rect 248616 326874 248644 338014
rect 248800 335354 248828 338014
rect 248708 335326 248828 335354
rect 248604 326868 248656 326874
rect 248604 326810 248656 326816
rect 248604 326664 248656 326670
rect 248604 326606 248656 326612
rect 248512 326392 248564 326398
rect 248512 326334 248564 326340
rect 248420 323604 248472 323610
rect 248420 323546 248472 323552
rect 247776 318164 247828 318170
rect 247776 318106 247828 318112
rect 247132 22772 247184 22778
rect 247132 22714 247184 22720
rect 248432 13190 248460 323546
rect 248524 17338 248552 326334
rect 248616 19990 248644 326606
rect 248708 323610 248736 335326
rect 249352 326398 249380 338014
rect 249340 326392 249392 326398
rect 249340 326334 249392 326340
rect 248696 323604 248748 323610
rect 248696 323546 248748 323552
rect 248604 19984 248656 19990
rect 248604 19926 248656 19932
rect 248512 17332 248564 17338
rect 248512 17274 248564 17280
rect 248420 13184 248472 13190
rect 248420 13126 248472 13132
rect 247040 11824 247092 11830
rect 247040 11766 247092 11772
rect 244372 10328 244424 10334
rect 244372 10270 244424 10276
rect 249812 9246 249840 338014
rect 250364 316034 250392 338014
rect 251088 335912 251140 335918
rect 251088 335854 251140 335860
rect 249904 316006 250392 316034
rect 249904 10402 249932 316006
rect 249892 10396 249944 10402
rect 249892 10338 249944 10344
rect 249800 9240 249852 9246
rect 249800 9182 249852 9188
rect 244280 6248 244332 6254
rect 244280 6190 244332 6196
rect 243084 6180 243136 6186
rect 243084 6122 243136 6128
rect 248788 4072 248840 4078
rect 248788 4014 248840 4020
rect 247592 4004 247644 4010
rect 247592 3946 247644 3952
rect 246396 3936 246448 3942
rect 246396 3878 246448 3884
rect 245200 3868 245252 3874
rect 245200 3810 245252 3816
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 241704 3392 241756 3398
rect 241704 3334 241756 3340
rect 242808 3392 242860 3398
rect 242808 3334 242860 3340
rect 241716 480 241744 3334
rect 242912 480 242940 3742
rect 244094 3632 244150 3641
rect 244094 3567 244150 3576
rect 244108 480 244136 3567
rect 245212 480 245240 3810
rect 246408 480 246436 3878
rect 247604 480 247632 3946
rect 248800 480 248828 4014
rect 251100 3398 251128 335854
rect 251180 323468 251232 323474
rect 251180 323410 251232 323416
rect 251192 4826 251220 323410
rect 251284 18698 251312 338028
rect 251468 338014 251850 338042
rect 252112 338014 252402 338042
rect 252572 338014 252954 338042
rect 253032 338014 253414 338042
rect 253966 338014 254164 338042
rect 251468 316034 251496 338014
rect 252112 323474 252140 338014
rect 252100 323468 252152 323474
rect 252100 323410 252152 323416
rect 251376 316006 251496 316034
rect 251376 21418 251404 316006
rect 251364 21412 251416 21418
rect 251364 21354 251416 21360
rect 251272 18692 251324 18698
rect 251272 18634 251324 18640
rect 252572 6322 252600 338014
rect 253032 316034 253060 338014
rect 253848 335844 253900 335850
rect 253848 335786 253900 335792
rect 252664 316006 253060 316034
rect 252664 11762 252692 316006
rect 252652 11756 252704 11762
rect 252652 11698 252704 11704
rect 253860 6914 253888 335786
rect 254136 328454 254164 338014
rect 254044 328426 254164 328454
rect 254228 338014 254518 338042
rect 254044 322402 254072 328426
rect 254044 322374 254164 322402
rect 254032 319524 254084 319530
rect 254032 319466 254084 319472
rect 253492 6886 253888 6914
rect 252560 6316 252612 6322
rect 252560 6258 252612 6264
rect 251180 4820 251232 4826
rect 251180 4762 251232 4768
rect 252376 4140 252428 4146
rect 252376 4082 252428 4088
rect 249984 3392 250036 3398
rect 249984 3334 250036 3340
rect 251088 3392 251140 3398
rect 251088 3334 251140 3340
rect 251180 3392 251232 3398
rect 251180 3334 251232 3340
rect 249996 480 250024 3334
rect 251192 480 251220 3334
rect 252388 480 252416 4082
rect 253492 480 253520 6886
rect 254044 6390 254072 319466
rect 254032 6384 254084 6390
rect 254032 6326 254084 6332
rect 254136 4894 254164 322374
rect 254228 319530 254256 338014
rect 254964 331974 254992 338028
rect 255332 338014 255530 338042
rect 255608 338014 256082 338042
rect 256344 338014 256634 338042
rect 256712 338014 257094 338042
rect 257172 338014 257646 338042
rect 254952 331968 255004 331974
rect 254952 331910 255004 331916
rect 254216 319524 254268 319530
rect 254216 319466 254268 319472
rect 255332 4962 255360 338014
rect 255608 335354 255636 338014
rect 255424 335326 255636 335354
rect 255424 6458 255452 335326
rect 256344 316034 256372 338014
rect 255516 316006 256372 316034
rect 255516 24138 255544 316006
rect 255504 24132 255556 24138
rect 255504 24074 255556 24080
rect 255412 6452 255464 6458
rect 255412 6394 255464 6400
rect 256712 5030 256740 338014
rect 257172 316034 257200 338014
rect 258184 334626 258212 338028
rect 258276 338014 258658 338042
rect 258920 338014 259210 338042
rect 258172 334620 258224 334626
rect 258172 334562 258224 334568
rect 258172 326392 258224 326398
rect 258172 326334 258224 326340
rect 256804 316006 257200 316034
rect 256804 6526 256832 316006
rect 258184 6594 258212 326334
rect 258172 6588 258224 6594
rect 258172 6530 258224 6536
rect 256792 6520 256844 6526
rect 256792 6462 256844 6468
rect 258276 5098 258304 338014
rect 258920 326398 258948 338014
rect 259368 335776 259420 335782
rect 259368 335718 259420 335724
rect 258908 326392 258960 326398
rect 258908 326334 258960 326340
rect 258264 5092 258316 5098
rect 258264 5034 258316 5040
rect 256700 5024 256752 5030
rect 256700 4966 256752 4972
rect 255320 4956 255372 4962
rect 255320 4898 255372 4904
rect 254124 4888 254176 4894
rect 254124 4830 254176 4836
rect 259380 3534 259408 335718
rect 259748 333402 259776 338028
rect 259932 338014 260314 338042
rect 260392 338014 260774 338042
rect 260852 338014 261326 338042
rect 261404 338014 261878 338042
rect 259736 333396 259788 333402
rect 259736 333338 259788 333344
rect 259552 326392 259604 326398
rect 259552 326334 259604 326340
rect 259564 31074 259592 326334
rect 259932 316034 259960 338014
rect 260392 326398 260420 338014
rect 260748 335640 260800 335646
rect 260748 335582 260800 335588
rect 260380 326392 260432 326398
rect 260380 326334 260432 326340
rect 259656 316006 259960 316034
rect 259552 31068 259604 31074
rect 259552 31010 259604 31016
rect 259656 5166 259684 316006
rect 260760 6914 260788 335582
rect 260668 6886 260788 6914
rect 259644 5160 259696 5166
rect 259644 5102 259696 5108
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 254676 3324 254728 3330
rect 254676 3266 254728 3272
rect 254688 480 254716 3266
rect 255872 3256 255924 3262
rect 255872 3198 255924 3204
rect 255884 480 255912 3198
rect 257068 3188 257120 3194
rect 257068 3130 257120 3136
rect 257080 480 257108 3130
rect 258276 480 258304 3470
rect 259460 3120 259512 3126
rect 259460 3062 259512 3068
rect 259472 480 259500 3062
rect 260668 480 260696 6886
rect 260852 3466 260880 338014
rect 261404 316034 261432 338014
rect 262324 336054 262352 338028
rect 262876 336190 262904 338028
rect 263060 338014 263442 338042
rect 262864 336184 262916 336190
rect 262864 336126 262916 336132
rect 262312 336048 262364 336054
rect 262312 335990 262364 335996
rect 263060 316034 263088 338014
rect 263980 336122 264008 338028
rect 264440 336326 264468 338028
rect 265006 338014 265112 338042
rect 264428 336320 264480 336326
rect 264428 336262 264480 336268
rect 263968 336116 264020 336122
rect 263968 336058 264020 336064
rect 264888 336048 264940 336054
rect 264888 335990 264940 335996
rect 260944 316006 261432 316034
rect 262324 316006 263088 316034
rect 260944 5234 260972 316006
rect 262324 5302 262352 316006
rect 262312 5296 262364 5302
rect 262312 5238 262364 5244
rect 260932 5228 260984 5234
rect 260932 5170 260984 5176
rect 264900 3534 264928 335990
rect 265084 5370 265112 338014
rect 265544 336258 265572 338028
rect 266096 336394 266124 338028
rect 266464 338014 266570 338042
rect 266084 336388 266136 336394
rect 266084 336330 266136 336336
rect 265532 336252 265584 336258
rect 265532 336194 265584 336200
rect 266464 5438 266492 338014
rect 267108 336462 267136 338028
rect 267660 336598 267688 338028
rect 267844 338014 268134 338042
rect 267648 336592 267700 336598
rect 267648 336534 267700 336540
rect 267096 336456 267148 336462
rect 267096 336398 267148 336404
rect 267844 5506 267872 338014
rect 268672 336530 268700 338028
rect 269238 338014 269344 338042
rect 268660 336524 268712 336530
rect 268660 336466 268712 336472
rect 269028 336116 269080 336122
rect 269028 336058 269080 336064
rect 267832 5500 267884 5506
rect 267832 5442 267884 5448
rect 266452 5432 266504 5438
rect 266452 5374 266504 5380
rect 265072 5364 265124 5370
rect 265072 5306 265124 5312
rect 269040 3534 269068 336058
rect 269212 330540 269264 330546
rect 269212 330482 269264 330488
rect 269224 8974 269252 330482
rect 269212 8968 269264 8974
rect 269212 8910 269264 8916
rect 269316 6914 269344 338014
rect 269408 338014 269790 338042
rect 269408 330546 269436 338014
rect 270236 336666 270264 338028
rect 270512 338014 270802 338042
rect 271064 338014 271354 338042
rect 271432 338014 271814 338042
rect 271892 338014 272366 338042
rect 270512 336734 270540 338014
rect 270500 336728 270552 336734
rect 270500 336670 270552 336676
rect 270684 336728 270736 336734
rect 270684 336670 270736 336676
rect 270224 336660 270276 336666
rect 270224 336602 270276 336608
rect 269396 330540 269448 330546
rect 269396 330482 269448 330488
rect 270592 330540 270644 330546
rect 270592 330482 270644 330488
rect 270604 14482 270632 330482
rect 270592 14476 270644 14482
rect 270592 14418 270644 14424
rect 269132 6886 269344 6914
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 267740 3528 267792 3534
rect 267740 3470 267792 3476
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 260840 3460 260892 3466
rect 260840 3402 260892 3408
rect 261760 3460 261812 3466
rect 261760 3402 261812 3408
rect 261772 480 261800 3402
rect 262956 3052 263008 3058
rect 262956 2994 263008 3000
rect 262968 480 262996 2994
rect 264164 480 264192 3470
rect 265348 2984 265400 2990
rect 265348 2926 265400 2932
rect 265360 480 265388 2926
rect 266544 2848 266596 2854
rect 266544 2790 266596 2796
rect 266556 480 266584 2790
rect 267752 480 267780 3470
rect 269132 3074 269160 6886
rect 270040 3800 270092 3806
rect 270040 3742 270092 3748
rect 268764 3046 269160 3074
rect 268764 2922 268792 3046
rect 268752 2916 268804 2922
rect 268752 2858 268804 2864
rect 268844 2916 268896 2922
rect 268844 2858 268896 2864
rect 268856 480 268884 2858
rect 270052 480 270080 3742
rect 270696 3602 270724 336670
rect 271064 330546 271092 338014
rect 271432 336734 271460 338014
rect 271420 336728 271472 336734
rect 271420 336670 271472 336676
rect 271788 336184 271840 336190
rect 271788 336126 271840 336132
rect 271052 330540 271104 330546
rect 271052 330482 271104 330488
rect 270684 3596 270736 3602
rect 270684 3538 270736 3544
rect 271800 3534 271828 336126
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271788 3528 271840 3534
rect 271788 3470 271840 3476
rect 271248 480 271276 3470
rect 271892 3369 271920 338014
rect 272904 329118 272932 338028
rect 273272 338014 273470 338042
rect 273548 338014 273930 338042
rect 274008 338014 274482 338042
rect 274836 338014 275034 338042
rect 272892 329112 272944 329118
rect 272892 329054 272944 329060
rect 272708 3528 272760 3534
rect 273272 3505 273300 338014
rect 273548 336682 273576 338014
rect 273364 336654 273576 336682
rect 273364 3602 273392 336654
rect 274008 335354 274036 338014
rect 273456 335326 274036 335354
rect 273456 7614 273484 335326
rect 273444 7608 273496 7614
rect 273444 7550 273496 7556
rect 274836 3738 274864 338014
rect 275572 335986 275600 338028
rect 276046 338014 276244 338042
rect 275560 335980 275612 335986
rect 275560 335922 275612 335928
rect 276216 330818 276244 338014
rect 276308 338014 276598 338042
rect 276768 338014 277150 338042
rect 277504 338014 277610 338042
rect 277780 338014 278162 338042
rect 278424 338014 278714 338042
rect 276204 330812 276256 330818
rect 276204 330754 276256 330760
rect 276308 330698 276336 338014
rect 276032 330670 276336 330698
rect 276032 3777 276060 330670
rect 276204 330608 276256 330614
rect 276204 330550 276256 330556
rect 276112 330540 276164 330546
rect 276112 330482 276164 330488
rect 276124 3806 276152 330482
rect 276216 4010 276244 330550
rect 276768 330546 276796 338014
rect 277216 336320 277268 336326
rect 277216 336262 277268 336268
rect 276756 330540 276808 330546
rect 276756 330482 276808 330488
rect 277228 6914 277256 336262
rect 277308 336252 277360 336258
rect 277308 336194 277360 336200
rect 277136 6886 277256 6914
rect 276204 4004 276256 4010
rect 276204 3946 276256 3952
rect 276112 3800 276164 3806
rect 276018 3768 276074 3777
rect 274824 3732 274876 3738
rect 276112 3742 276164 3748
rect 277032 3800 277084 3806
rect 277032 3742 277084 3748
rect 276018 3703 276074 3712
rect 274824 3674 274876 3680
rect 273352 3596 273404 3602
rect 273352 3538 273404 3544
rect 275008 3596 275060 3602
rect 275008 3538 275060 3544
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 273628 3528 273680 3534
rect 272708 3470 272760 3476
rect 273258 3496 273314 3505
rect 271878 3360 271934 3369
rect 271878 3295 271934 3304
rect 272720 1850 272748 3470
rect 273628 3470 273680 3476
rect 273258 3431 273314 3440
rect 272444 1822 272748 1850
rect 272444 480 272472 1822
rect 273640 480 273668 3470
rect 275020 1986 275048 3538
rect 274836 1958 275048 1986
rect 274836 480 274864 1958
rect 276032 480 276060 3538
rect 277044 3482 277072 3742
rect 277136 3602 277164 6886
rect 277216 4072 277268 4078
rect 277216 4014 277268 4020
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 277044 3454 277164 3482
rect 277136 480 277164 3454
rect 277228 3380 277256 4014
rect 277320 3806 277348 336194
rect 277400 330540 277452 330546
rect 277400 330482 277452 330488
rect 277412 3942 277440 330482
rect 277400 3936 277452 3942
rect 277400 3878 277452 3884
rect 277308 3800 277360 3806
rect 277308 3742 277360 3748
rect 277504 3670 277532 338014
rect 277780 316034 277808 338014
rect 278044 336456 278096 336462
rect 278044 336398 278096 336404
rect 277596 316006 277808 316034
rect 277492 3664 277544 3670
rect 277492 3606 277544 3612
rect 277596 3398 277624 316006
rect 278056 4010 278084 336398
rect 278424 330546 278452 338014
rect 279252 335918 279280 338028
rect 279344 338014 279726 338042
rect 280278 338014 280384 338042
rect 279240 335912 279292 335918
rect 279240 335854 279292 335860
rect 278412 330540 278464 330546
rect 278412 330482 278464 330488
rect 279344 316034 279372 338014
rect 280252 330540 280304 330546
rect 280252 330482 280304 330488
rect 278976 316006 279372 316034
rect 278044 4004 278096 4010
rect 278044 3946 278096 3952
rect 278976 3874 279004 316006
rect 278964 3868 279016 3874
rect 278964 3810 279016 3816
rect 279516 3732 279568 3738
rect 279516 3674 279568 3680
rect 277308 3392 277360 3398
rect 277228 3352 277308 3380
rect 277308 3334 277360 3340
rect 277584 3392 277636 3398
rect 277584 3334 277636 3340
rect 278320 3188 278372 3194
rect 278320 3130 278372 3136
rect 278332 480 278360 3130
rect 279528 480 279556 3674
rect 280264 3670 280292 330482
rect 280356 4146 280384 338014
rect 280816 335850 280844 338028
rect 281000 338014 281290 338042
rect 281736 338014 281842 338042
rect 282104 338014 282394 338042
rect 280896 336524 280948 336530
rect 280896 336466 280948 336472
rect 280804 335844 280856 335850
rect 280804 335786 280856 335792
rect 280908 316034 280936 336466
rect 281000 330546 281028 338014
rect 281448 336388 281500 336394
rect 281448 336330 281500 336336
rect 280988 330540 281040 330546
rect 280988 330482 281040 330488
rect 280816 316006 280936 316034
rect 280344 4140 280396 4146
rect 280344 4082 280396 4088
rect 280252 3664 280304 3670
rect 280252 3606 280304 3612
rect 280712 3460 280764 3466
rect 280712 3402 280764 3408
rect 280724 480 280752 3402
rect 280816 3194 280844 316006
rect 281460 3466 281488 336330
rect 281632 330540 281684 330546
rect 281632 330482 281684 330488
rect 281448 3460 281500 3466
rect 281448 3402 281500 3408
rect 281644 3262 281672 330482
rect 281736 3942 281764 338014
rect 282104 330546 282132 338014
rect 282828 336592 282880 336598
rect 282828 336534 282880 336540
rect 282092 330540 282144 330546
rect 282092 330482 282144 330488
rect 281724 3936 281776 3942
rect 281724 3878 281776 3884
rect 282840 3466 282868 336534
rect 282932 335782 282960 338028
rect 283116 338014 283406 338042
rect 282920 335776 282972 335782
rect 282920 335718 282972 335724
rect 283116 6914 283144 338014
rect 283944 335646 283972 338028
rect 284510 338014 284616 338042
rect 283932 335640 283984 335646
rect 283932 335582 283984 335588
rect 283564 335368 283616 335374
rect 283564 335310 283616 335316
rect 283024 6886 283144 6914
rect 281908 3460 281960 3466
rect 281908 3402 281960 3408
rect 282828 3460 282880 3466
rect 282828 3402 282880 3408
rect 281632 3256 281684 3262
rect 281632 3198 281684 3204
rect 280804 3188 280856 3194
rect 280804 3130 280856 3136
rect 281920 480 281948 3402
rect 283024 3126 283052 6886
rect 283576 3874 283604 335310
rect 284484 330540 284536 330546
rect 284484 330482 284536 330488
rect 283564 3868 283616 3874
rect 283564 3810 283616 3816
rect 283104 3800 283156 3806
rect 283104 3742 283156 3748
rect 283012 3120 283064 3126
rect 283012 3062 283064 3068
rect 283116 480 283144 3742
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 284312 480 284340 3606
rect 284496 3058 284524 330482
rect 284588 3330 284616 338014
rect 284680 338014 284970 338042
rect 285232 338014 285522 338042
rect 285784 338014 286074 338042
rect 286244 338014 286626 338042
rect 284680 330546 284708 338014
rect 285232 336054 285260 338014
rect 285588 336660 285640 336666
rect 285588 336602 285640 336608
rect 285220 336048 285272 336054
rect 285220 335990 285272 335996
rect 285496 336048 285548 336054
rect 285496 335990 285548 335996
rect 284668 330540 284720 330546
rect 284668 330482 284720 330488
rect 285508 3670 285536 335990
rect 285496 3664 285548 3670
rect 285496 3606 285548 3612
rect 285600 3516 285628 336602
rect 285416 3488 285628 3516
rect 284576 3324 284628 3330
rect 284576 3266 284628 3272
rect 284484 3052 284536 3058
rect 284484 2994 284536 3000
rect 285416 480 285444 3488
rect 285784 2990 285812 338014
rect 286244 316034 286272 338014
rect 286968 336728 287020 336734
rect 286968 336670 287020 336676
rect 285876 316006 286272 316034
rect 285772 2984 285824 2990
rect 285772 2926 285824 2932
rect 285876 2854 285904 316006
rect 286980 6914 287008 336670
rect 287072 336122 287100 338028
rect 287164 338014 287638 338042
rect 287716 338014 288190 338042
rect 287060 336116 287112 336122
rect 287060 336058 287112 336064
rect 286612 6886 287008 6914
rect 285864 2848 285916 2854
rect 285864 2790 285916 2796
rect 286612 480 286640 6886
rect 287164 2922 287192 338014
rect 287716 316034 287744 338014
rect 288728 336190 288756 338028
rect 288716 336184 288768 336190
rect 288716 336126 288768 336132
rect 289188 335374 289216 338028
rect 289372 338014 289754 338042
rect 289176 335368 289228 335374
rect 289176 335310 289228 335316
rect 289372 316034 289400 338014
rect 290292 336462 290320 338028
rect 290280 336456 290332 336462
rect 290280 336398 290332 336404
rect 290752 336326 290780 338028
rect 290740 336320 290792 336326
rect 290740 336262 290792 336268
rect 291304 336258 291332 338028
rect 291488 338014 291870 338042
rect 291948 338014 292422 338042
rect 291488 336530 291516 338014
rect 291948 336682 291976 338014
rect 291764 336654 291976 336682
rect 291476 336524 291528 336530
rect 291476 336466 291528 336472
rect 291292 336252 291344 336258
rect 291292 336194 291344 336200
rect 289728 336116 289780 336122
rect 289728 336058 289780 336064
rect 287348 316006 287744 316034
rect 288544 316006 289400 316034
rect 287348 3534 287376 316006
rect 288544 3602 288572 316006
rect 288532 3596 288584 3602
rect 288532 3538 288584 3544
rect 289740 3534 289768 336058
rect 291764 316034 291792 336654
rect 292868 336394 292896 338028
rect 293420 336598 293448 338028
rect 293986 338014 294092 338042
rect 293408 336592 293460 336598
rect 293408 336534 293460 336540
rect 292856 336388 292908 336394
rect 292856 336330 292908 336336
rect 292488 336184 292540 336190
rect 292488 336126 292540 336132
rect 291844 335640 291896 335646
rect 291844 335582 291896 335588
rect 291304 316006 291792 316034
rect 291304 3670 291332 316006
rect 291292 3664 291344 3670
rect 291292 3606 291344 3612
rect 287336 3528 287388 3534
rect 287336 3470 287388 3476
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 287796 3392 287848 3398
rect 287796 3334 287848 3340
rect 287152 2916 287204 2922
rect 287152 2858 287204 2864
rect 287808 480 287836 3334
rect 289004 480 289032 3470
rect 290188 3460 290240 3466
rect 290188 3402 290240 3408
rect 290200 480 290228 3402
rect 291396 480 291424 3470
rect 291856 3466 291884 335582
rect 292500 3534 292528 336126
rect 294064 3806 294092 338014
rect 294432 336054 294460 338028
rect 294984 336666 295012 338028
rect 295536 336734 295564 338028
rect 295628 338014 296102 338042
rect 295524 336728 295576 336734
rect 295524 336670 295576 336676
rect 294972 336660 295024 336666
rect 294972 336602 295024 336608
rect 294604 336388 294656 336394
rect 294604 336330 294656 336336
rect 294420 336048 294472 336054
rect 294420 335990 294472 335996
rect 294052 3800 294104 3806
rect 294052 3742 294104 3748
rect 294616 3534 294644 336330
rect 295628 316034 295656 338014
rect 296548 336122 296576 338028
rect 296536 336116 296588 336122
rect 296536 336058 296588 336064
rect 296628 336116 296680 336122
rect 296628 336058 296680 336064
rect 295444 316006 295656 316034
rect 294880 4072 294932 4078
rect 294880 4014 294932 4020
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 293684 3528 293736 3534
rect 293684 3470 293736 3476
rect 294604 3528 294656 3534
rect 294604 3470 294656 3476
rect 291844 3460 291896 3466
rect 291844 3402 291896 3408
rect 292580 3052 292632 3058
rect 292580 2994 292632 3000
rect 292592 480 292620 2994
rect 293696 480 293724 3470
rect 294892 480 294920 4014
rect 295444 3398 295472 316006
rect 296640 3534 296668 336058
rect 297100 335646 297128 338028
rect 297652 336190 297680 338028
rect 297640 336184 297692 336190
rect 297640 336126 297692 336132
rect 297088 335640 297140 335646
rect 297088 335582 297140 335588
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 296628 3528 296680 3534
rect 296628 3470 296680 3476
rect 295432 3392 295484 3398
rect 295432 3334 295484 3340
rect 296088 480 296116 3470
rect 297272 3188 297324 3194
rect 297272 3130 297324 3136
rect 297284 480 297312 3130
rect 298204 3058 298232 338028
rect 298664 336394 298692 338028
rect 298756 338014 299230 338042
rect 298652 336388 298704 336394
rect 298652 336330 298704 336336
rect 298756 316034 298784 338014
rect 299768 336122 299796 338028
rect 299860 338014 300242 338042
rect 299756 336116 299808 336122
rect 299756 336058 299808 336064
rect 299388 335640 299440 335646
rect 299388 335582 299440 335588
rect 298296 316006 298784 316034
rect 298296 4078 298324 316006
rect 298284 4072 298336 4078
rect 298284 4014 298336 4020
rect 299400 3534 299428 335582
rect 299860 316034 299888 338014
rect 300780 335646 300808 338028
rect 300964 338014 301346 338042
rect 301608 338014 301898 338042
rect 302252 338014 302358 338042
rect 302436 338014 302910 338042
rect 303462 338014 303568 338042
rect 300768 335640 300820 335646
rect 300768 335582 300820 335588
rect 300860 330540 300912 330546
rect 300860 330482 300912 330488
rect 299768 316006 299888 316034
rect 298468 3528 298520 3534
rect 298468 3470 298520 3476
rect 299388 3528 299440 3534
rect 299388 3470 299440 3476
rect 298192 3052 298244 3058
rect 298192 2994 298244 3000
rect 298480 480 298508 3470
rect 299664 3256 299716 3262
rect 299664 3198 299716 3204
rect 299676 480 299704 3198
rect 299768 3194 299796 316006
rect 300872 3482 300900 330482
rect 300780 3454 300900 3482
rect 299756 3188 299808 3194
rect 299756 3130 299808 3136
rect 300780 480 300808 3454
rect 300964 3262 300992 338014
rect 301608 330546 301636 338014
rect 301596 330540 301648 330546
rect 301596 330482 301648 330488
rect 302252 3482 302280 338014
rect 302436 316034 302464 338014
rect 303540 335354 303568 338014
rect 303908 336734 303936 338028
rect 303896 336728 303948 336734
rect 303896 336670 303948 336676
rect 304460 335714 304488 338028
rect 304908 336728 304960 336734
rect 304908 336670 304960 336676
rect 304448 335708 304500 335714
rect 304448 335650 304500 335656
rect 303540 335326 303844 335354
rect 302344 316006 302464 316034
rect 302344 3534 302372 316006
rect 303816 16574 303844 335326
rect 303816 16546 304396 16574
rect 301976 3454 302280 3482
rect 302332 3528 302384 3534
rect 302332 3470 302384 3476
rect 303160 3528 303212 3534
rect 303160 3470 303212 3476
rect 300952 3256 301004 3262
rect 300952 3198 301004 3204
rect 301976 480 302004 3454
rect 303172 480 303200 3470
rect 304368 480 304396 16546
rect 304920 3534 304948 336670
rect 305012 336190 305040 338028
rect 305578 338014 305960 338042
rect 305932 336274 305960 338014
rect 306024 336394 306052 338028
rect 306576 336734 306604 338028
rect 306564 336728 306616 336734
rect 306564 336670 306616 336676
rect 306012 336388 306064 336394
rect 306012 336330 306064 336336
rect 305932 336246 306328 336274
rect 305000 336184 305052 336190
rect 305000 336126 305052 336132
rect 306196 336184 306248 336190
rect 306196 336126 306248 336132
rect 306208 3602 306236 336126
rect 306300 4146 306328 336246
rect 306656 335708 306708 335714
rect 306656 335650 306708 335656
rect 306668 16574 306696 335650
rect 307128 335510 307156 338028
rect 307588 336258 307616 338028
rect 307668 336728 307720 336734
rect 307668 336670 307720 336676
rect 307576 336252 307628 336258
rect 307576 336194 307628 336200
rect 307116 335504 307168 335510
rect 307116 335446 307168 335452
rect 306668 16546 306788 16574
rect 306288 4140 306340 4146
rect 306288 4082 306340 4088
rect 306196 3596 306248 3602
rect 306196 3538 306248 3544
rect 304908 3528 304960 3534
rect 304908 3470 304960 3476
rect 305552 3528 305604 3534
rect 305552 3470 305604 3476
rect 305564 480 305592 3470
rect 306760 480 306788 16546
rect 307680 3262 307708 336670
rect 308140 336666 308168 338028
rect 308692 336734 308720 338028
rect 308680 336728 308732 336734
rect 308680 336670 308732 336676
rect 308128 336660 308180 336666
rect 308128 336602 308180 336608
rect 309244 335578 309272 338028
rect 309324 336388 309376 336394
rect 309324 336330 309376 336336
rect 309232 335572 309284 335578
rect 309232 335514 309284 335520
rect 309336 16574 309364 336330
rect 309704 335986 309732 338028
rect 309784 336728 309836 336734
rect 309784 336670 309836 336676
rect 309692 335980 309744 335986
rect 309692 335922 309744 335928
rect 309336 16546 309732 16574
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 307944 3596 307996 3602
rect 307944 3538 307996 3544
rect 307668 3256 307720 3262
rect 307668 3198 307720 3204
rect 307956 480 307984 3538
rect 309060 480 309088 4082
rect 309704 3584 309732 16546
rect 309796 4146 309824 336670
rect 310256 336394 310284 338028
rect 310808 336598 310836 338028
rect 311164 336660 311216 336666
rect 311164 336602 311216 336608
rect 310796 336592 310848 336598
rect 310796 336534 310848 336540
rect 310244 336388 310296 336394
rect 310244 336330 310296 336336
rect 310428 335572 310480 335578
rect 310428 335514 310480 335520
rect 309784 4140 309836 4146
rect 309784 4082 309836 4088
rect 310336 4140 310388 4146
rect 310336 4082 310388 4088
rect 309704 3556 310284 3584
rect 310256 480 310284 3556
rect 310348 3058 310376 4082
rect 310440 3398 310468 335514
rect 310428 3392 310480 3398
rect 310428 3334 310480 3340
rect 311176 3330 311204 336602
rect 311360 336326 311388 338028
rect 311820 336530 311848 338028
rect 312372 336666 312400 338028
rect 312924 336734 312952 338028
rect 312912 336728 312964 336734
rect 312912 336670 312964 336676
rect 312360 336660 312412 336666
rect 312360 336602 312412 336608
rect 313188 336660 313240 336666
rect 313188 336602 313240 336608
rect 311808 336524 311860 336530
rect 311808 336466 311860 336472
rect 311348 336320 311400 336326
rect 311348 336262 311400 336268
rect 312084 335504 312136 335510
rect 312084 335446 312136 335452
rect 312096 16574 312124 335446
rect 312096 16546 312676 16574
rect 311164 3324 311216 3330
rect 311164 3266 311216 3272
rect 311440 3256 311492 3262
rect 311440 3198 311492 3204
rect 310336 3052 310388 3058
rect 310336 2994 310388 3000
rect 311452 480 311480 3198
rect 312648 480 312676 16546
rect 313200 3534 313228 336602
rect 313384 336462 313412 338028
rect 313950 338014 314424 338042
rect 313372 336456 313424 336462
rect 313372 336398 313424 336404
rect 313924 336388 313976 336394
rect 313924 336330 313976 336336
rect 313372 336252 313424 336258
rect 313372 336194 313424 336200
rect 313384 16574 313412 336194
rect 313384 16546 313872 16574
rect 313188 3528 313240 3534
rect 313188 3470 313240 3476
rect 313844 480 313872 16546
rect 313936 3670 313964 336330
rect 314396 335354 314424 338014
rect 314488 336258 314516 338028
rect 314476 336252 314528 336258
rect 314476 336194 314528 336200
rect 315040 336122 315068 338028
rect 315514 338014 315988 338042
rect 315028 336116 315080 336122
rect 315028 336058 315080 336064
rect 314396 335326 314608 335354
rect 313924 3664 313976 3670
rect 313924 3606 313976 3612
rect 314580 3466 314608 335326
rect 315960 6254 315988 338014
rect 316052 336598 316080 338028
rect 316604 336734 316632 338028
rect 317078 338014 317184 338042
rect 316592 336728 316644 336734
rect 316592 336670 316644 336676
rect 316040 336592 316092 336598
rect 316040 336534 316092 336540
rect 317156 7682 317184 338014
rect 317328 336728 317380 336734
rect 317328 336670 317380 336676
rect 317236 336592 317288 336598
rect 317236 336534 317288 336540
rect 317144 7676 317196 7682
rect 317144 7618 317196 7624
rect 315948 6248 316000 6254
rect 315948 6190 316000 6196
rect 317248 4078 317276 336534
rect 317236 4072 317288 4078
rect 317236 4014 317288 4020
rect 317340 4010 317368 336670
rect 317616 336598 317644 338028
rect 318182 338014 318656 338042
rect 317604 336592 317656 336598
rect 317604 336534 317656 336540
rect 318064 336456 318116 336462
rect 318064 336398 318116 336404
rect 317512 335980 317564 335986
rect 317512 335922 317564 335928
rect 317524 16574 317552 335922
rect 317524 16546 318012 16574
rect 317328 4004 317380 4010
rect 317328 3946 317380 3952
rect 317984 3482 318012 16546
rect 318076 3942 318104 336398
rect 318628 4146 318656 338014
rect 318720 336734 318748 338028
rect 318708 336728 318760 336734
rect 318708 336670 318760 336676
rect 318708 336592 318760 336598
rect 318708 336534 318760 336540
rect 318616 4140 318668 4146
rect 318616 4082 318668 4088
rect 318064 3936 318116 3942
rect 318064 3878 318116 3884
rect 318720 3806 318748 336534
rect 319180 336462 319208 338028
rect 319444 336728 319496 336734
rect 319444 336670 319496 336676
rect 319168 336456 319220 336462
rect 319168 336398 319220 336404
rect 319456 10402 319484 336670
rect 319732 336190 319760 338028
rect 320284 336734 320312 338028
rect 320758 338014 321048 338042
rect 321310 338014 321508 338042
rect 320272 336728 320324 336734
rect 320272 336670 320324 336676
rect 320456 336660 320508 336666
rect 320456 336602 320508 336608
rect 320088 336456 320140 336462
rect 320088 336398 320140 336404
rect 319720 336184 319772 336190
rect 319720 336126 319772 336132
rect 320100 14482 320128 336398
rect 320468 16574 320496 336602
rect 321020 335354 321048 338014
rect 321376 336728 321428 336734
rect 321376 336670 321428 336676
rect 321020 335326 321324 335354
rect 320468 16546 320956 16574
rect 320088 14476 320140 14482
rect 320088 14418 320140 14424
rect 319444 10396 319496 10402
rect 319444 10338 319496 10344
rect 318708 3800 318760 3806
rect 318708 3742 318760 3748
rect 319720 3664 319772 3670
rect 319720 3606 319772 3612
rect 314568 3460 314620 3466
rect 317984 3454 318564 3482
rect 314568 3402 314620 3408
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 315028 3324 315080 3330
rect 315028 3266 315080 3272
rect 315040 480 315068 3266
rect 316224 3052 316276 3058
rect 316224 2994 316276 3000
rect 316236 480 316264 2994
rect 317340 480 317368 3334
rect 318536 480 318564 3454
rect 319732 480 319760 3606
rect 320928 480 320956 16546
rect 321296 13122 321324 335326
rect 321284 13116 321336 13122
rect 321284 13058 321336 13064
rect 321388 9042 321416 336670
rect 321376 9036 321428 9042
rect 321376 8978 321428 8984
rect 321480 3738 321508 338014
rect 321848 336734 321876 338028
rect 322414 338014 322796 338042
rect 321836 336728 321888 336734
rect 321836 336670 321888 336676
rect 322664 336728 322716 336734
rect 322664 336670 322716 336676
rect 321836 336320 321888 336326
rect 321836 336262 321888 336268
rect 321848 16574 321876 336262
rect 321848 16546 322152 16574
rect 321468 3732 321520 3738
rect 321468 3674 321520 3680
rect 322124 480 322152 16546
rect 322676 11830 322704 336670
rect 322664 11824 322716 11830
rect 322664 11766 322716 11772
rect 322768 6186 322796 338014
rect 322756 6180 322808 6186
rect 322756 6122 322808 6128
rect 322860 3874 322888 338028
rect 323426 338014 323900 338042
rect 323978 338014 324268 338042
rect 323124 336524 323176 336530
rect 323124 336466 323176 336472
rect 323136 16574 323164 336466
rect 323872 335354 323900 338014
rect 323872 335326 324176 335354
rect 323136 16546 323348 16574
rect 322848 3868 322900 3874
rect 322848 3810 322900 3816
rect 323320 480 323348 16546
rect 324148 15910 324176 335326
rect 324136 15904 324188 15910
rect 324136 15846 324188 15852
rect 324240 7614 324268 338014
rect 324412 336388 324464 336394
rect 324412 336330 324464 336336
rect 324424 335354 324452 336330
rect 324516 335986 324544 338028
rect 324504 335980 324556 335986
rect 324504 335922 324556 335928
rect 324424 335326 324544 335354
rect 324516 16574 324544 335326
rect 324976 334626 325004 338028
rect 325424 335980 325476 335986
rect 325424 335922 325476 335928
rect 324964 334620 325016 334626
rect 324964 334562 325016 334568
rect 324516 16546 325372 16574
rect 324228 7608 324280 7614
rect 324228 7550 324280 7556
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 325344 3482 325372 16546
rect 325436 3602 325464 335922
rect 325528 8974 325556 338028
rect 326080 336734 326108 338028
rect 326068 336728 326120 336734
rect 326068 336670 326120 336676
rect 326540 336054 326568 338028
rect 327092 336734 327120 338028
rect 327658 338014 328132 338042
rect 326988 336728 327040 336734
rect 326988 336670 327040 336676
rect 327080 336728 327132 336734
rect 327080 336670 327132 336676
rect 326528 336048 326580 336054
rect 326528 335990 326580 335996
rect 325516 8968 325568 8974
rect 325516 8910 325568 8916
rect 325516 4072 325568 4078
rect 325516 4014 325568 4020
rect 325528 3890 325556 4014
rect 326804 3936 326856 3942
rect 325528 3874 325648 3890
rect 326804 3878 326856 3884
rect 325528 3868 325660 3874
rect 325528 3862 325608 3868
rect 325608 3810 325660 3816
rect 325424 3596 325476 3602
rect 325424 3538 325476 3544
rect 324424 480 324452 3470
rect 325344 3454 325648 3482
rect 325620 480 325648 3454
rect 326816 480 326844 3878
rect 327000 3058 327028 336670
rect 327724 336252 327776 336258
rect 327724 336194 327776 336200
rect 327736 3398 327764 336194
rect 328104 325694 328132 338014
rect 328196 333266 328224 338028
rect 328276 336728 328328 336734
rect 328276 336670 328328 336676
rect 328184 333260 328236 333266
rect 328184 333202 328236 333208
rect 328104 325666 328224 325694
rect 328196 3466 328224 325666
rect 328288 17270 328316 336670
rect 328656 336258 328684 338028
rect 329208 336598 329236 338028
rect 329668 338014 329774 338042
rect 329196 336592 329248 336598
rect 329196 336534 329248 336540
rect 328644 336252 328696 336258
rect 328644 336194 328696 336200
rect 328276 17264 328328 17270
rect 328276 17206 328328 17212
rect 329668 4350 329696 338014
rect 329748 336592 329800 336598
rect 329748 336534 329800 336540
rect 329656 4344 329708 4350
rect 329656 4286 329708 4292
rect 328000 3460 328052 3466
rect 328000 3402 328052 3408
rect 328184 3460 328236 3466
rect 328184 3402 328236 3408
rect 327724 3392 327776 3398
rect 327724 3334 327776 3340
rect 326988 3052 327040 3058
rect 326988 2994 327040 3000
rect 328012 480 328040 3402
rect 329196 3392 329248 3398
rect 329196 3334 329248 3340
rect 329208 480 329236 3334
rect 329760 3126 329788 336534
rect 330220 336326 330248 338028
rect 330786 338014 331168 338042
rect 330208 336320 330260 336326
rect 330208 336262 330260 336268
rect 330024 336116 330076 336122
rect 330024 336058 330076 336064
rect 330036 16574 330064 336058
rect 330036 16546 330432 16574
rect 329748 3120 329800 3126
rect 329748 3062 329800 3068
rect 330404 480 330432 16546
rect 331140 3194 331168 338014
rect 331324 335782 331352 338028
rect 331890 338014 332272 338042
rect 332350 338014 332548 338042
rect 331312 335776 331364 335782
rect 331312 335718 331364 335724
rect 332244 335354 332272 338014
rect 332416 335776 332468 335782
rect 332416 335718 332468 335724
rect 332244 335326 332364 335354
rect 332336 18698 332364 335326
rect 332324 18692 332376 18698
rect 332324 18634 332376 18640
rect 331588 6248 331640 6254
rect 331588 6190 331640 6196
rect 331128 3188 331180 3194
rect 331128 3130 331180 3136
rect 331600 480 331628 6190
rect 332428 4418 332456 335718
rect 332416 4412 332468 4418
rect 332416 4354 332468 4360
rect 332520 3262 332548 338014
rect 332888 336734 332916 338028
rect 333454 338014 333836 338042
rect 332876 336728 332928 336734
rect 332876 336670 332928 336676
rect 333808 326398 333836 338014
rect 333888 336728 333940 336734
rect 333888 336670 333940 336676
rect 333796 326392 333848 326398
rect 333796 326334 333848 326340
rect 333900 4486 333928 336670
rect 333992 336666 334020 338028
rect 334452 336734 334480 338028
rect 335018 338014 335124 338042
rect 334440 336728 334492 336734
rect 334440 336670 334492 336676
rect 333980 336660 334032 336666
rect 333980 336602 334032 336608
rect 335096 10334 335124 338014
rect 335556 336734 335584 338028
rect 335176 336728 335228 336734
rect 335176 336670 335228 336676
rect 335544 336728 335596 336734
rect 335544 336670 335596 336676
rect 335084 10328 335136 10334
rect 335084 10270 335136 10276
rect 335084 7676 335136 7682
rect 335084 7618 335136 7624
rect 333888 4480 333940 4486
rect 333888 4422 333940 4428
rect 333888 4004 333940 4010
rect 333888 3946 333940 3952
rect 332692 3868 332744 3874
rect 332692 3810 332744 3816
rect 332508 3256 332560 3262
rect 332508 3198 332560 3204
rect 332704 480 332732 3810
rect 333900 480 333928 3946
rect 335096 480 335124 7618
rect 335188 4554 335216 336670
rect 335268 336660 335320 336666
rect 335268 336602 335320 336608
rect 335176 4548 335228 4554
rect 335176 4490 335228 4496
rect 335280 3330 335308 336602
rect 336016 336598 336044 338028
rect 336476 338014 336582 338042
rect 336004 336592 336056 336598
rect 336004 336534 336056 336540
rect 336476 20058 336504 338014
rect 337120 336734 337148 338028
rect 337686 338014 337976 338042
rect 336648 336728 336700 336734
rect 336648 336670 336700 336676
rect 337108 336728 337160 336734
rect 337108 336670 337160 336676
rect 336556 336592 336608 336598
rect 336556 336534 336608 336540
rect 336464 20052 336516 20058
rect 336464 19994 336516 20000
rect 336568 4622 336596 336534
rect 336556 4616 336608 4622
rect 336556 4558 336608 4564
rect 336280 3800 336332 3806
rect 336280 3742 336332 3748
rect 335268 3324 335320 3330
rect 335268 3266 335320 3272
rect 336292 480 336320 3742
rect 336660 3398 336688 336670
rect 337948 4690 337976 338014
rect 338132 336734 338160 338028
rect 338028 336728 338080 336734
rect 338028 336670 338080 336676
rect 338120 336728 338172 336734
rect 338120 336670 338172 336676
rect 337936 4684 337988 4690
rect 337936 4626 337988 4632
rect 338040 4146 338068 336670
rect 338684 336666 338712 338028
rect 339250 338014 339356 338042
rect 339224 336728 339276 336734
rect 339224 336670 339276 336676
rect 338672 336660 338724 336666
rect 338672 336602 338724 336608
rect 339236 11762 339264 336670
rect 339224 11756 339276 11762
rect 339224 11698 339276 11704
rect 338672 10396 338724 10402
rect 338672 10338 338724 10344
rect 338028 4140 338080 4146
rect 338028 4082 338080 4088
rect 337476 3732 337528 3738
rect 337476 3674 337528 3680
rect 336648 3392 336700 3398
rect 336648 3334 336700 3340
rect 337488 480 337516 3674
rect 338684 480 338712 10338
rect 339328 4758 339356 338014
rect 339696 336734 339724 338028
rect 339684 336728 339736 336734
rect 339684 336670 339736 336676
rect 339408 336660 339460 336666
rect 339408 336602 339460 336608
rect 339316 4752 339368 4758
rect 339316 4694 339368 4700
rect 339420 4078 339448 336602
rect 340248 335714 340276 338028
rect 340708 338014 340814 338042
rect 340604 336728 340656 336734
rect 340604 336670 340656 336676
rect 340236 335708 340288 335714
rect 340236 335650 340288 335656
rect 340616 14482 340644 336670
rect 339868 14476 339920 14482
rect 339868 14418 339920 14424
rect 340604 14476 340656 14482
rect 340604 14418 340656 14424
rect 339408 4072 339460 4078
rect 339408 4014 339460 4020
rect 339880 480 339908 14418
rect 340708 5438 340736 338014
rect 341352 336734 341380 338028
rect 341826 338014 342208 338042
rect 341340 336728 341392 336734
rect 341340 336670 341392 336676
rect 342076 336728 342128 336734
rect 342076 336670 342128 336676
rect 341064 336184 341116 336190
rect 341064 336126 341116 336132
rect 340788 335708 340840 335714
rect 340788 335650 340840 335656
rect 340696 5432 340748 5438
rect 340696 5374 340748 5380
rect 340800 4010 340828 335650
rect 341076 6914 341104 336126
rect 342088 13190 342116 336670
rect 342076 13184 342128 13190
rect 342076 13126 342128 13132
rect 342180 11778 342208 338014
rect 342364 336734 342392 338028
rect 342930 338014 343312 338042
rect 343390 338014 343588 338042
rect 342352 336728 342404 336734
rect 342352 336670 342404 336676
rect 343284 335354 343312 338014
rect 343456 336728 343508 336734
rect 343456 336670 343508 336676
rect 343284 335326 343404 335354
rect 343376 25634 343404 335326
rect 343364 25628 343416 25634
rect 343364 25570 343416 25576
rect 343364 13116 343416 13122
rect 343364 13058 343416 13064
rect 340984 6886 341104 6914
rect 342088 11750 342208 11778
rect 340788 4004 340840 4010
rect 340788 3946 340840 3952
rect 340984 480 341012 6886
rect 342088 3942 342116 11750
rect 342168 9036 342220 9042
rect 342168 8978 342220 8984
rect 342076 3936 342128 3942
rect 342076 3878 342128 3884
rect 342180 480 342208 8978
rect 343376 480 343404 13058
rect 343468 5506 343496 336670
rect 343456 5500 343508 5506
rect 343456 5442 343508 5448
rect 343560 3874 343588 338014
rect 343928 336734 343956 338028
rect 343916 336728 343968 336734
rect 343916 336670 343968 336676
rect 344480 336190 344508 338028
rect 344928 336728 344980 336734
rect 344928 336670 344980 336676
rect 344468 336184 344520 336190
rect 344468 336126 344520 336132
rect 344940 5370 344968 336670
rect 345032 335918 345060 338028
rect 345492 336734 345520 338028
rect 346058 338014 346164 338042
rect 345480 336728 345532 336734
rect 345480 336670 345532 336676
rect 345020 335912 345072 335918
rect 345020 335854 345072 335860
rect 346136 29646 346164 338014
rect 346216 336728 346268 336734
rect 346216 336670 346268 336676
rect 346124 29640 346176 29646
rect 346124 29582 346176 29588
rect 345756 11824 345808 11830
rect 345756 11766 345808 11772
rect 344928 5364 344980 5370
rect 344928 5306 344980 5312
rect 343548 3868 343600 3874
rect 343548 3810 343600 3816
rect 344560 3664 344612 3670
rect 344560 3606 344612 3612
rect 344572 480 344600 3606
rect 345768 480 345796 11766
rect 346228 5302 346256 336670
rect 346308 335912 346360 335918
rect 346308 335854 346360 335860
rect 346216 5296 346268 5302
rect 346216 5238 346268 5244
rect 346320 3806 346348 335854
rect 346596 335578 346624 338028
rect 347148 336734 347176 338028
rect 347516 338014 347622 338042
rect 347136 336728 347188 336734
rect 347136 336670 347188 336676
rect 346584 335572 346636 335578
rect 346584 335514 346636 335520
rect 347516 324970 347544 338014
rect 348160 336734 348188 338028
rect 348726 338014 349016 338042
rect 347596 336728 347648 336734
rect 347596 336670 347648 336676
rect 348148 336728 348200 336734
rect 348148 336670 348200 336676
rect 347504 324964 347556 324970
rect 347504 324906 347556 324912
rect 346952 6180 347004 6186
rect 346952 6122 347004 6128
rect 346308 3800 346360 3806
rect 346308 3742 346360 3748
rect 346964 480 346992 6122
rect 347608 5234 347636 336670
rect 347688 335572 347740 335578
rect 347688 335514 347740 335520
rect 347596 5228 347648 5234
rect 347596 5170 347648 5176
rect 347700 3738 347728 335514
rect 348988 5166 349016 338014
rect 349068 336728 349120 336734
rect 349068 336670 349120 336676
rect 348976 5160 349028 5166
rect 348976 5102 349028 5108
rect 347688 3732 347740 3738
rect 347688 3674 347740 3680
rect 349080 3670 349108 336670
rect 349172 336122 349200 338028
rect 349724 336666 349752 338028
rect 350290 338014 350488 338042
rect 349712 336660 349764 336666
rect 349712 336602 349764 336608
rect 349804 336252 349856 336258
rect 349804 336194 349856 336200
rect 349160 336116 349212 336122
rect 349160 336058 349212 336064
rect 349816 15910 349844 336194
rect 350356 336116 350408 336122
rect 350356 336058 350408 336064
rect 349252 15904 349304 15910
rect 349252 15846 349304 15852
rect 349804 15904 349856 15910
rect 349804 15846 349856 15852
rect 349068 3664 349120 3670
rect 349068 3606 349120 3612
rect 348056 3596 348108 3602
rect 348056 3538 348108 3544
rect 348068 480 348096 3538
rect 349264 480 349292 15846
rect 350368 10402 350396 336058
rect 350356 10396 350408 10402
rect 350356 10338 350408 10344
rect 350356 7608 350408 7614
rect 350356 7550 350408 7556
rect 350368 3482 350396 7550
rect 350460 5098 350488 338014
rect 350828 330614 350856 338028
rect 351288 336598 351316 338028
rect 351748 338014 351854 338042
rect 351276 336592 351328 336598
rect 351276 336534 351328 336540
rect 350816 330608 350868 330614
rect 350816 330550 350868 330556
rect 350448 5092 350500 5098
rect 350448 5034 350500 5040
rect 351748 5030 351776 338014
rect 352392 336734 352420 338028
rect 352380 336728 352432 336734
rect 352380 336670 352432 336676
rect 352852 336666 352880 338028
rect 353404 336734 353432 338028
rect 353970 338014 354444 338042
rect 354522 338014 354628 338042
rect 353208 336728 353260 336734
rect 353208 336670 353260 336676
rect 353392 336728 353444 336734
rect 353392 336670 353444 336676
rect 352840 336660 352892 336666
rect 352840 336602 352892 336608
rect 351828 336592 351880 336598
rect 351828 336534 351880 336540
rect 351736 5024 351788 5030
rect 351736 4966 351788 4972
rect 351840 3602 351868 336534
rect 352564 336320 352616 336326
rect 352564 336262 352616 336268
rect 351920 334620 351972 334626
rect 351920 334562 351972 334568
rect 351932 16574 351960 334562
rect 351932 16546 352512 16574
rect 351828 3596 351880 3602
rect 351828 3538 351880 3544
rect 351644 3528 351696 3534
rect 350368 3454 350488 3482
rect 351644 3470 351696 3476
rect 352484 3482 352512 16546
rect 352576 6186 352604 336262
rect 353220 28286 353248 336670
rect 354416 31074 354444 338014
rect 354496 336728 354548 336734
rect 354496 336670 354548 336676
rect 354404 31068 354456 31074
rect 354404 31010 354456 31016
rect 353208 28280 353260 28286
rect 353208 28222 353260 28228
rect 354036 8968 354088 8974
rect 354036 8910 354088 8916
rect 352564 6180 352616 6186
rect 352564 6122 352616 6128
rect 350460 480 350488 3454
rect 351656 480 351684 3470
rect 352484 3454 352880 3482
rect 352852 480 352880 3454
rect 354048 480 354076 8910
rect 354508 4962 354536 336670
rect 354496 4956 354548 4962
rect 354496 4898 354548 4904
rect 354600 3534 354628 338014
rect 354968 336734 354996 338028
rect 355534 338014 355916 338042
rect 354956 336728 355008 336734
rect 354956 336670 355008 336676
rect 355888 323678 355916 338014
rect 355968 336728 356020 336734
rect 355968 336670 356020 336676
rect 355876 323672 355928 323678
rect 355876 323614 355928 323620
rect 355980 4894 356008 336670
rect 356072 336462 356100 338028
rect 356532 336734 356560 338028
rect 357098 338014 357296 338042
rect 356520 336728 356572 336734
rect 356520 336670 356572 336676
rect 356060 336456 356112 336462
rect 356060 336398 356112 336404
rect 356152 335980 356204 335986
rect 356152 335922 356204 335928
rect 356164 16574 356192 335922
rect 357268 19990 357296 338014
rect 357636 336734 357664 338028
rect 357348 336728 357400 336734
rect 357348 336670 357400 336676
rect 357624 336728 357676 336734
rect 357624 336670 357676 336676
rect 357256 19984 357308 19990
rect 357256 19926 357308 19932
rect 356164 16546 356376 16574
rect 355968 4888 356020 4894
rect 355968 4830 356020 4836
rect 354588 3528 354640 3534
rect 354588 3470 354640 3476
rect 355232 3052 355284 3058
rect 355232 2994 355284 3000
rect 355244 480 355272 2994
rect 356348 480 356376 16546
rect 357360 4826 357388 336670
rect 358084 336184 358136 336190
rect 358084 336126 358136 336132
rect 358096 26926 358124 336126
rect 358188 336054 358216 338028
rect 358176 336048 358228 336054
rect 358176 335990 358228 335996
rect 358084 26920 358136 26926
rect 358084 26862 358136 26868
rect 357532 17264 357584 17270
rect 357532 17206 357584 17212
rect 357348 4820 357400 4826
rect 357348 4762 357400 4768
rect 357544 480 357572 17206
rect 358648 7206 358676 338028
rect 359200 336734 359228 338028
rect 359766 338014 360056 338042
rect 358728 336728 358780 336734
rect 358728 336670 358780 336676
rect 359188 336728 359240 336734
rect 359188 336670 359240 336676
rect 358636 7200 358688 7206
rect 358636 7142 358688 7148
rect 358740 3618 358768 336670
rect 358820 333260 358872 333266
rect 358820 333202 358872 333208
rect 358832 16574 358860 333202
rect 360028 232558 360056 338014
rect 360108 336728 360160 336734
rect 360108 336670 360160 336676
rect 360016 232552 360068 232558
rect 360016 232494 360068 232500
rect 358832 16546 359964 16574
rect 358740 3590 358860 3618
rect 358832 3466 358860 3590
rect 358728 3460 358780 3466
rect 358728 3402 358780 3408
rect 358820 3460 358872 3466
rect 358820 3402 358872 3408
rect 358740 480 358768 3402
rect 359936 480 359964 16546
rect 360120 2854 360148 336670
rect 360304 335646 360332 338028
rect 360764 336734 360792 338028
rect 360752 336728 360804 336734
rect 360752 336670 360804 336676
rect 360292 335640 360344 335646
rect 360292 335582 360344 335588
rect 361316 15910 361344 338028
rect 361868 336734 361896 338028
rect 361488 336728 361540 336734
rect 361488 336670 361540 336676
rect 361856 336728 361908 336734
rect 361856 336670 361908 336676
rect 361396 335640 361448 335646
rect 361396 335582 361448 335588
rect 361120 15904 361172 15910
rect 361120 15846 361172 15852
rect 361304 15904 361356 15910
rect 361304 15846 361356 15852
rect 360108 2848 360160 2854
rect 360108 2790 360160 2796
rect 361132 480 361160 15846
rect 361408 7274 361436 335582
rect 361396 7268 361448 7274
rect 361396 7210 361448 7216
rect 361500 2922 361528 336670
rect 362328 336462 362356 338028
rect 362788 338014 362894 338042
rect 362316 336456 362368 336462
rect 362316 336398 362368 336404
rect 362788 329186 362816 338014
rect 363432 336734 363460 338028
rect 363998 338014 364288 338042
rect 362868 336728 362920 336734
rect 362868 336670 362920 336676
rect 363420 336728 363472 336734
rect 363420 336670 363472 336676
rect 364156 336728 364208 336734
rect 364156 336670 364208 336676
rect 362776 329180 362828 329186
rect 362776 329122 362828 329128
rect 362880 326466 362908 336670
rect 362868 326460 362920 326466
rect 362868 326402 362920 326408
rect 364168 44878 364196 336670
rect 364156 44872 364208 44878
rect 364156 44814 364208 44820
rect 363512 4344 363564 4350
rect 363512 4286 363564 4292
rect 362316 3120 362368 3126
rect 362316 3062 362368 3068
rect 361488 2916 361540 2922
rect 361488 2858 361540 2864
rect 362328 480 362356 3062
rect 363524 480 363552 4286
rect 364260 2990 364288 338014
rect 364444 336734 364472 338028
rect 365010 338014 365392 338042
rect 364432 336728 364484 336734
rect 364432 336670 364484 336676
rect 365364 335354 365392 338014
rect 365548 336258 365576 338028
rect 366008 336734 366036 338028
rect 366574 338014 366956 338042
rect 365628 336728 365680 336734
rect 365628 336670 365680 336676
rect 365996 336728 366048 336734
rect 365996 336670 366048 336676
rect 365536 336252 365588 336258
rect 365536 336194 365588 336200
rect 365364 335326 365576 335354
rect 365548 174554 365576 335326
rect 365536 174548 365588 174554
rect 365536 174490 365588 174496
rect 365640 17270 365668 336670
rect 366928 322250 366956 338014
rect 367112 336734 367140 338028
rect 367678 338014 368060 338042
rect 368138 338014 368336 338042
rect 367008 336728 367060 336734
rect 367008 336670 367060 336676
rect 367100 336728 367152 336734
rect 367100 336670 367152 336676
rect 366916 322244 366968 322250
rect 366916 322186 366968 322192
rect 367020 18630 367048 336670
rect 368032 327826 368060 338014
rect 368020 327820 368072 327826
rect 368020 327762 368072 327768
rect 368308 35222 368336 338014
rect 368388 336728 368440 336734
rect 368388 336670 368440 336676
rect 368296 35216 368348 35222
rect 368296 35158 368348 35164
rect 367100 18692 367152 18698
rect 367100 18634 367152 18640
rect 367008 18624 367060 18630
rect 367008 18566 367060 18572
rect 365628 17264 365680 17270
rect 365628 17206 365680 17212
rect 367112 16574 367140 18634
rect 367112 16546 368244 16574
rect 364616 6180 364668 6186
rect 364616 6122 364668 6128
rect 364248 2984 364300 2990
rect 364248 2926 364300 2932
rect 364628 480 364656 6122
rect 367008 4412 367060 4418
rect 367008 4354 367060 4360
rect 365812 3188 365864 3194
rect 365812 3130 365864 3136
rect 365824 480 365852 3130
rect 367020 480 367048 4354
rect 368216 480 368244 16546
rect 368400 3058 368428 336670
rect 368676 336190 368704 338028
rect 369228 336394 369256 338028
rect 369216 336388 369268 336394
rect 369216 336330 369268 336336
rect 368664 336184 368716 336190
rect 368664 336126 368716 336132
rect 369780 320890 369808 338028
rect 370240 336734 370268 338028
rect 370806 338014 371096 338042
rect 370228 336728 370280 336734
rect 370228 336670 370280 336676
rect 370504 336388 370556 336394
rect 370504 336330 370556 336336
rect 369768 320884 369820 320890
rect 369768 320826 369820 320832
rect 370516 21418 370544 336330
rect 371068 22778 371096 338014
rect 371344 336734 371372 338028
rect 371148 336728 371200 336734
rect 371148 336670 371200 336676
rect 371332 336728 371384 336734
rect 371332 336670 371384 336676
rect 371056 22772 371108 22778
rect 371056 22714 371108 22720
rect 370504 21412 370556 21418
rect 370504 21354 370556 21360
rect 370596 4412 370648 4418
rect 370596 4354 370648 4360
rect 369400 3256 369452 3262
rect 369400 3198 369452 3204
rect 368388 3052 368440 3058
rect 368388 2994 368440 3000
rect 369412 480 369440 3198
rect 370608 480 370636 4354
rect 371160 3126 371188 336670
rect 371804 336258 371832 338028
rect 372370 338014 372568 338042
rect 372436 336728 372488 336734
rect 372436 336670 372488 336676
rect 371792 336252 371844 336258
rect 371792 336194 371844 336200
rect 371240 326392 371292 326398
rect 371240 326334 371292 326340
rect 371252 16574 371280 326334
rect 372448 175982 372476 336670
rect 372436 175976 372488 175982
rect 372436 175918 372488 175924
rect 372540 24138 372568 338014
rect 372908 333334 372936 338028
rect 373474 338014 373764 338042
rect 372896 333328 372948 333334
rect 372896 333270 372948 333276
rect 372528 24132 372580 24138
rect 372528 24074 372580 24080
rect 371252 16546 371740 16574
rect 371148 3120 371200 3126
rect 371148 3062 371200 3068
rect 371712 480 371740 16546
rect 372896 3324 372948 3330
rect 372896 3266 372948 3272
rect 372908 480 372936 3266
rect 373736 3194 373764 338014
rect 373828 338014 373934 338042
rect 373828 5710 373856 338014
rect 374472 336734 374500 338028
rect 374460 336728 374512 336734
rect 374460 336670 374512 336676
rect 375024 336054 375052 338028
rect 375484 336734 375512 338028
rect 376050 338014 376524 338042
rect 376602 338014 376708 338042
rect 375288 336728 375340 336734
rect 375288 336670 375340 336676
rect 375472 336728 375524 336734
rect 375472 336670 375524 336676
rect 374644 336048 374696 336054
rect 374644 335990 374696 335996
rect 375012 336048 375064 336054
rect 375012 335990 375064 335996
rect 374000 10328 374052 10334
rect 374000 10270 374052 10276
rect 373816 5704 373868 5710
rect 373816 5646 373868 5652
rect 374012 3330 374040 10270
rect 374656 9042 374684 335990
rect 375300 319462 375328 336670
rect 375288 319456 375340 319462
rect 375288 319398 375340 319404
rect 376496 316742 376524 338014
rect 376576 336728 376628 336734
rect 376576 336670 376628 336676
rect 376484 316736 376536 316742
rect 376484 316678 376536 316684
rect 374644 9036 374696 9042
rect 374644 8978 374696 8984
rect 376588 5778 376616 336670
rect 376576 5772 376628 5778
rect 376576 5714 376628 5720
rect 374092 4480 374144 4486
rect 374092 4422 374144 4428
rect 374000 3324 374052 3330
rect 374000 3266 374052 3272
rect 373724 3188 373776 3194
rect 373724 3130 373776 3136
rect 374104 480 374132 4422
rect 376484 3392 376536 3398
rect 376484 3334 376536 3340
rect 375288 3324 375340 3330
rect 375288 3266 375340 3272
rect 375300 480 375328 3266
rect 376496 480 376524 3334
rect 376680 3262 376708 338014
rect 377140 336734 377168 338028
rect 377614 338014 377996 338042
rect 377128 336728 377180 336734
rect 377128 336670 377180 336676
rect 377968 318102 377996 338014
rect 378048 336728 378100 336734
rect 378048 336670 378100 336676
rect 377956 318096 378008 318102
rect 377956 318038 378008 318044
rect 378060 5846 378088 336670
rect 378152 336122 378180 338028
rect 378704 336734 378732 338028
rect 379178 338014 379376 338042
rect 378692 336728 378744 336734
rect 378692 336670 378744 336676
rect 378140 336116 378192 336122
rect 378140 336058 378192 336064
rect 379348 25566 379376 338014
rect 379428 336728 379480 336734
rect 379428 336670 379480 336676
rect 379336 25560 379388 25566
rect 379336 25502 379388 25508
rect 378140 20052 378192 20058
rect 378140 19994 378192 20000
rect 378152 16574 378180 19994
rect 378152 16546 378916 16574
rect 378048 5840 378100 5846
rect 378048 5782 378100 5788
rect 377680 4616 377732 4622
rect 377680 4558 377732 4564
rect 376668 3256 376720 3262
rect 376668 3198 376720 3204
rect 377692 480 377720 4558
rect 378888 480 378916 16546
rect 379440 5914 379468 336670
rect 379716 336190 379744 338028
rect 380282 338014 380756 338042
rect 380624 336728 380676 336734
rect 380624 336670 380676 336676
rect 379704 336184 379756 336190
rect 379704 336126 379756 336132
rect 380636 329118 380664 336670
rect 380624 329112 380676 329118
rect 380624 329054 380676 329060
rect 380728 5982 380756 338014
rect 380820 336734 380848 338028
rect 380808 336728 380860 336734
rect 380808 336670 380860 336676
rect 380808 336184 380860 336190
rect 380808 336126 380860 336132
rect 380716 5976 380768 5982
rect 380716 5918 380768 5924
rect 379428 5908 379480 5914
rect 379428 5850 379480 5856
rect 379980 4140 380032 4146
rect 379980 4082 380032 4088
rect 379992 480 380020 4082
rect 380820 3330 380848 336126
rect 381280 336054 381308 338028
rect 381846 338014 382228 338042
rect 381268 336048 381320 336054
rect 381268 335990 381320 335996
rect 382200 8974 382228 338014
rect 382384 336734 382412 338028
rect 382950 338014 383332 338042
rect 382372 336728 382424 336734
rect 382372 336670 382424 336676
rect 383304 325694 383332 338014
rect 383396 331974 383424 338028
rect 383568 336728 383620 336734
rect 383568 336670 383620 336676
rect 383384 331968 383436 331974
rect 383384 331910 383436 331916
rect 383304 325666 383516 325694
rect 383488 315314 383516 325666
rect 383476 315308 383528 315314
rect 383476 315250 383528 315256
rect 382372 11756 382424 11762
rect 382372 11698 382424 11704
rect 382188 8968 382240 8974
rect 382188 8910 382240 8916
rect 381176 4684 381228 4690
rect 381176 4626 381228 4632
rect 380808 3324 380860 3330
rect 380808 3266 380860 3272
rect 381188 480 381216 4626
rect 382384 480 382412 11698
rect 383580 6050 383608 336670
rect 383948 335374 383976 338028
rect 384514 338014 384896 338042
rect 383936 335368 383988 335374
rect 383936 335310 383988 335316
rect 384868 311166 384896 338014
rect 384960 336734 384988 338028
rect 384948 336728 385000 336734
rect 384948 336670 385000 336676
rect 385512 335986 385540 338028
rect 386078 338014 386276 338042
rect 385684 336728 385736 336734
rect 385684 336670 385736 336676
rect 385500 335980 385552 335986
rect 385500 335922 385552 335928
rect 384948 335232 385000 335238
rect 384948 335174 385000 335180
rect 384856 311160 384908 311166
rect 384856 311102 384908 311108
rect 384960 6118 384988 335174
rect 385696 10334 385724 336670
rect 386248 251870 386276 338014
rect 386328 335980 386380 335986
rect 386328 335922 386380 335928
rect 386236 251864 386288 251870
rect 386236 251806 386288 251812
rect 385960 14476 386012 14482
rect 385960 14418 386012 14424
rect 385684 10328 385736 10334
rect 385684 10270 385736 10276
rect 384948 6112 385000 6118
rect 384948 6054 385000 6060
rect 383568 6044 383620 6050
rect 383568 5986 383620 5992
rect 384764 4752 384816 4758
rect 384764 4694 384816 4700
rect 383568 4072 383620 4078
rect 383568 4014 383620 4020
rect 383580 480 383608 4014
rect 384776 480 384804 4694
rect 385972 480 386000 14418
rect 386340 6866 386368 335922
rect 386616 334694 386644 338028
rect 387090 338014 387564 338042
rect 386604 334688 386656 334694
rect 386604 334630 386656 334636
rect 386328 6860 386380 6866
rect 386328 6802 386380 6808
rect 387536 6798 387564 338014
rect 387628 326398 387656 338028
rect 388180 336734 388208 338028
rect 388654 338014 389128 338042
rect 388168 336728 388220 336734
rect 388168 336670 388220 336676
rect 388996 336728 389048 336734
rect 388996 336670 389048 336676
rect 387616 326392 387668 326398
rect 387616 326334 387668 326340
rect 389008 13122 389036 336670
rect 388996 13116 389048 13122
rect 388996 13058 389048 13064
rect 387524 6792 387576 6798
rect 387524 6734 387576 6740
rect 389100 6730 389128 338014
rect 389192 335986 389220 338028
rect 389758 338014 390232 338042
rect 390310 338014 390508 338042
rect 390204 336682 390232 338014
rect 390204 336654 390416 336682
rect 389180 335980 389232 335986
rect 389180 335922 389232 335928
rect 390284 335980 390336 335986
rect 390284 335922 390336 335928
rect 390296 313954 390324 335922
rect 390284 313948 390336 313954
rect 390284 313890 390336 313896
rect 390388 14482 390416 336654
rect 390376 14476 390428 14482
rect 390376 14418 390428 14424
rect 389456 13184 389508 13190
rect 389456 13126 389508 13132
rect 389088 6724 389140 6730
rect 389088 6666 389140 6672
rect 388260 5432 388312 5438
rect 388260 5374 388312 5380
rect 387156 4004 387208 4010
rect 387156 3946 387208 3952
rect 387168 480 387196 3946
rect 388272 480 388300 5374
rect 389468 480 389496 13126
rect 390480 6662 390508 338014
rect 390756 336734 390784 338028
rect 390744 336728 390796 336734
rect 390744 336670 390796 336676
rect 391308 330546 391336 338028
rect 391756 336728 391808 336734
rect 391756 336670 391808 336676
rect 391296 330540 391348 330546
rect 391296 330482 391348 330488
rect 391768 323610 391796 336670
rect 391756 323604 391808 323610
rect 391756 323546 391808 323552
rect 390468 6656 390520 6662
rect 390468 6598 390520 6604
rect 391860 6594 391888 338028
rect 392320 336734 392348 338028
rect 392886 338014 393268 338042
rect 392308 336728 392360 336734
rect 392308 336670 392360 336676
rect 393136 336728 393188 336734
rect 393136 336670 393188 336676
rect 393148 309806 393176 336670
rect 393136 309800 393188 309806
rect 393136 309742 393188 309748
rect 391940 25628 391992 25634
rect 391940 25570 391992 25576
rect 391952 16574 391980 25570
rect 391952 16546 393084 16574
rect 391848 6588 391900 6594
rect 391848 6530 391900 6536
rect 391848 5500 391900 5506
rect 391848 5442 391900 5448
rect 390652 3936 390704 3942
rect 390652 3878 390704 3884
rect 390664 480 390692 3878
rect 391860 480 391888 5442
rect 393056 480 393084 16546
rect 393240 11762 393268 338014
rect 393424 335986 393452 338028
rect 393990 338014 394372 338042
rect 394450 338014 394648 338042
rect 394344 336682 394372 338014
rect 394344 336654 394556 336682
rect 393412 335980 393464 335986
rect 393412 335922 393464 335928
rect 394424 335980 394476 335986
rect 394424 335922 394476 335928
rect 393228 11756 393280 11762
rect 393228 11698 393280 11704
rect 394436 6526 394464 335922
rect 394528 307086 394556 336654
rect 394620 333266 394648 338014
rect 394988 336734 395016 338028
rect 395554 338014 395936 338042
rect 394976 336728 395028 336734
rect 394976 336670 395028 336676
rect 394608 333260 394660 333266
rect 394608 333202 394660 333208
rect 395908 308446 395936 338014
rect 395988 336728 396040 336734
rect 395988 336670 396040 336676
rect 395896 308440 395948 308446
rect 395896 308382 395948 308388
rect 394516 307080 394568 307086
rect 394516 307022 394568 307028
rect 394424 6520 394476 6526
rect 394424 6462 394476 6468
rect 396000 6458 396028 336670
rect 396092 335986 396120 338028
rect 396552 336734 396580 338028
rect 397118 338014 397224 338042
rect 396540 336728 396592 336734
rect 396540 336670 396592 336676
rect 396080 335980 396132 335986
rect 396080 335922 396132 335928
rect 397196 305658 397224 338014
rect 397276 336728 397328 336734
rect 397276 336670 397328 336676
rect 397184 305652 397236 305658
rect 397184 305594 397236 305600
rect 396080 26920 396132 26926
rect 396080 26862 396132 26868
rect 396092 16574 396120 26862
rect 396092 16546 396580 16574
rect 395988 6452 396040 6458
rect 395988 6394 396040 6400
rect 395344 5364 395396 5370
rect 395344 5306 395396 5312
rect 394240 3868 394292 3874
rect 394240 3810 394292 3816
rect 394252 480 394280 3810
rect 395356 480 395384 5306
rect 396552 480 396580 16546
rect 397288 6390 397316 336670
rect 397656 335986 397684 338028
rect 398116 336734 398144 338028
rect 398576 338014 398682 338042
rect 398104 336728 398156 336734
rect 398104 336670 398156 336676
rect 397368 335980 397420 335986
rect 397368 335922 397420 335928
rect 397644 335980 397696 335986
rect 397644 335922 397696 335928
rect 397276 6384 397328 6390
rect 397276 6326 397328 6332
rect 397380 4282 397408 335922
rect 398576 327758 398604 338014
rect 399220 336734 399248 338028
rect 399786 338014 400076 338042
rect 398656 336728 398708 336734
rect 398656 336670 398708 336676
rect 399208 336728 399260 336734
rect 399208 336670 399260 336676
rect 398564 327752 398616 327758
rect 398564 327694 398616 327700
rect 398668 6322 398696 336670
rect 398748 335980 398800 335986
rect 398748 335922 398800 335928
rect 398656 6316 398708 6322
rect 398656 6258 398708 6264
rect 398760 4350 398788 335922
rect 398840 29640 398892 29646
rect 398840 29582 398892 29588
rect 398748 4344 398800 4350
rect 398748 4286 398800 4292
rect 397368 4276 397420 4282
rect 397368 4218 397420 4224
rect 397736 3800 397788 3806
rect 397736 3742 397788 3748
rect 397748 480 397776 3742
rect 398852 3398 398880 29582
rect 400048 6254 400076 338014
rect 400232 336734 400260 338028
rect 400128 336728 400180 336734
rect 400128 336670 400180 336676
rect 400220 336728 400272 336734
rect 400220 336670 400272 336676
rect 400036 6248 400088 6254
rect 400036 6190 400088 6196
rect 398932 5296 398984 5302
rect 398932 5238 398984 5244
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 5238
rect 400140 4418 400168 336670
rect 400784 335986 400812 338028
rect 401350 338014 401456 338042
rect 401324 336728 401376 336734
rect 401324 336670 401376 336676
rect 400772 335980 400824 335986
rect 400772 335922 400824 335928
rect 401336 302938 401364 336670
rect 401324 302932 401376 302938
rect 401324 302874 401376 302880
rect 401428 6186 401456 338014
rect 401508 335980 401560 335986
rect 401508 335922 401560 335928
rect 401416 6180 401468 6186
rect 401416 6122 401468 6128
rect 401520 4486 401548 335922
rect 401796 331906 401824 338028
rect 402348 336734 402376 338028
rect 402808 338014 402914 338042
rect 403466 338014 403848 338042
rect 403926 338014 404308 338042
rect 402336 336728 402388 336734
rect 402336 336670 402388 336676
rect 401784 331900 401836 331906
rect 401784 331842 401836 331848
rect 402808 7342 402836 338014
rect 402888 336728 402940 336734
rect 402888 336670 402940 336676
rect 402796 7336 402848 7342
rect 402796 7278 402848 7284
rect 402520 5228 402572 5234
rect 402520 5170 402572 5176
rect 401508 4480 401560 4486
rect 401508 4422 401560 4428
rect 400128 4412 400180 4418
rect 400128 4354 400180 4360
rect 401324 3732 401376 3738
rect 401324 3674 401376 3680
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 401336 480 401364 3674
rect 402532 480 402560 5170
rect 402900 4554 402928 336670
rect 403820 335354 403848 338014
rect 403820 335326 404216 335354
rect 402980 324964 403032 324970
rect 402980 324906 403032 324912
rect 402992 16574 403020 324906
rect 404188 301510 404216 335326
rect 404176 301504 404228 301510
rect 404176 301446 404228 301452
rect 402992 16546 403664 16574
rect 402888 4548 402940 4554
rect 402888 4490 402940 4496
rect 403636 480 403664 16546
rect 404280 4622 404308 338014
rect 404464 336734 404492 338028
rect 404452 336728 404504 336734
rect 404452 336670 404504 336676
rect 405016 334626 405044 338028
rect 405476 338014 405582 338042
rect 405004 334620 405056 334626
rect 405004 334562 405056 334568
rect 405476 4690 405504 338014
rect 406028 336734 406056 338028
rect 406594 338014 406976 338042
rect 405556 336728 405608 336734
rect 405556 336670 405608 336676
rect 406016 336728 406068 336734
rect 406016 336670 406068 336676
rect 405568 7410 405596 336670
rect 406948 304298 406976 338014
rect 407132 336734 407160 338028
rect 407606 338014 408080 338042
rect 408158 338014 408448 338042
rect 407028 336728 407080 336734
rect 407028 336670 407080 336676
rect 407120 336728 407172 336734
rect 407120 336670 407172 336676
rect 406936 304292 406988 304298
rect 406936 304234 406988 304240
rect 407040 7478 407068 336670
rect 407396 336660 407448 336666
rect 407396 336602 407448 336608
rect 407212 10396 407264 10402
rect 407212 10338 407264 10344
rect 407028 7472 407080 7478
rect 407028 7414 407080 7420
rect 405556 7404 405608 7410
rect 405556 7346 405608 7352
rect 406016 5160 406068 5166
rect 406016 5102 406068 5108
rect 405464 4684 405516 4690
rect 405464 4626 405516 4632
rect 404268 4616 404320 4622
rect 404268 4558 404320 4564
rect 404820 3664 404872 3670
rect 404820 3606 404872 3612
rect 404832 480 404860 3606
rect 406028 480 406056 5102
rect 407224 480 407252 10338
rect 407408 6914 407436 336602
rect 408052 335354 408080 338014
rect 408316 336728 408368 336734
rect 408316 336670 408368 336676
rect 408052 335326 408264 335354
rect 408236 7546 408264 335326
rect 408224 7540 408276 7546
rect 408224 7482 408276 7488
rect 407408 6886 408264 6914
rect 408236 3482 408264 6886
rect 408328 4758 408356 336670
rect 408316 4752 408368 4758
rect 408316 4694 408368 4700
rect 408420 3618 408448 338014
rect 408696 336734 408724 338028
rect 409262 338014 409644 338042
rect 409722 338014 409828 338042
rect 408684 336728 408736 336734
rect 408684 336670 408736 336676
rect 409616 8294 409644 338014
rect 409696 336728 409748 336734
rect 409696 336670 409748 336676
rect 409604 8288 409656 8294
rect 409604 8230 409656 8236
rect 409708 5506 409736 336670
rect 409696 5500 409748 5506
rect 409696 5442 409748 5448
rect 409604 5092 409656 5098
rect 409604 5034 409656 5040
rect 408420 3590 408540 3618
rect 408236 3454 408448 3482
rect 408420 480 408448 3454
rect 408512 3398 408540 3590
rect 408500 3392 408552 3398
rect 408500 3334 408552 3340
rect 409616 480 409644 5034
rect 409800 4146 409828 338014
rect 410260 336734 410288 338028
rect 410826 338014 411116 338042
rect 410248 336728 410300 336734
rect 410248 336670 410300 336676
rect 409880 330608 409932 330614
rect 409880 330550 409932 330556
rect 409892 16574 409920 330550
rect 409892 16546 410840 16574
rect 409788 4140 409840 4146
rect 409788 4082 409840 4088
rect 410812 480 410840 16546
rect 411088 8226 411116 338014
rect 411168 336728 411220 336734
rect 411168 336670 411220 336676
rect 411076 8220 411128 8226
rect 411076 8162 411128 8168
rect 411180 5438 411208 336670
rect 411272 335578 411300 338028
rect 411824 336734 411852 338028
rect 411812 336728 411864 336734
rect 411812 336670 411864 336676
rect 411260 335572 411312 335578
rect 411260 335514 411312 335520
rect 412376 8158 412404 338028
rect 412456 336728 412508 336734
rect 412456 336670 412508 336676
rect 412364 8152 412416 8158
rect 412364 8094 412416 8100
rect 411168 5432 411220 5438
rect 411168 5374 411220 5380
rect 412468 5370 412496 336670
rect 412548 335572 412600 335578
rect 412548 335514 412600 335520
rect 412456 5364 412508 5370
rect 412456 5306 412508 5312
rect 412560 4078 412588 335514
rect 412928 335374 412956 338028
rect 413388 336734 413416 338028
rect 413756 338014 413954 338042
rect 413376 336728 413428 336734
rect 413376 336670 413428 336676
rect 412916 335368 412968 335374
rect 412916 335310 412968 335316
rect 413756 8090 413784 338014
rect 414492 336734 414520 338028
rect 414966 338014 415256 338042
rect 413836 336728 413888 336734
rect 413836 336670 413888 336676
rect 414480 336728 414532 336734
rect 414480 336670 414532 336676
rect 413744 8084 413796 8090
rect 413744 8026 413796 8032
rect 413848 5302 413876 336670
rect 413928 335232 413980 335238
rect 413928 335174 413980 335180
rect 413836 5296 413888 5302
rect 413836 5238 413888 5244
rect 413100 5024 413152 5030
rect 413100 4966 413152 4972
rect 412548 4072 412600 4078
rect 412548 4014 412600 4020
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 411916 480 411944 3538
rect 413112 480 413140 4966
rect 413940 4010 413968 335174
rect 414020 28280 414072 28286
rect 414020 28222 414072 28228
rect 414032 16574 414060 28222
rect 414032 16546 414336 16574
rect 413928 4004 413980 4010
rect 413928 3946 413980 3952
rect 414308 480 414336 16546
rect 415228 5234 415256 338014
rect 415504 336734 415532 338028
rect 415308 336728 415360 336734
rect 415308 336670 415360 336676
rect 415492 336728 415544 336734
rect 415492 336670 415544 336676
rect 415216 5228 415268 5234
rect 415216 5170 415268 5176
rect 415320 3942 415348 336670
rect 416056 336666 416084 338028
rect 416504 336728 416556 336734
rect 416504 336670 416556 336676
rect 416044 336660 416096 336666
rect 416044 336602 416096 336608
rect 415676 336592 415728 336598
rect 415676 336534 415728 336540
rect 415688 6914 415716 336534
rect 416516 8022 416544 336670
rect 416504 8016 416556 8022
rect 416504 7958 416556 7964
rect 415504 6886 415716 6914
rect 415308 3936 415360 3942
rect 415308 3878 415360 3884
rect 415504 480 415532 6886
rect 416608 5166 416636 338028
rect 417068 336666 417096 338028
rect 417634 338014 418108 338042
rect 416688 336660 416740 336666
rect 416688 336602 416740 336608
rect 417056 336660 417108 336666
rect 417056 336602 417108 336608
rect 417976 336660 418028 336666
rect 417976 336602 418028 336608
rect 416596 5160 416648 5166
rect 416596 5102 416648 5108
rect 416700 4978 416728 336602
rect 416780 31068 416832 31074
rect 416780 31010 416832 31016
rect 416792 16574 416820 31010
rect 416792 16546 417924 16574
rect 416504 4956 416556 4962
rect 416504 4898 416556 4904
rect 416608 4950 416728 4978
rect 416516 2530 416544 4898
rect 416608 3874 416636 4950
rect 416596 3868 416648 3874
rect 416596 3810 416648 3816
rect 416516 2502 416728 2530
rect 416700 480 416728 2502
rect 417896 480 417924 16546
rect 417988 7954 418016 336602
rect 417976 7948 418028 7954
rect 417976 7890 418028 7896
rect 418080 3806 418108 338014
rect 418172 336734 418200 338028
rect 418738 338014 419120 338042
rect 419198 338014 419488 338042
rect 418160 336728 418212 336734
rect 418160 336670 418212 336676
rect 419092 335354 419120 338014
rect 419356 336728 419408 336734
rect 419356 336670 419408 336676
rect 419092 335326 419304 335354
rect 419276 7138 419304 335326
rect 419264 7132 419316 7138
rect 419264 7074 419316 7080
rect 419368 5098 419396 336670
rect 419356 5092 419408 5098
rect 419356 5034 419408 5040
rect 418068 3800 418120 3806
rect 418068 3742 418120 3748
rect 419460 3738 419488 338014
rect 419736 336734 419764 338028
rect 420302 338014 420684 338042
rect 420762 338014 420868 338042
rect 419724 336728 419776 336734
rect 419724 336670 419776 336676
rect 420656 7886 420684 338014
rect 420736 336728 420788 336734
rect 420736 336670 420788 336676
rect 420644 7880 420696 7886
rect 420644 7822 420696 7828
rect 420748 5030 420776 336670
rect 420736 5024 420788 5030
rect 420736 4966 420788 4972
rect 420184 4888 420236 4894
rect 420184 4830 420236 4836
rect 419448 3732 419500 3738
rect 419448 3674 419500 3680
rect 418988 3528 419040 3534
rect 418988 3470 419040 3476
rect 419000 480 419028 3470
rect 420196 480 420224 4830
rect 420840 3670 420868 338014
rect 421300 336666 421328 338028
rect 421866 338014 422156 338042
rect 421288 336660 421340 336666
rect 421288 336602 421340 336608
rect 420920 323672 420972 323678
rect 420920 323614 420972 323620
rect 420932 16574 420960 323614
rect 420932 16546 421420 16574
rect 420828 3664 420880 3670
rect 420828 3606 420880 3612
rect 421392 480 421420 16546
rect 422128 7818 422156 338014
rect 422404 336666 422432 338028
rect 422864 336734 422892 338028
rect 422852 336728 422904 336734
rect 422852 336670 422904 336676
rect 422208 336660 422260 336666
rect 422208 336602 422260 336608
rect 422392 336660 422444 336666
rect 422392 336602 422444 336608
rect 422116 7812 422168 7818
rect 422116 7754 422168 7760
rect 422220 4962 422248 336602
rect 422576 336524 422628 336530
rect 422576 336466 422628 336472
rect 422208 4956 422260 4962
rect 422208 4898 422260 4904
rect 422588 480 422616 336466
rect 423416 7750 423444 338028
rect 423496 336728 423548 336734
rect 423496 336670 423548 336676
rect 423404 7744 423456 7750
rect 423404 7686 423456 7692
rect 423508 4894 423536 336670
rect 423588 336660 423640 336666
rect 423588 336602 423640 336608
rect 423496 4888 423548 4894
rect 423496 4830 423548 4836
rect 423600 3602 423628 336602
rect 423968 335374 423996 338028
rect 424428 336734 424456 338028
rect 424796 338014 424994 338042
rect 425546 338014 425928 338042
rect 426098 338014 426388 338042
rect 424416 336728 424468 336734
rect 424416 336670 424468 336676
rect 423956 335368 424008 335374
rect 423956 335310 424008 335316
rect 423680 19984 423732 19990
rect 423680 19926 423732 19932
rect 423692 7614 423720 19926
rect 424692 8356 424744 8362
rect 424692 8298 424744 8304
rect 423680 7608 423732 7614
rect 423680 7550 423732 7556
rect 423772 4820 423824 4826
rect 423772 4762 423824 4768
rect 423588 3596 423640 3602
rect 423588 3538 423640 3544
rect 423784 480 423812 4762
rect 424704 3534 424732 8298
rect 424796 7682 424824 338014
rect 424876 336728 424928 336734
rect 424876 336670 424928 336676
rect 424784 7676 424836 7682
rect 424784 7618 424836 7624
rect 424888 4826 424916 336670
rect 425900 335354 425928 338014
rect 425900 335326 426296 335354
rect 424968 335232 425020 335238
rect 424968 335174 425020 335180
rect 424980 8362 425008 335174
rect 424968 8356 425020 8362
rect 424968 8298 425020 8304
rect 424968 7608 425020 7614
rect 424968 7550 425020 7556
rect 424876 4820 424928 4826
rect 424876 4762 424928 4768
rect 424692 3528 424744 3534
rect 424692 3470 424744 3476
rect 424980 480 425008 7550
rect 426268 3466 426296 335326
rect 426360 3777 426388 338014
rect 426544 336598 426572 338028
rect 427110 338014 427492 338042
rect 427662 338014 427768 338042
rect 427464 336682 427492 338014
rect 427464 336654 427676 336682
rect 426532 336592 426584 336598
rect 426532 336534 426584 336540
rect 427544 336592 427596 336598
rect 427544 336534 427596 336540
rect 427268 9036 427320 9042
rect 427268 8978 427320 8984
rect 426346 3768 426402 3777
rect 426346 3703 426402 3712
rect 426164 3460 426216 3466
rect 426164 3402 426216 3408
rect 426256 3460 426308 3466
rect 426256 3402 426308 3408
rect 426176 480 426204 3402
rect 427280 480 427308 8978
rect 427556 3505 427584 336534
rect 427648 3641 427676 336654
rect 427634 3632 427690 3641
rect 427634 3567 427690 3576
rect 427542 3496 427598 3505
rect 427542 3431 427598 3440
rect 427740 3369 427768 338014
rect 429212 299470 429240 405855
rect 429566 402792 429622 402801
rect 429566 402727 429568 402736
rect 429620 402727 429622 402736
rect 429568 402698 429620 402704
rect 429290 399800 429346 399809
rect 429290 399735 429346 399744
rect 429200 299464 429252 299470
rect 429200 299406 429252 299412
rect 429304 273222 429332 399735
rect 429382 396808 429438 396817
rect 429382 396743 429438 396752
rect 429292 273216 429344 273222
rect 429292 273158 429344 273164
rect 429396 259418 429424 396743
rect 429474 393816 429530 393825
rect 429474 393751 429530 393760
rect 429384 259412 429436 259418
rect 429384 259354 429436 259360
rect 429488 245614 429516 393751
rect 429566 390824 429622 390833
rect 429566 390759 429568 390768
rect 429620 390759 429622 390768
rect 429568 390730 429620 390736
rect 429568 387864 429620 387870
rect 429566 387832 429568 387841
rect 429620 387832 429622 387841
rect 429566 387767 429622 387776
rect 429566 384704 429622 384713
rect 429566 384639 429622 384648
rect 429476 245608 429528 245614
rect 429476 245550 429528 245556
rect 429580 206990 429608 384639
rect 429658 381712 429714 381721
rect 429658 381647 429714 381656
rect 429568 206984 429620 206990
rect 429568 206926 429620 206932
rect 429672 193186 429700 381647
rect 429750 378720 429806 378729
rect 429750 378655 429806 378664
rect 429660 193180 429712 193186
rect 429660 193122 429712 193128
rect 429764 179382 429792 378655
rect 429856 364334 429884 417823
rect 429948 373994 429976 420951
rect 430040 379506 430068 423943
rect 430132 391950 430160 426935
rect 430224 405686 430252 429927
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 433984 414860 434036 414866
rect 433984 414802 434036 414808
rect 430212 405680 430264 405686
rect 430212 405622 430264 405628
rect 432604 402756 432656 402762
rect 432604 402698 432656 402704
rect 430120 391944 430172 391950
rect 430120 391886 430172 391892
rect 431224 390788 431276 390794
rect 431224 390730 431276 390736
rect 430028 379500 430080 379506
rect 430028 379442 430080 379448
rect 430486 375728 430542 375737
rect 430486 375663 430542 375672
rect 429948 373966 430068 373994
rect 429934 369608 429990 369617
rect 429934 369543 429990 369552
rect 429948 368558 429976 369543
rect 429936 368552 429988 368558
rect 429936 368494 429988 368500
rect 430040 365702 430068 373966
rect 430394 372736 430450 372745
rect 430394 372671 430450 372680
rect 430302 366616 430358 366625
rect 430302 366551 430358 366560
rect 430028 365696 430080 365702
rect 430028 365638 430080 365644
rect 429856 364306 429976 364334
rect 429842 354512 429898 354521
rect 429842 354447 429898 354456
rect 429856 353138 429884 354447
rect 429948 353258 429976 364306
rect 430210 363624 430266 363633
rect 430210 363559 430266 363568
rect 430118 360632 430174 360641
rect 430118 360567 430174 360576
rect 430026 357640 430082 357649
rect 430026 357575 430082 357584
rect 429936 353252 429988 353258
rect 429936 353194 429988 353200
rect 429856 353110 429976 353138
rect 429842 351520 429898 351529
rect 429842 351455 429898 351464
rect 429856 350606 429884 351455
rect 429844 350600 429896 350606
rect 429844 350542 429896 350548
rect 429842 348528 429898 348537
rect 429842 348463 429898 348472
rect 429856 347818 429884 348463
rect 429844 347812 429896 347818
rect 429844 347754 429896 347760
rect 429842 345536 429898 345545
rect 429842 345471 429898 345480
rect 429752 179376 429804 179382
rect 429752 179318 429804 179324
rect 429856 33114 429884 345471
rect 429948 73166 429976 353110
rect 430040 86970 430068 357575
rect 430132 100706 430160 360567
rect 430224 113150 430252 363559
rect 430316 126954 430344 366551
rect 430408 153202 430436 372671
rect 430500 167006 430528 375663
rect 431236 233238 431264 390730
rect 432616 285666 432644 402698
rect 433996 339454 434024 414802
rect 435364 411324 435416 411330
rect 435364 411266 435416 411272
rect 433984 339448 434036 339454
rect 433984 339390 434036 339396
rect 434720 326460 434772 326466
rect 434720 326402 434772 326408
rect 432604 285660 432656 285666
rect 432604 285602 432656 285608
rect 431224 233232 431276 233238
rect 431224 233174 431276 233180
rect 430580 232552 430632 232558
rect 430580 232494 430632 232500
rect 430488 167000 430540 167006
rect 430488 166942 430540 166948
rect 430396 153196 430448 153202
rect 430396 153138 430448 153144
rect 430304 126948 430356 126954
rect 430304 126890 430356 126896
rect 430212 113144 430264 113150
rect 430212 113086 430264 113092
rect 430120 100700 430172 100706
rect 430120 100642 430172 100648
rect 430028 86964 430080 86970
rect 430028 86906 430080 86912
rect 429936 73160 429988 73166
rect 429936 73102 429988 73108
rect 429844 33108 429896 33114
rect 429844 33050 429896 33056
rect 430592 16574 430620 232494
rect 434732 16574 434760 326402
rect 435376 325650 435404 411266
rect 461584 408536 461636 408542
rect 461584 408478 461636 408484
rect 454684 387864 454736 387870
rect 454684 387806 454736 387812
rect 447784 368552 447836 368558
rect 447784 368494 447836 368500
rect 442264 350600 442316 350606
rect 442264 350542 442316 350548
rect 439504 347812 439556 347818
rect 439504 347754 439556 347760
rect 436100 336456 436152 336462
rect 436100 336398 436152 336404
rect 435364 325644 435416 325650
rect 435364 325586 435416 325592
rect 436112 16574 436140 336398
rect 437480 329180 437532 329186
rect 437480 329122 437532 329128
rect 437492 16574 437520 329122
rect 439516 46918 439544 347754
rect 441620 174548 441672 174554
rect 441620 174490 441672 174496
rect 439504 46912 439556 46918
rect 439504 46854 439556 46860
rect 438860 44872 438912 44878
rect 438860 44814 438912 44820
rect 438872 16574 438900 44814
rect 440332 17264 440384 17270
rect 440332 17206 440384 17212
rect 430592 16546 430896 16574
rect 434732 16546 435588 16574
rect 436112 16546 436784 16574
rect 437492 16546 437980 16574
rect 438872 16546 439176 16574
rect 428464 7200 428516 7206
rect 428464 7142 428516 7148
rect 427726 3360 427782 3369
rect 427726 3295 427782 3304
rect 428476 480 428504 7142
rect 429660 2848 429712 2854
rect 429660 2790 429712 2796
rect 429672 480 429700 2790
rect 430868 480 430896 16546
rect 434444 15904 434496 15910
rect 434444 15846 434496 15852
rect 432052 7268 432104 7274
rect 432052 7210 432104 7216
rect 432064 480 432092 7210
rect 433248 2916 433300 2922
rect 433248 2858 433300 2864
rect 433260 480 433288 2858
rect 434456 480 434484 15846
rect 435560 480 435588 16546
rect 436756 480 436784 16546
rect 437952 480 437980 16546
rect 439148 480 439176 16546
rect 440344 2990 440372 17206
rect 441632 16574 441660 174490
rect 442276 60722 442304 350542
rect 443000 336388 443052 336394
rect 443000 336330 443052 336336
rect 442264 60716 442316 60722
rect 442264 60658 442316 60664
rect 443012 16574 443040 336330
rect 445760 322244 445812 322250
rect 445760 322186 445812 322192
rect 444380 18624 444432 18630
rect 444380 18566 444432 18572
rect 444392 16574 444420 18566
rect 445772 16574 445800 322186
rect 447796 139398 447824 368494
rect 449900 336320 449952 336326
rect 449900 336262 449952 336268
rect 448520 327820 448572 327826
rect 448520 327762 448572 327768
rect 447784 139392 447836 139398
rect 447784 139334 447836 139340
rect 441632 16546 442672 16574
rect 443012 16546 443868 16574
rect 444392 16546 445064 16574
rect 445772 16546 446260 16574
rect 440240 2984 440292 2990
rect 440240 2926 440292 2932
rect 440332 2984 440384 2990
rect 440332 2926 440384 2932
rect 441528 2984 441580 2990
rect 441528 2926 441580 2932
rect 440252 1578 440280 2926
rect 440252 1550 440372 1578
rect 440344 480 440372 1550
rect 441540 480 441568 2926
rect 442644 480 442672 16546
rect 443840 480 443868 16546
rect 445036 480 445064 16546
rect 446232 480 446260 16546
rect 448532 3482 448560 327762
rect 448612 35216 448664 35222
rect 448612 35158 448664 35164
rect 448624 4214 448652 35158
rect 449912 16574 449940 336262
rect 452660 320884 452712 320890
rect 452660 320826 452712 320832
rect 451280 21412 451332 21418
rect 451280 21354 451332 21360
rect 451292 16574 451320 21354
rect 452672 16574 452700 320826
rect 454696 219434 454724 387806
rect 456800 336252 456852 336258
rect 456800 336194 456852 336200
rect 454684 219428 454736 219434
rect 454684 219370 454736 219376
rect 455420 22772 455472 22778
rect 455420 22714 455472 22720
rect 455432 16574 455460 22714
rect 449912 16546 450952 16574
rect 451292 16546 452148 16574
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 448612 4208 448664 4214
rect 448612 4150 448664 4156
rect 449808 4208 449860 4214
rect 449808 4150 449860 4156
rect 448532 3454 448652 3482
rect 447416 3052 447468 3058
rect 447416 2994 447468 3000
rect 447428 480 447456 2994
rect 448624 480 448652 3454
rect 449820 480 449848 4150
rect 450924 480 450952 16546
rect 452120 480 452148 16546
rect 453316 480 453344 16546
rect 454500 3120 454552 3126
rect 454500 3062 454552 3068
rect 454512 480 454540 3062
rect 455708 480 455736 16546
rect 456812 3126 456840 336194
rect 459560 333328 459612 333334
rect 459560 333270 459612 333276
rect 456892 175976 456944 175982
rect 456892 175918 456944 175924
rect 456800 3120 456852 3126
rect 456800 3062 456852 3068
rect 456904 480 456932 175918
rect 458180 24132 458232 24138
rect 458180 24074 458232 24080
rect 458192 16574 458220 24074
rect 459572 16574 459600 333270
rect 461596 313274 461624 408478
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 391944 580224 391950
rect 580172 391886 580224 391892
rect 580184 391785 580212 391886
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 489184 339516 489236 339522
rect 489184 339458 489236 339464
rect 465080 336184 465132 336190
rect 465080 336126 465132 336132
rect 463700 319456 463752 319462
rect 463700 319398 463752 319404
rect 461584 313268 461636 313274
rect 461584 313210 461636 313216
rect 463712 16574 463740 319398
rect 465092 16574 465120 336126
rect 471980 336116 472032 336122
rect 471980 336058 472032 336064
rect 470600 318096 470652 318102
rect 470600 318038 470652 318044
rect 466460 316736 466512 316742
rect 466460 316678 466512 316684
rect 466472 16574 466500 316678
rect 470612 16574 470640 318038
rect 471992 16574 472020 336058
rect 478880 336048 478932 336054
rect 478880 335990 478932 335996
rect 477500 329112 477552 329118
rect 477500 329054 477552 329060
rect 473360 25560 473412 25566
rect 473360 25502 473412 25508
rect 458192 16546 459232 16574
rect 459572 16546 460428 16574
rect 463712 16546 464016 16574
rect 465092 16546 465212 16574
rect 466472 16546 467512 16574
rect 470612 16546 471100 16574
rect 471992 16546 472296 16574
rect 458088 3120 458140 3126
rect 458088 3062 458140 3068
rect 458100 480 458128 3062
rect 459204 480 459232 16546
rect 460400 480 460428 16546
rect 462780 5704 462832 5710
rect 462780 5646 462832 5652
rect 461584 3188 461636 3194
rect 461584 3130 461636 3136
rect 461596 480 461624 3130
rect 462792 480 462820 5646
rect 463988 480 464016 16546
rect 465184 480 465212 16546
rect 466276 5772 466328 5778
rect 466276 5714 466328 5720
rect 466288 480 466316 5714
rect 467484 480 467512 16546
rect 469864 5840 469916 5846
rect 469864 5782 469916 5788
rect 468668 3256 468720 3262
rect 468668 3198 468720 3204
rect 468680 480 468708 3198
rect 469876 480 469904 5782
rect 471072 480 471100 16546
rect 472268 480 472296 16546
rect 473372 3330 473400 25502
rect 477512 16574 477540 329054
rect 478892 16574 478920 335990
rect 483020 331968 483072 331974
rect 483020 331910 483072 331916
rect 481640 315308 481692 315314
rect 481640 315250 481692 315256
rect 477512 16546 478184 16574
rect 478892 16546 479380 16574
rect 476948 5976 477000 5982
rect 476948 5918 477000 5924
rect 473452 5908 473504 5914
rect 473452 5850 473504 5856
rect 473360 3324 473412 3330
rect 473360 3266 473412 3272
rect 473464 480 473492 5850
rect 474556 3324 474608 3330
rect 474556 3266 474608 3272
rect 474568 480 474596 3266
rect 475752 3256 475804 3262
rect 475752 3198 475804 3204
rect 475764 480 475792 3198
rect 476960 480 476988 5918
rect 478156 480 478184 16546
rect 479352 480 479380 16546
rect 480536 8968 480588 8974
rect 480536 8910 480588 8916
rect 480548 480 480576 8910
rect 481652 3330 481680 315250
rect 483032 16574 483060 331910
rect 485780 311160 485832 311166
rect 485780 311102 485832 311108
rect 485792 16574 485820 311102
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 481732 6044 481784 6050
rect 481732 5986 481784 5992
rect 481640 3324 481692 3330
rect 481640 3266 481692 3272
rect 481744 480 481772 5986
rect 482836 3324 482888 3330
rect 482836 3266 482888 3272
rect 482848 480 482876 3266
rect 484044 480 484072 16546
rect 485228 6112 485280 6118
rect 485228 6054 485280 6060
rect 485240 480 485268 6054
rect 486436 480 486464 16546
rect 489196 11830 489224 339458
rect 579988 339448 580040 339454
rect 579988 339390 580040 339396
rect 580000 338609 580028 339390
rect 579986 338600 580042 338609
rect 579986 338535 580042 338544
rect 489920 334688 489972 334694
rect 489920 334630 489972 334636
rect 489184 11824 489236 11830
rect 489184 11766 489236 11772
rect 487620 10328 487672 10334
rect 487620 10270 487672 10276
rect 487632 480 487660 10270
rect 488816 6860 488868 6866
rect 488816 6802 488868 6808
rect 488828 480 488856 6802
rect 489932 3330 489960 334630
rect 531320 334620 531372 334626
rect 531320 334562 531372 334568
rect 507860 333260 507912 333266
rect 507860 333202 507912 333208
rect 500960 330540 501012 330546
rect 500960 330482 501012 330488
rect 492680 326392 492732 326398
rect 492680 326334 492732 326340
rect 490012 251864 490064 251870
rect 490012 251806 490064 251812
rect 489920 3324 489972 3330
rect 489920 3266 489972 3272
rect 490024 1442 490052 251806
rect 492692 16574 492720 326334
rect 499580 323604 499632 323610
rect 499580 323546 499632 323552
rect 496820 313948 496872 313954
rect 496820 313890 496872 313896
rect 496832 16574 496860 313890
rect 499592 16574 499620 323546
rect 500972 16574 501000 330482
rect 503720 309800 503772 309806
rect 503720 309742 503772 309748
rect 503732 16574 503760 309742
rect 506480 307080 506532 307086
rect 506480 307022 506532 307028
rect 492692 16546 493548 16574
rect 496832 16546 497136 16574
rect 499592 16546 500632 16574
rect 500972 16546 501828 16574
rect 503732 16546 504220 16574
rect 492312 6792 492364 6798
rect 492312 6734 492364 6740
rect 491116 3324 491168 3330
rect 491116 3266 491168 3272
rect 489932 1414 490052 1442
rect 489932 480 489960 1414
rect 491128 480 491156 3266
rect 492324 480 492352 6734
rect 493520 480 493548 16546
rect 494704 13116 494756 13122
rect 494704 13058 494756 13064
rect 494716 480 494744 13058
rect 495900 6724 495952 6730
rect 495900 6666 495952 6672
rect 495912 480 495940 6666
rect 497108 480 497136 16546
rect 498200 14476 498252 14482
rect 498200 14418 498252 14424
rect 498212 480 498240 14418
rect 499396 6656 499448 6662
rect 499396 6598 499448 6604
rect 499408 480 499436 6598
rect 500604 480 500632 16546
rect 501800 480 501828 16546
rect 502984 6588 503036 6594
rect 502984 6530 503036 6536
rect 502996 480 503024 6530
rect 504192 480 504220 16546
rect 505376 11756 505428 11762
rect 505376 11698 505428 11704
rect 505388 480 505416 11698
rect 506492 3330 506520 307022
rect 507872 16574 507900 333202
rect 524420 331900 524472 331906
rect 524420 331842 524472 331848
rect 517520 327752 517572 327758
rect 517520 327694 517572 327700
rect 510620 308440 510672 308446
rect 510620 308382 510672 308388
rect 510632 16574 510660 308382
rect 514760 305652 514812 305658
rect 514760 305594 514812 305600
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 506572 6520 506624 6526
rect 506572 6462 506624 6468
rect 506480 3324 506532 3330
rect 506480 3266 506532 3272
rect 506584 3210 506612 6462
rect 507676 3324 507728 3330
rect 507676 3266 507728 3272
rect 506492 3182 506612 3210
rect 506492 480 506520 3182
rect 507688 480 507716 3266
rect 508884 480 508912 16546
rect 510068 6452 510120 6458
rect 510068 6394 510120 6400
rect 510080 480 510108 6394
rect 511276 480 511304 16546
rect 513564 6384 513616 6390
rect 513564 6326 513616 6332
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 513576 480 513604 6326
rect 514772 480 514800 305594
rect 517532 16574 517560 327694
rect 521660 302932 521712 302938
rect 521660 302874 521712 302880
rect 521672 16574 521700 302874
rect 524432 16574 524460 331842
rect 528560 301504 528612 301510
rect 528560 301446 528612 301452
rect 528572 16574 528600 301446
rect 517532 16546 518388 16574
rect 521672 16546 521884 16574
rect 524432 16546 525472 16574
rect 528572 16546 529060 16574
rect 517152 6316 517204 6322
rect 517152 6258 517204 6264
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517164 480 517192 6258
rect 518360 480 518388 16546
rect 520740 6248 520792 6254
rect 520740 6190 520792 6196
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 519556 480 519584 4354
rect 520752 480 520780 6190
rect 521856 480 521884 16546
rect 524236 6180 524288 6186
rect 524236 6122 524288 6128
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 523052 480 523080 4422
rect 524248 480 524276 6122
rect 525444 480 525472 16546
rect 527824 7336 527876 7342
rect 527824 7278 527876 7284
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526640 480 526668 4490
rect 527836 480 527864 7278
rect 529032 480 529060 16546
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 530136 480 530164 4558
rect 531332 3330 531360 334562
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 535460 304292 535512 304298
rect 535460 304234 535512 304240
rect 535472 16574 535500 304234
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 285660 580224 285666
rect 580172 285602 580224 285608
rect 580184 285433 580212 285602
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 535472 16546 536144 16574
rect 534908 7472 534960 7478
rect 534908 7414 534960 7420
rect 531412 7404 531464 7410
rect 531412 7346 531464 7352
rect 531320 3324 531372 3330
rect 531320 3266 531372 3272
rect 531424 1442 531452 7346
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 532516 3324 532568 3330
rect 532516 3266 532568 3272
rect 531332 1414 531452 1442
rect 531332 480 531360 1414
rect 532528 480 532556 3266
rect 533724 480 533752 4626
rect 534920 480 534948 7414
rect 536116 480 536144 16546
rect 580264 11824 580316 11830
rect 580264 11766 580316 11772
rect 541992 8288 542044 8294
rect 541992 8230 542044 8236
rect 538404 7540 538456 7546
rect 538404 7482 538456 7488
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 538416 480 538444 7482
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3392 539652 3398
rect 539600 3334 539652 3340
rect 539612 480 539640 3334
rect 540808 480 540836 5442
rect 542004 480 542032 8230
rect 545488 8220 545540 8226
rect 545488 8162 545540 8168
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 4140 543240 4146
rect 543188 4082 543240 4088
rect 543200 480 543228 4082
rect 544396 480 544424 5374
rect 545500 480 545528 8162
rect 549076 8152 549128 8158
rect 549076 8094 549128 8100
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 4072 546736 4078
rect 546684 4014 546736 4020
rect 546696 480 546724 4014
rect 547892 480 547920 5306
rect 549088 480 549116 8094
rect 552664 8084 552716 8090
rect 552664 8026 552716 8032
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 4004 550324 4010
rect 550272 3946 550324 3952
rect 550284 480 550312 3946
rect 551480 480 551508 5238
rect 552676 480 552704 8026
rect 556160 8016 556212 8022
rect 556160 7958 556212 7964
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3936 553820 3942
rect 553768 3878 553820 3884
rect 553780 480 553808 3878
rect 554976 480 555004 5170
rect 556172 480 556200 7958
rect 559748 7948 559800 7954
rect 559748 7890 559800 7896
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3868 557408 3874
rect 557356 3810 557408 3816
rect 557368 480 557396 3810
rect 558564 480 558592 5102
rect 559760 480 559788 7890
rect 563244 7880 563296 7886
rect 563244 7822 563296 7828
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 560852 3800 560904 3806
rect 560852 3742 560904 3748
rect 560864 480 560892 3742
rect 562060 480 562088 5034
rect 563256 480 563284 7822
rect 566832 7812 566884 7818
rect 566832 7754 566884 7760
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 564440 3732 564492 3738
rect 564440 3674 564492 3680
rect 564452 480 564480 3674
rect 565648 480 565676 4966
rect 566844 480 566872 7754
rect 570328 7744 570380 7750
rect 570328 7686 570380 7692
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3664 568080 3670
rect 568028 3606 568080 3612
rect 568040 480 568068 3606
rect 569144 480 569172 4898
rect 570340 480 570368 7686
rect 573916 7676 573968 7682
rect 573916 7618 573968 7624
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 571524 3596 571576 3602
rect 571524 3538 571576 3544
rect 571536 480 571564 3538
rect 572732 480 572760 4830
rect 573928 480 573956 7618
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 575112 3528 575164 3534
rect 575112 3470 575164 3476
rect 575124 480 575152 3470
rect 576320 480 576348 4762
rect 577424 480 577452 7550
rect 580276 6633 580304 11766
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 579802 3768 579858 3777
rect 579802 3703 579858 3712
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 578620 480 578648 3402
rect 579816 480 579844 3703
rect 582194 3632 582250 3641
rect 582194 3567 582250 3576
rect 580998 3496 581054 3505
rect 580998 3431 581054 3440
rect 581012 480 581040 3431
rect 582208 480 582236 3567
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3146 553832 3202 553888
rect 3054 540776 3110 540832
rect 2962 527856 3018 527912
rect 2870 514800 2926 514856
rect 2778 501744 2834 501800
rect 3514 671200 3570 671256
rect 3606 658144 3662 658200
rect 3422 488688 3478 488744
rect 3698 645088 3754 645144
rect 3790 632032 3846 632088
rect 3882 619112 3938 619168
rect 3974 606056 4030 606112
rect 4066 593000 4122 593056
rect 3514 475632 3570 475688
rect 580170 697176 580226 697232
rect 165618 493312 165674 493368
rect 165618 490320 165674 490376
rect 165618 487328 165674 487384
rect 429382 487328 429438 487384
rect 165618 484472 165674 484528
rect 165618 481480 165674 481536
rect 165618 478488 165674 478544
rect 165618 475496 165674 475552
rect 429474 475224 429530 475280
rect 165618 472640 165674 472696
rect 165618 469648 165674 469704
rect 165618 466656 165674 466712
rect 165618 463664 165674 463720
rect 429198 463120 429254 463176
rect 3606 462576 3662 462632
rect 165618 460672 165674 460728
rect 165618 457816 165674 457872
rect 580170 683848 580226 683904
rect 429842 496304 429898 496360
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 429934 493312 429990 493368
rect 580170 670656 580226 670692
rect 580262 657328 580318 657384
rect 580170 644000 580226 644056
rect 430026 490320 430082 490376
rect 579986 630808 580042 630864
rect 429750 466112 429806 466168
rect 429658 460128 429714 460184
rect 429566 457136 429622 457192
rect 165618 454824 165674 454880
rect 429198 454144 429254 454200
rect 165618 451832 165674 451888
rect 429566 451016 429622 451072
rect 3698 449520 3754 449576
rect 165618 448840 165674 448896
rect 430118 484336 430174 484392
rect 580170 617480 580226 617536
rect 430210 481208 430266 481264
rect 579618 590960 579674 591016
rect 430302 478216 430358 478272
rect 579618 577632 579674 577688
rect 430394 472232 430450 472288
rect 429842 448024 429898 448080
rect 165618 445984 165674 446040
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580354 604152 580410 604208
rect 579618 484608 579674 484664
rect 580446 551112 580502 551168
rect 579618 471416 579674 471472
rect 430486 469240 430542 469296
rect 580538 511264 580594 511320
rect 580170 458088 580226 458144
rect 429934 445032 429990 445088
rect 165618 442992 165674 443048
rect 165618 440000 165674 440056
rect 580630 497936 580686 497992
rect 580170 444760 580226 444816
rect 430026 442040 430082 442096
rect 429842 439048 429898 439104
rect 165618 437008 165674 437064
rect 3422 436600 3478 436656
rect 429934 436056 429990 436112
rect 165618 434016 165674 434072
rect 429842 432928 429898 432984
rect 165618 431160 165674 431216
rect 3422 423544 3478 423600
rect 3054 332288 3110 332344
rect 3054 319232 3110 319288
rect 3146 306176 3202 306232
rect 3330 384376 3386 384432
rect 3238 293120 3294 293176
rect 3238 280100 3240 280120
rect 3240 280100 3292 280120
rect 3292 280100 3294 280120
rect 3238 280064 3294 280100
rect 3054 267144 3110 267200
rect 3238 254088 3294 254144
rect 3238 241032 3294 241088
rect 3238 227976 3294 228032
rect 3238 214920 3294 214976
rect 165618 428168 165674 428224
rect 166262 425176 166318 425232
rect 165618 422184 165674 422240
rect 165618 419328 165674 419384
rect 165618 416336 165674 416392
rect 3790 410488 3846 410544
rect 165618 407360 165674 407416
rect 165618 404504 165674 404560
rect 3698 397432 3754 397488
rect 165618 395528 165674 395584
rect 3606 371320 3662 371376
rect 3514 358400 3570 358456
rect 3422 345344 3478 345400
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3330 175888 3386 175944
rect 3330 149776 3386 149832
rect 3146 123664 3202 123720
rect 3146 84632 3202 84688
rect 2870 58520 2926 58576
rect 4066 162832 4122 162888
rect 3974 136720 4030 136776
rect 3882 110608 3938 110664
rect 3790 97552 3846 97608
rect 3698 71576 3754 71632
rect 3606 45464 3662 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 6458 3304 6514 3360
rect 15934 3576 15990 3632
rect 14738 3440 14794 3496
rect 165618 392672 165674 392728
rect 579802 431568 579858 431624
rect 430210 429936 430266 429992
rect 430118 426944 430174 427000
rect 430026 423952 430082 424008
rect 429934 420960 429990 421016
rect 429842 417832 429898 417888
rect 429566 414860 429622 414896
rect 429566 414840 429568 414860
rect 429568 414840 429620 414860
rect 429620 414840 429622 414860
rect 166906 413344 166962 413400
rect 166814 410352 166870 410408
rect 166722 401512 166778 401568
rect 166630 398520 166686 398576
rect 166538 389680 166594 389736
rect 166446 386688 166502 386744
rect 165618 383716 165674 383752
rect 165618 383696 165620 383716
rect 165620 383696 165672 383716
rect 165672 383696 165674 383716
rect 165618 380704 165674 380760
rect 166354 377848 166410 377904
rect 165618 374856 165674 374912
rect 165618 371864 165674 371920
rect 165618 368872 165674 368928
rect 166262 366016 166318 366072
rect 165618 363024 165674 363080
rect 165618 360032 165674 360088
rect 165618 357040 165674 357096
rect 165618 354048 165674 354104
rect 165618 351192 165674 351248
rect 24214 3712 24270 3768
rect 165618 348200 165674 348256
rect 165618 345208 165674 345264
rect 165618 342252 165620 342272
rect 165620 342252 165672 342272
rect 165672 342252 165674 342272
rect 165618 342216 165674 342252
rect 165618 339360 165674 339416
rect 429566 411848 429622 411904
rect 429474 408856 429530 408912
rect 429198 405864 429254 405920
rect 429106 339516 429162 339552
rect 429106 339496 429108 339516
rect 429108 339496 429160 339516
rect 429160 339496 429162 339516
rect 169942 3304 169998 3360
rect 174082 3576 174138 3632
rect 173990 3440 174046 3496
rect 178038 3712 178094 3768
rect 234618 3304 234674 3360
rect 237010 3440 237066 3496
rect 244094 3576 244150 3632
rect 276018 3712 276074 3768
rect 271878 3304 271934 3360
rect 273258 3440 273314 3496
rect 426346 3712 426402 3768
rect 427634 3576 427690 3632
rect 427542 3440 427598 3496
rect 429566 402756 429622 402792
rect 429566 402736 429568 402756
rect 429568 402736 429620 402756
rect 429620 402736 429622 402756
rect 429290 399744 429346 399800
rect 429382 396752 429438 396808
rect 429474 393760 429530 393816
rect 429566 390788 429622 390824
rect 429566 390768 429568 390788
rect 429568 390768 429620 390788
rect 429620 390768 429622 390788
rect 429566 387812 429568 387832
rect 429568 387812 429620 387832
rect 429620 387812 429622 387832
rect 429566 387776 429622 387812
rect 429566 384648 429622 384704
rect 429658 381656 429714 381712
rect 429750 378664 429806 378720
rect 580170 418240 580226 418296
rect 430486 375672 430542 375728
rect 429934 369552 429990 369608
rect 430394 372680 430450 372736
rect 430302 366560 430358 366616
rect 429842 354456 429898 354512
rect 430210 363568 430266 363624
rect 430118 360576 430174 360632
rect 430026 357584 430082 357640
rect 429842 351464 429898 351520
rect 429842 348472 429898 348528
rect 429842 345480 429898 345536
rect 427726 3304 427782 3360
rect 580170 404912 580226 404968
rect 580170 391720 580226 391776
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579986 338544 580042 338600
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 285368 580226 285424
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580262 6568 580318 6624
rect 579802 3712 579858 3768
rect 582194 3576 582250 3632
rect 580998 3440 581054 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3366 697370 3372 697372
rect -960 697310 3372 697370
rect -960 697220 480 697310
rect 3366 697308 3372 697310
rect 3436 697308 3442 697372
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3601 658202 3667 658205
rect -960 658200 3667 658202
rect -960 658144 3606 658200
rect 3662 658144 3667 658200
rect -960 658142 3667 658144
rect -960 658052 480 658142
rect 3601 658139 3667 658142
rect 580257 657386 580323 657389
rect 583520 657386 584960 657476
rect 580257 657384 584960 657386
rect 580257 657328 580262 657384
rect 580318 657328 584960 657384
rect 580257 657326 584960 657328
rect 580257 657323 580323 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 3693 645146 3759 645149
rect -960 645144 3759 645146
rect -960 645088 3698 645144
rect 3754 645088 3759 645144
rect -960 645086 3759 645088
rect -960 644996 480 645086
rect 3693 645083 3759 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3785 632090 3851 632093
rect -960 632088 3851 632090
rect -960 632032 3790 632088
rect 3846 632032 3851 632088
rect -960 632030 3851 632032
rect -960 631940 480 632030
rect 3785 632027 3851 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3877 619170 3943 619173
rect -960 619168 3943 619170
rect -960 619112 3882 619168
rect 3938 619112 3943 619168
rect -960 619110 3943 619112
rect -960 619020 480 619110
rect 3877 619107 3943 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3969 606114 4035 606117
rect -960 606112 4035 606114
rect -960 606056 3974 606112
rect 4030 606056 4035 606112
rect -960 606054 4035 606056
rect -960 605964 480 606054
rect 3969 606051 4035 606054
rect 580349 604210 580415 604213
rect 583520 604210 584960 604300
rect 580349 604208 584960 604210
rect 580349 604152 580354 604208
rect 580410 604152 584960 604208
rect 580349 604150 584960 604152
rect 580349 604147 580415 604150
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 4061 593058 4127 593061
rect -960 593056 4127 593058
rect -960 593000 4066 593056
rect 4122 593000 4127 593056
rect -960 592998 4127 593000
rect -960 592908 480 592998
rect 4061 592995 4127 592998
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect 580441 551170 580507 551173
rect 583520 551170 584960 551260
rect 580441 551168 584960 551170
rect 580441 551112 580446 551168
rect 580502 551112 584960 551168
rect 580441 551110 584960 551112
rect 580441 551107 580507 551110
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3049 540834 3115 540837
rect -960 540832 3115 540834
rect -960 540776 3054 540832
rect 3110 540776 3115 540832
rect -960 540774 3115 540776
rect -960 540684 480 540774
rect 3049 540771 3115 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2865 514858 2931 514861
rect -960 514856 2931 514858
rect -960 514800 2870 514856
rect 2926 514800 2931 514856
rect -960 514798 2931 514800
rect -960 514708 480 514798
rect 2865 514795 2931 514798
rect 580533 511322 580599 511325
rect 583520 511322 584960 511412
rect 580533 511320 584960 511322
rect 580533 511264 580538 511320
rect 580594 511264 584960 511320
rect 580533 511262 584960 511264
rect 580533 511259 580599 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 580625 497994 580691 497997
rect 583520 497994 584960 498084
rect 580625 497992 584960 497994
rect 580625 497936 580630 497992
rect 580686 497936 584960 497992
rect 580625 497934 584960 497936
rect 580625 497931 580691 497934
rect 583520 497844 584960 497934
rect 429837 496362 429903 496365
rect 427892 496360 429903 496362
rect 3366 495484 3372 495548
rect 3436 495546 3442 495548
rect 168054 495546 168114 496332
rect 427892 496304 429842 496360
rect 429898 496304 429903 496360
rect 427892 496302 429903 496304
rect 429837 496299 429903 496302
rect 3436 495486 168114 495546
rect 3436 495484 3442 495486
rect 165613 493370 165679 493373
rect 429929 493370 429995 493373
rect 165613 493368 168084 493370
rect 165613 493312 165618 493368
rect 165674 493312 168084 493368
rect 165613 493310 168084 493312
rect 427892 493368 429995 493370
rect 427892 493312 429934 493368
rect 429990 493312 429995 493368
rect 427892 493310 429995 493312
rect 165613 493307 165679 493310
rect 429929 493307 429995 493310
rect 165613 490378 165679 490381
rect 430021 490378 430087 490381
rect 165613 490376 168084 490378
rect 165613 490320 165618 490376
rect 165674 490320 168084 490376
rect 165613 490318 168084 490320
rect 427892 490376 430087 490378
rect 427892 490320 430026 490376
rect 430082 490320 430087 490376
rect 427892 490318 430087 490320
rect 165613 490315 165679 490318
rect 430021 490315 430087 490318
rect -960 488746 480 488836
rect 3417 488746 3483 488749
rect -960 488744 3483 488746
rect -960 488688 3422 488744
rect 3478 488688 3483 488744
rect -960 488686 3483 488688
rect -960 488596 480 488686
rect 3417 488683 3483 488686
rect 165613 487386 165679 487389
rect 429377 487386 429443 487389
rect 165613 487384 168084 487386
rect 165613 487328 165618 487384
rect 165674 487328 168084 487384
rect 165613 487326 168084 487328
rect 427892 487384 429443 487386
rect 427892 487328 429382 487384
rect 429438 487328 429443 487384
rect 427892 487326 429443 487328
rect 165613 487323 165679 487326
rect 429377 487323 429443 487326
rect 579613 484666 579679 484669
rect 583520 484666 584960 484756
rect 579613 484664 584960 484666
rect 579613 484608 579618 484664
rect 579674 484608 584960 484664
rect 579613 484606 584960 484608
rect 579613 484603 579679 484606
rect 165613 484530 165679 484533
rect 165613 484528 168084 484530
rect 165613 484472 165618 484528
rect 165674 484472 168084 484528
rect 583520 484516 584960 484606
rect 165613 484470 168084 484472
rect 165613 484467 165679 484470
rect 430113 484394 430179 484397
rect 427892 484392 430179 484394
rect 427892 484336 430118 484392
rect 430174 484336 430179 484392
rect 427892 484334 430179 484336
rect 430113 484331 430179 484334
rect 165613 481538 165679 481541
rect 165613 481536 168084 481538
rect 165613 481480 165618 481536
rect 165674 481480 168084 481536
rect 165613 481478 168084 481480
rect 165613 481475 165679 481478
rect 430205 481266 430271 481269
rect 427892 481264 430271 481266
rect 427892 481208 430210 481264
rect 430266 481208 430271 481264
rect 427892 481206 430271 481208
rect 430205 481203 430271 481206
rect 165613 478546 165679 478549
rect 165613 478544 168084 478546
rect 165613 478488 165618 478544
rect 165674 478488 168084 478544
rect 165613 478486 168084 478488
rect 165613 478483 165679 478486
rect 430297 478274 430363 478277
rect 427892 478272 430363 478274
rect 427892 478216 430302 478272
rect 430358 478216 430363 478272
rect 427892 478214 430363 478216
rect 430297 478211 430363 478214
rect -960 475690 480 475780
rect 3509 475690 3575 475693
rect -960 475688 3575 475690
rect -960 475632 3514 475688
rect 3570 475632 3575 475688
rect -960 475630 3575 475632
rect -960 475540 480 475630
rect 3509 475627 3575 475630
rect 165613 475554 165679 475557
rect 165613 475552 168084 475554
rect 165613 475496 165618 475552
rect 165674 475496 168084 475552
rect 165613 475494 168084 475496
rect 165613 475491 165679 475494
rect 429469 475282 429535 475285
rect 427892 475280 429535 475282
rect 427892 475224 429474 475280
rect 429530 475224 429535 475280
rect 427892 475222 429535 475224
rect 429469 475219 429535 475222
rect 165613 472698 165679 472701
rect 165613 472696 168084 472698
rect 165613 472640 165618 472696
rect 165674 472640 168084 472696
rect 165613 472638 168084 472640
rect 165613 472635 165679 472638
rect 430389 472290 430455 472293
rect 427892 472288 430455 472290
rect 427892 472232 430394 472288
rect 430450 472232 430455 472288
rect 427892 472230 430455 472232
rect 430389 472227 430455 472230
rect 579613 471474 579679 471477
rect 583520 471474 584960 471564
rect 579613 471472 584960 471474
rect 579613 471416 579618 471472
rect 579674 471416 584960 471472
rect 579613 471414 584960 471416
rect 579613 471411 579679 471414
rect 583520 471324 584960 471414
rect 165613 469706 165679 469709
rect 165613 469704 168084 469706
rect 165613 469648 165618 469704
rect 165674 469648 168084 469704
rect 165613 469646 168084 469648
rect 165613 469643 165679 469646
rect 430481 469298 430547 469301
rect 427892 469296 430547 469298
rect 427892 469240 430486 469296
rect 430542 469240 430547 469296
rect 427892 469238 430547 469240
rect 430481 469235 430547 469238
rect 165613 466714 165679 466717
rect 165613 466712 168084 466714
rect 165613 466656 165618 466712
rect 165674 466656 168084 466712
rect 165613 466654 168084 466656
rect 165613 466651 165679 466654
rect 429745 466170 429811 466173
rect 427892 466168 429811 466170
rect 427892 466112 429750 466168
rect 429806 466112 429811 466168
rect 427892 466110 429811 466112
rect 429745 466107 429811 466110
rect 165613 463722 165679 463725
rect 165613 463720 168084 463722
rect 165613 463664 165618 463720
rect 165674 463664 168084 463720
rect 165613 463662 168084 463664
rect 165613 463659 165679 463662
rect 429193 463178 429259 463181
rect 427892 463176 429259 463178
rect 427892 463120 429198 463176
rect 429254 463120 429259 463176
rect 427892 463118 429259 463120
rect 429193 463115 429259 463118
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 165613 460730 165679 460733
rect 165613 460728 168084 460730
rect 165613 460672 165618 460728
rect 165674 460672 168084 460728
rect 165613 460670 168084 460672
rect 165613 460667 165679 460670
rect 429653 460186 429719 460189
rect 427892 460184 429719 460186
rect 427892 460128 429658 460184
rect 429714 460128 429719 460184
rect 427892 460126 429719 460128
rect 429653 460123 429719 460126
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 165613 457874 165679 457877
rect 165613 457872 168084 457874
rect 165613 457816 165618 457872
rect 165674 457816 168084 457872
rect 165613 457814 168084 457816
rect 165613 457811 165679 457814
rect 429561 457194 429627 457197
rect 427892 457192 429627 457194
rect 427892 457136 429566 457192
rect 429622 457136 429627 457192
rect 427892 457134 429627 457136
rect 429561 457131 429627 457134
rect 165613 454882 165679 454885
rect 165613 454880 168084 454882
rect 165613 454824 165618 454880
rect 165674 454824 168084 454880
rect 165613 454822 168084 454824
rect 165613 454819 165679 454822
rect 429193 454202 429259 454205
rect 427892 454200 429259 454202
rect 427892 454144 429198 454200
rect 429254 454144 429259 454200
rect 427892 454142 429259 454144
rect 429193 454139 429259 454142
rect 165613 451890 165679 451893
rect 165613 451888 168084 451890
rect 165613 451832 165618 451888
rect 165674 451832 168084 451888
rect 165613 451830 168084 451832
rect 165613 451827 165679 451830
rect 429561 451074 429627 451077
rect 427892 451072 429627 451074
rect 427892 451016 429566 451072
rect 429622 451016 429627 451072
rect 427892 451014 429627 451016
rect 429561 451011 429627 451014
rect -960 449578 480 449668
rect 3693 449578 3759 449581
rect -960 449576 3759 449578
rect -960 449520 3698 449576
rect 3754 449520 3759 449576
rect -960 449518 3759 449520
rect -960 449428 480 449518
rect 3693 449515 3759 449518
rect 165613 448898 165679 448901
rect 165613 448896 168084 448898
rect 165613 448840 165618 448896
rect 165674 448840 168084 448896
rect 165613 448838 168084 448840
rect 165613 448835 165679 448838
rect 429837 448082 429903 448085
rect 427892 448080 429903 448082
rect 427892 448024 429842 448080
rect 429898 448024 429903 448080
rect 427892 448022 429903 448024
rect 429837 448019 429903 448022
rect 165613 446042 165679 446045
rect 165613 446040 168084 446042
rect 165613 445984 165618 446040
rect 165674 445984 168084 446040
rect 165613 445982 168084 445984
rect 165613 445979 165679 445982
rect 429929 445090 429995 445093
rect 427892 445088 429995 445090
rect 427892 445032 429934 445088
rect 429990 445032 429995 445088
rect 427892 445030 429995 445032
rect 429929 445027 429995 445030
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 165613 443050 165679 443053
rect 165613 443048 168084 443050
rect 165613 442992 165618 443048
rect 165674 442992 168084 443048
rect 165613 442990 168084 442992
rect 165613 442987 165679 442990
rect 430021 442098 430087 442101
rect 427892 442096 430087 442098
rect 427892 442040 430026 442096
rect 430082 442040 430087 442096
rect 427892 442038 430087 442040
rect 430021 442035 430087 442038
rect 165613 440058 165679 440061
rect 165613 440056 168084 440058
rect 165613 440000 165618 440056
rect 165674 440000 168084 440056
rect 165613 439998 168084 440000
rect 165613 439995 165679 439998
rect 429837 439106 429903 439109
rect 427892 439104 429903 439106
rect 427892 439048 429842 439104
rect 429898 439048 429903 439104
rect 427892 439046 429903 439048
rect 429837 439043 429903 439046
rect 165613 437066 165679 437069
rect 165613 437064 168084 437066
rect 165613 437008 165618 437064
rect 165674 437008 168084 437064
rect 165613 437006 168084 437008
rect 165613 437003 165679 437006
rect -960 436658 480 436748
rect 3417 436658 3483 436661
rect -960 436656 3483 436658
rect -960 436600 3422 436656
rect 3478 436600 3483 436656
rect -960 436598 3483 436600
rect -960 436508 480 436598
rect 3417 436595 3483 436598
rect 429929 436114 429995 436117
rect 427892 436112 429995 436114
rect 427892 436056 429934 436112
rect 429990 436056 429995 436112
rect 427892 436054 429995 436056
rect 429929 436051 429995 436054
rect 165613 434074 165679 434077
rect 165613 434072 168084 434074
rect 165613 434016 165618 434072
rect 165674 434016 168084 434072
rect 165613 434014 168084 434016
rect 165613 434011 165679 434014
rect 429837 432986 429903 432989
rect 427892 432984 429903 432986
rect 427892 432928 429842 432984
rect 429898 432928 429903 432984
rect 427892 432926 429903 432928
rect 429837 432923 429903 432926
rect 579797 431626 579863 431629
rect 583520 431626 584960 431716
rect 579797 431624 584960 431626
rect 579797 431568 579802 431624
rect 579858 431568 584960 431624
rect 579797 431566 584960 431568
rect 579797 431563 579863 431566
rect 583520 431476 584960 431566
rect 165613 431218 165679 431221
rect 165613 431216 168084 431218
rect 165613 431160 165618 431216
rect 165674 431160 168084 431216
rect 165613 431158 168084 431160
rect 165613 431155 165679 431158
rect 430205 429994 430271 429997
rect 427892 429992 430271 429994
rect 427892 429936 430210 429992
rect 430266 429936 430271 429992
rect 427892 429934 430271 429936
rect 430205 429931 430271 429934
rect 165613 428226 165679 428229
rect 165613 428224 168084 428226
rect 165613 428168 165618 428224
rect 165674 428168 168084 428224
rect 165613 428166 168084 428168
rect 165613 428163 165679 428166
rect 430113 427002 430179 427005
rect 427892 427000 430179 427002
rect 427892 426944 430118 427000
rect 430174 426944 430179 427000
rect 427892 426942 430179 426944
rect 430113 426939 430179 426942
rect 166257 425234 166323 425237
rect 166257 425232 168084 425234
rect 166257 425176 166262 425232
rect 166318 425176 168084 425232
rect 166257 425174 168084 425176
rect 166257 425171 166323 425174
rect 430021 424010 430087 424013
rect 427892 424008 430087 424010
rect 427892 423952 430026 424008
rect 430082 423952 430087 424008
rect 427892 423950 430087 423952
rect 430021 423947 430087 423950
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 165613 422242 165679 422245
rect 165613 422240 168084 422242
rect 165613 422184 165618 422240
rect 165674 422184 168084 422240
rect 165613 422182 168084 422184
rect 165613 422179 165679 422182
rect 429929 421018 429995 421021
rect 427892 421016 429995 421018
rect 427892 420960 429934 421016
rect 429990 420960 429995 421016
rect 427892 420958 429995 420960
rect 429929 420955 429995 420958
rect 165613 419386 165679 419389
rect 165613 419384 168084 419386
rect 165613 419328 165618 419384
rect 165674 419328 168084 419384
rect 165613 419326 168084 419328
rect 165613 419323 165679 419326
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 429837 417890 429903 417893
rect 427892 417888 429903 417890
rect 427892 417832 429842 417888
rect 429898 417832 429903 417888
rect 427892 417830 429903 417832
rect 429837 417827 429903 417830
rect 165613 416394 165679 416397
rect 165613 416392 168084 416394
rect 165613 416336 165618 416392
rect 165674 416336 168084 416392
rect 165613 416334 168084 416336
rect 165613 416331 165679 416334
rect 429561 414898 429627 414901
rect 427892 414896 429627 414898
rect 427892 414840 429566 414896
rect 429622 414840 429627 414896
rect 427892 414838 429627 414840
rect 429561 414835 429627 414838
rect 166901 413402 166967 413405
rect 166901 413400 168084 413402
rect 166901 413344 166906 413400
rect 166962 413344 168084 413400
rect 166901 413342 168084 413344
rect 166901 413339 166967 413342
rect 429561 411906 429627 411909
rect 427892 411904 429627 411906
rect 427892 411848 429566 411904
rect 429622 411848 429627 411904
rect 427892 411846 429627 411848
rect 429561 411843 429627 411846
rect -960 410546 480 410636
rect 3785 410546 3851 410549
rect -960 410544 3851 410546
rect -960 410488 3790 410544
rect 3846 410488 3851 410544
rect -960 410486 3851 410488
rect -960 410396 480 410486
rect 3785 410483 3851 410486
rect 166809 410410 166875 410413
rect 166809 410408 168084 410410
rect 166809 410352 166814 410408
rect 166870 410352 168084 410408
rect 166809 410350 168084 410352
rect 166809 410347 166875 410350
rect 429469 408914 429535 408917
rect 427892 408912 429535 408914
rect 427892 408856 429474 408912
rect 429530 408856 429535 408912
rect 427892 408854 429535 408856
rect 429469 408851 429535 408854
rect 165613 407418 165679 407421
rect 165613 407416 168084 407418
rect 165613 407360 165618 407416
rect 165674 407360 168084 407416
rect 165613 407358 168084 407360
rect 165613 407355 165679 407358
rect 429193 405922 429259 405925
rect 427892 405920 429259 405922
rect 427892 405864 429198 405920
rect 429254 405864 429259 405920
rect 427892 405862 429259 405864
rect 429193 405859 429259 405862
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 165613 404562 165679 404565
rect 165613 404560 168084 404562
rect 165613 404504 165618 404560
rect 165674 404504 168084 404560
rect 165613 404502 168084 404504
rect 165613 404499 165679 404502
rect 429561 402794 429627 402797
rect 427892 402792 429627 402794
rect 427892 402736 429566 402792
rect 429622 402736 429627 402792
rect 427892 402734 429627 402736
rect 429561 402731 429627 402734
rect 166717 401570 166783 401573
rect 166717 401568 168084 401570
rect 166717 401512 166722 401568
rect 166778 401512 168084 401568
rect 166717 401510 168084 401512
rect 166717 401507 166783 401510
rect 429285 399802 429351 399805
rect 427892 399800 429351 399802
rect 427892 399744 429290 399800
rect 429346 399744 429351 399800
rect 427892 399742 429351 399744
rect 429285 399739 429351 399742
rect 166625 398578 166691 398581
rect 166625 398576 168084 398578
rect 166625 398520 166630 398576
rect 166686 398520 168084 398576
rect 166625 398518 168084 398520
rect 166625 398515 166691 398518
rect -960 397490 480 397580
rect 3693 397490 3759 397493
rect -960 397488 3759 397490
rect -960 397432 3698 397488
rect 3754 397432 3759 397488
rect -960 397430 3759 397432
rect -960 397340 480 397430
rect 3693 397427 3759 397430
rect 429377 396810 429443 396813
rect 427892 396808 429443 396810
rect 427892 396752 429382 396808
rect 429438 396752 429443 396808
rect 427892 396750 429443 396752
rect 429377 396747 429443 396750
rect 165613 395586 165679 395589
rect 165613 395584 168084 395586
rect 165613 395528 165618 395584
rect 165674 395528 168084 395584
rect 165613 395526 168084 395528
rect 165613 395523 165679 395526
rect 429469 393818 429535 393821
rect 427892 393816 429535 393818
rect 427892 393760 429474 393816
rect 429530 393760 429535 393816
rect 427892 393758 429535 393760
rect 429469 393755 429535 393758
rect 165613 392730 165679 392733
rect 165613 392728 168084 392730
rect 165613 392672 165618 392728
rect 165674 392672 168084 392728
rect 165613 392670 168084 392672
rect 165613 392667 165679 392670
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect 429561 390826 429627 390829
rect 427892 390824 429627 390826
rect 427892 390768 429566 390824
rect 429622 390768 429627 390824
rect 427892 390766 429627 390768
rect 429561 390763 429627 390766
rect 166533 389738 166599 389741
rect 166533 389736 168084 389738
rect 166533 389680 166538 389736
rect 166594 389680 168084 389736
rect 166533 389678 168084 389680
rect 166533 389675 166599 389678
rect 429561 387834 429627 387837
rect 427892 387832 429627 387834
rect 427892 387776 429566 387832
rect 429622 387776 429627 387832
rect 427892 387774 429627 387776
rect 429561 387771 429627 387774
rect 166441 386746 166507 386749
rect 166441 386744 168084 386746
rect 166441 386688 166446 386744
rect 166502 386688 168084 386744
rect 166441 386686 168084 386688
rect 166441 386683 166507 386686
rect 429561 384706 429627 384709
rect 427892 384704 429627 384706
rect 427892 384648 429566 384704
rect 429622 384648 429627 384704
rect 427892 384646 429627 384648
rect 429561 384643 429627 384646
rect -960 384434 480 384524
rect 3325 384434 3391 384437
rect -960 384432 3391 384434
rect -960 384376 3330 384432
rect 3386 384376 3391 384432
rect -960 384374 3391 384376
rect -960 384284 480 384374
rect 3325 384371 3391 384374
rect 165613 383754 165679 383757
rect 165613 383752 168084 383754
rect 165613 383696 165618 383752
rect 165674 383696 168084 383752
rect 165613 383694 168084 383696
rect 165613 383691 165679 383694
rect 429653 381714 429719 381717
rect 427892 381712 429719 381714
rect 427892 381656 429658 381712
rect 429714 381656 429719 381712
rect 427892 381654 429719 381656
rect 429653 381651 429719 381654
rect 165613 380762 165679 380765
rect 165613 380760 168084 380762
rect 165613 380704 165618 380760
rect 165674 380704 168084 380760
rect 165613 380702 168084 380704
rect 165613 380699 165679 380702
rect 429745 378722 429811 378725
rect 427892 378720 429811 378722
rect 427892 378664 429750 378720
rect 429806 378664 429811 378720
rect 427892 378662 429811 378664
rect 429745 378659 429811 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 166349 377906 166415 377909
rect 166349 377904 168084 377906
rect 166349 377848 166354 377904
rect 166410 377848 168084 377904
rect 166349 377846 168084 377848
rect 166349 377843 166415 377846
rect 430481 375730 430547 375733
rect 427892 375728 430547 375730
rect 427892 375672 430486 375728
rect 430542 375672 430547 375728
rect 427892 375670 430547 375672
rect 430481 375667 430547 375670
rect 165613 374914 165679 374917
rect 165613 374912 168084 374914
rect 165613 374856 165618 374912
rect 165674 374856 168084 374912
rect 165613 374854 168084 374856
rect 165613 374851 165679 374854
rect 430389 372738 430455 372741
rect 427892 372736 430455 372738
rect 427892 372680 430394 372736
rect 430450 372680 430455 372736
rect 427892 372678 430455 372680
rect 430389 372675 430455 372678
rect 165613 371922 165679 371925
rect 165613 371920 168084 371922
rect 165613 371864 165618 371920
rect 165674 371864 168084 371920
rect 165613 371862 168084 371864
rect 165613 371859 165679 371862
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 429929 369610 429995 369613
rect 427892 369608 429995 369610
rect 427892 369552 429934 369608
rect 429990 369552 429995 369608
rect 427892 369550 429995 369552
rect 429929 369547 429995 369550
rect 165613 368930 165679 368933
rect 165613 368928 168084 368930
rect 165613 368872 165618 368928
rect 165674 368872 168084 368928
rect 165613 368870 168084 368872
rect 165613 368867 165679 368870
rect 430297 366618 430363 366621
rect 427892 366616 430363 366618
rect 427892 366560 430302 366616
rect 430358 366560 430363 366616
rect 427892 366558 430363 366560
rect 430297 366555 430363 366558
rect 166257 366074 166323 366077
rect 166257 366072 168084 366074
rect 166257 366016 166262 366072
rect 166318 366016 168084 366072
rect 166257 366014 168084 366016
rect 166257 366011 166323 366014
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 430205 363626 430271 363629
rect 427892 363624 430271 363626
rect 427892 363568 430210 363624
rect 430266 363568 430271 363624
rect 427892 363566 430271 363568
rect 430205 363563 430271 363566
rect 165613 363082 165679 363085
rect 165613 363080 168084 363082
rect 165613 363024 165618 363080
rect 165674 363024 168084 363080
rect 165613 363022 168084 363024
rect 165613 363019 165679 363022
rect 430113 360634 430179 360637
rect 427892 360632 430179 360634
rect 427892 360576 430118 360632
rect 430174 360576 430179 360632
rect 427892 360574 430179 360576
rect 430113 360571 430179 360574
rect 165613 360090 165679 360093
rect 165613 360088 168084 360090
rect 165613 360032 165618 360088
rect 165674 360032 168084 360088
rect 165613 360030 168084 360032
rect 165613 360027 165679 360030
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 430021 357642 430087 357645
rect 427892 357640 430087 357642
rect 427892 357584 430026 357640
rect 430082 357584 430087 357640
rect 427892 357582 430087 357584
rect 430021 357579 430087 357582
rect 165613 357098 165679 357101
rect 165613 357096 168084 357098
rect 165613 357040 165618 357096
rect 165674 357040 168084 357096
rect 165613 357038 168084 357040
rect 165613 357035 165679 357038
rect 429837 354514 429903 354517
rect 427892 354512 429903 354514
rect 427892 354456 429842 354512
rect 429898 354456 429903 354512
rect 427892 354454 429903 354456
rect 429837 354451 429903 354454
rect 165613 354106 165679 354109
rect 165613 354104 168084 354106
rect 165613 354048 165618 354104
rect 165674 354048 168084 354104
rect 165613 354046 168084 354048
rect 165613 354043 165679 354046
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 429837 351522 429903 351525
rect 427892 351520 429903 351522
rect 427892 351464 429842 351520
rect 429898 351464 429903 351520
rect 427892 351462 429903 351464
rect 429837 351459 429903 351462
rect 165613 351250 165679 351253
rect 165613 351248 168084 351250
rect 165613 351192 165618 351248
rect 165674 351192 168084 351248
rect 165613 351190 168084 351192
rect 165613 351187 165679 351190
rect 429837 348530 429903 348533
rect 427892 348528 429903 348530
rect 427892 348472 429842 348528
rect 429898 348472 429903 348528
rect 427892 348470 429903 348472
rect 429837 348467 429903 348470
rect 165613 348258 165679 348261
rect 165613 348256 168084 348258
rect 165613 348200 165618 348256
rect 165674 348200 168084 348256
rect 165613 348198 168084 348200
rect 165613 348195 165679 348198
rect 429837 345538 429903 345541
rect 427892 345536 429903 345538
rect -960 345402 480 345492
rect 427892 345480 429842 345536
rect 429898 345480 429903 345536
rect 427892 345478 429903 345480
rect 429837 345475 429903 345478
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 165613 345266 165679 345269
rect 165613 345264 168084 345266
rect 165613 345208 165618 345264
rect 165674 345208 168084 345264
rect 165613 345206 168084 345208
rect 165613 345203 165679 345206
rect 429694 342546 429700 342548
rect 427892 342486 429700 342546
rect 429694 342484 429700 342486
rect 429764 342484 429770 342548
rect 165613 342274 165679 342277
rect 165613 342272 168084 342274
rect 165613 342216 165618 342272
rect 165674 342216 168084 342272
rect 165613 342214 168084 342216
rect 165613 342211 165679 342214
rect 429101 339554 429167 339557
rect 427892 339552 429167 339554
rect 427892 339496 429106 339552
rect 429162 339496 429167 339552
rect 427892 339494 429167 339496
rect 429101 339491 429167 339494
rect 165613 339418 165679 339421
rect 165613 339416 168084 339418
rect 165613 339360 165618 339416
rect 165674 339360 168084 339416
rect 165613 339358 168084 339360
rect 165613 339355 165679 339358
rect 579981 338602 580047 338605
rect 583520 338602 584960 338692
rect 579981 338600 584960 338602
rect 579981 338544 579986 338600
rect 580042 338544 584960 338600
rect 579981 338542 584960 338544
rect 579981 338539 580047 338542
rect 583520 338452 584960 338542
rect -960 332346 480 332436
rect 3049 332346 3115 332349
rect -960 332344 3115 332346
rect -960 332288 3054 332344
rect 3110 332288 3115 332344
rect -960 332286 3115 332288
rect -960 332196 480 332286
rect 3049 332283 3115 332286
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3049 319290 3115 319293
rect -960 319288 3115 319290
rect -960 319232 3054 319288
rect 3110 319232 3115 319288
rect -960 319230 3115 319232
rect -960 319140 480 319230
rect 3049 319227 3115 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3141 306234 3207 306237
rect -960 306232 3207 306234
rect -960 306176 3146 306232
rect 3202 306176 3207 306232
rect -960 306174 3207 306176
rect -960 306084 480 306174
rect 3141 306171 3207 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3233 293178 3299 293181
rect -960 293176 3299 293178
rect -960 293120 3238 293176
rect 3294 293120 3299 293176
rect -960 293118 3299 293120
rect -960 293028 480 293118
rect 3233 293115 3299 293118
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect -960 280122 480 280212
rect 3233 280122 3299 280125
rect -960 280120 3299 280122
rect -960 280064 3238 280120
rect 3294 280064 3299 280120
rect -960 280062 3299 280064
rect -960 279972 480 280062
rect 3233 280059 3299 280062
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3233 254146 3299 254149
rect -960 254144 3299 254146
rect -960 254088 3238 254144
rect 3294 254088 3299 254144
rect -960 254086 3299 254088
rect -960 253996 480 254086
rect 3233 254083 3299 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3233 228034 3299 228037
rect -960 228032 3299 228034
rect -960 227976 3238 228032
rect 3294 227976 3299 228032
rect -960 227974 3299 227976
rect -960 227884 480 227974
rect 3233 227971 3299 227974
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3233 214978 3299 214981
rect -960 214976 3299 214978
rect -960 214920 3238 214976
rect 3294 214920 3299 214976
rect -960 214918 3299 214920
rect -960 214828 480 214918
rect 3233 214915 3299 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 3325 175946 3391 175949
rect -960 175944 3391 175946
rect -960 175888 3330 175944
rect 3386 175888 3391 175944
rect -960 175886 3391 175888
rect -960 175796 480 175886
rect 3325 175883 3391 175886
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 4061 162890 4127 162893
rect -960 162888 4127 162890
rect -960 162832 4066 162888
rect 4122 162832 4127 162888
rect -960 162830 4127 162832
rect -960 162740 480 162830
rect 4061 162827 4127 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3969 136778 4035 136781
rect -960 136776 4035 136778
rect -960 136720 3974 136776
rect 4030 136720 4035 136776
rect -960 136718 4035 136720
rect -960 136628 480 136718
rect 3969 136715 4035 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3141 123722 3207 123725
rect -960 123720 3207 123722
rect -960 123664 3146 123720
rect 3202 123664 3207 123720
rect -960 123662 3207 123664
rect -960 123572 480 123662
rect 3141 123659 3207 123662
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3877 110666 3943 110669
rect -960 110664 3943 110666
rect -960 110608 3882 110664
rect 3938 110608 3943 110664
rect -960 110606 3943 110608
rect -960 110516 480 110606
rect 3877 110603 3943 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3785 97610 3851 97613
rect -960 97608 3851 97610
rect -960 97552 3790 97608
rect 3846 97552 3851 97608
rect -960 97550 3851 97552
rect -960 97460 480 97550
rect 3785 97547 3851 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3693 71634 3759 71637
rect -960 71632 3759 71634
rect -960 71576 3698 71632
rect 3754 71576 3759 71632
rect -960 71574 3759 71576
rect -960 71484 480 71574
rect 3693 71571 3759 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2865 58578 2931 58581
rect -960 58576 2931 58578
rect -960 58520 2870 58576
rect 2926 58520 2931 58576
rect -960 58518 2931 58520
rect -960 58428 480 58518
rect 2865 58515 2931 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 583520 19818 584960 19908
rect 567150 19758 584960 19818
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 429694 19348 429700 19412
rect 429764 19410 429770 19412
rect 567150 19410 567210 19758
rect 583520 19668 584960 19758
rect 429764 19350 567210 19410
rect 429764 19348 429770 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 24209 3770 24275 3773
rect 178033 3770 178099 3773
rect 276013 3770 276079 3773
rect 24209 3768 178099 3770
rect 24209 3712 24214 3768
rect 24270 3712 178038 3768
rect 178094 3712 178099 3768
rect 24209 3710 178099 3712
rect 24209 3707 24275 3710
rect 178033 3707 178099 3710
rect 258030 3768 276079 3770
rect 258030 3712 276018 3768
rect 276074 3712 276079 3768
rect 258030 3710 276079 3712
rect 15929 3634 15995 3637
rect 174077 3634 174143 3637
rect 15929 3632 174143 3634
rect 15929 3576 15934 3632
rect 15990 3576 174082 3632
rect 174138 3576 174143 3632
rect 15929 3574 174143 3576
rect 15929 3571 15995 3574
rect 174077 3571 174143 3574
rect 244089 3634 244155 3637
rect 258030 3634 258090 3710
rect 276013 3707 276079 3710
rect 426341 3770 426407 3773
rect 579797 3770 579863 3773
rect 426341 3768 579863 3770
rect 426341 3712 426346 3768
rect 426402 3712 579802 3768
rect 579858 3712 579863 3768
rect 426341 3710 579863 3712
rect 426341 3707 426407 3710
rect 579797 3707 579863 3710
rect 244089 3632 258090 3634
rect 244089 3576 244094 3632
rect 244150 3576 258090 3632
rect 244089 3574 258090 3576
rect 427629 3634 427695 3637
rect 582189 3634 582255 3637
rect 427629 3632 582255 3634
rect 427629 3576 427634 3632
rect 427690 3576 582194 3632
rect 582250 3576 582255 3632
rect 427629 3574 582255 3576
rect 244089 3571 244155 3574
rect 427629 3571 427695 3574
rect 582189 3571 582255 3574
rect 14733 3498 14799 3501
rect 173985 3498 174051 3501
rect 14733 3496 174051 3498
rect 14733 3440 14738 3496
rect 14794 3440 173990 3496
rect 174046 3440 174051 3496
rect 14733 3438 174051 3440
rect 14733 3435 14799 3438
rect 173985 3435 174051 3438
rect 237005 3498 237071 3501
rect 273253 3498 273319 3501
rect 237005 3496 273319 3498
rect 237005 3440 237010 3496
rect 237066 3440 273258 3496
rect 273314 3440 273319 3496
rect 237005 3438 273319 3440
rect 237005 3435 237071 3438
rect 273253 3435 273319 3438
rect 427537 3498 427603 3501
rect 580993 3498 581059 3501
rect 427537 3496 581059 3498
rect 427537 3440 427542 3496
rect 427598 3440 580998 3496
rect 581054 3440 581059 3496
rect 427537 3438 581059 3440
rect 427537 3435 427603 3438
rect 580993 3435 581059 3438
rect 6453 3362 6519 3365
rect 169937 3362 170003 3365
rect 6453 3360 170003 3362
rect 6453 3304 6458 3360
rect 6514 3304 169942 3360
rect 169998 3304 170003 3360
rect 6453 3302 170003 3304
rect 6453 3299 6519 3302
rect 169937 3299 170003 3302
rect 234613 3362 234679 3365
rect 271873 3362 271939 3365
rect 234613 3360 271939 3362
rect 234613 3304 234618 3360
rect 234674 3304 271878 3360
rect 271934 3304 271939 3360
rect 234613 3302 271939 3304
rect 234613 3299 234679 3302
rect 271873 3299 271939 3302
rect 427721 3362 427787 3365
rect 583385 3362 583451 3365
rect 427721 3360 583451 3362
rect 427721 3304 427726 3360
rect 427782 3304 583390 3360
rect 583446 3304 583451 3360
rect 427721 3302 583451 3304
rect 427721 3299 427787 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 3372 697308 3436 697372
rect 3372 495484 3436 495548
rect 429700 342484 429764 342548
rect 429700 19348 429764 19412
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 680254 -7976 710862
rect -8576 680018 -8394 680254
rect -8158 680018 -7976 680254
rect -8576 679934 -7976 680018
rect -8576 679698 -8394 679934
rect -8158 679698 -7976 679934
rect -8576 644254 -7976 679698
rect -8576 644018 -8394 644254
rect -8158 644018 -7976 644254
rect -8576 643934 -7976 644018
rect -8576 643698 -8394 643934
rect -8158 643698 -7976 643934
rect -8576 608254 -7976 643698
rect -8576 608018 -8394 608254
rect -8158 608018 -7976 608254
rect -8576 607934 -7976 608018
rect -8576 607698 -8394 607934
rect -8158 607698 -7976 607934
rect -8576 572254 -7976 607698
rect -8576 572018 -8394 572254
rect -8158 572018 -7976 572254
rect -8576 571934 -7976 572018
rect -8576 571698 -8394 571934
rect -8158 571698 -7976 571934
rect -8576 536254 -7976 571698
rect -8576 536018 -8394 536254
rect -8158 536018 -7976 536254
rect -8576 535934 -7976 536018
rect -8576 535698 -8394 535934
rect -8158 535698 -7976 535934
rect -8576 500254 -7976 535698
rect -8576 500018 -8394 500254
rect -8158 500018 -7976 500254
rect -8576 499934 -7976 500018
rect -8576 499698 -8394 499934
rect -8158 499698 -7976 499934
rect -8576 464254 -7976 499698
rect -8576 464018 -8394 464254
rect -8158 464018 -7976 464254
rect -8576 463934 -7976 464018
rect -8576 463698 -8394 463934
rect -8158 463698 -7976 463934
rect -8576 428254 -7976 463698
rect -8576 428018 -8394 428254
rect -8158 428018 -7976 428254
rect -8576 427934 -7976 428018
rect -8576 427698 -8394 427934
rect -8158 427698 -7976 427934
rect -8576 392254 -7976 427698
rect -8576 392018 -8394 392254
rect -8158 392018 -7976 392254
rect -8576 391934 -7976 392018
rect -8576 391698 -8394 391934
rect -8158 391698 -7976 391934
rect -8576 356254 -7976 391698
rect -8576 356018 -8394 356254
rect -8158 356018 -7976 356254
rect -8576 355934 -7976 356018
rect -8576 355698 -8394 355934
rect -8158 355698 -7976 355934
rect -8576 320254 -7976 355698
rect -8576 320018 -8394 320254
rect -8158 320018 -7976 320254
rect -8576 319934 -7976 320018
rect -8576 319698 -8394 319934
rect -8158 319698 -7976 319934
rect -8576 284254 -7976 319698
rect -8576 284018 -8394 284254
rect -8158 284018 -7976 284254
rect -8576 283934 -7976 284018
rect -8576 283698 -8394 283934
rect -8158 283698 -7976 283934
rect -8576 248254 -7976 283698
rect -8576 248018 -8394 248254
rect -8158 248018 -7976 248254
rect -8576 247934 -7976 248018
rect -8576 247698 -8394 247934
rect -8158 247698 -7976 247934
rect -8576 212254 -7976 247698
rect -8576 212018 -8394 212254
rect -8158 212018 -7976 212254
rect -8576 211934 -7976 212018
rect -8576 211698 -8394 211934
rect -8158 211698 -7976 211934
rect -8576 176254 -7976 211698
rect -8576 176018 -8394 176254
rect -8158 176018 -7976 176254
rect -8576 175934 -7976 176018
rect -8576 175698 -8394 175934
rect -8158 175698 -7976 175934
rect -8576 140254 -7976 175698
rect -8576 140018 -8394 140254
rect -8158 140018 -7976 140254
rect -8576 139934 -7976 140018
rect -8576 139698 -8394 139934
rect -8158 139698 -7976 139934
rect -8576 104254 -7976 139698
rect -8576 104018 -8394 104254
rect -8158 104018 -7976 104254
rect -8576 103934 -7976 104018
rect -8576 103698 -8394 103934
rect -8158 103698 -7976 103934
rect -8576 68254 -7976 103698
rect -8576 68018 -8394 68254
rect -8158 68018 -7976 68254
rect -8576 67934 -7976 68018
rect -8576 67698 -8394 67934
rect -8158 67698 -7976 67934
rect -8576 32254 -7976 67698
rect -8576 32018 -8394 32254
rect -8158 32018 -7976 32254
rect -8576 31934 -7976 32018
rect -8576 31698 -8394 31934
rect -8158 31698 -7976 31934
rect -8576 -6926 -7976 31698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 698254 -7036 709922
rect 12604 710478 13204 711440
rect 12604 710242 12786 710478
rect 13022 710242 13204 710478
rect 12604 710158 13204 710242
rect 12604 709922 12786 710158
rect 13022 709922 13204 710158
rect -7636 698018 -7454 698254
rect -7218 698018 -7036 698254
rect -7636 697934 -7036 698018
rect -7636 697698 -7454 697934
rect -7218 697698 -7036 697934
rect -7636 662254 -7036 697698
rect -7636 662018 -7454 662254
rect -7218 662018 -7036 662254
rect -7636 661934 -7036 662018
rect -7636 661698 -7454 661934
rect -7218 661698 -7036 661934
rect -7636 626254 -7036 661698
rect -7636 626018 -7454 626254
rect -7218 626018 -7036 626254
rect -7636 625934 -7036 626018
rect -7636 625698 -7454 625934
rect -7218 625698 -7036 625934
rect -7636 590254 -7036 625698
rect -7636 590018 -7454 590254
rect -7218 590018 -7036 590254
rect -7636 589934 -7036 590018
rect -7636 589698 -7454 589934
rect -7218 589698 -7036 589934
rect -7636 554254 -7036 589698
rect -7636 554018 -7454 554254
rect -7218 554018 -7036 554254
rect -7636 553934 -7036 554018
rect -7636 553698 -7454 553934
rect -7218 553698 -7036 553934
rect -7636 518254 -7036 553698
rect -7636 518018 -7454 518254
rect -7218 518018 -7036 518254
rect -7636 517934 -7036 518018
rect -7636 517698 -7454 517934
rect -7218 517698 -7036 517934
rect -7636 482254 -7036 517698
rect -7636 482018 -7454 482254
rect -7218 482018 -7036 482254
rect -7636 481934 -7036 482018
rect -7636 481698 -7454 481934
rect -7218 481698 -7036 481934
rect -7636 446254 -7036 481698
rect -7636 446018 -7454 446254
rect -7218 446018 -7036 446254
rect -7636 445934 -7036 446018
rect -7636 445698 -7454 445934
rect -7218 445698 -7036 445934
rect -7636 410254 -7036 445698
rect -7636 410018 -7454 410254
rect -7218 410018 -7036 410254
rect -7636 409934 -7036 410018
rect -7636 409698 -7454 409934
rect -7218 409698 -7036 409934
rect -7636 374254 -7036 409698
rect -7636 374018 -7454 374254
rect -7218 374018 -7036 374254
rect -7636 373934 -7036 374018
rect -7636 373698 -7454 373934
rect -7218 373698 -7036 373934
rect -7636 338254 -7036 373698
rect -7636 338018 -7454 338254
rect -7218 338018 -7036 338254
rect -7636 337934 -7036 338018
rect -7636 337698 -7454 337934
rect -7218 337698 -7036 337934
rect -7636 302254 -7036 337698
rect -7636 302018 -7454 302254
rect -7218 302018 -7036 302254
rect -7636 301934 -7036 302018
rect -7636 301698 -7454 301934
rect -7218 301698 -7036 301934
rect -7636 266254 -7036 301698
rect -7636 266018 -7454 266254
rect -7218 266018 -7036 266254
rect -7636 265934 -7036 266018
rect -7636 265698 -7454 265934
rect -7218 265698 -7036 265934
rect -7636 230254 -7036 265698
rect -7636 230018 -7454 230254
rect -7218 230018 -7036 230254
rect -7636 229934 -7036 230018
rect -7636 229698 -7454 229934
rect -7218 229698 -7036 229934
rect -7636 194254 -7036 229698
rect -7636 194018 -7454 194254
rect -7218 194018 -7036 194254
rect -7636 193934 -7036 194018
rect -7636 193698 -7454 193934
rect -7218 193698 -7036 193934
rect -7636 158254 -7036 193698
rect -7636 158018 -7454 158254
rect -7218 158018 -7036 158254
rect -7636 157934 -7036 158018
rect -7636 157698 -7454 157934
rect -7218 157698 -7036 157934
rect -7636 122254 -7036 157698
rect -7636 122018 -7454 122254
rect -7218 122018 -7036 122254
rect -7636 121934 -7036 122018
rect -7636 121698 -7454 121934
rect -7218 121698 -7036 121934
rect -7636 86254 -7036 121698
rect -7636 86018 -7454 86254
rect -7218 86018 -7036 86254
rect -7636 85934 -7036 86018
rect -7636 85698 -7454 85934
rect -7218 85698 -7036 85934
rect -7636 50254 -7036 85698
rect -7636 50018 -7454 50254
rect -7218 50018 -7036 50254
rect -7636 49934 -7036 50018
rect -7636 49698 -7454 49934
rect -7218 49698 -7036 49934
rect -7636 14254 -7036 49698
rect -7636 14018 -7454 14254
rect -7218 14018 -7036 14254
rect -7636 13934 -7036 14018
rect -7636 13698 -7454 13934
rect -7218 13698 -7036 13934
rect -7636 -5986 -7036 13698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 676654 -6096 708982
rect -6696 676418 -6514 676654
rect -6278 676418 -6096 676654
rect -6696 676334 -6096 676418
rect -6696 676098 -6514 676334
rect -6278 676098 -6096 676334
rect -6696 640654 -6096 676098
rect -6696 640418 -6514 640654
rect -6278 640418 -6096 640654
rect -6696 640334 -6096 640418
rect -6696 640098 -6514 640334
rect -6278 640098 -6096 640334
rect -6696 604654 -6096 640098
rect -6696 604418 -6514 604654
rect -6278 604418 -6096 604654
rect -6696 604334 -6096 604418
rect -6696 604098 -6514 604334
rect -6278 604098 -6096 604334
rect -6696 568654 -6096 604098
rect -6696 568418 -6514 568654
rect -6278 568418 -6096 568654
rect -6696 568334 -6096 568418
rect -6696 568098 -6514 568334
rect -6278 568098 -6096 568334
rect -6696 532654 -6096 568098
rect -6696 532418 -6514 532654
rect -6278 532418 -6096 532654
rect -6696 532334 -6096 532418
rect -6696 532098 -6514 532334
rect -6278 532098 -6096 532334
rect -6696 496654 -6096 532098
rect -6696 496418 -6514 496654
rect -6278 496418 -6096 496654
rect -6696 496334 -6096 496418
rect -6696 496098 -6514 496334
rect -6278 496098 -6096 496334
rect -6696 460654 -6096 496098
rect -6696 460418 -6514 460654
rect -6278 460418 -6096 460654
rect -6696 460334 -6096 460418
rect -6696 460098 -6514 460334
rect -6278 460098 -6096 460334
rect -6696 424654 -6096 460098
rect -6696 424418 -6514 424654
rect -6278 424418 -6096 424654
rect -6696 424334 -6096 424418
rect -6696 424098 -6514 424334
rect -6278 424098 -6096 424334
rect -6696 388654 -6096 424098
rect -6696 388418 -6514 388654
rect -6278 388418 -6096 388654
rect -6696 388334 -6096 388418
rect -6696 388098 -6514 388334
rect -6278 388098 -6096 388334
rect -6696 352654 -6096 388098
rect -6696 352418 -6514 352654
rect -6278 352418 -6096 352654
rect -6696 352334 -6096 352418
rect -6696 352098 -6514 352334
rect -6278 352098 -6096 352334
rect -6696 316654 -6096 352098
rect -6696 316418 -6514 316654
rect -6278 316418 -6096 316654
rect -6696 316334 -6096 316418
rect -6696 316098 -6514 316334
rect -6278 316098 -6096 316334
rect -6696 280654 -6096 316098
rect -6696 280418 -6514 280654
rect -6278 280418 -6096 280654
rect -6696 280334 -6096 280418
rect -6696 280098 -6514 280334
rect -6278 280098 -6096 280334
rect -6696 244654 -6096 280098
rect -6696 244418 -6514 244654
rect -6278 244418 -6096 244654
rect -6696 244334 -6096 244418
rect -6696 244098 -6514 244334
rect -6278 244098 -6096 244334
rect -6696 208654 -6096 244098
rect -6696 208418 -6514 208654
rect -6278 208418 -6096 208654
rect -6696 208334 -6096 208418
rect -6696 208098 -6514 208334
rect -6278 208098 -6096 208334
rect -6696 172654 -6096 208098
rect -6696 172418 -6514 172654
rect -6278 172418 -6096 172654
rect -6696 172334 -6096 172418
rect -6696 172098 -6514 172334
rect -6278 172098 -6096 172334
rect -6696 136654 -6096 172098
rect -6696 136418 -6514 136654
rect -6278 136418 -6096 136654
rect -6696 136334 -6096 136418
rect -6696 136098 -6514 136334
rect -6278 136098 -6096 136334
rect -6696 100654 -6096 136098
rect -6696 100418 -6514 100654
rect -6278 100418 -6096 100654
rect -6696 100334 -6096 100418
rect -6696 100098 -6514 100334
rect -6278 100098 -6096 100334
rect -6696 64654 -6096 100098
rect -6696 64418 -6514 64654
rect -6278 64418 -6096 64654
rect -6696 64334 -6096 64418
rect -6696 64098 -6514 64334
rect -6278 64098 -6096 64334
rect -6696 28654 -6096 64098
rect -6696 28418 -6514 28654
rect -6278 28418 -6096 28654
rect -6696 28334 -6096 28418
rect -6696 28098 -6514 28334
rect -6278 28098 -6096 28334
rect -6696 -5046 -6096 28098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 694654 -5156 708042
rect 9004 708598 9604 709560
rect 9004 708362 9186 708598
rect 9422 708362 9604 708598
rect 9004 708278 9604 708362
rect 9004 708042 9186 708278
rect 9422 708042 9604 708278
rect -5756 694418 -5574 694654
rect -5338 694418 -5156 694654
rect -5756 694334 -5156 694418
rect -5756 694098 -5574 694334
rect -5338 694098 -5156 694334
rect -5756 658654 -5156 694098
rect -5756 658418 -5574 658654
rect -5338 658418 -5156 658654
rect -5756 658334 -5156 658418
rect -5756 658098 -5574 658334
rect -5338 658098 -5156 658334
rect -5756 622654 -5156 658098
rect -5756 622418 -5574 622654
rect -5338 622418 -5156 622654
rect -5756 622334 -5156 622418
rect -5756 622098 -5574 622334
rect -5338 622098 -5156 622334
rect -5756 586654 -5156 622098
rect -5756 586418 -5574 586654
rect -5338 586418 -5156 586654
rect -5756 586334 -5156 586418
rect -5756 586098 -5574 586334
rect -5338 586098 -5156 586334
rect -5756 550654 -5156 586098
rect -5756 550418 -5574 550654
rect -5338 550418 -5156 550654
rect -5756 550334 -5156 550418
rect -5756 550098 -5574 550334
rect -5338 550098 -5156 550334
rect -5756 514654 -5156 550098
rect -5756 514418 -5574 514654
rect -5338 514418 -5156 514654
rect -5756 514334 -5156 514418
rect -5756 514098 -5574 514334
rect -5338 514098 -5156 514334
rect -5756 478654 -5156 514098
rect -5756 478418 -5574 478654
rect -5338 478418 -5156 478654
rect -5756 478334 -5156 478418
rect -5756 478098 -5574 478334
rect -5338 478098 -5156 478334
rect -5756 442654 -5156 478098
rect -5756 442418 -5574 442654
rect -5338 442418 -5156 442654
rect -5756 442334 -5156 442418
rect -5756 442098 -5574 442334
rect -5338 442098 -5156 442334
rect -5756 406654 -5156 442098
rect -5756 406418 -5574 406654
rect -5338 406418 -5156 406654
rect -5756 406334 -5156 406418
rect -5756 406098 -5574 406334
rect -5338 406098 -5156 406334
rect -5756 370654 -5156 406098
rect -5756 370418 -5574 370654
rect -5338 370418 -5156 370654
rect -5756 370334 -5156 370418
rect -5756 370098 -5574 370334
rect -5338 370098 -5156 370334
rect -5756 334654 -5156 370098
rect -5756 334418 -5574 334654
rect -5338 334418 -5156 334654
rect -5756 334334 -5156 334418
rect -5756 334098 -5574 334334
rect -5338 334098 -5156 334334
rect -5756 298654 -5156 334098
rect -5756 298418 -5574 298654
rect -5338 298418 -5156 298654
rect -5756 298334 -5156 298418
rect -5756 298098 -5574 298334
rect -5338 298098 -5156 298334
rect -5756 262654 -5156 298098
rect -5756 262418 -5574 262654
rect -5338 262418 -5156 262654
rect -5756 262334 -5156 262418
rect -5756 262098 -5574 262334
rect -5338 262098 -5156 262334
rect -5756 226654 -5156 262098
rect -5756 226418 -5574 226654
rect -5338 226418 -5156 226654
rect -5756 226334 -5156 226418
rect -5756 226098 -5574 226334
rect -5338 226098 -5156 226334
rect -5756 190654 -5156 226098
rect -5756 190418 -5574 190654
rect -5338 190418 -5156 190654
rect -5756 190334 -5156 190418
rect -5756 190098 -5574 190334
rect -5338 190098 -5156 190334
rect -5756 154654 -5156 190098
rect -5756 154418 -5574 154654
rect -5338 154418 -5156 154654
rect -5756 154334 -5156 154418
rect -5756 154098 -5574 154334
rect -5338 154098 -5156 154334
rect -5756 118654 -5156 154098
rect -5756 118418 -5574 118654
rect -5338 118418 -5156 118654
rect -5756 118334 -5156 118418
rect -5756 118098 -5574 118334
rect -5338 118098 -5156 118334
rect -5756 82654 -5156 118098
rect -5756 82418 -5574 82654
rect -5338 82418 -5156 82654
rect -5756 82334 -5156 82418
rect -5756 82098 -5574 82334
rect -5338 82098 -5156 82334
rect -5756 46654 -5156 82098
rect -5756 46418 -5574 46654
rect -5338 46418 -5156 46654
rect -5756 46334 -5156 46418
rect -5756 46098 -5574 46334
rect -5338 46098 -5156 46334
rect -5756 10654 -5156 46098
rect -5756 10418 -5574 10654
rect -5338 10418 -5156 10654
rect -5756 10334 -5156 10418
rect -5756 10098 -5574 10334
rect -5338 10098 -5156 10334
rect -5756 -4106 -5156 10098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 673054 -4216 707102
rect -4816 672818 -4634 673054
rect -4398 672818 -4216 673054
rect -4816 672734 -4216 672818
rect -4816 672498 -4634 672734
rect -4398 672498 -4216 672734
rect -4816 637054 -4216 672498
rect -4816 636818 -4634 637054
rect -4398 636818 -4216 637054
rect -4816 636734 -4216 636818
rect -4816 636498 -4634 636734
rect -4398 636498 -4216 636734
rect -4816 601054 -4216 636498
rect -4816 600818 -4634 601054
rect -4398 600818 -4216 601054
rect -4816 600734 -4216 600818
rect -4816 600498 -4634 600734
rect -4398 600498 -4216 600734
rect -4816 565054 -4216 600498
rect -4816 564818 -4634 565054
rect -4398 564818 -4216 565054
rect -4816 564734 -4216 564818
rect -4816 564498 -4634 564734
rect -4398 564498 -4216 564734
rect -4816 529054 -4216 564498
rect -4816 528818 -4634 529054
rect -4398 528818 -4216 529054
rect -4816 528734 -4216 528818
rect -4816 528498 -4634 528734
rect -4398 528498 -4216 528734
rect -4816 493054 -4216 528498
rect -4816 492818 -4634 493054
rect -4398 492818 -4216 493054
rect -4816 492734 -4216 492818
rect -4816 492498 -4634 492734
rect -4398 492498 -4216 492734
rect -4816 457054 -4216 492498
rect -4816 456818 -4634 457054
rect -4398 456818 -4216 457054
rect -4816 456734 -4216 456818
rect -4816 456498 -4634 456734
rect -4398 456498 -4216 456734
rect -4816 421054 -4216 456498
rect -4816 420818 -4634 421054
rect -4398 420818 -4216 421054
rect -4816 420734 -4216 420818
rect -4816 420498 -4634 420734
rect -4398 420498 -4216 420734
rect -4816 385054 -4216 420498
rect -4816 384818 -4634 385054
rect -4398 384818 -4216 385054
rect -4816 384734 -4216 384818
rect -4816 384498 -4634 384734
rect -4398 384498 -4216 384734
rect -4816 349054 -4216 384498
rect -4816 348818 -4634 349054
rect -4398 348818 -4216 349054
rect -4816 348734 -4216 348818
rect -4816 348498 -4634 348734
rect -4398 348498 -4216 348734
rect -4816 313054 -4216 348498
rect -4816 312818 -4634 313054
rect -4398 312818 -4216 313054
rect -4816 312734 -4216 312818
rect -4816 312498 -4634 312734
rect -4398 312498 -4216 312734
rect -4816 277054 -4216 312498
rect -4816 276818 -4634 277054
rect -4398 276818 -4216 277054
rect -4816 276734 -4216 276818
rect -4816 276498 -4634 276734
rect -4398 276498 -4216 276734
rect -4816 241054 -4216 276498
rect -4816 240818 -4634 241054
rect -4398 240818 -4216 241054
rect -4816 240734 -4216 240818
rect -4816 240498 -4634 240734
rect -4398 240498 -4216 240734
rect -4816 205054 -4216 240498
rect -4816 204818 -4634 205054
rect -4398 204818 -4216 205054
rect -4816 204734 -4216 204818
rect -4816 204498 -4634 204734
rect -4398 204498 -4216 204734
rect -4816 169054 -4216 204498
rect -4816 168818 -4634 169054
rect -4398 168818 -4216 169054
rect -4816 168734 -4216 168818
rect -4816 168498 -4634 168734
rect -4398 168498 -4216 168734
rect -4816 133054 -4216 168498
rect -4816 132818 -4634 133054
rect -4398 132818 -4216 133054
rect -4816 132734 -4216 132818
rect -4816 132498 -4634 132734
rect -4398 132498 -4216 132734
rect -4816 97054 -4216 132498
rect -4816 96818 -4634 97054
rect -4398 96818 -4216 97054
rect -4816 96734 -4216 96818
rect -4816 96498 -4634 96734
rect -4398 96498 -4216 96734
rect -4816 61054 -4216 96498
rect -4816 60818 -4634 61054
rect -4398 60818 -4216 61054
rect -4816 60734 -4216 60818
rect -4816 60498 -4634 60734
rect -4398 60498 -4216 60734
rect -4816 25054 -4216 60498
rect -4816 24818 -4634 25054
rect -4398 24818 -4216 25054
rect -4816 24734 -4216 24818
rect -4816 24498 -4634 24734
rect -4398 24498 -4216 24734
rect -4816 -3166 -4216 24498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 691054 -3276 706162
rect 5404 706718 6004 707680
rect 5404 706482 5586 706718
rect 5822 706482 6004 706718
rect 5404 706398 6004 706482
rect 5404 706162 5586 706398
rect 5822 706162 6004 706398
rect -3876 690818 -3694 691054
rect -3458 690818 -3276 691054
rect -3876 690734 -3276 690818
rect -3876 690498 -3694 690734
rect -3458 690498 -3276 690734
rect -3876 655054 -3276 690498
rect -3876 654818 -3694 655054
rect -3458 654818 -3276 655054
rect -3876 654734 -3276 654818
rect -3876 654498 -3694 654734
rect -3458 654498 -3276 654734
rect -3876 619054 -3276 654498
rect -3876 618818 -3694 619054
rect -3458 618818 -3276 619054
rect -3876 618734 -3276 618818
rect -3876 618498 -3694 618734
rect -3458 618498 -3276 618734
rect -3876 583054 -3276 618498
rect -3876 582818 -3694 583054
rect -3458 582818 -3276 583054
rect -3876 582734 -3276 582818
rect -3876 582498 -3694 582734
rect -3458 582498 -3276 582734
rect -3876 547054 -3276 582498
rect -3876 546818 -3694 547054
rect -3458 546818 -3276 547054
rect -3876 546734 -3276 546818
rect -3876 546498 -3694 546734
rect -3458 546498 -3276 546734
rect -3876 511054 -3276 546498
rect -3876 510818 -3694 511054
rect -3458 510818 -3276 511054
rect -3876 510734 -3276 510818
rect -3876 510498 -3694 510734
rect -3458 510498 -3276 510734
rect -3876 475054 -3276 510498
rect -3876 474818 -3694 475054
rect -3458 474818 -3276 475054
rect -3876 474734 -3276 474818
rect -3876 474498 -3694 474734
rect -3458 474498 -3276 474734
rect -3876 439054 -3276 474498
rect -3876 438818 -3694 439054
rect -3458 438818 -3276 439054
rect -3876 438734 -3276 438818
rect -3876 438498 -3694 438734
rect -3458 438498 -3276 438734
rect -3876 403054 -3276 438498
rect -3876 402818 -3694 403054
rect -3458 402818 -3276 403054
rect -3876 402734 -3276 402818
rect -3876 402498 -3694 402734
rect -3458 402498 -3276 402734
rect -3876 367054 -3276 402498
rect -3876 366818 -3694 367054
rect -3458 366818 -3276 367054
rect -3876 366734 -3276 366818
rect -3876 366498 -3694 366734
rect -3458 366498 -3276 366734
rect -3876 331054 -3276 366498
rect -3876 330818 -3694 331054
rect -3458 330818 -3276 331054
rect -3876 330734 -3276 330818
rect -3876 330498 -3694 330734
rect -3458 330498 -3276 330734
rect -3876 295054 -3276 330498
rect -3876 294818 -3694 295054
rect -3458 294818 -3276 295054
rect -3876 294734 -3276 294818
rect -3876 294498 -3694 294734
rect -3458 294498 -3276 294734
rect -3876 259054 -3276 294498
rect -3876 258818 -3694 259054
rect -3458 258818 -3276 259054
rect -3876 258734 -3276 258818
rect -3876 258498 -3694 258734
rect -3458 258498 -3276 258734
rect -3876 223054 -3276 258498
rect -3876 222818 -3694 223054
rect -3458 222818 -3276 223054
rect -3876 222734 -3276 222818
rect -3876 222498 -3694 222734
rect -3458 222498 -3276 222734
rect -3876 187054 -3276 222498
rect -3876 186818 -3694 187054
rect -3458 186818 -3276 187054
rect -3876 186734 -3276 186818
rect -3876 186498 -3694 186734
rect -3458 186498 -3276 186734
rect -3876 151054 -3276 186498
rect -3876 150818 -3694 151054
rect -3458 150818 -3276 151054
rect -3876 150734 -3276 150818
rect -3876 150498 -3694 150734
rect -3458 150498 -3276 150734
rect -3876 115054 -3276 150498
rect -3876 114818 -3694 115054
rect -3458 114818 -3276 115054
rect -3876 114734 -3276 114818
rect -3876 114498 -3694 114734
rect -3458 114498 -3276 114734
rect -3876 79054 -3276 114498
rect -3876 78818 -3694 79054
rect -3458 78818 -3276 79054
rect -3876 78734 -3276 78818
rect -3876 78498 -3694 78734
rect -3458 78498 -3276 78734
rect -3876 43054 -3276 78498
rect -3876 42818 -3694 43054
rect -3458 42818 -3276 43054
rect -3876 42734 -3276 42818
rect -3876 42498 -3694 42734
rect -3458 42498 -3276 42734
rect -3876 7054 -3276 42498
rect -3876 6818 -3694 7054
rect -3458 6818 -3276 7054
rect -3876 6734 -3276 6818
rect -3876 6498 -3694 6734
rect -3458 6498 -3276 6734
rect -3876 -2226 -3276 6498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 669454 -2336 705222
rect -2936 669218 -2754 669454
rect -2518 669218 -2336 669454
rect -2936 669134 -2336 669218
rect -2936 668898 -2754 669134
rect -2518 668898 -2336 669134
rect -2936 633454 -2336 668898
rect -2936 633218 -2754 633454
rect -2518 633218 -2336 633454
rect -2936 633134 -2336 633218
rect -2936 632898 -2754 633134
rect -2518 632898 -2336 633134
rect -2936 597454 -2336 632898
rect -2936 597218 -2754 597454
rect -2518 597218 -2336 597454
rect -2936 597134 -2336 597218
rect -2936 596898 -2754 597134
rect -2518 596898 -2336 597134
rect -2936 561454 -2336 596898
rect -2936 561218 -2754 561454
rect -2518 561218 -2336 561454
rect -2936 561134 -2336 561218
rect -2936 560898 -2754 561134
rect -2518 560898 -2336 561134
rect -2936 525454 -2336 560898
rect -2936 525218 -2754 525454
rect -2518 525218 -2336 525454
rect -2936 525134 -2336 525218
rect -2936 524898 -2754 525134
rect -2518 524898 -2336 525134
rect -2936 489454 -2336 524898
rect -2936 489218 -2754 489454
rect -2518 489218 -2336 489454
rect -2936 489134 -2336 489218
rect -2936 488898 -2754 489134
rect -2518 488898 -2336 489134
rect -2936 453454 -2336 488898
rect -2936 453218 -2754 453454
rect -2518 453218 -2336 453454
rect -2936 453134 -2336 453218
rect -2936 452898 -2754 453134
rect -2518 452898 -2336 453134
rect -2936 417454 -2336 452898
rect -2936 417218 -2754 417454
rect -2518 417218 -2336 417454
rect -2936 417134 -2336 417218
rect -2936 416898 -2754 417134
rect -2518 416898 -2336 417134
rect -2936 381454 -2336 416898
rect -2936 381218 -2754 381454
rect -2518 381218 -2336 381454
rect -2936 381134 -2336 381218
rect -2936 380898 -2754 381134
rect -2518 380898 -2336 381134
rect -2936 345454 -2336 380898
rect -2936 345218 -2754 345454
rect -2518 345218 -2336 345454
rect -2936 345134 -2336 345218
rect -2936 344898 -2754 345134
rect -2518 344898 -2336 345134
rect -2936 309454 -2336 344898
rect -2936 309218 -2754 309454
rect -2518 309218 -2336 309454
rect -2936 309134 -2336 309218
rect -2936 308898 -2754 309134
rect -2518 308898 -2336 309134
rect -2936 273454 -2336 308898
rect -2936 273218 -2754 273454
rect -2518 273218 -2336 273454
rect -2936 273134 -2336 273218
rect -2936 272898 -2754 273134
rect -2518 272898 -2336 273134
rect -2936 237454 -2336 272898
rect -2936 237218 -2754 237454
rect -2518 237218 -2336 237454
rect -2936 237134 -2336 237218
rect -2936 236898 -2754 237134
rect -2518 236898 -2336 237134
rect -2936 201454 -2336 236898
rect -2936 201218 -2754 201454
rect -2518 201218 -2336 201454
rect -2936 201134 -2336 201218
rect -2936 200898 -2754 201134
rect -2518 200898 -2336 201134
rect -2936 165454 -2336 200898
rect -2936 165218 -2754 165454
rect -2518 165218 -2336 165454
rect -2936 165134 -2336 165218
rect -2936 164898 -2754 165134
rect -2518 164898 -2336 165134
rect -2936 129454 -2336 164898
rect -2936 129218 -2754 129454
rect -2518 129218 -2336 129454
rect -2936 129134 -2336 129218
rect -2936 128898 -2754 129134
rect -2518 128898 -2336 129134
rect -2936 93454 -2336 128898
rect -2936 93218 -2754 93454
rect -2518 93218 -2336 93454
rect -2936 93134 -2336 93218
rect -2936 92898 -2754 93134
rect -2518 92898 -2336 93134
rect -2936 57454 -2336 92898
rect -2936 57218 -2754 57454
rect -2518 57218 -2336 57454
rect -2936 57134 -2336 57218
rect -2936 56898 -2754 57134
rect -2518 56898 -2336 57134
rect -2936 21454 -2336 56898
rect -2936 21218 -2754 21454
rect -2518 21218 -2336 21454
rect -2936 21134 -2336 21218
rect -2936 20898 -2754 21134
rect -2518 20898 -2336 21134
rect -2936 -1286 -2336 20898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 687454 -1396 704282
rect -1996 687218 -1814 687454
rect -1578 687218 -1396 687454
rect -1996 687134 -1396 687218
rect -1996 686898 -1814 687134
rect -1578 686898 -1396 687134
rect -1996 651454 -1396 686898
rect -1996 651218 -1814 651454
rect -1578 651218 -1396 651454
rect -1996 651134 -1396 651218
rect -1996 650898 -1814 651134
rect -1578 650898 -1396 651134
rect -1996 615454 -1396 650898
rect -1996 615218 -1814 615454
rect -1578 615218 -1396 615454
rect -1996 615134 -1396 615218
rect -1996 614898 -1814 615134
rect -1578 614898 -1396 615134
rect -1996 579454 -1396 614898
rect -1996 579218 -1814 579454
rect -1578 579218 -1396 579454
rect -1996 579134 -1396 579218
rect -1996 578898 -1814 579134
rect -1578 578898 -1396 579134
rect -1996 543454 -1396 578898
rect -1996 543218 -1814 543454
rect -1578 543218 -1396 543454
rect -1996 543134 -1396 543218
rect -1996 542898 -1814 543134
rect -1578 542898 -1396 543134
rect -1996 507454 -1396 542898
rect -1996 507218 -1814 507454
rect -1578 507218 -1396 507454
rect -1996 507134 -1396 507218
rect -1996 506898 -1814 507134
rect -1578 506898 -1396 507134
rect -1996 471454 -1396 506898
rect -1996 471218 -1814 471454
rect -1578 471218 -1396 471454
rect -1996 471134 -1396 471218
rect -1996 470898 -1814 471134
rect -1578 470898 -1396 471134
rect -1996 435454 -1396 470898
rect -1996 435218 -1814 435454
rect -1578 435218 -1396 435454
rect -1996 435134 -1396 435218
rect -1996 434898 -1814 435134
rect -1578 434898 -1396 435134
rect -1996 399454 -1396 434898
rect -1996 399218 -1814 399454
rect -1578 399218 -1396 399454
rect -1996 399134 -1396 399218
rect -1996 398898 -1814 399134
rect -1578 398898 -1396 399134
rect -1996 363454 -1396 398898
rect -1996 363218 -1814 363454
rect -1578 363218 -1396 363454
rect -1996 363134 -1396 363218
rect -1996 362898 -1814 363134
rect -1578 362898 -1396 363134
rect -1996 327454 -1396 362898
rect -1996 327218 -1814 327454
rect -1578 327218 -1396 327454
rect -1996 327134 -1396 327218
rect -1996 326898 -1814 327134
rect -1578 326898 -1396 327134
rect -1996 291454 -1396 326898
rect -1996 291218 -1814 291454
rect -1578 291218 -1396 291454
rect -1996 291134 -1396 291218
rect -1996 290898 -1814 291134
rect -1578 290898 -1396 291134
rect -1996 255454 -1396 290898
rect -1996 255218 -1814 255454
rect -1578 255218 -1396 255454
rect -1996 255134 -1396 255218
rect -1996 254898 -1814 255134
rect -1578 254898 -1396 255134
rect -1996 219454 -1396 254898
rect -1996 219218 -1814 219454
rect -1578 219218 -1396 219454
rect -1996 219134 -1396 219218
rect -1996 218898 -1814 219134
rect -1578 218898 -1396 219134
rect -1996 183454 -1396 218898
rect -1996 183218 -1814 183454
rect -1578 183218 -1396 183454
rect -1996 183134 -1396 183218
rect -1996 182898 -1814 183134
rect -1578 182898 -1396 183134
rect -1996 147454 -1396 182898
rect -1996 147218 -1814 147454
rect -1578 147218 -1396 147454
rect -1996 147134 -1396 147218
rect -1996 146898 -1814 147134
rect -1578 146898 -1396 147134
rect -1996 111454 -1396 146898
rect -1996 111218 -1814 111454
rect -1578 111218 -1396 111454
rect -1996 111134 -1396 111218
rect -1996 110898 -1814 111134
rect -1578 110898 -1396 111134
rect -1996 75454 -1396 110898
rect -1996 75218 -1814 75454
rect -1578 75218 -1396 75454
rect -1996 75134 -1396 75218
rect -1996 74898 -1814 75134
rect -1578 74898 -1396 75134
rect -1996 39454 -1396 74898
rect -1996 39218 -1814 39454
rect -1578 39218 -1396 39454
rect -1996 39134 -1396 39218
rect -1996 38898 -1814 39134
rect -1578 38898 -1396 39134
rect -1996 3454 -1396 38898
rect -1996 3218 -1814 3454
rect -1578 3218 -1396 3454
rect -1996 3134 -1396 3218
rect -1996 2898 -1814 3134
rect -1578 2898 -1396 3134
rect -1996 -346 -1396 2898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 1804 704838 2404 705800
rect 1804 704602 1986 704838
rect 2222 704602 2404 704838
rect 1804 704518 2404 704602
rect 1804 704282 1986 704518
rect 2222 704282 2404 704518
rect 1804 687454 2404 704282
rect 3371 697372 3437 697373
rect 3371 697308 3372 697372
rect 3436 697308 3437 697372
rect 3371 697307 3437 697308
rect 1804 687218 1986 687454
rect 2222 687218 2404 687454
rect 1804 687134 2404 687218
rect 1804 686898 1986 687134
rect 2222 686898 2404 687134
rect 1804 651454 2404 686898
rect 1804 651218 1986 651454
rect 2222 651218 2404 651454
rect 1804 651134 2404 651218
rect 1804 650898 1986 651134
rect 2222 650898 2404 651134
rect 1804 615454 2404 650898
rect 1804 615218 1986 615454
rect 2222 615218 2404 615454
rect 1804 615134 2404 615218
rect 1804 614898 1986 615134
rect 2222 614898 2404 615134
rect 1804 579454 2404 614898
rect 1804 579218 1986 579454
rect 2222 579218 2404 579454
rect 1804 579134 2404 579218
rect 1804 578898 1986 579134
rect 2222 578898 2404 579134
rect 1804 543454 2404 578898
rect 1804 543218 1986 543454
rect 2222 543218 2404 543454
rect 1804 543134 2404 543218
rect 1804 542898 1986 543134
rect 2222 542898 2404 543134
rect 1804 507454 2404 542898
rect 1804 507218 1986 507454
rect 2222 507218 2404 507454
rect 1804 507134 2404 507218
rect 1804 506898 1986 507134
rect 2222 506898 2404 507134
rect 1804 471454 2404 506898
rect 3374 495549 3434 697307
rect 5404 691054 6004 706162
rect 5404 690818 5586 691054
rect 5822 690818 6004 691054
rect 5404 690734 6004 690818
rect 5404 690498 5586 690734
rect 5822 690498 6004 690734
rect 5404 655054 6004 690498
rect 5404 654818 5586 655054
rect 5822 654818 6004 655054
rect 5404 654734 6004 654818
rect 5404 654498 5586 654734
rect 5822 654498 6004 654734
rect 5404 619054 6004 654498
rect 5404 618818 5586 619054
rect 5822 618818 6004 619054
rect 5404 618734 6004 618818
rect 5404 618498 5586 618734
rect 5822 618498 6004 618734
rect 5404 583054 6004 618498
rect 5404 582818 5586 583054
rect 5822 582818 6004 583054
rect 5404 582734 6004 582818
rect 5404 582498 5586 582734
rect 5822 582498 6004 582734
rect 5404 547054 6004 582498
rect 5404 546818 5586 547054
rect 5822 546818 6004 547054
rect 5404 546734 6004 546818
rect 5404 546498 5586 546734
rect 5822 546498 6004 546734
rect 5404 511054 6004 546498
rect 5404 510818 5586 511054
rect 5822 510818 6004 511054
rect 5404 510734 6004 510818
rect 5404 510498 5586 510734
rect 5822 510498 6004 510734
rect 3371 495548 3437 495549
rect 3371 495484 3372 495548
rect 3436 495484 3437 495548
rect 3371 495483 3437 495484
rect 1804 471218 1986 471454
rect 2222 471218 2404 471454
rect 1804 471134 2404 471218
rect 1804 470898 1986 471134
rect 2222 470898 2404 471134
rect 1804 435454 2404 470898
rect 1804 435218 1986 435454
rect 2222 435218 2404 435454
rect 1804 435134 2404 435218
rect 1804 434898 1986 435134
rect 2222 434898 2404 435134
rect 1804 399454 2404 434898
rect 1804 399218 1986 399454
rect 2222 399218 2404 399454
rect 1804 399134 2404 399218
rect 1804 398898 1986 399134
rect 2222 398898 2404 399134
rect 1804 363454 2404 398898
rect 1804 363218 1986 363454
rect 2222 363218 2404 363454
rect 1804 363134 2404 363218
rect 1804 362898 1986 363134
rect 2222 362898 2404 363134
rect 1804 327454 2404 362898
rect 1804 327218 1986 327454
rect 2222 327218 2404 327454
rect 1804 327134 2404 327218
rect 1804 326898 1986 327134
rect 2222 326898 2404 327134
rect 1804 291454 2404 326898
rect 1804 291218 1986 291454
rect 2222 291218 2404 291454
rect 1804 291134 2404 291218
rect 1804 290898 1986 291134
rect 2222 290898 2404 291134
rect 1804 255454 2404 290898
rect 1804 255218 1986 255454
rect 2222 255218 2404 255454
rect 1804 255134 2404 255218
rect 1804 254898 1986 255134
rect 2222 254898 2404 255134
rect 1804 219454 2404 254898
rect 1804 219218 1986 219454
rect 2222 219218 2404 219454
rect 1804 219134 2404 219218
rect 1804 218898 1986 219134
rect 2222 218898 2404 219134
rect 1804 183454 2404 218898
rect 1804 183218 1986 183454
rect 2222 183218 2404 183454
rect 1804 183134 2404 183218
rect 1804 182898 1986 183134
rect 2222 182898 2404 183134
rect 1804 147454 2404 182898
rect 1804 147218 1986 147454
rect 2222 147218 2404 147454
rect 1804 147134 2404 147218
rect 1804 146898 1986 147134
rect 2222 146898 2404 147134
rect 1804 111454 2404 146898
rect 1804 111218 1986 111454
rect 2222 111218 2404 111454
rect 1804 111134 2404 111218
rect 1804 110898 1986 111134
rect 2222 110898 2404 111134
rect 1804 75454 2404 110898
rect 1804 75218 1986 75454
rect 2222 75218 2404 75454
rect 1804 75134 2404 75218
rect 1804 74898 1986 75134
rect 2222 74898 2404 75134
rect 1804 39454 2404 74898
rect 1804 39218 1986 39454
rect 2222 39218 2404 39454
rect 1804 39134 2404 39218
rect 1804 38898 1986 39134
rect 2222 38898 2404 39134
rect 1804 3454 2404 38898
rect 1804 3218 1986 3454
rect 2222 3218 2404 3454
rect 1804 3134 2404 3218
rect 1804 2898 1986 3134
rect 2222 2898 2404 3134
rect 1804 -346 2404 2898
rect 1804 -582 1986 -346
rect 2222 -582 2404 -346
rect 1804 -666 2404 -582
rect 1804 -902 1986 -666
rect 2222 -902 2404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 1804 -1864 2404 -902
rect 5404 475054 6004 510498
rect 5404 474818 5586 475054
rect 5822 474818 6004 475054
rect 5404 474734 6004 474818
rect 5404 474498 5586 474734
rect 5822 474498 6004 474734
rect 5404 439054 6004 474498
rect 5404 438818 5586 439054
rect 5822 438818 6004 439054
rect 5404 438734 6004 438818
rect 5404 438498 5586 438734
rect 5822 438498 6004 438734
rect 5404 403054 6004 438498
rect 5404 402818 5586 403054
rect 5822 402818 6004 403054
rect 5404 402734 6004 402818
rect 5404 402498 5586 402734
rect 5822 402498 6004 402734
rect 5404 367054 6004 402498
rect 5404 366818 5586 367054
rect 5822 366818 6004 367054
rect 5404 366734 6004 366818
rect 5404 366498 5586 366734
rect 5822 366498 6004 366734
rect 5404 331054 6004 366498
rect 5404 330818 5586 331054
rect 5822 330818 6004 331054
rect 5404 330734 6004 330818
rect 5404 330498 5586 330734
rect 5822 330498 6004 330734
rect 5404 295054 6004 330498
rect 5404 294818 5586 295054
rect 5822 294818 6004 295054
rect 5404 294734 6004 294818
rect 5404 294498 5586 294734
rect 5822 294498 6004 294734
rect 5404 259054 6004 294498
rect 5404 258818 5586 259054
rect 5822 258818 6004 259054
rect 5404 258734 6004 258818
rect 5404 258498 5586 258734
rect 5822 258498 6004 258734
rect 5404 223054 6004 258498
rect 5404 222818 5586 223054
rect 5822 222818 6004 223054
rect 5404 222734 6004 222818
rect 5404 222498 5586 222734
rect 5822 222498 6004 222734
rect 5404 187054 6004 222498
rect 5404 186818 5586 187054
rect 5822 186818 6004 187054
rect 5404 186734 6004 186818
rect 5404 186498 5586 186734
rect 5822 186498 6004 186734
rect 5404 151054 6004 186498
rect 5404 150818 5586 151054
rect 5822 150818 6004 151054
rect 5404 150734 6004 150818
rect 5404 150498 5586 150734
rect 5822 150498 6004 150734
rect 5404 115054 6004 150498
rect 5404 114818 5586 115054
rect 5822 114818 6004 115054
rect 5404 114734 6004 114818
rect 5404 114498 5586 114734
rect 5822 114498 6004 114734
rect 5404 79054 6004 114498
rect 5404 78818 5586 79054
rect 5822 78818 6004 79054
rect 5404 78734 6004 78818
rect 5404 78498 5586 78734
rect 5822 78498 6004 78734
rect 5404 43054 6004 78498
rect 5404 42818 5586 43054
rect 5822 42818 6004 43054
rect 5404 42734 6004 42818
rect 5404 42498 5586 42734
rect 5822 42498 6004 42734
rect 5404 7054 6004 42498
rect 5404 6818 5586 7054
rect 5822 6818 6004 7054
rect 5404 6734 6004 6818
rect 5404 6498 5586 6734
rect 5822 6498 6004 6734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 5404 -2226 6004 6498
rect 5404 -2462 5586 -2226
rect 5822 -2462 6004 -2226
rect 5404 -2546 6004 -2462
rect 5404 -2782 5586 -2546
rect 5822 -2782 6004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 5404 -3744 6004 -2782
rect 9004 694654 9604 708042
rect 9004 694418 9186 694654
rect 9422 694418 9604 694654
rect 9004 694334 9604 694418
rect 9004 694098 9186 694334
rect 9422 694098 9604 694334
rect 9004 658654 9604 694098
rect 9004 658418 9186 658654
rect 9422 658418 9604 658654
rect 9004 658334 9604 658418
rect 9004 658098 9186 658334
rect 9422 658098 9604 658334
rect 9004 622654 9604 658098
rect 9004 622418 9186 622654
rect 9422 622418 9604 622654
rect 9004 622334 9604 622418
rect 9004 622098 9186 622334
rect 9422 622098 9604 622334
rect 9004 586654 9604 622098
rect 9004 586418 9186 586654
rect 9422 586418 9604 586654
rect 9004 586334 9604 586418
rect 9004 586098 9186 586334
rect 9422 586098 9604 586334
rect 9004 550654 9604 586098
rect 9004 550418 9186 550654
rect 9422 550418 9604 550654
rect 9004 550334 9604 550418
rect 9004 550098 9186 550334
rect 9422 550098 9604 550334
rect 9004 514654 9604 550098
rect 9004 514418 9186 514654
rect 9422 514418 9604 514654
rect 9004 514334 9604 514418
rect 9004 514098 9186 514334
rect 9422 514098 9604 514334
rect 9004 478654 9604 514098
rect 9004 478418 9186 478654
rect 9422 478418 9604 478654
rect 9004 478334 9604 478418
rect 9004 478098 9186 478334
rect 9422 478098 9604 478334
rect 9004 442654 9604 478098
rect 9004 442418 9186 442654
rect 9422 442418 9604 442654
rect 9004 442334 9604 442418
rect 9004 442098 9186 442334
rect 9422 442098 9604 442334
rect 9004 406654 9604 442098
rect 9004 406418 9186 406654
rect 9422 406418 9604 406654
rect 9004 406334 9604 406418
rect 9004 406098 9186 406334
rect 9422 406098 9604 406334
rect 9004 370654 9604 406098
rect 9004 370418 9186 370654
rect 9422 370418 9604 370654
rect 9004 370334 9604 370418
rect 9004 370098 9186 370334
rect 9422 370098 9604 370334
rect 9004 334654 9604 370098
rect 9004 334418 9186 334654
rect 9422 334418 9604 334654
rect 9004 334334 9604 334418
rect 9004 334098 9186 334334
rect 9422 334098 9604 334334
rect 9004 298654 9604 334098
rect 9004 298418 9186 298654
rect 9422 298418 9604 298654
rect 9004 298334 9604 298418
rect 9004 298098 9186 298334
rect 9422 298098 9604 298334
rect 9004 262654 9604 298098
rect 9004 262418 9186 262654
rect 9422 262418 9604 262654
rect 9004 262334 9604 262418
rect 9004 262098 9186 262334
rect 9422 262098 9604 262334
rect 9004 226654 9604 262098
rect 9004 226418 9186 226654
rect 9422 226418 9604 226654
rect 9004 226334 9604 226418
rect 9004 226098 9186 226334
rect 9422 226098 9604 226334
rect 9004 190654 9604 226098
rect 9004 190418 9186 190654
rect 9422 190418 9604 190654
rect 9004 190334 9604 190418
rect 9004 190098 9186 190334
rect 9422 190098 9604 190334
rect 9004 154654 9604 190098
rect 9004 154418 9186 154654
rect 9422 154418 9604 154654
rect 9004 154334 9604 154418
rect 9004 154098 9186 154334
rect 9422 154098 9604 154334
rect 9004 118654 9604 154098
rect 9004 118418 9186 118654
rect 9422 118418 9604 118654
rect 9004 118334 9604 118418
rect 9004 118098 9186 118334
rect 9422 118098 9604 118334
rect 9004 82654 9604 118098
rect 9004 82418 9186 82654
rect 9422 82418 9604 82654
rect 9004 82334 9604 82418
rect 9004 82098 9186 82334
rect 9422 82098 9604 82334
rect 9004 46654 9604 82098
rect 9004 46418 9186 46654
rect 9422 46418 9604 46654
rect 9004 46334 9604 46418
rect 9004 46098 9186 46334
rect 9422 46098 9604 46334
rect 9004 10654 9604 46098
rect 9004 10418 9186 10654
rect 9422 10418 9604 10654
rect 9004 10334 9604 10418
rect 9004 10098 9186 10334
rect 9422 10098 9604 10334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 9004 -4106 9604 10098
rect 9004 -4342 9186 -4106
rect 9422 -4342 9604 -4106
rect 9004 -4426 9604 -4342
rect 9004 -4662 9186 -4426
rect 9422 -4662 9604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 9004 -5624 9604 -4662
rect 12604 698254 13204 709922
rect 30604 711418 31204 711440
rect 30604 711182 30786 711418
rect 31022 711182 31204 711418
rect 30604 711098 31204 711182
rect 30604 710862 30786 711098
rect 31022 710862 31204 711098
rect 27004 709538 27604 709560
rect 27004 709302 27186 709538
rect 27422 709302 27604 709538
rect 27004 709218 27604 709302
rect 27004 708982 27186 709218
rect 27422 708982 27604 709218
rect 23404 707658 24004 707680
rect 23404 707422 23586 707658
rect 23822 707422 24004 707658
rect 23404 707338 24004 707422
rect 23404 707102 23586 707338
rect 23822 707102 24004 707338
rect 12604 698018 12786 698254
rect 13022 698018 13204 698254
rect 12604 697934 13204 698018
rect 12604 697698 12786 697934
rect 13022 697698 13204 697934
rect 12604 662254 13204 697698
rect 12604 662018 12786 662254
rect 13022 662018 13204 662254
rect 12604 661934 13204 662018
rect 12604 661698 12786 661934
rect 13022 661698 13204 661934
rect 12604 626254 13204 661698
rect 12604 626018 12786 626254
rect 13022 626018 13204 626254
rect 12604 625934 13204 626018
rect 12604 625698 12786 625934
rect 13022 625698 13204 625934
rect 12604 590254 13204 625698
rect 12604 590018 12786 590254
rect 13022 590018 13204 590254
rect 12604 589934 13204 590018
rect 12604 589698 12786 589934
rect 13022 589698 13204 589934
rect 12604 554254 13204 589698
rect 12604 554018 12786 554254
rect 13022 554018 13204 554254
rect 12604 553934 13204 554018
rect 12604 553698 12786 553934
rect 13022 553698 13204 553934
rect 12604 518254 13204 553698
rect 12604 518018 12786 518254
rect 13022 518018 13204 518254
rect 12604 517934 13204 518018
rect 12604 517698 12786 517934
rect 13022 517698 13204 517934
rect 12604 482254 13204 517698
rect 12604 482018 12786 482254
rect 13022 482018 13204 482254
rect 12604 481934 13204 482018
rect 12604 481698 12786 481934
rect 13022 481698 13204 481934
rect 12604 446254 13204 481698
rect 12604 446018 12786 446254
rect 13022 446018 13204 446254
rect 12604 445934 13204 446018
rect 12604 445698 12786 445934
rect 13022 445698 13204 445934
rect 12604 410254 13204 445698
rect 12604 410018 12786 410254
rect 13022 410018 13204 410254
rect 12604 409934 13204 410018
rect 12604 409698 12786 409934
rect 13022 409698 13204 409934
rect 12604 374254 13204 409698
rect 12604 374018 12786 374254
rect 13022 374018 13204 374254
rect 12604 373934 13204 374018
rect 12604 373698 12786 373934
rect 13022 373698 13204 373934
rect 12604 338254 13204 373698
rect 12604 338018 12786 338254
rect 13022 338018 13204 338254
rect 12604 337934 13204 338018
rect 12604 337698 12786 337934
rect 13022 337698 13204 337934
rect 12604 302254 13204 337698
rect 12604 302018 12786 302254
rect 13022 302018 13204 302254
rect 12604 301934 13204 302018
rect 12604 301698 12786 301934
rect 13022 301698 13204 301934
rect 12604 266254 13204 301698
rect 12604 266018 12786 266254
rect 13022 266018 13204 266254
rect 12604 265934 13204 266018
rect 12604 265698 12786 265934
rect 13022 265698 13204 265934
rect 12604 230254 13204 265698
rect 12604 230018 12786 230254
rect 13022 230018 13204 230254
rect 12604 229934 13204 230018
rect 12604 229698 12786 229934
rect 13022 229698 13204 229934
rect 12604 194254 13204 229698
rect 12604 194018 12786 194254
rect 13022 194018 13204 194254
rect 12604 193934 13204 194018
rect 12604 193698 12786 193934
rect 13022 193698 13204 193934
rect 12604 158254 13204 193698
rect 12604 158018 12786 158254
rect 13022 158018 13204 158254
rect 12604 157934 13204 158018
rect 12604 157698 12786 157934
rect 13022 157698 13204 157934
rect 12604 122254 13204 157698
rect 12604 122018 12786 122254
rect 13022 122018 13204 122254
rect 12604 121934 13204 122018
rect 12604 121698 12786 121934
rect 13022 121698 13204 121934
rect 12604 86254 13204 121698
rect 12604 86018 12786 86254
rect 13022 86018 13204 86254
rect 12604 85934 13204 86018
rect 12604 85698 12786 85934
rect 13022 85698 13204 85934
rect 12604 50254 13204 85698
rect 12604 50018 12786 50254
rect 13022 50018 13204 50254
rect 12604 49934 13204 50018
rect 12604 49698 12786 49934
rect 13022 49698 13204 49934
rect 12604 14254 13204 49698
rect 12604 14018 12786 14254
rect 13022 14018 13204 14254
rect 12604 13934 13204 14018
rect 12604 13698 12786 13934
rect 13022 13698 13204 13934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 12604 -5986 13204 13698
rect 19804 705778 20404 705800
rect 19804 705542 19986 705778
rect 20222 705542 20404 705778
rect 19804 705458 20404 705542
rect 19804 705222 19986 705458
rect 20222 705222 20404 705458
rect 19804 669454 20404 705222
rect 19804 669218 19986 669454
rect 20222 669218 20404 669454
rect 19804 669134 20404 669218
rect 19804 668898 19986 669134
rect 20222 668898 20404 669134
rect 19804 633454 20404 668898
rect 19804 633218 19986 633454
rect 20222 633218 20404 633454
rect 19804 633134 20404 633218
rect 19804 632898 19986 633134
rect 20222 632898 20404 633134
rect 19804 597454 20404 632898
rect 19804 597218 19986 597454
rect 20222 597218 20404 597454
rect 19804 597134 20404 597218
rect 19804 596898 19986 597134
rect 20222 596898 20404 597134
rect 19804 561454 20404 596898
rect 19804 561218 19986 561454
rect 20222 561218 20404 561454
rect 19804 561134 20404 561218
rect 19804 560898 19986 561134
rect 20222 560898 20404 561134
rect 19804 525454 20404 560898
rect 19804 525218 19986 525454
rect 20222 525218 20404 525454
rect 19804 525134 20404 525218
rect 19804 524898 19986 525134
rect 20222 524898 20404 525134
rect 19804 489454 20404 524898
rect 19804 489218 19986 489454
rect 20222 489218 20404 489454
rect 19804 489134 20404 489218
rect 19804 488898 19986 489134
rect 20222 488898 20404 489134
rect 19804 453454 20404 488898
rect 19804 453218 19986 453454
rect 20222 453218 20404 453454
rect 19804 453134 20404 453218
rect 19804 452898 19986 453134
rect 20222 452898 20404 453134
rect 19804 417454 20404 452898
rect 19804 417218 19986 417454
rect 20222 417218 20404 417454
rect 19804 417134 20404 417218
rect 19804 416898 19986 417134
rect 20222 416898 20404 417134
rect 19804 381454 20404 416898
rect 19804 381218 19986 381454
rect 20222 381218 20404 381454
rect 19804 381134 20404 381218
rect 19804 380898 19986 381134
rect 20222 380898 20404 381134
rect 19804 345454 20404 380898
rect 19804 345218 19986 345454
rect 20222 345218 20404 345454
rect 19804 345134 20404 345218
rect 19804 344898 19986 345134
rect 20222 344898 20404 345134
rect 19804 309454 20404 344898
rect 19804 309218 19986 309454
rect 20222 309218 20404 309454
rect 19804 309134 20404 309218
rect 19804 308898 19986 309134
rect 20222 308898 20404 309134
rect 19804 273454 20404 308898
rect 19804 273218 19986 273454
rect 20222 273218 20404 273454
rect 19804 273134 20404 273218
rect 19804 272898 19986 273134
rect 20222 272898 20404 273134
rect 19804 237454 20404 272898
rect 19804 237218 19986 237454
rect 20222 237218 20404 237454
rect 19804 237134 20404 237218
rect 19804 236898 19986 237134
rect 20222 236898 20404 237134
rect 19804 201454 20404 236898
rect 19804 201218 19986 201454
rect 20222 201218 20404 201454
rect 19804 201134 20404 201218
rect 19804 200898 19986 201134
rect 20222 200898 20404 201134
rect 19804 165454 20404 200898
rect 19804 165218 19986 165454
rect 20222 165218 20404 165454
rect 19804 165134 20404 165218
rect 19804 164898 19986 165134
rect 20222 164898 20404 165134
rect 19804 129454 20404 164898
rect 19804 129218 19986 129454
rect 20222 129218 20404 129454
rect 19804 129134 20404 129218
rect 19804 128898 19986 129134
rect 20222 128898 20404 129134
rect 19804 93454 20404 128898
rect 19804 93218 19986 93454
rect 20222 93218 20404 93454
rect 19804 93134 20404 93218
rect 19804 92898 19986 93134
rect 20222 92898 20404 93134
rect 19804 57454 20404 92898
rect 19804 57218 19986 57454
rect 20222 57218 20404 57454
rect 19804 57134 20404 57218
rect 19804 56898 19986 57134
rect 20222 56898 20404 57134
rect 19804 21454 20404 56898
rect 19804 21218 19986 21454
rect 20222 21218 20404 21454
rect 19804 21134 20404 21218
rect 19804 20898 19986 21134
rect 20222 20898 20404 21134
rect 19804 -1286 20404 20898
rect 19804 -1522 19986 -1286
rect 20222 -1522 20404 -1286
rect 19804 -1606 20404 -1522
rect 19804 -1842 19986 -1606
rect 20222 -1842 20404 -1606
rect 19804 -1864 20404 -1842
rect 23404 673054 24004 707102
rect 23404 672818 23586 673054
rect 23822 672818 24004 673054
rect 23404 672734 24004 672818
rect 23404 672498 23586 672734
rect 23822 672498 24004 672734
rect 23404 637054 24004 672498
rect 23404 636818 23586 637054
rect 23822 636818 24004 637054
rect 23404 636734 24004 636818
rect 23404 636498 23586 636734
rect 23822 636498 24004 636734
rect 23404 601054 24004 636498
rect 23404 600818 23586 601054
rect 23822 600818 24004 601054
rect 23404 600734 24004 600818
rect 23404 600498 23586 600734
rect 23822 600498 24004 600734
rect 23404 565054 24004 600498
rect 23404 564818 23586 565054
rect 23822 564818 24004 565054
rect 23404 564734 24004 564818
rect 23404 564498 23586 564734
rect 23822 564498 24004 564734
rect 23404 529054 24004 564498
rect 23404 528818 23586 529054
rect 23822 528818 24004 529054
rect 23404 528734 24004 528818
rect 23404 528498 23586 528734
rect 23822 528498 24004 528734
rect 23404 493054 24004 528498
rect 23404 492818 23586 493054
rect 23822 492818 24004 493054
rect 23404 492734 24004 492818
rect 23404 492498 23586 492734
rect 23822 492498 24004 492734
rect 23404 457054 24004 492498
rect 23404 456818 23586 457054
rect 23822 456818 24004 457054
rect 23404 456734 24004 456818
rect 23404 456498 23586 456734
rect 23822 456498 24004 456734
rect 23404 421054 24004 456498
rect 23404 420818 23586 421054
rect 23822 420818 24004 421054
rect 23404 420734 24004 420818
rect 23404 420498 23586 420734
rect 23822 420498 24004 420734
rect 23404 385054 24004 420498
rect 23404 384818 23586 385054
rect 23822 384818 24004 385054
rect 23404 384734 24004 384818
rect 23404 384498 23586 384734
rect 23822 384498 24004 384734
rect 23404 349054 24004 384498
rect 23404 348818 23586 349054
rect 23822 348818 24004 349054
rect 23404 348734 24004 348818
rect 23404 348498 23586 348734
rect 23822 348498 24004 348734
rect 23404 313054 24004 348498
rect 23404 312818 23586 313054
rect 23822 312818 24004 313054
rect 23404 312734 24004 312818
rect 23404 312498 23586 312734
rect 23822 312498 24004 312734
rect 23404 277054 24004 312498
rect 23404 276818 23586 277054
rect 23822 276818 24004 277054
rect 23404 276734 24004 276818
rect 23404 276498 23586 276734
rect 23822 276498 24004 276734
rect 23404 241054 24004 276498
rect 23404 240818 23586 241054
rect 23822 240818 24004 241054
rect 23404 240734 24004 240818
rect 23404 240498 23586 240734
rect 23822 240498 24004 240734
rect 23404 205054 24004 240498
rect 23404 204818 23586 205054
rect 23822 204818 24004 205054
rect 23404 204734 24004 204818
rect 23404 204498 23586 204734
rect 23822 204498 24004 204734
rect 23404 169054 24004 204498
rect 23404 168818 23586 169054
rect 23822 168818 24004 169054
rect 23404 168734 24004 168818
rect 23404 168498 23586 168734
rect 23822 168498 24004 168734
rect 23404 133054 24004 168498
rect 23404 132818 23586 133054
rect 23822 132818 24004 133054
rect 23404 132734 24004 132818
rect 23404 132498 23586 132734
rect 23822 132498 24004 132734
rect 23404 97054 24004 132498
rect 23404 96818 23586 97054
rect 23822 96818 24004 97054
rect 23404 96734 24004 96818
rect 23404 96498 23586 96734
rect 23822 96498 24004 96734
rect 23404 61054 24004 96498
rect 23404 60818 23586 61054
rect 23822 60818 24004 61054
rect 23404 60734 24004 60818
rect 23404 60498 23586 60734
rect 23822 60498 24004 60734
rect 23404 25054 24004 60498
rect 23404 24818 23586 25054
rect 23822 24818 24004 25054
rect 23404 24734 24004 24818
rect 23404 24498 23586 24734
rect 23822 24498 24004 24734
rect 23404 -3166 24004 24498
rect 23404 -3402 23586 -3166
rect 23822 -3402 24004 -3166
rect 23404 -3486 24004 -3402
rect 23404 -3722 23586 -3486
rect 23822 -3722 24004 -3486
rect 23404 -3744 24004 -3722
rect 27004 676654 27604 708982
rect 27004 676418 27186 676654
rect 27422 676418 27604 676654
rect 27004 676334 27604 676418
rect 27004 676098 27186 676334
rect 27422 676098 27604 676334
rect 27004 640654 27604 676098
rect 27004 640418 27186 640654
rect 27422 640418 27604 640654
rect 27004 640334 27604 640418
rect 27004 640098 27186 640334
rect 27422 640098 27604 640334
rect 27004 604654 27604 640098
rect 27004 604418 27186 604654
rect 27422 604418 27604 604654
rect 27004 604334 27604 604418
rect 27004 604098 27186 604334
rect 27422 604098 27604 604334
rect 27004 568654 27604 604098
rect 27004 568418 27186 568654
rect 27422 568418 27604 568654
rect 27004 568334 27604 568418
rect 27004 568098 27186 568334
rect 27422 568098 27604 568334
rect 27004 532654 27604 568098
rect 27004 532418 27186 532654
rect 27422 532418 27604 532654
rect 27004 532334 27604 532418
rect 27004 532098 27186 532334
rect 27422 532098 27604 532334
rect 27004 496654 27604 532098
rect 27004 496418 27186 496654
rect 27422 496418 27604 496654
rect 27004 496334 27604 496418
rect 27004 496098 27186 496334
rect 27422 496098 27604 496334
rect 27004 460654 27604 496098
rect 27004 460418 27186 460654
rect 27422 460418 27604 460654
rect 27004 460334 27604 460418
rect 27004 460098 27186 460334
rect 27422 460098 27604 460334
rect 27004 424654 27604 460098
rect 27004 424418 27186 424654
rect 27422 424418 27604 424654
rect 27004 424334 27604 424418
rect 27004 424098 27186 424334
rect 27422 424098 27604 424334
rect 27004 388654 27604 424098
rect 27004 388418 27186 388654
rect 27422 388418 27604 388654
rect 27004 388334 27604 388418
rect 27004 388098 27186 388334
rect 27422 388098 27604 388334
rect 27004 352654 27604 388098
rect 27004 352418 27186 352654
rect 27422 352418 27604 352654
rect 27004 352334 27604 352418
rect 27004 352098 27186 352334
rect 27422 352098 27604 352334
rect 27004 316654 27604 352098
rect 27004 316418 27186 316654
rect 27422 316418 27604 316654
rect 27004 316334 27604 316418
rect 27004 316098 27186 316334
rect 27422 316098 27604 316334
rect 27004 280654 27604 316098
rect 27004 280418 27186 280654
rect 27422 280418 27604 280654
rect 27004 280334 27604 280418
rect 27004 280098 27186 280334
rect 27422 280098 27604 280334
rect 27004 244654 27604 280098
rect 27004 244418 27186 244654
rect 27422 244418 27604 244654
rect 27004 244334 27604 244418
rect 27004 244098 27186 244334
rect 27422 244098 27604 244334
rect 27004 208654 27604 244098
rect 27004 208418 27186 208654
rect 27422 208418 27604 208654
rect 27004 208334 27604 208418
rect 27004 208098 27186 208334
rect 27422 208098 27604 208334
rect 27004 172654 27604 208098
rect 27004 172418 27186 172654
rect 27422 172418 27604 172654
rect 27004 172334 27604 172418
rect 27004 172098 27186 172334
rect 27422 172098 27604 172334
rect 27004 136654 27604 172098
rect 27004 136418 27186 136654
rect 27422 136418 27604 136654
rect 27004 136334 27604 136418
rect 27004 136098 27186 136334
rect 27422 136098 27604 136334
rect 27004 100654 27604 136098
rect 27004 100418 27186 100654
rect 27422 100418 27604 100654
rect 27004 100334 27604 100418
rect 27004 100098 27186 100334
rect 27422 100098 27604 100334
rect 27004 64654 27604 100098
rect 27004 64418 27186 64654
rect 27422 64418 27604 64654
rect 27004 64334 27604 64418
rect 27004 64098 27186 64334
rect 27422 64098 27604 64334
rect 27004 28654 27604 64098
rect 27004 28418 27186 28654
rect 27422 28418 27604 28654
rect 27004 28334 27604 28418
rect 27004 28098 27186 28334
rect 27422 28098 27604 28334
rect 27004 -5046 27604 28098
rect 27004 -5282 27186 -5046
rect 27422 -5282 27604 -5046
rect 27004 -5366 27604 -5282
rect 27004 -5602 27186 -5366
rect 27422 -5602 27604 -5366
rect 27004 -5624 27604 -5602
rect 30604 680254 31204 710862
rect 48604 710478 49204 711440
rect 48604 710242 48786 710478
rect 49022 710242 49204 710478
rect 48604 710158 49204 710242
rect 48604 709922 48786 710158
rect 49022 709922 49204 710158
rect 45004 708598 45604 709560
rect 45004 708362 45186 708598
rect 45422 708362 45604 708598
rect 45004 708278 45604 708362
rect 45004 708042 45186 708278
rect 45422 708042 45604 708278
rect 41404 706718 42004 707680
rect 41404 706482 41586 706718
rect 41822 706482 42004 706718
rect 41404 706398 42004 706482
rect 41404 706162 41586 706398
rect 41822 706162 42004 706398
rect 30604 680018 30786 680254
rect 31022 680018 31204 680254
rect 30604 679934 31204 680018
rect 30604 679698 30786 679934
rect 31022 679698 31204 679934
rect 30604 644254 31204 679698
rect 30604 644018 30786 644254
rect 31022 644018 31204 644254
rect 30604 643934 31204 644018
rect 30604 643698 30786 643934
rect 31022 643698 31204 643934
rect 30604 608254 31204 643698
rect 30604 608018 30786 608254
rect 31022 608018 31204 608254
rect 30604 607934 31204 608018
rect 30604 607698 30786 607934
rect 31022 607698 31204 607934
rect 30604 572254 31204 607698
rect 30604 572018 30786 572254
rect 31022 572018 31204 572254
rect 30604 571934 31204 572018
rect 30604 571698 30786 571934
rect 31022 571698 31204 571934
rect 30604 536254 31204 571698
rect 30604 536018 30786 536254
rect 31022 536018 31204 536254
rect 30604 535934 31204 536018
rect 30604 535698 30786 535934
rect 31022 535698 31204 535934
rect 30604 500254 31204 535698
rect 30604 500018 30786 500254
rect 31022 500018 31204 500254
rect 30604 499934 31204 500018
rect 30604 499698 30786 499934
rect 31022 499698 31204 499934
rect 30604 464254 31204 499698
rect 30604 464018 30786 464254
rect 31022 464018 31204 464254
rect 30604 463934 31204 464018
rect 30604 463698 30786 463934
rect 31022 463698 31204 463934
rect 30604 428254 31204 463698
rect 30604 428018 30786 428254
rect 31022 428018 31204 428254
rect 30604 427934 31204 428018
rect 30604 427698 30786 427934
rect 31022 427698 31204 427934
rect 30604 392254 31204 427698
rect 30604 392018 30786 392254
rect 31022 392018 31204 392254
rect 30604 391934 31204 392018
rect 30604 391698 30786 391934
rect 31022 391698 31204 391934
rect 30604 356254 31204 391698
rect 30604 356018 30786 356254
rect 31022 356018 31204 356254
rect 30604 355934 31204 356018
rect 30604 355698 30786 355934
rect 31022 355698 31204 355934
rect 30604 320254 31204 355698
rect 30604 320018 30786 320254
rect 31022 320018 31204 320254
rect 30604 319934 31204 320018
rect 30604 319698 30786 319934
rect 31022 319698 31204 319934
rect 30604 284254 31204 319698
rect 30604 284018 30786 284254
rect 31022 284018 31204 284254
rect 30604 283934 31204 284018
rect 30604 283698 30786 283934
rect 31022 283698 31204 283934
rect 30604 248254 31204 283698
rect 30604 248018 30786 248254
rect 31022 248018 31204 248254
rect 30604 247934 31204 248018
rect 30604 247698 30786 247934
rect 31022 247698 31204 247934
rect 30604 212254 31204 247698
rect 30604 212018 30786 212254
rect 31022 212018 31204 212254
rect 30604 211934 31204 212018
rect 30604 211698 30786 211934
rect 31022 211698 31204 211934
rect 30604 176254 31204 211698
rect 30604 176018 30786 176254
rect 31022 176018 31204 176254
rect 30604 175934 31204 176018
rect 30604 175698 30786 175934
rect 31022 175698 31204 175934
rect 30604 140254 31204 175698
rect 30604 140018 30786 140254
rect 31022 140018 31204 140254
rect 30604 139934 31204 140018
rect 30604 139698 30786 139934
rect 31022 139698 31204 139934
rect 30604 104254 31204 139698
rect 30604 104018 30786 104254
rect 31022 104018 31204 104254
rect 30604 103934 31204 104018
rect 30604 103698 30786 103934
rect 31022 103698 31204 103934
rect 30604 68254 31204 103698
rect 30604 68018 30786 68254
rect 31022 68018 31204 68254
rect 30604 67934 31204 68018
rect 30604 67698 30786 67934
rect 31022 67698 31204 67934
rect 30604 32254 31204 67698
rect 30604 32018 30786 32254
rect 31022 32018 31204 32254
rect 30604 31934 31204 32018
rect 30604 31698 30786 31934
rect 31022 31698 31204 31934
rect 12604 -6222 12786 -5986
rect 13022 -6222 13204 -5986
rect 12604 -6306 13204 -6222
rect 12604 -6542 12786 -6306
rect 13022 -6542 13204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 12604 -7504 13204 -6542
rect 30604 -6926 31204 31698
rect 37804 704838 38404 705800
rect 37804 704602 37986 704838
rect 38222 704602 38404 704838
rect 37804 704518 38404 704602
rect 37804 704282 37986 704518
rect 38222 704282 38404 704518
rect 37804 687454 38404 704282
rect 37804 687218 37986 687454
rect 38222 687218 38404 687454
rect 37804 687134 38404 687218
rect 37804 686898 37986 687134
rect 38222 686898 38404 687134
rect 37804 651454 38404 686898
rect 37804 651218 37986 651454
rect 38222 651218 38404 651454
rect 37804 651134 38404 651218
rect 37804 650898 37986 651134
rect 38222 650898 38404 651134
rect 37804 615454 38404 650898
rect 37804 615218 37986 615454
rect 38222 615218 38404 615454
rect 37804 615134 38404 615218
rect 37804 614898 37986 615134
rect 38222 614898 38404 615134
rect 37804 579454 38404 614898
rect 37804 579218 37986 579454
rect 38222 579218 38404 579454
rect 37804 579134 38404 579218
rect 37804 578898 37986 579134
rect 38222 578898 38404 579134
rect 37804 543454 38404 578898
rect 37804 543218 37986 543454
rect 38222 543218 38404 543454
rect 37804 543134 38404 543218
rect 37804 542898 37986 543134
rect 38222 542898 38404 543134
rect 37804 507454 38404 542898
rect 37804 507218 37986 507454
rect 38222 507218 38404 507454
rect 37804 507134 38404 507218
rect 37804 506898 37986 507134
rect 38222 506898 38404 507134
rect 37804 471454 38404 506898
rect 37804 471218 37986 471454
rect 38222 471218 38404 471454
rect 37804 471134 38404 471218
rect 37804 470898 37986 471134
rect 38222 470898 38404 471134
rect 37804 435454 38404 470898
rect 37804 435218 37986 435454
rect 38222 435218 38404 435454
rect 37804 435134 38404 435218
rect 37804 434898 37986 435134
rect 38222 434898 38404 435134
rect 37804 399454 38404 434898
rect 37804 399218 37986 399454
rect 38222 399218 38404 399454
rect 37804 399134 38404 399218
rect 37804 398898 37986 399134
rect 38222 398898 38404 399134
rect 37804 363454 38404 398898
rect 37804 363218 37986 363454
rect 38222 363218 38404 363454
rect 37804 363134 38404 363218
rect 37804 362898 37986 363134
rect 38222 362898 38404 363134
rect 37804 327454 38404 362898
rect 37804 327218 37986 327454
rect 38222 327218 38404 327454
rect 37804 327134 38404 327218
rect 37804 326898 37986 327134
rect 38222 326898 38404 327134
rect 37804 291454 38404 326898
rect 37804 291218 37986 291454
rect 38222 291218 38404 291454
rect 37804 291134 38404 291218
rect 37804 290898 37986 291134
rect 38222 290898 38404 291134
rect 37804 255454 38404 290898
rect 37804 255218 37986 255454
rect 38222 255218 38404 255454
rect 37804 255134 38404 255218
rect 37804 254898 37986 255134
rect 38222 254898 38404 255134
rect 37804 219454 38404 254898
rect 37804 219218 37986 219454
rect 38222 219218 38404 219454
rect 37804 219134 38404 219218
rect 37804 218898 37986 219134
rect 38222 218898 38404 219134
rect 37804 183454 38404 218898
rect 37804 183218 37986 183454
rect 38222 183218 38404 183454
rect 37804 183134 38404 183218
rect 37804 182898 37986 183134
rect 38222 182898 38404 183134
rect 37804 147454 38404 182898
rect 37804 147218 37986 147454
rect 38222 147218 38404 147454
rect 37804 147134 38404 147218
rect 37804 146898 37986 147134
rect 38222 146898 38404 147134
rect 37804 111454 38404 146898
rect 37804 111218 37986 111454
rect 38222 111218 38404 111454
rect 37804 111134 38404 111218
rect 37804 110898 37986 111134
rect 38222 110898 38404 111134
rect 37804 75454 38404 110898
rect 37804 75218 37986 75454
rect 38222 75218 38404 75454
rect 37804 75134 38404 75218
rect 37804 74898 37986 75134
rect 38222 74898 38404 75134
rect 37804 39454 38404 74898
rect 37804 39218 37986 39454
rect 38222 39218 38404 39454
rect 37804 39134 38404 39218
rect 37804 38898 37986 39134
rect 38222 38898 38404 39134
rect 37804 3454 38404 38898
rect 37804 3218 37986 3454
rect 38222 3218 38404 3454
rect 37804 3134 38404 3218
rect 37804 2898 37986 3134
rect 38222 2898 38404 3134
rect 37804 -346 38404 2898
rect 37804 -582 37986 -346
rect 38222 -582 38404 -346
rect 37804 -666 38404 -582
rect 37804 -902 37986 -666
rect 38222 -902 38404 -666
rect 37804 -1864 38404 -902
rect 41404 691054 42004 706162
rect 41404 690818 41586 691054
rect 41822 690818 42004 691054
rect 41404 690734 42004 690818
rect 41404 690498 41586 690734
rect 41822 690498 42004 690734
rect 41404 655054 42004 690498
rect 41404 654818 41586 655054
rect 41822 654818 42004 655054
rect 41404 654734 42004 654818
rect 41404 654498 41586 654734
rect 41822 654498 42004 654734
rect 41404 619054 42004 654498
rect 41404 618818 41586 619054
rect 41822 618818 42004 619054
rect 41404 618734 42004 618818
rect 41404 618498 41586 618734
rect 41822 618498 42004 618734
rect 41404 583054 42004 618498
rect 41404 582818 41586 583054
rect 41822 582818 42004 583054
rect 41404 582734 42004 582818
rect 41404 582498 41586 582734
rect 41822 582498 42004 582734
rect 41404 547054 42004 582498
rect 41404 546818 41586 547054
rect 41822 546818 42004 547054
rect 41404 546734 42004 546818
rect 41404 546498 41586 546734
rect 41822 546498 42004 546734
rect 41404 511054 42004 546498
rect 41404 510818 41586 511054
rect 41822 510818 42004 511054
rect 41404 510734 42004 510818
rect 41404 510498 41586 510734
rect 41822 510498 42004 510734
rect 41404 475054 42004 510498
rect 41404 474818 41586 475054
rect 41822 474818 42004 475054
rect 41404 474734 42004 474818
rect 41404 474498 41586 474734
rect 41822 474498 42004 474734
rect 41404 439054 42004 474498
rect 41404 438818 41586 439054
rect 41822 438818 42004 439054
rect 41404 438734 42004 438818
rect 41404 438498 41586 438734
rect 41822 438498 42004 438734
rect 41404 403054 42004 438498
rect 41404 402818 41586 403054
rect 41822 402818 42004 403054
rect 41404 402734 42004 402818
rect 41404 402498 41586 402734
rect 41822 402498 42004 402734
rect 41404 367054 42004 402498
rect 41404 366818 41586 367054
rect 41822 366818 42004 367054
rect 41404 366734 42004 366818
rect 41404 366498 41586 366734
rect 41822 366498 42004 366734
rect 41404 331054 42004 366498
rect 41404 330818 41586 331054
rect 41822 330818 42004 331054
rect 41404 330734 42004 330818
rect 41404 330498 41586 330734
rect 41822 330498 42004 330734
rect 41404 295054 42004 330498
rect 41404 294818 41586 295054
rect 41822 294818 42004 295054
rect 41404 294734 42004 294818
rect 41404 294498 41586 294734
rect 41822 294498 42004 294734
rect 41404 259054 42004 294498
rect 41404 258818 41586 259054
rect 41822 258818 42004 259054
rect 41404 258734 42004 258818
rect 41404 258498 41586 258734
rect 41822 258498 42004 258734
rect 41404 223054 42004 258498
rect 41404 222818 41586 223054
rect 41822 222818 42004 223054
rect 41404 222734 42004 222818
rect 41404 222498 41586 222734
rect 41822 222498 42004 222734
rect 41404 187054 42004 222498
rect 41404 186818 41586 187054
rect 41822 186818 42004 187054
rect 41404 186734 42004 186818
rect 41404 186498 41586 186734
rect 41822 186498 42004 186734
rect 41404 151054 42004 186498
rect 41404 150818 41586 151054
rect 41822 150818 42004 151054
rect 41404 150734 42004 150818
rect 41404 150498 41586 150734
rect 41822 150498 42004 150734
rect 41404 115054 42004 150498
rect 41404 114818 41586 115054
rect 41822 114818 42004 115054
rect 41404 114734 42004 114818
rect 41404 114498 41586 114734
rect 41822 114498 42004 114734
rect 41404 79054 42004 114498
rect 41404 78818 41586 79054
rect 41822 78818 42004 79054
rect 41404 78734 42004 78818
rect 41404 78498 41586 78734
rect 41822 78498 42004 78734
rect 41404 43054 42004 78498
rect 41404 42818 41586 43054
rect 41822 42818 42004 43054
rect 41404 42734 42004 42818
rect 41404 42498 41586 42734
rect 41822 42498 42004 42734
rect 41404 7054 42004 42498
rect 41404 6818 41586 7054
rect 41822 6818 42004 7054
rect 41404 6734 42004 6818
rect 41404 6498 41586 6734
rect 41822 6498 42004 6734
rect 41404 -2226 42004 6498
rect 41404 -2462 41586 -2226
rect 41822 -2462 42004 -2226
rect 41404 -2546 42004 -2462
rect 41404 -2782 41586 -2546
rect 41822 -2782 42004 -2546
rect 41404 -3744 42004 -2782
rect 45004 694654 45604 708042
rect 45004 694418 45186 694654
rect 45422 694418 45604 694654
rect 45004 694334 45604 694418
rect 45004 694098 45186 694334
rect 45422 694098 45604 694334
rect 45004 658654 45604 694098
rect 45004 658418 45186 658654
rect 45422 658418 45604 658654
rect 45004 658334 45604 658418
rect 45004 658098 45186 658334
rect 45422 658098 45604 658334
rect 45004 622654 45604 658098
rect 45004 622418 45186 622654
rect 45422 622418 45604 622654
rect 45004 622334 45604 622418
rect 45004 622098 45186 622334
rect 45422 622098 45604 622334
rect 45004 586654 45604 622098
rect 45004 586418 45186 586654
rect 45422 586418 45604 586654
rect 45004 586334 45604 586418
rect 45004 586098 45186 586334
rect 45422 586098 45604 586334
rect 45004 550654 45604 586098
rect 45004 550418 45186 550654
rect 45422 550418 45604 550654
rect 45004 550334 45604 550418
rect 45004 550098 45186 550334
rect 45422 550098 45604 550334
rect 45004 514654 45604 550098
rect 45004 514418 45186 514654
rect 45422 514418 45604 514654
rect 45004 514334 45604 514418
rect 45004 514098 45186 514334
rect 45422 514098 45604 514334
rect 45004 478654 45604 514098
rect 45004 478418 45186 478654
rect 45422 478418 45604 478654
rect 45004 478334 45604 478418
rect 45004 478098 45186 478334
rect 45422 478098 45604 478334
rect 45004 442654 45604 478098
rect 45004 442418 45186 442654
rect 45422 442418 45604 442654
rect 45004 442334 45604 442418
rect 45004 442098 45186 442334
rect 45422 442098 45604 442334
rect 45004 406654 45604 442098
rect 45004 406418 45186 406654
rect 45422 406418 45604 406654
rect 45004 406334 45604 406418
rect 45004 406098 45186 406334
rect 45422 406098 45604 406334
rect 45004 370654 45604 406098
rect 45004 370418 45186 370654
rect 45422 370418 45604 370654
rect 45004 370334 45604 370418
rect 45004 370098 45186 370334
rect 45422 370098 45604 370334
rect 45004 334654 45604 370098
rect 45004 334418 45186 334654
rect 45422 334418 45604 334654
rect 45004 334334 45604 334418
rect 45004 334098 45186 334334
rect 45422 334098 45604 334334
rect 45004 298654 45604 334098
rect 45004 298418 45186 298654
rect 45422 298418 45604 298654
rect 45004 298334 45604 298418
rect 45004 298098 45186 298334
rect 45422 298098 45604 298334
rect 45004 262654 45604 298098
rect 45004 262418 45186 262654
rect 45422 262418 45604 262654
rect 45004 262334 45604 262418
rect 45004 262098 45186 262334
rect 45422 262098 45604 262334
rect 45004 226654 45604 262098
rect 45004 226418 45186 226654
rect 45422 226418 45604 226654
rect 45004 226334 45604 226418
rect 45004 226098 45186 226334
rect 45422 226098 45604 226334
rect 45004 190654 45604 226098
rect 45004 190418 45186 190654
rect 45422 190418 45604 190654
rect 45004 190334 45604 190418
rect 45004 190098 45186 190334
rect 45422 190098 45604 190334
rect 45004 154654 45604 190098
rect 45004 154418 45186 154654
rect 45422 154418 45604 154654
rect 45004 154334 45604 154418
rect 45004 154098 45186 154334
rect 45422 154098 45604 154334
rect 45004 118654 45604 154098
rect 45004 118418 45186 118654
rect 45422 118418 45604 118654
rect 45004 118334 45604 118418
rect 45004 118098 45186 118334
rect 45422 118098 45604 118334
rect 45004 82654 45604 118098
rect 45004 82418 45186 82654
rect 45422 82418 45604 82654
rect 45004 82334 45604 82418
rect 45004 82098 45186 82334
rect 45422 82098 45604 82334
rect 45004 46654 45604 82098
rect 45004 46418 45186 46654
rect 45422 46418 45604 46654
rect 45004 46334 45604 46418
rect 45004 46098 45186 46334
rect 45422 46098 45604 46334
rect 45004 10654 45604 46098
rect 45004 10418 45186 10654
rect 45422 10418 45604 10654
rect 45004 10334 45604 10418
rect 45004 10098 45186 10334
rect 45422 10098 45604 10334
rect 45004 -4106 45604 10098
rect 45004 -4342 45186 -4106
rect 45422 -4342 45604 -4106
rect 45004 -4426 45604 -4342
rect 45004 -4662 45186 -4426
rect 45422 -4662 45604 -4426
rect 45004 -5624 45604 -4662
rect 48604 698254 49204 709922
rect 66604 711418 67204 711440
rect 66604 711182 66786 711418
rect 67022 711182 67204 711418
rect 66604 711098 67204 711182
rect 66604 710862 66786 711098
rect 67022 710862 67204 711098
rect 63004 709538 63604 709560
rect 63004 709302 63186 709538
rect 63422 709302 63604 709538
rect 63004 709218 63604 709302
rect 63004 708982 63186 709218
rect 63422 708982 63604 709218
rect 59404 707658 60004 707680
rect 59404 707422 59586 707658
rect 59822 707422 60004 707658
rect 59404 707338 60004 707422
rect 59404 707102 59586 707338
rect 59822 707102 60004 707338
rect 48604 698018 48786 698254
rect 49022 698018 49204 698254
rect 48604 697934 49204 698018
rect 48604 697698 48786 697934
rect 49022 697698 49204 697934
rect 48604 662254 49204 697698
rect 48604 662018 48786 662254
rect 49022 662018 49204 662254
rect 48604 661934 49204 662018
rect 48604 661698 48786 661934
rect 49022 661698 49204 661934
rect 48604 626254 49204 661698
rect 48604 626018 48786 626254
rect 49022 626018 49204 626254
rect 48604 625934 49204 626018
rect 48604 625698 48786 625934
rect 49022 625698 49204 625934
rect 48604 590254 49204 625698
rect 48604 590018 48786 590254
rect 49022 590018 49204 590254
rect 48604 589934 49204 590018
rect 48604 589698 48786 589934
rect 49022 589698 49204 589934
rect 48604 554254 49204 589698
rect 48604 554018 48786 554254
rect 49022 554018 49204 554254
rect 48604 553934 49204 554018
rect 48604 553698 48786 553934
rect 49022 553698 49204 553934
rect 48604 518254 49204 553698
rect 48604 518018 48786 518254
rect 49022 518018 49204 518254
rect 48604 517934 49204 518018
rect 48604 517698 48786 517934
rect 49022 517698 49204 517934
rect 48604 482254 49204 517698
rect 48604 482018 48786 482254
rect 49022 482018 49204 482254
rect 48604 481934 49204 482018
rect 48604 481698 48786 481934
rect 49022 481698 49204 481934
rect 48604 446254 49204 481698
rect 48604 446018 48786 446254
rect 49022 446018 49204 446254
rect 48604 445934 49204 446018
rect 48604 445698 48786 445934
rect 49022 445698 49204 445934
rect 48604 410254 49204 445698
rect 48604 410018 48786 410254
rect 49022 410018 49204 410254
rect 48604 409934 49204 410018
rect 48604 409698 48786 409934
rect 49022 409698 49204 409934
rect 48604 374254 49204 409698
rect 48604 374018 48786 374254
rect 49022 374018 49204 374254
rect 48604 373934 49204 374018
rect 48604 373698 48786 373934
rect 49022 373698 49204 373934
rect 48604 338254 49204 373698
rect 48604 338018 48786 338254
rect 49022 338018 49204 338254
rect 48604 337934 49204 338018
rect 48604 337698 48786 337934
rect 49022 337698 49204 337934
rect 48604 302254 49204 337698
rect 48604 302018 48786 302254
rect 49022 302018 49204 302254
rect 48604 301934 49204 302018
rect 48604 301698 48786 301934
rect 49022 301698 49204 301934
rect 48604 266254 49204 301698
rect 48604 266018 48786 266254
rect 49022 266018 49204 266254
rect 48604 265934 49204 266018
rect 48604 265698 48786 265934
rect 49022 265698 49204 265934
rect 48604 230254 49204 265698
rect 48604 230018 48786 230254
rect 49022 230018 49204 230254
rect 48604 229934 49204 230018
rect 48604 229698 48786 229934
rect 49022 229698 49204 229934
rect 48604 194254 49204 229698
rect 48604 194018 48786 194254
rect 49022 194018 49204 194254
rect 48604 193934 49204 194018
rect 48604 193698 48786 193934
rect 49022 193698 49204 193934
rect 48604 158254 49204 193698
rect 48604 158018 48786 158254
rect 49022 158018 49204 158254
rect 48604 157934 49204 158018
rect 48604 157698 48786 157934
rect 49022 157698 49204 157934
rect 48604 122254 49204 157698
rect 48604 122018 48786 122254
rect 49022 122018 49204 122254
rect 48604 121934 49204 122018
rect 48604 121698 48786 121934
rect 49022 121698 49204 121934
rect 48604 86254 49204 121698
rect 48604 86018 48786 86254
rect 49022 86018 49204 86254
rect 48604 85934 49204 86018
rect 48604 85698 48786 85934
rect 49022 85698 49204 85934
rect 48604 50254 49204 85698
rect 48604 50018 48786 50254
rect 49022 50018 49204 50254
rect 48604 49934 49204 50018
rect 48604 49698 48786 49934
rect 49022 49698 49204 49934
rect 48604 14254 49204 49698
rect 48604 14018 48786 14254
rect 49022 14018 49204 14254
rect 48604 13934 49204 14018
rect 48604 13698 48786 13934
rect 49022 13698 49204 13934
rect 30604 -7162 30786 -6926
rect 31022 -7162 31204 -6926
rect 30604 -7246 31204 -7162
rect 30604 -7482 30786 -7246
rect 31022 -7482 31204 -7246
rect 30604 -7504 31204 -7482
rect 48604 -5986 49204 13698
rect 55804 705778 56404 705800
rect 55804 705542 55986 705778
rect 56222 705542 56404 705778
rect 55804 705458 56404 705542
rect 55804 705222 55986 705458
rect 56222 705222 56404 705458
rect 55804 669454 56404 705222
rect 55804 669218 55986 669454
rect 56222 669218 56404 669454
rect 55804 669134 56404 669218
rect 55804 668898 55986 669134
rect 56222 668898 56404 669134
rect 55804 633454 56404 668898
rect 55804 633218 55986 633454
rect 56222 633218 56404 633454
rect 55804 633134 56404 633218
rect 55804 632898 55986 633134
rect 56222 632898 56404 633134
rect 55804 597454 56404 632898
rect 55804 597218 55986 597454
rect 56222 597218 56404 597454
rect 55804 597134 56404 597218
rect 55804 596898 55986 597134
rect 56222 596898 56404 597134
rect 55804 561454 56404 596898
rect 55804 561218 55986 561454
rect 56222 561218 56404 561454
rect 55804 561134 56404 561218
rect 55804 560898 55986 561134
rect 56222 560898 56404 561134
rect 55804 525454 56404 560898
rect 55804 525218 55986 525454
rect 56222 525218 56404 525454
rect 55804 525134 56404 525218
rect 55804 524898 55986 525134
rect 56222 524898 56404 525134
rect 55804 489454 56404 524898
rect 55804 489218 55986 489454
rect 56222 489218 56404 489454
rect 55804 489134 56404 489218
rect 55804 488898 55986 489134
rect 56222 488898 56404 489134
rect 55804 453454 56404 488898
rect 55804 453218 55986 453454
rect 56222 453218 56404 453454
rect 55804 453134 56404 453218
rect 55804 452898 55986 453134
rect 56222 452898 56404 453134
rect 55804 417454 56404 452898
rect 55804 417218 55986 417454
rect 56222 417218 56404 417454
rect 55804 417134 56404 417218
rect 55804 416898 55986 417134
rect 56222 416898 56404 417134
rect 55804 381454 56404 416898
rect 55804 381218 55986 381454
rect 56222 381218 56404 381454
rect 55804 381134 56404 381218
rect 55804 380898 55986 381134
rect 56222 380898 56404 381134
rect 55804 345454 56404 380898
rect 55804 345218 55986 345454
rect 56222 345218 56404 345454
rect 55804 345134 56404 345218
rect 55804 344898 55986 345134
rect 56222 344898 56404 345134
rect 55804 309454 56404 344898
rect 55804 309218 55986 309454
rect 56222 309218 56404 309454
rect 55804 309134 56404 309218
rect 55804 308898 55986 309134
rect 56222 308898 56404 309134
rect 55804 273454 56404 308898
rect 55804 273218 55986 273454
rect 56222 273218 56404 273454
rect 55804 273134 56404 273218
rect 55804 272898 55986 273134
rect 56222 272898 56404 273134
rect 55804 237454 56404 272898
rect 55804 237218 55986 237454
rect 56222 237218 56404 237454
rect 55804 237134 56404 237218
rect 55804 236898 55986 237134
rect 56222 236898 56404 237134
rect 55804 201454 56404 236898
rect 55804 201218 55986 201454
rect 56222 201218 56404 201454
rect 55804 201134 56404 201218
rect 55804 200898 55986 201134
rect 56222 200898 56404 201134
rect 55804 165454 56404 200898
rect 55804 165218 55986 165454
rect 56222 165218 56404 165454
rect 55804 165134 56404 165218
rect 55804 164898 55986 165134
rect 56222 164898 56404 165134
rect 55804 129454 56404 164898
rect 55804 129218 55986 129454
rect 56222 129218 56404 129454
rect 55804 129134 56404 129218
rect 55804 128898 55986 129134
rect 56222 128898 56404 129134
rect 55804 93454 56404 128898
rect 55804 93218 55986 93454
rect 56222 93218 56404 93454
rect 55804 93134 56404 93218
rect 55804 92898 55986 93134
rect 56222 92898 56404 93134
rect 55804 57454 56404 92898
rect 55804 57218 55986 57454
rect 56222 57218 56404 57454
rect 55804 57134 56404 57218
rect 55804 56898 55986 57134
rect 56222 56898 56404 57134
rect 55804 21454 56404 56898
rect 55804 21218 55986 21454
rect 56222 21218 56404 21454
rect 55804 21134 56404 21218
rect 55804 20898 55986 21134
rect 56222 20898 56404 21134
rect 55804 -1286 56404 20898
rect 55804 -1522 55986 -1286
rect 56222 -1522 56404 -1286
rect 55804 -1606 56404 -1522
rect 55804 -1842 55986 -1606
rect 56222 -1842 56404 -1606
rect 55804 -1864 56404 -1842
rect 59404 673054 60004 707102
rect 59404 672818 59586 673054
rect 59822 672818 60004 673054
rect 59404 672734 60004 672818
rect 59404 672498 59586 672734
rect 59822 672498 60004 672734
rect 59404 637054 60004 672498
rect 59404 636818 59586 637054
rect 59822 636818 60004 637054
rect 59404 636734 60004 636818
rect 59404 636498 59586 636734
rect 59822 636498 60004 636734
rect 59404 601054 60004 636498
rect 59404 600818 59586 601054
rect 59822 600818 60004 601054
rect 59404 600734 60004 600818
rect 59404 600498 59586 600734
rect 59822 600498 60004 600734
rect 59404 565054 60004 600498
rect 59404 564818 59586 565054
rect 59822 564818 60004 565054
rect 59404 564734 60004 564818
rect 59404 564498 59586 564734
rect 59822 564498 60004 564734
rect 59404 529054 60004 564498
rect 59404 528818 59586 529054
rect 59822 528818 60004 529054
rect 59404 528734 60004 528818
rect 59404 528498 59586 528734
rect 59822 528498 60004 528734
rect 59404 493054 60004 528498
rect 59404 492818 59586 493054
rect 59822 492818 60004 493054
rect 59404 492734 60004 492818
rect 59404 492498 59586 492734
rect 59822 492498 60004 492734
rect 59404 457054 60004 492498
rect 59404 456818 59586 457054
rect 59822 456818 60004 457054
rect 59404 456734 60004 456818
rect 59404 456498 59586 456734
rect 59822 456498 60004 456734
rect 59404 421054 60004 456498
rect 59404 420818 59586 421054
rect 59822 420818 60004 421054
rect 59404 420734 60004 420818
rect 59404 420498 59586 420734
rect 59822 420498 60004 420734
rect 59404 385054 60004 420498
rect 59404 384818 59586 385054
rect 59822 384818 60004 385054
rect 59404 384734 60004 384818
rect 59404 384498 59586 384734
rect 59822 384498 60004 384734
rect 59404 349054 60004 384498
rect 59404 348818 59586 349054
rect 59822 348818 60004 349054
rect 59404 348734 60004 348818
rect 59404 348498 59586 348734
rect 59822 348498 60004 348734
rect 59404 313054 60004 348498
rect 59404 312818 59586 313054
rect 59822 312818 60004 313054
rect 59404 312734 60004 312818
rect 59404 312498 59586 312734
rect 59822 312498 60004 312734
rect 59404 277054 60004 312498
rect 59404 276818 59586 277054
rect 59822 276818 60004 277054
rect 59404 276734 60004 276818
rect 59404 276498 59586 276734
rect 59822 276498 60004 276734
rect 59404 241054 60004 276498
rect 59404 240818 59586 241054
rect 59822 240818 60004 241054
rect 59404 240734 60004 240818
rect 59404 240498 59586 240734
rect 59822 240498 60004 240734
rect 59404 205054 60004 240498
rect 59404 204818 59586 205054
rect 59822 204818 60004 205054
rect 59404 204734 60004 204818
rect 59404 204498 59586 204734
rect 59822 204498 60004 204734
rect 59404 169054 60004 204498
rect 59404 168818 59586 169054
rect 59822 168818 60004 169054
rect 59404 168734 60004 168818
rect 59404 168498 59586 168734
rect 59822 168498 60004 168734
rect 59404 133054 60004 168498
rect 59404 132818 59586 133054
rect 59822 132818 60004 133054
rect 59404 132734 60004 132818
rect 59404 132498 59586 132734
rect 59822 132498 60004 132734
rect 59404 97054 60004 132498
rect 59404 96818 59586 97054
rect 59822 96818 60004 97054
rect 59404 96734 60004 96818
rect 59404 96498 59586 96734
rect 59822 96498 60004 96734
rect 59404 61054 60004 96498
rect 59404 60818 59586 61054
rect 59822 60818 60004 61054
rect 59404 60734 60004 60818
rect 59404 60498 59586 60734
rect 59822 60498 60004 60734
rect 59404 25054 60004 60498
rect 59404 24818 59586 25054
rect 59822 24818 60004 25054
rect 59404 24734 60004 24818
rect 59404 24498 59586 24734
rect 59822 24498 60004 24734
rect 59404 -3166 60004 24498
rect 59404 -3402 59586 -3166
rect 59822 -3402 60004 -3166
rect 59404 -3486 60004 -3402
rect 59404 -3722 59586 -3486
rect 59822 -3722 60004 -3486
rect 59404 -3744 60004 -3722
rect 63004 676654 63604 708982
rect 63004 676418 63186 676654
rect 63422 676418 63604 676654
rect 63004 676334 63604 676418
rect 63004 676098 63186 676334
rect 63422 676098 63604 676334
rect 63004 640654 63604 676098
rect 63004 640418 63186 640654
rect 63422 640418 63604 640654
rect 63004 640334 63604 640418
rect 63004 640098 63186 640334
rect 63422 640098 63604 640334
rect 63004 604654 63604 640098
rect 63004 604418 63186 604654
rect 63422 604418 63604 604654
rect 63004 604334 63604 604418
rect 63004 604098 63186 604334
rect 63422 604098 63604 604334
rect 63004 568654 63604 604098
rect 63004 568418 63186 568654
rect 63422 568418 63604 568654
rect 63004 568334 63604 568418
rect 63004 568098 63186 568334
rect 63422 568098 63604 568334
rect 63004 532654 63604 568098
rect 63004 532418 63186 532654
rect 63422 532418 63604 532654
rect 63004 532334 63604 532418
rect 63004 532098 63186 532334
rect 63422 532098 63604 532334
rect 63004 496654 63604 532098
rect 63004 496418 63186 496654
rect 63422 496418 63604 496654
rect 63004 496334 63604 496418
rect 63004 496098 63186 496334
rect 63422 496098 63604 496334
rect 63004 460654 63604 496098
rect 63004 460418 63186 460654
rect 63422 460418 63604 460654
rect 63004 460334 63604 460418
rect 63004 460098 63186 460334
rect 63422 460098 63604 460334
rect 63004 424654 63604 460098
rect 63004 424418 63186 424654
rect 63422 424418 63604 424654
rect 63004 424334 63604 424418
rect 63004 424098 63186 424334
rect 63422 424098 63604 424334
rect 63004 388654 63604 424098
rect 63004 388418 63186 388654
rect 63422 388418 63604 388654
rect 63004 388334 63604 388418
rect 63004 388098 63186 388334
rect 63422 388098 63604 388334
rect 63004 352654 63604 388098
rect 63004 352418 63186 352654
rect 63422 352418 63604 352654
rect 63004 352334 63604 352418
rect 63004 352098 63186 352334
rect 63422 352098 63604 352334
rect 63004 316654 63604 352098
rect 63004 316418 63186 316654
rect 63422 316418 63604 316654
rect 63004 316334 63604 316418
rect 63004 316098 63186 316334
rect 63422 316098 63604 316334
rect 63004 280654 63604 316098
rect 63004 280418 63186 280654
rect 63422 280418 63604 280654
rect 63004 280334 63604 280418
rect 63004 280098 63186 280334
rect 63422 280098 63604 280334
rect 63004 244654 63604 280098
rect 63004 244418 63186 244654
rect 63422 244418 63604 244654
rect 63004 244334 63604 244418
rect 63004 244098 63186 244334
rect 63422 244098 63604 244334
rect 63004 208654 63604 244098
rect 63004 208418 63186 208654
rect 63422 208418 63604 208654
rect 63004 208334 63604 208418
rect 63004 208098 63186 208334
rect 63422 208098 63604 208334
rect 63004 172654 63604 208098
rect 63004 172418 63186 172654
rect 63422 172418 63604 172654
rect 63004 172334 63604 172418
rect 63004 172098 63186 172334
rect 63422 172098 63604 172334
rect 63004 136654 63604 172098
rect 63004 136418 63186 136654
rect 63422 136418 63604 136654
rect 63004 136334 63604 136418
rect 63004 136098 63186 136334
rect 63422 136098 63604 136334
rect 63004 100654 63604 136098
rect 63004 100418 63186 100654
rect 63422 100418 63604 100654
rect 63004 100334 63604 100418
rect 63004 100098 63186 100334
rect 63422 100098 63604 100334
rect 63004 64654 63604 100098
rect 63004 64418 63186 64654
rect 63422 64418 63604 64654
rect 63004 64334 63604 64418
rect 63004 64098 63186 64334
rect 63422 64098 63604 64334
rect 63004 28654 63604 64098
rect 63004 28418 63186 28654
rect 63422 28418 63604 28654
rect 63004 28334 63604 28418
rect 63004 28098 63186 28334
rect 63422 28098 63604 28334
rect 63004 -5046 63604 28098
rect 63004 -5282 63186 -5046
rect 63422 -5282 63604 -5046
rect 63004 -5366 63604 -5282
rect 63004 -5602 63186 -5366
rect 63422 -5602 63604 -5366
rect 63004 -5624 63604 -5602
rect 66604 680254 67204 710862
rect 84604 710478 85204 711440
rect 84604 710242 84786 710478
rect 85022 710242 85204 710478
rect 84604 710158 85204 710242
rect 84604 709922 84786 710158
rect 85022 709922 85204 710158
rect 81004 708598 81604 709560
rect 81004 708362 81186 708598
rect 81422 708362 81604 708598
rect 81004 708278 81604 708362
rect 81004 708042 81186 708278
rect 81422 708042 81604 708278
rect 77404 706718 78004 707680
rect 77404 706482 77586 706718
rect 77822 706482 78004 706718
rect 77404 706398 78004 706482
rect 77404 706162 77586 706398
rect 77822 706162 78004 706398
rect 66604 680018 66786 680254
rect 67022 680018 67204 680254
rect 66604 679934 67204 680018
rect 66604 679698 66786 679934
rect 67022 679698 67204 679934
rect 66604 644254 67204 679698
rect 66604 644018 66786 644254
rect 67022 644018 67204 644254
rect 66604 643934 67204 644018
rect 66604 643698 66786 643934
rect 67022 643698 67204 643934
rect 66604 608254 67204 643698
rect 66604 608018 66786 608254
rect 67022 608018 67204 608254
rect 66604 607934 67204 608018
rect 66604 607698 66786 607934
rect 67022 607698 67204 607934
rect 66604 572254 67204 607698
rect 66604 572018 66786 572254
rect 67022 572018 67204 572254
rect 66604 571934 67204 572018
rect 66604 571698 66786 571934
rect 67022 571698 67204 571934
rect 66604 536254 67204 571698
rect 66604 536018 66786 536254
rect 67022 536018 67204 536254
rect 66604 535934 67204 536018
rect 66604 535698 66786 535934
rect 67022 535698 67204 535934
rect 66604 500254 67204 535698
rect 66604 500018 66786 500254
rect 67022 500018 67204 500254
rect 66604 499934 67204 500018
rect 66604 499698 66786 499934
rect 67022 499698 67204 499934
rect 66604 464254 67204 499698
rect 66604 464018 66786 464254
rect 67022 464018 67204 464254
rect 66604 463934 67204 464018
rect 66604 463698 66786 463934
rect 67022 463698 67204 463934
rect 66604 428254 67204 463698
rect 66604 428018 66786 428254
rect 67022 428018 67204 428254
rect 66604 427934 67204 428018
rect 66604 427698 66786 427934
rect 67022 427698 67204 427934
rect 66604 392254 67204 427698
rect 66604 392018 66786 392254
rect 67022 392018 67204 392254
rect 66604 391934 67204 392018
rect 66604 391698 66786 391934
rect 67022 391698 67204 391934
rect 66604 356254 67204 391698
rect 66604 356018 66786 356254
rect 67022 356018 67204 356254
rect 66604 355934 67204 356018
rect 66604 355698 66786 355934
rect 67022 355698 67204 355934
rect 66604 320254 67204 355698
rect 66604 320018 66786 320254
rect 67022 320018 67204 320254
rect 66604 319934 67204 320018
rect 66604 319698 66786 319934
rect 67022 319698 67204 319934
rect 66604 284254 67204 319698
rect 66604 284018 66786 284254
rect 67022 284018 67204 284254
rect 66604 283934 67204 284018
rect 66604 283698 66786 283934
rect 67022 283698 67204 283934
rect 66604 248254 67204 283698
rect 66604 248018 66786 248254
rect 67022 248018 67204 248254
rect 66604 247934 67204 248018
rect 66604 247698 66786 247934
rect 67022 247698 67204 247934
rect 66604 212254 67204 247698
rect 66604 212018 66786 212254
rect 67022 212018 67204 212254
rect 66604 211934 67204 212018
rect 66604 211698 66786 211934
rect 67022 211698 67204 211934
rect 66604 176254 67204 211698
rect 66604 176018 66786 176254
rect 67022 176018 67204 176254
rect 66604 175934 67204 176018
rect 66604 175698 66786 175934
rect 67022 175698 67204 175934
rect 66604 140254 67204 175698
rect 66604 140018 66786 140254
rect 67022 140018 67204 140254
rect 66604 139934 67204 140018
rect 66604 139698 66786 139934
rect 67022 139698 67204 139934
rect 66604 104254 67204 139698
rect 66604 104018 66786 104254
rect 67022 104018 67204 104254
rect 66604 103934 67204 104018
rect 66604 103698 66786 103934
rect 67022 103698 67204 103934
rect 66604 68254 67204 103698
rect 66604 68018 66786 68254
rect 67022 68018 67204 68254
rect 66604 67934 67204 68018
rect 66604 67698 66786 67934
rect 67022 67698 67204 67934
rect 66604 32254 67204 67698
rect 66604 32018 66786 32254
rect 67022 32018 67204 32254
rect 66604 31934 67204 32018
rect 66604 31698 66786 31934
rect 67022 31698 67204 31934
rect 48604 -6222 48786 -5986
rect 49022 -6222 49204 -5986
rect 48604 -6306 49204 -6222
rect 48604 -6542 48786 -6306
rect 49022 -6542 49204 -6306
rect 48604 -7504 49204 -6542
rect 66604 -6926 67204 31698
rect 73804 704838 74404 705800
rect 73804 704602 73986 704838
rect 74222 704602 74404 704838
rect 73804 704518 74404 704602
rect 73804 704282 73986 704518
rect 74222 704282 74404 704518
rect 73804 687454 74404 704282
rect 73804 687218 73986 687454
rect 74222 687218 74404 687454
rect 73804 687134 74404 687218
rect 73804 686898 73986 687134
rect 74222 686898 74404 687134
rect 73804 651454 74404 686898
rect 73804 651218 73986 651454
rect 74222 651218 74404 651454
rect 73804 651134 74404 651218
rect 73804 650898 73986 651134
rect 74222 650898 74404 651134
rect 73804 615454 74404 650898
rect 73804 615218 73986 615454
rect 74222 615218 74404 615454
rect 73804 615134 74404 615218
rect 73804 614898 73986 615134
rect 74222 614898 74404 615134
rect 73804 579454 74404 614898
rect 73804 579218 73986 579454
rect 74222 579218 74404 579454
rect 73804 579134 74404 579218
rect 73804 578898 73986 579134
rect 74222 578898 74404 579134
rect 73804 543454 74404 578898
rect 73804 543218 73986 543454
rect 74222 543218 74404 543454
rect 73804 543134 74404 543218
rect 73804 542898 73986 543134
rect 74222 542898 74404 543134
rect 73804 507454 74404 542898
rect 73804 507218 73986 507454
rect 74222 507218 74404 507454
rect 73804 507134 74404 507218
rect 73804 506898 73986 507134
rect 74222 506898 74404 507134
rect 73804 471454 74404 506898
rect 73804 471218 73986 471454
rect 74222 471218 74404 471454
rect 73804 471134 74404 471218
rect 73804 470898 73986 471134
rect 74222 470898 74404 471134
rect 73804 435454 74404 470898
rect 73804 435218 73986 435454
rect 74222 435218 74404 435454
rect 73804 435134 74404 435218
rect 73804 434898 73986 435134
rect 74222 434898 74404 435134
rect 73804 399454 74404 434898
rect 73804 399218 73986 399454
rect 74222 399218 74404 399454
rect 73804 399134 74404 399218
rect 73804 398898 73986 399134
rect 74222 398898 74404 399134
rect 73804 363454 74404 398898
rect 73804 363218 73986 363454
rect 74222 363218 74404 363454
rect 73804 363134 74404 363218
rect 73804 362898 73986 363134
rect 74222 362898 74404 363134
rect 73804 327454 74404 362898
rect 73804 327218 73986 327454
rect 74222 327218 74404 327454
rect 73804 327134 74404 327218
rect 73804 326898 73986 327134
rect 74222 326898 74404 327134
rect 73804 291454 74404 326898
rect 73804 291218 73986 291454
rect 74222 291218 74404 291454
rect 73804 291134 74404 291218
rect 73804 290898 73986 291134
rect 74222 290898 74404 291134
rect 73804 255454 74404 290898
rect 73804 255218 73986 255454
rect 74222 255218 74404 255454
rect 73804 255134 74404 255218
rect 73804 254898 73986 255134
rect 74222 254898 74404 255134
rect 73804 219454 74404 254898
rect 73804 219218 73986 219454
rect 74222 219218 74404 219454
rect 73804 219134 74404 219218
rect 73804 218898 73986 219134
rect 74222 218898 74404 219134
rect 73804 183454 74404 218898
rect 73804 183218 73986 183454
rect 74222 183218 74404 183454
rect 73804 183134 74404 183218
rect 73804 182898 73986 183134
rect 74222 182898 74404 183134
rect 73804 147454 74404 182898
rect 73804 147218 73986 147454
rect 74222 147218 74404 147454
rect 73804 147134 74404 147218
rect 73804 146898 73986 147134
rect 74222 146898 74404 147134
rect 73804 111454 74404 146898
rect 73804 111218 73986 111454
rect 74222 111218 74404 111454
rect 73804 111134 74404 111218
rect 73804 110898 73986 111134
rect 74222 110898 74404 111134
rect 73804 75454 74404 110898
rect 73804 75218 73986 75454
rect 74222 75218 74404 75454
rect 73804 75134 74404 75218
rect 73804 74898 73986 75134
rect 74222 74898 74404 75134
rect 73804 39454 74404 74898
rect 73804 39218 73986 39454
rect 74222 39218 74404 39454
rect 73804 39134 74404 39218
rect 73804 38898 73986 39134
rect 74222 38898 74404 39134
rect 73804 3454 74404 38898
rect 73804 3218 73986 3454
rect 74222 3218 74404 3454
rect 73804 3134 74404 3218
rect 73804 2898 73986 3134
rect 74222 2898 74404 3134
rect 73804 -346 74404 2898
rect 73804 -582 73986 -346
rect 74222 -582 74404 -346
rect 73804 -666 74404 -582
rect 73804 -902 73986 -666
rect 74222 -902 74404 -666
rect 73804 -1864 74404 -902
rect 77404 691054 78004 706162
rect 77404 690818 77586 691054
rect 77822 690818 78004 691054
rect 77404 690734 78004 690818
rect 77404 690498 77586 690734
rect 77822 690498 78004 690734
rect 77404 655054 78004 690498
rect 77404 654818 77586 655054
rect 77822 654818 78004 655054
rect 77404 654734 78004 654818
rect 77404 654498 77586 654734
rect 77822 654498 78004 654734
rect 77404 619054 78004 654498
rect 77404 618818 77586 619054
rect 77822 618818 78004 619054
rect 77404 618734 78004 618818
rect 77404 618498 77586 618734
rect 77822 618498 78004 618734
rect 77404 583054 78004 618498
rect 77404 582818 77586 583054
rect 77822 582818 78004 583054
rect 77404 582734 78004 582818
rect 77404 582498 77586 582734
rect 77822 582498 78004 582734
rect 77404 547054 78004 582498
rect 77404 546818 77586 547054
rect 77822 546818 78004 547054
rect 77404 546734 78004 546818
rect 77404 546498 77586 546734
rect 77822 546498 78004 546734
rect 77404 511054 78004 546498
rect 77404 510818 77586 511054
rect 77822 510818 78004 511054
rect 77404 510734 78004 510818
rect 77404 510498 77586 510734
rect 77822 510498 78004 510734
rect 77404 475054 78004 510498
rect 77404 474818 77586 475054
rect 77822 474818 78004 475054
rect 77404 474734 78004 474818
rect 77404 474498 77586 474734
rect 77822 474498 78004 474734
rect 77404 439054 78004 474498
rect 77404 438818 77586 439054
rect 77822 438818 78004 439054
rect 77404 438734 78004 438818
rect 77404 438498 77586 438734
rect 77822 438498 78004 438734
rect 77404 403054 78004 438498
rect 77404 402818 77586 403054
rect 77822 402818 78004 403054
rect 77404 402734 78004 402818
rect 77404 402498 77586 402734
rect 77822 402498 78004 402734
rect 77404 367054 78004 402498
rect 77404 366818 77586 367054
rect 77822 366818 78004 367054
rect 77404 366734 78004 366818
rect 77404 366498 77586 366734
rect 77822 366498 78004 366734
rect 77404 331054 78004 366498
rect 77404 330818 77586 331054
rect 77822 330818 78004 331054
rect 77404 330734 78004 330818
rect 77404 330498 77586 330734
rect 77822 330498 78004 330734
rect 77404 295054 78004 330498
rect 77404 294818 77586 295054
rect 77822 294818 78004 295054
rect 77404 294734 78004 294818
rect 77404 294498 77586 294734
rect 77822 294498 78004 294734
rect 77404 259054 78004 294498
rect 77404 258818 77586 259054
rect 77822 258818 78004 259054
rect 77404 258734 78004 258818
rect 77404 258498 77586 258734
rect 77822 258498 78004 258734
rect 77404 223054 78004 258498
rect 77404 222818 77586 223054
rect 77822 222818 78004 223054
rect 77404 222734 78004 222818
rect 77404 222498 77586 222734
rect 77822 222498 78004 222734
rect 77404 187054 78004 222498
rect 77404 186818 77586 187054
rect 77822 186818 78004 187054
rect 77404 186734 78004 186818
rect 77404 186498 77586 186734
rect 77822 186498 78004 186734
rect 77404 151054 78004 186498
rect 77404 150818 77586 151054
rect 77822 150818 78004 151054
rect 77404 150734 78004 150818
rect 77404 150498 77586 150734
rect 77822 150498 78004 150734
rect 77404 115054 78004 150498
rect 77404 114818 77586 115054
rect 77822 114818 78004 115054
rect 77404 114734 78004 114818
rect 77404 114498 77586 114734
rect 77822 114498 78004 114734
rect 77404 79054 78004 114498
rect 77404 78818 77586 79054
rect 77822 78818 78004 79054
rect 77404 78734 78004 78818
rect 77404 78498 77586 78734
rect 77822 78498 78004 78734
rect 77404 43054 78004 78498
rect 77404 42818 77586 43054
rect 77822 42818 78004 43054
rect 77404 42734 78004 42818
rect 77404 42498 77586 42734
rect 77822 42498 78004 42734
rect 77404 7054 78004 42498
rect 77404 6818 77586 7054
rect 77822 6818 78004 7054
rect 77404 6734 78004 6818
rect 77404 6498 77586 6734
rect 77822 6498 78004 6734
rect 77404 -2226 78004 6498
rect 77404 -2462 77586 -2226
rect 77822 -2462 78004 -2226
rect 77404 -2546 78004 -2462
rect 77404 -2782 77586 -2546
rect 77822 -2782 78004 -2546
rect 77404 -3744 78004 -2782
rect 81004 694654 81604 708042
rect 81004 694418 81186 694654
rect 81422 694418 81604 694654
rect 81004 694334 81604 694418
rect 81004 694098 81186 694334
rect 81422 694098 81604 694334
rect 81004 658654 81604 694098
rect 81004 658418 81186 658654
rect 81422 658418 81604 658654
rect 81004 658334 81604 658418
rect 81004 658098 81186 658334
rect 81422 658098 81604 658334
rect 81004 622654 81604 658098
rect 81004 622418 81186 622654
rect 81422 622418 81604 622654
rect 81004 622334 81604 622418
rect 81004 622098 81186 622334
rect 81422 622098 81604 622334
rect 81004 586654 81604 622098
rect 81004 586418 81186 586654
rect 81422 586418 81604 586654
rect 81004 586334 81604 586418
rect 81004 586098 81186 586334
rect 81422 586098 81604 586334
rect 81004 550654 81604 586098
rect 81004 550418 81186 550654
rect 81422 550418 81604 550654
rect 81004 550334 81604 550418
rect 81004 550098 81186 550334
rect 81422 550098 81604 550334
rect 81004 514654 81604 550098
rect 81004 514418 81186 514654
rect 81422 514418 81604 514654
rect 81004 514334 81604 514418
rect 81004 514098 81186 514334
rect 81422 514098 81604 514334
rect 81004 478654 81604 514098
rect 81004 478418 81186 478654
rect 81422 478418 81604 478654
rect 81004 478334 81604 478418
rect 81004 478098 81186 478334
rect 81422 478098 81604 478334
rect 81004 442654 81604 478098
rect 81004 442418 81186 442654
rect 81422 442418 81604 442654
rect 81004 442334 81604 442418
rect 81004 442098 81186 442334
rect 81422 442098 81604 442334
rect 81004 406654 81604 442098
rect 81004 406418 81186 406654
rect 81422 406418 81604 406654
rect 81004 406334 81604 406418
rect 81004 406098 81186 406334
rect 81422 406098 81604 406334
rect 81004 370654 81604 406098
rect 81004 370418 81186 370654
rect 81422 370418 81604 370654
rect 81004 370334 81604 370418
rect 81004 370098 81186 370334
rect 81422 370098 81604 370334
rect 81004 334654 81604 370098
rect 81004 334418 81186 334654
rect 81422 334418 81604 334654
rect 81004 334334 81604 334418
rect 81004 334098 81186 334334
rect 81422 334098 81604 334334
rect 81004 298654 81604 334098
rect 81004 298418 81186 298654
rect 81422 298418 81604 298654
rect 81004 298334 81604 298418
rect 81004 298098 81186 298334
rect 81422 298098 81604 298334
rect 81004 262654 81604 298098
rect 81004 262418 81186 262654
rect 81422 262418 81604 262654
rect 81004 262334 81604 262418
rect 81004 262098 81186 262334
rect 81422 262098 81604 262334
rect 81004 226654 81604 262098
rect 81004 226418 81186 226654
rect 81422 226418 81604 226654
rect 81004 226334 81604 226418
rect 81004 226098 81186 226334
rect 81422 226098 81604 226334
rect 81004 190654 81604 226098
rect 81004 190418 81186 190654
rect 81422 190418 81604 190654
rect 81004 190334 81604 190418
rect 81004 190098 81186 190334
rect 81422 190098 81604 190334
rect 81004 154654 81604 190098
rect 81004 154418 81186 154654
rect 81422 154418 81604 154654
rect 81004 154334 81604 154418
rect 81004 154098 81186 154334
rect 81422 154098 81604 154334
rect 81004 118654 81604 154098
rect 81004 118418 81186 118654
rect 81422 118418 81604 118654
rect 81004 118334 81604 118418
rect 81004 118098 81186 118334
rect 81422 118098 81604 118334
rect 81004 82654 81604 118098
rect 81004 82418 81186 82654
rect 81422 82418 81604 82654
rect 81004 82334 81604 82418
rect 81004 82098 81186 82334
rect 81422 82098 81604 82334
rect 81004 46654 81604 82098
rect 81004 46418 81186 46654
rect 81422 46418 81604 46654
rect 81004 46334 81604 46418
rect 81004 46098 81186 46334
rect 81422 46098 81604 46334
rect 81004 10654 81604 46098
rect 81004 10418 81186 10654
rect 81422 10418 81604 10654
rect 81004 10334 81604 10418
rect 81004 10098 81186 10334
rect 81422 10098 81604 10334
rect 81004 -4106 81604 10098
rect 81004 -4342 81186 -4106
rect 81422 -4342 81604 -4106
rect 81004 -4426 81604 -4342
rect 81004 -4662 81186 -4426
rect 81422 -4662 81604 -4426
rect 81004 -5624 81604 -4662
rect 84604 698254 85204 709922
rect 102604 711418 103204 711440
rect 102604 711182 102786 711418
rect 103022 711182 103204 711418
rect 102604 711098 103204 711182
rect 102604 710862 102786 711098
rect 103022 710862 103204 711098
rect 99004 709538 99604 709560
rect 99004 709302 99186 709538
rect 99422 709302 99604 709538
rect 99004 709218 99604 709302
rect 99004 708982 99186 709218
rect 99422 708982 99604 709218
rect 95404 707658 96004 707680
rect 95404 707422 95586 707658
rect 95822 707422 96004 707658
rect 95404 707338 96004 707422
rect 95404 707102 95586 707338
rect 95822 707102 96004 707338
rect 84604 698018 84786 698254
rect 85022 698018 85204 698254
rect 84604 697934 85204 698018
rect 84604 697698 84786 697934
rect 85022 697698 85204 697934
rect 84604 662254 85204 697698
rect 84604 662018 84786 662254
rect 85022 662018 85204 662254
rect 84604 661934 85204 662018
rect 84604 661698 84786 661934
rect 85022 661698 85204 661934
rect 84604 626254 85204 661698
rect 84604 626018 84786 626254
rect 85022 626018 85204 626254
rect 84604 625934 85204 626018
rect 84604 625698 84786 625934
rect 85022 625698 85204 625934
rect 84604 590254 85204 625698
rect 84604 590018 84786 590254
rect 85022 590018 85204 590254
rect 84604 589934 85204 590018
rect 84604 589698 84786 589934
rect 85022 589698 85204 589934
rect 84604 554254 85204 589698
rect 84604 554018 84786 554254
rect 85022 554018 85204 554254
rect 84604 553934 85204 554018
rect 84604 553698 84786 553934
rect 85022 553698 85204 553934
rect 84604 518254 85204 553698
rect 84604 518018 84786 518254
rect 85022 518018 85204 518254
rect 84604 517934 85204 518018
rect 84604 517698 84786 517934
rect 85022 517698 85204 517934
rect 84604 482254 85204 517698
rect 84604 482018 84786 482254
rect 85022 482018 85204 482254
rect 84604 481934 85204 482018
rect 84604 481698 84786 481934
rect 85022 481698 85204 481934
rect 84604 446254 85204 481698
rect 84604 446018 84786 446254
rect 85022 446018 85204 446254
rect 84604 445934 85204 446018
rect 84604 445698 84786 445934
rect 85022 445698 85204 445934
rect 84604 410254 85204 445698
rect 84604 410018 84786 410254
rect 85022 410018 85204 410254
rect 84604 409934 85204 410018
rect 84604 409698 84786 409934
rect 85022 409698 85204 409934
rect 84604 374254 85204 409698
rect 84604 374018 84786 374254
rect 85022 374018 85204 374254
rect 84604 373934 85204 374018
rect 84604 373698 84786 373934
rect 85022 373698 85204 373934
rect 84604 338254 85204 373698
rect 84604 338018 84786 338254
rect 85022 338018 85204 338254
rect 84604 337934 85204 338018
rect 84604 337698 84786 337934
rect 85022 337698 85204 337934
rect 84604 302254 85204 337698
rect 84604 302018 84786 302254
rect 85022 302018 85204 302254
rect 84604 301934 85204 302018
rect 84604 301698 84786 301934
rect 85022 301698 85204 301934
rect 84604 266254 85204 301698
rect 84604 266018 84786 266254
rect 85022 266018 85204 266254
rect 84604 265934 85204 266018
rect 84604 265698 84786 265934
rect 85022 265698 85204 265934
rect 84604 230254 85204 265698
rect 84604 230018 84786 230254
rect 85022 230018 85204 230254
rect 84604 229934 85204 230018
rect 84604 229698 84786 229934
rect 85022 229698 85204 229934
rect 84604 194254 85204 229698
rect 84604 194018 84786 194254
rect 85022 194018 85204 194254
rect 84604 193934 85204 194018
rect 84604 193698 84786 193934
rect 85022 193698 85204 193934
rect 84604 158254 85204 193698
rect 84604 158018 84786 158254
rect 85022 158018 85204 158254
rect 84604 157934 85204 158018
rect 84604 157698 84786 157934
rect 85022 157698 85204 157934
rect 84604 122254 85204 157698
rect 84604 122018 84786 122254
rect 85022 122018 85204 122254
rect 84604 121934 85204 122018
rect 84604 121698 84786 121934
rect 85022 121698 85204 121934
rect 84604 86254 85204 121698
rect 84604 86018 84786 86254
rect 85022 86018 85204 86254
rect 84604 85934 85204 86018
rect 84604 85698 84786 85934
rect 85022 85698 85204 85934
rect 84604 50254 85204 85698
rect 84604 50018 84786 50254
rect 85022 50018 85204 50254
rect 84604 49934 85204 50018
rect 84604 49698 84786 49934
rect 85022 49698 85204 49934
rect 84604 14254 85204 49698
rect 84604 14018 84786 14254
rect 85022 14018 85204 14254
rect 84604 13934 85204 14018
rect 84604 13698 84786 13934
rect 85022 13698 85204 13934
rect 66604 -7162 66786 -6926
rect 67022 -7162 67204 -6926
rect 66604 -7246 67204 -7162
rect 66604 -7482 66786 -7246
rect 67022 -7482 67204 -7246
rect 66604 -7504 67204 -7482
rect 84604 -5986 85204 13698
rect 91804 705778 92404 705800
rect 91804 705542 91986 705778
rect 92222 705542 92404 705778
rect 91804 705458 92404 705542
rect 91804 705222 91986 705458
rect 92222 705222 92404 705458
rect 91804 669454 92404 705222
rect 91804 669218 91986 669454
rect 92222 669218 92404 669454
rect 91804 669134 92404 669218
rect 91804 668898 91986 669134
rect 92222 668898 92404 669134
rect 91804 633454 92404 668898
rect 91804 633218 91986 633454
rect 92222 633218 92404 633454
rect 91804 633134 92404 633218
rect 91804 632898 91986 633134
rect 92222 632898 92404 633134
rect 91804 597454 92404 632898
rect 91804 597218 91986 597454
rect 92222 597218 92404 597454
rect 91804 597134 92404 597218
rect 91804 596898 91986 597134
rect 92222 596898 92404 597134
rect 91804 561454 92404 596898
rect 91804 561218 91986 561454
rect 92222 561218 92404 561454
rect 91804 561134 92404 561218
rect 91804 560898 91986 561134
rect 92222 560898 92404 561134
rect 91804 525454 92404 560898
rect 91804 525218 91986 525454
rect 92222 525218 92404 525454
rect 91804 525134 92404 525218
rect 91804 524898 91986 525134
rect 92222 524898 92404 525134
rect 91804 489454 92404 524898
rect 91804 489218 91986 489454
rect 92222 489218 92404 489454
rect 91804 489134 92404 489218
rect 91804 488898 91986 489134
rect 92222 488898 92404 489134
rect 91804 453454 92404 488898
rect 91804 453218 91986 453454
rect 92222 453218 92404 453454
rect 91804 453134 92404 453218
rect 91804 452898 91986 453134
rect 92222 452898 92404 453134
rect 91804 417454 92404 452898
rect 91804 417218 91986 417454
rect 92222 417218 92404 417454
rect 91804 417134 92404 417218
rect 91804 416898 91986 417134
rect 92222 416898 92404 417134
rect 91804 381454 92404 416898
rect 91804 381218 91986 381454
rect 92222 381218 92404 381454
rect 91804 381134 92404 381218
rect 91804 380898 91986 381134
rect 92222 380898 92404 381134
rect 91804 345454 92404 380898
rect 91804 345218 91986 345454
rect 92222 345218 92404 345454
rect 91804 345134 92404 345218
rect 91804 344898 91986 345134
rect 92222 344898 92404 345134
rect 91804 309454 92404 344898
rect 91804 309218 91986 309454
rect 92222 309218 92404 309454
rect 91804 309134 92404 309218
rect 91804 308898 91986 309134
rect 92222 308898 92404 309134
rect 91804 273454 92404 308898
rect 91804 273218 91986 273454
rect 92222 273218 92404 273454
rect 91804 273134 92404 273218
rect 91804 272898 91986 273134
rect 92222 272898 92404 273134
rect 91804 237454 92404 272898
rect 91804 237218 91986 237454
rect 92222 237218 92404 237454
rect 91804 237134 92404 237218
rect 91804 236898 91986 237134
rect 92222 236898 92404 237134
rect 91804 201454 92404 236898
rect 91804 201218 91986 201454
rect 92222 201218 92404 201454
rect 91804 201134 92404 201218
rect 91804 200898 91986 201134
rect 92222 200898 92404 201134
rect 91804 165454 92404 200898
rect 91804 165218 91986 165454
rect 92222 165218 92404 165454
rect 91804 165134 92404 165218
rect 91804 164898 91986 165134
rect 92222 164898 92404 165134
rect 91804 129454 92404 164898
rect 91804 129218 91986 129454
rect 92222 129218 92404 129454
rect 91804 129134 92404 129218
rect 91804 128898 91986 129134
rect 92222 128898 92404 129134
rect 91804 93454 92404 128898
rect 91804 93218 91986 93454
rect 92222 93218 92404 93454
rect 91804 93134 92404 93218
rect 91804 92898 91986 93134
rect 92222 92898 92404 93134
rect 91804 57454 92404 92898
rect 91804 57218 91986 57454
rect 92222 57218 92404 57454
rect 91804 57134 92404 57218
rect 91804 56898 91986 57134
rect 92222 56898 92404 57134
rect 91804 21454 92404 56898
rect 91804 21218 91986 21454
rect 92222 21218 92404 21454
rect 91804 21134 92404 21218
rect 91804 20898 91986 21134
rect 92222 20898 92404 21134
rect 91804 -1286 92404 20898
rect 91804 -1522 91986 -1286
rect 92222 -1522 92404 -1286
rect 91804 -1606 92404 -1522
rect 91804 -1842 91986 -1606
rect 92222 -1842 92404 -1606
rect 91804 -1864 92404 -1842
rect 95404 673054 96004 707102
rect 95404 672818 95586 673054
rect 95822 672818 96004 673054
rect 95404 672734 96004 672818
rect 95404 672498 95586 672734
rect 95822 672498 96004 672734
rect 95404 637054 96004 672498
rect 95404 636818 95586 637054
rect 95822 636818 96004 637054
rect 95404 636734 96004 636818
rect 95404 636498 95586 636734
rect 95822 636498 96004 636734
rect 95404 601054 96004 636498
rect 95404 600818 95586 601054
rect 95822 600818 96004 601054
rect 95404 600734 96004 600818
rect 95404 600498 95586 600734
rect 95822 600498 96004 600734
rect 95404 565054 96004 600498
rect 95404 564818 95586 565054
rect 95822 564818 96004 565054
rect 95404 564734 96004 564818
rect 95404 564498 95586 564734
rect 95822 564498 96004 564734
rect 95404 529054 96004 564498
rect 95404 528818 95586 529054
rect 95822 528818 96004 529054
rect 95404 528734 96004 528818
rect 95404 528498 95586 528734
rect 95822 528498 96004 528734
rect 95404 493054 96004 528498
rect 95404 492818 95586 493054
rect 95822 492818 96004 493054
rect 95404 492734 96004 492818
rect 95404 492498 95586 492734
rect 95822 492498 96004 492734
rect 95404 457054 96004 492498
rect 95404 456818 95586 457054
rect 95822 456818 96004 457054
rect 95404 456734 96004 456818
rect 95404 456498 95586 456734
rect 95822 456498 96004 456734
rect 95404 421054 96004 456498
rect 95404 420818 95586 421054
rect 95822 420818 96004 421054
rect 95404 420734 96004 420818
rect 95404 420498 95586 420734
rect 95822 420498 96004 420734
rect 95404 385054 96004 420498
rect 95404 384818 95586 385054
rect 95822 384818 96004 385054
rect 95404 384734 96004 384818
rect 95404 384498 95586 384734
rect 95822 384498 96004 384734
rect 95404 349054 96004 384498
rect 95404 348818 95586 349054
rect 95822 348818 96004 349054
rect 95404 348734 96004 348818
rect 95404 348498 95586 348734
rect 95822 348498 96004 348734
rect 95404 313054 96004 348498
rect 95404 312818 95586 313054
rect 95822 312818 96004 313054
rect 95404 312734 96004 312818
rect 95404 312498 95586 312734
rect 95822 312498 96004 312734
rect 95404 277054 96004 312498
rect 95404 276818 95586 277054
rect 95822 276818 96004 277054
rect 95404 276734 96004 276818
rect 95404 276498 95586 276734
rect 95822 276498 96004 276734
rect 95404 241054 96004 276498
rect 95404 240818 95586 241054
rect 95822 240818 96004 241054
rect 95404 240734 96004 240818
rect 95404 240498 95586 240734
rect 95822 240498 96004 240734
rect 95404 205054 96004 240498
rect 95404 204818 95586 205054
rect 95822 204818 96004 205054
rect 95404 204734 96004 204818
rect 95404 204498 95586 204734
rect 95822 204498 96004 204734
rect 95404 169054 96004 204498
rect 95404 168818 95586 169054
rect 95822 168818 96004 169054
rect 95404 168734 96004 168818
rect 95404 168498 95586 168734
rect 95822 168498 96004 168734
rect 95404 133054 96004 168498
rect 95404 132818 95586 133054
rect 95822 132818 96004 133054
rect 95404 132734 96004 132818
rect 95404 132498 95586 132734
rect 95822 132498 96004 132734
rect 95404 97054 96004 132498
rect 95404 96818 95586 97054
rect 95822 96818 96004 97054
rect 95404 96734 96004 96818
rect 95404 96498 95586 96734
rect 95822 96498 96004 96734
rect 95404 61054 96004 96498
rect 95404 60818 95586 61054
rect 95822 60818 96004 61054
rect 95404 60734 96004 60818
rect 95404 60498 95586 60734
rect 95822 60498 96004 60734
rect 95404 25054 96004 60498
rect 95404 24818 95586 25054
rect 95822 24818 96004 25054
rect 95404 24734 96004 24818
rect 95404 24498 95586 24734
rect 95822 24498 96004 24734
rect 95404 -3166 96004 24498
rect 95404 -3402 95586 -3166
rect 95822 -3402 96004 -3166
rect 95404 -3486 96004 -3402
rect 95404 -3722 95586 -3486
rect 95822 -3722 96004 -3486
rect 95404 -3744 96004 -3722
rect 99004 676654 99604 708982
rect 99004 676418 99186 676654
rect 99422 676418 99604 676654
rect 99004 676334 99604 676418
rect 99004 676098 99186 676334
rect 99422 676098 99604 676334
rect 99004 640654 99604 676098
rect 99004 640418 99186 640654
rect 99422 640418 99604 640654
rect 99004 640334 99604 640418
rect 99004 640098 99186 640334
rect 99422 640098 99604 640334
rect 99004 604654 99604 640098
rect 99004 604418 99186 604654
rect 99422 604418 99604 604654
rect 99004 604334 99604 604418
rect 99004 604098 99186 604334
rect 99422 604098 99604 604334
rect 99004 568654 99604 604098
rect 99004 568418 99186 568654
rect 99422 568418 99604 568654
rect 99004 568334 99604 568418
rect 99004 568098 99186 568334
rect 99422 568098 99604 568334
rect 99004 532654 99604 568098
rect 99004 532418 99186 532654
rect 99422 532418 99604 532654
rect 99004 532334 99604 532418
rect 99004 532098 99186 532334
rect 99422 532098 99604 532334
rect 99004 496654 99604 532098
rect 99004 496418 99186 496654
rect 99422 496418 99604 496654
rect 99004 496334 99604 496418
rect 99004 496098 99186 496334
rect 99422 496098 99604 496334
rect 99004 460654 99604 496098
rect 99004 460418 99186 460654
rect 99422 460418 99604 460654
rect 99004 460334 99604 460418
rect 99004 460098 99186 460334
rect 99422 460098 99604 460334
rect 99004 424654 99604 460098
rect 99004 424418 99186 424654
rect 99422 424418 99604 424654
rect 99004 424334 99604 424418
rect 99004 424098 99186 424334
rect 99422 424098 99604 424334
rect 99004 388654 99604 424098
rect 99004 388418 99186 388654
rect 99422 388418 99604 388654
rect 99004 388334 99604 388418
rect 99004 388098 99186 388334
rect 99422 388098 99604 388334
rect 99004 352654 99604 388098
rect 99004 352418 99186 352654
rect 99422 352418 99604 352654
rect 99004 352334 99604 352418
rect 99004 352098 99186 352334
rect 99422 352098 99604 352334
rect 99004 316654 99604 352098
rect 99004 316418 99186 316654
rect 99422 316418 99604 316654
rect 99004 316334 99604 316418
rect 99004 316098 99186 316334
rect 99422 316098 99604 316334
rect 99004 280654 99604 316098
rect 99004 280418 99186 280654
rect 99422 280418 99604 280654
rect 99004 280334 99604 280418
rect 99004 280098 99186 280334
rect 99422 280098 99604 280334
rect 99004 244654 99604 280098
rect 99004 244418 99186 244654
rect 99422 244418 99604 244654
rect 99004 244334 99604 244418
rect 99004 244098 99186 244334
rect 99422 244098 99604 244334
rect 99004 208654 99604 244098
rect 99004 208418 99186 208654
rect 99422 208418 99604 208654
rect 99004 208334 99604 208418
rect 99004 208098 99186 208334
rect 99422 208098 99604 208334
rect 99004 172654 99604 208098
rect 99004 172418 99186 172654
rect 99422 172418 99604 172654
rect 99004 172334 99604 172418
rect 99004 172098 99186 172334
rect 99422 172098 99604 172334
rect 99004 136654 99604 172098
rect 99004 136418 99186 136654
rect 99422 136418 99604 136654
rect 99004 136334 99604 136418
rect 99004 136098 99186 136334
rect 99422 136098 99604 136334
rect 99004 100654 99604 136098
rect 99004 100418 99186 100654
rect 99422 100418 99604 100654
rect 99004 100334 99604 100418
rect 99004 100098 99186 100334
rect 99422 100098 99604 100334
rect 99004 64654 99604 100098
rect 99004 64418 99186 64654
rect 99422 64418 99604 64654
rect 99004 64334 99604 64418
rect 99004 64098 99186 64334
rect 99422 64098 99604 64334
rect 99004 28654 99604 64098
rect 99004 28418 99186 28654
rect 99422 28418 99604 28654
rect 99004 28334 99604 28418
rect 99004 28098 99186 28334
rect 99422 28098 99604 28334
rect 99004 -5046 99604 28098
rect 99004 -5282 99186 -5046
rect 99422 -5282 99604 -5046
rect 99004 -5366 99604 -5282
rect 99004 -5602 99186 -5366
rect 99422 -5602 99604 -5366
rect 99004 -5624 99604 -5602
rect 102604 680254 103204 710862
rect 120604 710478 121204 711440
rect 120604 710242 120786 710478
rect 121022 710242 121204 710478
rect 120604 710158 121204 710242
rect 120604 709922 120786 710158
rect 121022 709922 121204 710158
rect 117004 708598 117604 709560
rect 117004 708362 117186 708598
rect 117422 708362 117604 708598
rect 117004 708278 117604 708362
rect 117004 708042 117186 708278
rect 117422 708042 117604 708278
rect 113404 706718 114004 707680
rect 113404 706482 113586 706718
rect 113822 706482 114004 706718
rect 113404 706398 114004 706482
rect 113404 706162 113586 706398
rect 113822 706162 114004 706398
rect 102604 680018 102786 680254
rect 103022 680018 103204 680254
rect 102604 679934 103204 680018
rect 102604 679698 102786 679934
rect 103022 679698 103204 679934
rect 102604 644254 103204 679698
rect 102604 644018 102786 644254
rect 103022 644018 103204 644254
rect 102604 643934 103204 644018
rect 102604 643698 102786 643934
rect 103022 643698 103204 643934
rect 102604 608254 103204 643698
rect 102604 608018 102786 608254
rect 103022 608018 103204 608254
rect 102604 607934 103204 608018
rect 102604 607698 102786 607934
rect 103022 607698 103204 607934
rect 102604 572254 103204 607698
rect 102604 572018 102786 572254
rect 103022 572018 103204 572254
rect 102604 571934 103204 572018
rect 102604 571698 102786 571934
rect 103022 571698 103204 571934
rect 102604 536254 103204 571698
rect 102604 536018 102786 536254
rect 103022 536018 103204 536254
rect 102604 535934 103204 536018
rect 102604 535698 102786 535934
rect 103022 535698 103204 535934
rect 102604 500254 103204 535698
rect 102604 500018 102786 500254
rect 103022 500018 103204 500254
rect 102604 499934 103204 500018
rect 102604 499698 102786 499934
rect 103022 499698 103204 499934
rect 102604 464254 103204 499698
rect 102604 464018 102786 464254
rect 103022 464018 103204 464254
rect 102604 463934 103204 464018
rect 102604 463698 102786 463934
rect 103022 463698 103204 463934
rect 102604 428254 103204 463698
rect 102604 428018 102786 428254
rect 103022 428018 103204 428254
rect 102604 427934 103204 428018
rect 102604 427698 102786 427934
rect 103022 427698 103204 427934
rect 102604 392254 103204 427698
rect 102604 392018 102786 392254
rect 103022 392018 103204 392254
rect 102604 391934 103204 392018
rect 102604 391698 102786 391934
rect 103022 391698 103204 391934
rect 102604 356254 103204 391698
rect 102604 356018 102786 356254
rect 103022 356018 103204 356254
rect 102604 355934 103204 356018
rect 102604 355698 102786 355934
rect 103022 355698 103204 355934
rect 102604 320254 103204 355698
rect 102604 320018 102786 320254
rect 103022 320018 103204 320254
rect 102604 319934 103204 320018
rect 102604 319698 102786 319934
rect 103022 319698 103204 319934
rect 102604 284254 103204 319698
rect 102604 284018 102786 284254
rect 103022 284018 103204 284254
rect 102604 283934 103204 284018
rect 102604 283698 102786 283934
rect 103022 283698 103204 283934
rect 102604 248254 103204 283698
rect 102604 248018 102786 248254
rect 103022 248018 103204 248254
rect 102604 247934 103204 248018
rect 102604 247698 102786 247934
rect 103022 247698 103204 247934
rect 102604 212254 103204 247698
rect 102604 212018 102786 212254
rect 103022 212018 103204 212254
rect 102604 211934 103204 212018
rect 102604 211698 102786 211934
rect 103022 211698 103204 211934
rect 102604 176254 103204 211698
rect 102604 176018 102786 176254
rect 103022 176018 103204 176254
rect 102604 175934 103204 176018
rect 102604 175698 102786 175934
rect 103022 175698 103204 175934
rect 102604 140254 103204 175698
rect 102604 140018 102786 140254
rect 103022 140018 103204 140254
rect 102604 139934 103204 140018
rect 102604 139698 102786 139934
rect 103022 139698 103204 139934
rect 102604 104254 103204 139698
rect 102604 104018 102786 104254
rect 103022 104018 103204 104254
rect 102604 103934 103204 104018
rect 102604 103698 102786 103934
rect 103022 103698 103204 103934
rect 102604 68254 103204 103698
rect 102604 68018 102786 68254
rect 103022 68018 103204 68254
rect 102604 67934 103204 68018
rect 102604 67698 102786 67934
rect 103022 67698 103204 67934
rect 102604 32254 103204 67698
rect 102604 32018 102786 32254
rect 103022 32018 103204 32254
rect 102604 31934 103204 32018
rect 102604 31698 102786 31934
rect 103022 31698 103204 31934
rect 84604 -6222 84786 -5986
rect 85022 -6222 85204 -5986
rect 84604 -6306 85204 -6222
rect 84604 -6542 84786 -6306
rect 85022 -6542 85204 -6306
rect 84604 -7504 85204 -6542
rect 102604 -6926 103204 31698
rect 109804 704838 110404 705800
rect 109804 704602 109986 704838
rect 110222 704602 110404 704838
rect 109804 704518 110404 704602
rect 109804 704282 109986 704518
rect 110222 704282 110404 704518
rect 109804 687454 110404 704282
rect 109804 687218 109986 687454
rect 110222 687218 110404 687454
rect 109804 687134 110404 687218
rect 109804 686898 109986 687134
rect 110222 686898 110404 687134
rect 109804 651454 110404 686898
rect 109804 651218 109986 651454
rect 110222 651218 110404 651454
rect 109804 651134 110404 651218
rect 109804 650898 109986 651134
rect 110222 650898 110404 651134
rect 109804 615454 110404 650898
rect 109804 615218 109986 615454
rect 110222 615218 110404 615454
rect 109804 615134 110404 615218
rect 109804 614898 109986 615134
rect 110222 614898 110404 615134
rect 109804 579454 110404 614898
rect 109804 579218 109986 579454
rect 110222 579218 110404 579454
rect 109804 579134 110404 579218
rect 109804 578898 109986 579134
rect 110222 578898 110404 579134
rect 109804 543454 110404 578898
rect 109804 543218 109986 543454
rect 110222 543218 110404 543454
rect 109804 543134 110404 543218
rect 109804 542898 109986 543134
rect 110222 542898 110404 543134
rect 109804 507454 110404 542898
rect 109804 507218 109986 507454
rect 110222 507218 110404 507454
rect 109804 507134 110404 507218
rect 109804 506898 109986 507134
rect 110222 506898 110404 507134
rect 109804 471454 110404 506898
rect 109804 471218 109986 471454
rect 110222 471218 110404 471454
rect 109804 471134 110404 471218
rect 109804 470898 109986 471134
rect 110222 470898 110404 471134
rect 109804 435454 110404 470898
rect 109804 435218 109986 435454
rect 110222 435218 110404 435454
rect 109804 435134 110404 435218
rect 109804 434898 109986 435134
rect 110222 434898 110404 435134
rect 109804 399454 110404 434898
rect 109804 399218 109986 399454
rect 110222 399218 110404 399454
rect 109804 399134 110404 399218
rect 109804 398898 109986 399134
rect 110222 398898 110404 399134
rect 109804 363454 110404 398898
rect 109804 363218 109986 363454
rect 110222 363218 110404 363454
rect 109804 363134 110404 363218
rect 109804 362898 109986 363134
rect 110222 362898 110404 363134
rect 109804 327454 110404 362898
rect 109804 327218 109986 327454
rect 110222 327218 110404 327454
rect 109804 327134 110404 327218
rect 109804 326898 109986 327134
rect 110222 326898 110404 327134
rect 109804 291454 110404 326898
rect 109804 291218 109986 291454
rect 110222 291218 110404 291454
rect 109804 291134 110404 291218
rect 109804 290898 109986 291134
rect 110222 290898 110404 291134
rect 109804 255454 110404 290898
rect 109804 255218 109986 255454
rect 110222 255218 110404 255454
rect 109804 255134 110404 255218
rect 109804 254898 109986 255134
rect 110222 254898 110404 255134
rect 109804 219454 110404 254898
rect 109804 219218 109986 219454
rect 110222 219218 110404 219454
rect 109804 219134 110404 219218
rect 109804 218898 109986 219134
rect 110222 218898 110404 219134
rect 109804 183454 110404 218898
rect 109804 183218 109986 183454
rect 110222 183218 110404 183454
rect 109804 183134 110404 183218
rect 109804 182898 109986 183134
rect 110222 182898 110404 183134
rect 109804 147454 110404 182898
rect 109804 147218 109986 147454
rect 110222 147218 110404 147454
rect 109804 147134 110404 147218
rect 109804 146898 109986 147134
rect 110222 146898 110404 147134
rect 109804 111454 110404 146898
rect 109804 111218 109986 111454
rect 110222 111218 110404 111454
rect 109804 111134 110404 111218
rect 109804 110898 109986 111134
rect 110222 110898 110404 111134
rect 109804 75454 110404 110898
rect 109804 75218 109986 75454
rect 110222 75218 110404 75454
rect 109804 75134 110404 75218
rect 109804 74898 109986 75134
rect 110222 74898 110404 75134
rect 109804 39454 110404 74898
rect 109804 39218 109986 39454
rect 110222 39218 110404 39454
rect 109804 39134 110404 39218
rect 109804 38898 109986 39134
rect 110222 38898 110404 39134
rect 109804 3454 110404 38898
rect 109804 3218 109986 3454
rect 110222 3218 110404 3454
rect 109804 3134 110404 3218
rect 109804 2898 109986 3134
rect 110222 2898 110404 3134
rect 109804 -346 110404 2898
rect 109804 -582 109986 -346
rect 110222 -582 110404 -346
rect 109804 -666 110404 -582
rect 109804 -902 109986 -666
rect 110222 -902 110404 -666
rect 109804 -1864 110404 -902
rect 113404 691054 114004 706162
rect 113404 690818 113586 691054
rect 113822 690818 114004 691054
rect 113404 690734 114004 690818
rect 113404 690498 113586 690734
rect 113822 690498 114004 690734
rect 113404 655054 114004 690498
rect 113404 654818 113586 655054
rect 113822 654818 114004 655054
rect 113404 654734 114004 654818
rect 113404 654498 113586 654734
rect 113822 654498 114004 654734
rect 113404 619054 114004 654498
rect 113404 618818 113586 619054
rect 113822 618818 114004 619054
rect 113404 618734 114004 618818
rect 113404 618498 113586 618734
rect 113822 618498 114004 618734
rect 113404 583054 114004 618498
rect 113404 582818 113586 583054
rect 113822 582818 114004 583054
rect 113404 582734 114004 582818
rect 113404 582498 113586 582734
rect 113822 582498 114004 582734
rect 113404 547054 114004 582498
rect 113404 546818 113586 547054
rect 113822 546818 114004 547054
rect 113404 546734 114004 546818
rect 113404 546498 113586 546734
rect 113822 546498 114004 546734
rect 113404 511054 114004 546498
rect 113404 510818 113586 511054
rect 113822 510818 114004 511054
rect 113404 510734 114004 510818
rect 113404 510498 113586 510734
rect 113822 510498 114004 510734
rect 113404 475054 114004 510498
rect 113404 474818 113586 475054
rect 113822 474818 114004 475054
rect 113404 474734 114004 474818
rect 113404 474498 113586 474734
rect 113822 474498 114004 474734
rect 113404 439054 114004 474498
rect 113404 438818 113586 439054
rect 113822 438818 114004 439054
rect 113404 438734 114004 438818
rect 113404 438498 113586 438734
rect 113822 438498 114004 438734
rect 113404 403054 114004 438498
rect 113404 402818 113586 403054
rect 113822 402818 114004 403054
rect 113404 402734 114004 402818
rect 113404 402498 113586 402734
rect 113822 402498 114004 402734
rect 113404 367054 114004 402498
rect 113404 366818 113586 367054
rect 113822 366818 114004 367054
rect 113404 366734 114004 366818
rect 113404 366498 113586 366734
rect 113822 366498 114004 366734
rect 113404 331054 114004 366498
rect 113404 330818 113586 331054
rect 113822 330818 114004 331054
rect 113404 330734 114004 330818
rect 113404 330498 113586 330734
rect 113822 330498 114004 330734
rect 113404 295054 114004 330498
rect 113404 294818 113586 295054
rect 113822 294818 114004 295054
rect 113404 294734 114004 294818
rect 113404 294498 113586 294734
rect 113822 294498 114004 294734
rect 113404 259054 114004 294498
rect 113404 258818 113586 259054
rect 113822 258818 114004 259054
rect 113404 258734 114004 258818
rect 113404 258498 113586 258734
rect 113822 258498 114004 258734
rect 113404 223054 114004 258498
rect 113404 222818 113586 223054
rect 113822 222818 114004 223054
rect 113404 222734 114004 222818
rect 113404 222498 113586 222734
rect 113822 222498 114004 222734
rect 113404 187054 114004 222498
rect 113404 186818 113586 187054
rect 113822 186818 114004 187054
rect 113404 186734 114004 186818
rect 113404 186498 113586 186734
rect 113822 186498 114004 186734
rect 113404 151054 114004 186498
rect 113404 150818 113586 151054
rect 113822 150818 114004 151054
rect 113404 150734 114004 150818
rect 113404 150498 113586 150734
rect 113822 150498 114004 150734
rect 113404 115054 114004 150498
rect 113404 114818 113586 115054
rect 113822 114818 114004 115054
rect 113404 114734 114004 114818
rect 113404 114498 113586 114734
rect 113822 114498 114004 114734
rect 113404 79054 114004 114498
rect 113404 78818 113586 79054
rect 113822 78818 114004 79054
rect 113404 78734 114004 78818
rect 113404 78498 113586 78734
rect 113822 78498 114004 78734
rect 113404 43054 114004 78498
rect 113404 42818 113586 43054
rect 113822 42818 114004 43054
rect 113404 42734 114004 42818
rect 113404 42498 113586 42734
rect 113822 42498 114004 42734
rect 113404 7054 114004 42498
rect 113404 6818 113586 7054
rect 113822 6818 114004 7054
rect 113404 6734 114004 6818
rect 113404 6498 113586 6734
rect 113822 6498 114004 6734
rect 113404 -2226 114004 6498
rect 113404 -2462 113586 -2226
rect 113822 -2462 114004 -2226
rect 113404 -2546 114004 -2462
rect 113404 -2782 113586 -2546
rect 113822 -2782 114004 -2546
rect 113404 -3744 114004 -2782
rect 117004 694654 117604 708042
rect 117004 694418 117186 694654
rect 117422 694418 117604 694654
rect 117004 694334 117604 694418
rect 117004 694098 117186 694334
rect 117422 694098 117604 694334
rect 117004 658654 117604 694098
rect 117004 658418 117186 658654
rect 117422 658418 117604 658654
rect 117004 658334 117604 658418
rect 117004 658098 117186 658334
rect 117422 658098 117604 658334
rect 117004 622654 117604 658098
rect 117004 622418 117186 622654
rect 117422 622418 117604 622654
rect 117004 622334 117604 622418
rect 117004 622098 117186 622334
rect 117422 622098 117604 622334
rect 117004 586654 117604 622098
rect 117004 586418 117186 586654
rect 117422 586418 117604 586654
rect 117004 586334 117604 586418
rect 117004 586098 117186 586334
rect 117422 586098 117604 586334
rect 117004 550654 117604 586098
rect 117004 550418 117186 550654
rect 117422 550418 117604 550654
rect 117004 550334 117604 550418
rect 117004 550098 117186 550334
rect 117422 550098 117604 550334
rect 117004 514654 117604 550098
rect 117004 514418 117186 514654
rect 117422 514418 117604 514654
rect 117004 514334 117604 514418
rect 117004 514098 117186 514334
rect 117422 514098 117604 514334
rect 117004 478654 117604 514098
rect 117004 478418 117186 478654
rect 117422 478418 117604 478654
rect 117004 478334 117604 478418
rect 117004 478098 117186 478334
rect 117422 478098 117604 478334
rect 117004 442654 117604 478098
rect 117004 442418 117186 442654
rect 117422 442418 117604 442654
rect 117004 442334 117604 442418
rect 117004 442098 117186 442334
rect 117422 442098 117604 442334
rect 117004 406654 117604 442098
rect 117004 406418 117186 406654
rect 117422 406418 117604 406654
rect 117004 406334 117604 406418
rect 117004 406098 117186 406334
rect 117422 406098 117604 406334
rect 117004 370654 117604 406098
rect 117004 370418 117186 370654
rect 117422 370418 117604 370654
rect 117004 370334 117604 370418
rect 117004 370098 117186 370334
rect 117422 370098 117604 370334
rect 117004 334654 117604 370098
rect 117004 334418 117186 334654
rect 117422 334418 117604 334654
rect 117004 334334 117604 334418
rect 117004 334098 117186 334334
rect 117422 334098 117604 334334
rect 117004 298654 117604 334098
rect 117004 298418 117186 298654
rect 117422 298418 117604 298654
rect 117004 298334 117604 298418
rect 117004 298098 117186 298334
rect 117422 298098 117604 298334
rect 117004 262654 117604 298098
rect 117004 262418 117186 262654
rect 117422 262418 117604 262654
rect 117004 262334 117604 262418
rect 117004 262098 117186 262334
rect 117422 262098 117604 262334
rect 117004 226654 117604 262098
rect 117004 226418 117186 226654
rect 117422 226418 117604 226654
rect 117004 226334 117604 226418
rect 117004 226098 117186 226334
rect 117422 226098 117604 226334
rect 117004 190654 117604 226098
rect 117004 190418 117186 190654
rect 117422 190418 117604 190654
rect 117004 190334 117604 190418
rect 117004 190098 117186 190334
rect 117422 190098 117604 190334
rect 117004 154654 117604 190098
rect 117004 154418 117186 154654
rect 117422 154418 117604 154654
rect 117004 154334 117604 154418
rect 117004 154098 117186 154334
rect 117422 154098 117604 154334
rect 117004 118654 117604 154098
rect 117004 118418 117186 118654
rect 117422 118418 117604 118654
rect 117004 118334 117604 118418
rect 117004 118098 117186 118334
rect 117422 118098 117604 118334
rect 117004 82654 117604 118098
rect 117004 82418 117186 82654
rect 117422 82418 117604 82654
rect 117004 82334 117604 82418
rect 117004 82098 117186 82334
rect 117422 82098 117604 82334
rect 117004 46654 117604 82098
rect 117004 46418 117186 46654
rect 117422 46418 117604 46654
rect 117004 46334 117604 46418
rect 117004 46098 117186 46334
rect 117422 46098 117604 46334
rect 117004 10654 117604 46098
rect 117004 10418 117186 10654
rect 117422 10418 117604 10654
rect 117004 10334 117604 10418
rect 117004 10098 117186 10334
rect 117422 10098 117604 10334
rect 117004 -4106 117604 10098
rect 117004 -4342 117186 -4106
rect 117422 -4342 117604 -4106
rect 117004 -4426 117604 -4342
rect 117004 -4662 117186 -4426
rect 117422 -4662 117604 -4426
rect 117004 -5624 117604 -4662
rect 120604 698254 121204 709922
rect 138604 711418 139204 711440
rect 138604 711182 138786 711418
rect 139022 711182 139204 711418
rect 138604 711098 139204 711182
rect 138604 710862 138786 711098
rect 139022 710862 139204 711098
rect 135004 709538 135604 709560
rect 135004 709302 135186 709538
rect 135422 709302 135604 709538
rect 135004 709218 135604 709302
rect 135004 708982 135186 709218
rect 135422 708982 135604 709218
rect 131404 707658 132004 707680
rect 131404 707422 131586 707658
rect 131822 707422 132004 707658
rect 131404 707338 132004 707422
rect 131404 707102 131586 707338
rect 131822 707102 132004 707338
rect 120604 698018 120786 698254
rect 121022 698018 121204 698254
rect 120604 697934 121204 698018
rect 120604 697698 120786 697934
rect 121022 697698 121204 697934
rect 120604 662254 121204 697698
rect 120604 662018 120786 662254
rect 121022 662018 121204 662254
rect 120604 661934 121204 662018
rect 120604 661698 120786 661934
rect 121022 661698 121204 661934
rect 120604 626254 121204 661698
rect 120604 626018 120786 626254
rect 121022 626018 121204 626254
rect 120604 625934 121204 626018
rect 120604 625698 120786 625934
rect 121022 625698 121204 625934
rect 120604 590254 121204 625698
rect 120604 590018 120786 590254
rect 121022 590018 121204 590254
rect 120604 589934 121204 590018
rect 120604 589698 120786 589934
rect 121022 589698 121204 589934
rect 120604 554254 121204 589698
rect 120604 554018 120786 554254
rect 121022 554018 121204 554254
rect 120604 553934 121204 554018
rect 120604 553698 120786 553934
rect 121022 553698 121204 553934
rect 120604 518254 121204 553698
rect 120604 518018 120786 518254
rect 121022 518018 121204 518254
rect 120604 517934 121204 518018
rect 120604 517698 120786 517934
rect 121022 517698 121204 517934
rect 120604 482254 121204 517698
rect 120604 482018 120786 482254
rect 121022 482018 121204 482254
rect 120604 481934 121204 482018
rect 120604 481698 120786 481934
rect 121022 481698 121204 481934
rect 120604 446254 121204 481698
rect 120604 446018 120786 446254
rect 121022 446018 121204 446254
rect 120604 445934 121204 446018
rect 120604 445698 120786 445934
rect 121022 445698 121204 445934
rect 120604 410254 121204 445698
rect 120604 410018 120786 410254
rect 121022 410018 121204 410254
rect 120604 409934 121204 410018
rect 120604 409698 120786 409934
rect 121022 409698 121204 409934
rect 120604 374254 121204 409698
rect 120604 374018 120786 374254
rect 121022 374018 121204 374254
rect 120604 373934 121204 374018
rect 120604 373698 120786 373934
rect 121022 373698 121204 373934
rect 120604 338254 121204 373698
rect 120604 338018 120786 338254
rect 121022 338018 121204 338254
rect 120604 337934 121204 338018
rect 120604 337698 120786 337934
rect 121022 337698 121204 337934
rect 120604 302254 121204 337698
rect 120604 302018 120786 302254
rect 121022 302018 121204 302254
rect 120604 301934 121204 302018
rect 120604 301698 120786 301934
rect 121022 301698 121204 301934
rect 120604 266254 121204 301698
rect 120604 266018 120786 266254
rect 121022 266018 121204 266254
rect 120604 265934 121204 266018
rect 120604 265698 120786 265934
rect 121022 265698 121204 265934
rect 120604 230254 121204 265698
rect 120604 230018 120786 230254
rect 121022 230018 121204 230254
rect 120604 229934 121204 230018
rect 120604 229698 120786 229934
rect 121022 229698 121204 229934
rect 120604 194254 121204 229698
rect 120604 194018 120786 194254
rect 121022 194018 121204 194254
rect 120604 193934 121204 194018
rect 120604 193698 120786 193934
rect 121022 193698 121204 193934
rect 120604 158254 121204 193698
rect 120604 158018 120786 158254
rect 121022 158018 121204 158254
rect 120604 157934 121204 158018
rect 120604 157698 120786 157934
rect 121022 157698 121204 157934
rect 120604 122254 121204 157698
rect 120604 122018 120786 122254
rect 121022 122018 121204 122254
rect 120604 121934 121204 122018
rect 120604 121698 120786 121934
rect 121022 121698 121204 121934
rect 120604 86254 121204 121698
rect 120604 86018 120786 86254
rect 121022 86018 121204 86254
rect 120604 85934 121204 86018
rect 120604 85698 120786 85934
rect 121022 85698 121204 85934
rect 120604 50254 121204 85698
rect 120604 50018 120786 50254
rect 121022 50018 121204 50254
rect 120604 49934 121204 50018
rect 120604 49698 120786 49934
rect 121022 49698 121204 49934
rect 120604 14254 121204 49698
rect 120604 14018 120786 14254
rect 121022 14018 121204 14254
rect 120604 13934 121204 14018
rect 120604 13698 120786 13934
rect 121022 13698 121204 13934
rect 102604 -7162 102786 -6926
rect 103022 -7162 103204 -6926
rect 102604 -7246 103204 -7162
rect 102604 -7482 102786 -7246
rect 103022 -7482 103204 -7246
rect 102604 -7504 103204 -7482
rect 120604 -5986 121204 13698
rect 127804 705778 128404 705800
rect 127804 705542 127986 705778
rect 128222 705542 128404 705778
rect 127804 705458 128404 705542
rect 127804 705222 127986 705458
rect 128222 705222 128404 705458
rect 127804 669454 128404 705222
rect 127804 669218 127986 669454
rect 128222 669218 128404 669454
rect 127804 669134 128404 669218
rect 127804 668898 127986 669134
rect 128222 668898 128404 669134
rect 127804 633454 128404 668898
rect 127804 633218 127986 633454
rect 128222 633218 128404 633454
rect 127804 633134 128404 633218
rect 127804 632898 127986 633134
rect 128222 632898 128404 633134
rect 127804 597454 128404 632898
rect 127804 597218 127986 597454
rect 128222 597218 128404 597454
rect 127804 597134 128404 597218
rect 127804 596898 127986 597134
rect 128222 596898 128404 597134
rect 127804 561454 128404 596898
rect 127804 561218 127986 561454
rect 128222 561218 128404 561454
rect 127804 561134 128404 561218
rect 127804 560898 127986 561134
rect 128222 560898 128404 561134
rect 127804 525454 128404 560898
rect 127804 525218 127986 525454
rect 128222 525218 128404 525454
rect 127804 525134 128404 525218
rect 127804 524898 127986 525134
rect 128222 524898 128404 525134
rect 127804 489454 128404 524898
rect 127804 489218 127986 489454
rect 128222 489218 128404 489454
rect 127804 489134 128404 489218
rect 127804 488898 127986 489134
rect 128222 488898 128404 489134
rect 127804 453454 128404 488898
rect 127804 453218 127986 453454
rect 128222 453218 128404 453454
rect 127804 453134 128404 453218
rect 127804 452898 127986 453134
rect 128222 452898 128404 453134
rect 127804 417454 128404 452898
rect 127804 417218 127986 417454
rect 128222 417218 128404 417454
rect 127804 417134 128404 417218
rect 127804 416898 127986 417134
rect 128222 416898 128404 417134
rect 127804 381454 128404 416898
rect 127804 381218 127986 381454
rect 128222 381218 128404 381454
rect 127804 381134 128404 381218
rect 127804 380898 127986 381134
rect 128222 380898 128404 381134
rect 127804 345454 128404 380898
rect 127804 345218 127986 345454
rect 128222 345218 128404 345454
rect 127804 345134 128404 345218
rect 127804 344898 127986 345134
rect 128222 344898 128404 345134
rect 127804 309454 128404 344898
rect 127804 309218 127986 309454
rect 128222 309218 128404 309454
rect 127804 309134 128404 309218
rect 127804 308898 127986 309134
rect 128222 308898 128404 309134
rect 127804 273454 128404 308898
rect 127804 273218 127986 273454
rect 128222 273218 128404 273454
rect 127804 273134 128404 273218
rect 127804 272898 127986 273134
rect 128222 272898 128404 273134
rect 127804 237454 128404 272898
rect 127804 237218 127986 237454
rect 128222 237218 128404 237454
rect 127804 237134 128404 237218
rect 127804 236898 127986 237134
rect 128222 236898 128404 237134
rect 127804 201454 128404 236898
rect 127804 201218 127986 201454
rect 128222 201218 128404 201454
rect 127804 201134 128404 201218
rect 127804 200898 127986 201134
rect 128222 200898 128404 201134
rect 127804 165454 128404 200898
rect 127804 165218 127986 165454
rect 128222 165218 128404 165454
rect 127804 165134 128404 165218
rect 127804 164898 127986 165134
rect 128222 164898 128404 165134
rect 127804 129454 128404 164898
rect 127804 129218 127986 129454
rect 128222 129218 128404 129454
rect 127804 129134 128404 129218
rect 127804 128898 127986 129134
rect 128222 128898 128404 129134
rect 127804 93454 128404 128898
rect 127804 93218 127986 93454
rect 128222 93218 128404 93454
rect 127804 93134 128404 93218
rect 127804 92898 127986 93134
rect 128222 92898 128404 93134
rect 127804 57454 128404 92898
rect 127804 57218 127986 57454
rect 128222 57218 128404 57454
rect 127804 57134 128404 57218
rect 127804 56898 127986 57134
rect 128222 56898 128404 57134
rect 127804 21454 128404 56898
rect 127804 21218 127986 21454
rect 128222 21218 128404 21454
rect 127804 21134 128404 21218
rect 127804 20898 127986 21134
rect 128222 20898 128404 21134
rect 127804 -1286 128404 20898
rect 127804 -1522 127986 -1286
rect 128222 -1522 128404 -1286
rect 127804 -1606 128404 -1522
rect 127804 -1842 127986 -1606
rect 128222 -1842 128404 -1606
rect 127804 -1864 128404 -1842
rect 131404 673054 132004 707102
rect 131404 672818 131586 673054
rect 131822 672818 132004 673054
rect 131404 672734 132004 672818
rect 131404 672498 131586 672734
rect 131822 672498 132004 672734
rect 131404 637054 132004 672498
rect 131404 636818 131586 637054
rect 131822 636818 132004 637054
rect 131404 636734 132004 636818
rect 131404 636498 131586 636734
rect 131822 636498 132004 636734
rect 131404 601054 132004 636498
rect 131404 600818 131586 601054
rect 131822 600818 132004 601054
rect 131404 600734 132004 600818
rect 131404 600498 131586 600734
rect 131822 600498 132004 600734
rect 131404 565054 132004 600498
rect 131404 564818 131586 565054
rect 131822 564818 132004 565054
rect 131404 564734 132004 564818
rect 131404 564498 131586 564734
rect 131822 564498 132004 564734
rect 131404 529054 132004 564498
rect 131404 528818 131586 529054
rect 131822 528818 132004 529054
rect 131404 528734 132004 528818
rect 131404 528498 131586 528734
rect 131822 528498 132004 528734
rect 131404 493054 132004 528498
rect 131404 492818 131586 493054
rect 131822 492818 132004 493054
rect 131404 492734 132004 492818
rect 131404 492498 131586 492734
rect 131822 492498 132004 492734
rect 131404 457054 132004 492498
rect 131404 456818 131586 457054
rect 131822 456818 132004 457054
rect 131404 456734 132004 456818
rect 131404 456498 131586 456734
rect 131822 456498 132004 456734
rect 131404 421054 132004 456498
rect 131404 420818 131586 421054
rect 131822 420818 132004 421054
rect 131404 420734 132004 420818
rect 131404 420498 131586 420734
rect 131822 420498 132004 420734
rect 131404 385054 132004 420498
rect 131404 384818 131586 385054
rect 131822 384818 132004 385054
rect 131404 384734 132004 384818
rect 131404 384498 131586 384734
rect 131822 384498 132004 384734
rect 131404 349054 132004 384498
rect 131404 348818 131586 349054
rect 131822 348818 132004 349054
rect 131404 348734 132004 348818
rect 131404 348498 131586 348734
rect 131822 348498 132004 348734
rect 131404 313054 132004 348498
rect 131404 312818 131586 313054
rect 131822 312818 132004 313054
rect 131404 312734 132004 312818
rect 131404 312498 131586 312734
rect 131822 312498 132004 312734
rect 131404 277054 132004 312498
rect 131404 276818 131586 277054
rect 131822 276818 132004 277054
rect 131404 276734 132004 276818
rect 131404 276498 131586 276734
rect 131822 276498 132004 276734
rect 131404 241054 132004 276498
rect 131404 240818 131586 241054
rect 131822 240818 132004 241054
rect 131404 240734 132004 240818
rect 131404 240498 131586 240734
rect 131822 240498 132004 240734
rect 131404 205054 132004 240498
rect 131404 204818 131586 205054
rect 131822 204818 132004 205054
rect 131404 204734 132004 204818
rect 131404 204498 131586 204734
rect 131822 204498 132004 204734
rect 131404 169054 132004 204498
rect 131404 168818 131586 169054
rect 131822 168818 132004 169054
rect 131404 168734 132004 168818
rect 131404 168498 131586 168734
rect 131822 168498 132004 168734
rect 131404 133054 132004 168498
rect 131404 132818 131586 133054
rect 131822 132818 132004 133054
rect 131404 132734 132004 132818
rect 131404 132498 131586 132734
rect 131822 132498 132004 132734
rect 131404 97054 132004 132498
rect 131404 96818 131586 97054
rect 131822 96818 132004 97054
rect 131404 96734 132004 96818
rect 131404 96498 131586 96734
rect 131822 96498 132004 96734
rect 131404 61054 132004 96498
rect 131404 60818 131586 61054
rect 131822 60818 132004 61054
rect 131404 60734 132004 60818
rect 131404 60498 131586 60734
rect 131822 60498 132004 60734
rect 131404 25054 132004 60498
rect 131404 24818 131586 25054
rect 131822 24818 132004 25054
rect 131404 24734 132004 24818
rect 131404 24498 131586 24734
rect 131822 24498 132004 24734
rect 131404 -3166 132004 24498
rect 131404 -3402 131586 -3166
rect 131822 -3402 132004 -3166
rect 131404 -3486 132004 -3402
rect 131404 -3722 131586 -3486
rect 131822 -3722 132004 -3486
rect 131404 -3744 132004 -3722
rect 135004 676654 135604 708982
rect 135004 676418 135186 676654
rect 135422 676418 135604 676654
rect 135004 676334 135604 676418
rect 135004 676098 135186 676334
rect 135422 676098 135604 676334
rect 135004 640654 135604 676098
rect 135004 640418 135186 640654
rect 135422 640418 135604 640654
rect 135004 640334 135604 640418
rect 135004 640098 135186 640334
rect 135422 640098 135604 640334
rect 135004 604654 135604 640098
rect 135004 604418 135186 604654
rect 135422 604418 135604 604654
rect 135004 604334 135604 604418
rect 135004 604098 135186 604334
rect 135422 604098 135604 604334
rect 135004 568654 135604 604098
rect 135004 568418 135186 568654
rect 135422 568418 135604 568654
rect 135004 568334 135604 568418
rect 135004 568098 135186 568334
rect 135422 568098 135604 568334
rect 135004 532654 135604 568098
rect 135004 532418 135186 532654
rect 135422 532418 135604 532654
rect 135004 532334 135604 532418
rect 135004 532098 135186 532334
rect 135422 532098 135604 532334
rect 135004 496654 135604 532098
rect 135004 496418 135186 496654
rect 135422 496418 135604 496654
rect 135004 496334 135604 496418
rect 135004 496098 135186 496334
rect 135422 496098 135604 496334
rect 135004 460654 135604 496098
rect 135004 460418 135186 460654
rect 135422 460418 135604 460654
rect 135004 460334 135604 460418
rect 135004 460098 135186 460334
rect 135422 460098 135604 460334
rect 135004 424654 135604 460098
rect 135004 424418 135186 424654
rect 135422 424418 135604 424654
rect 135004 424334 135604 424418
rect 135004 424098 135186 424334
rect 135422 424098 135604 424334
rect 135004 388654 135604 424098
rect 135004 388418 135186 388654
rect 135422 388418 135604 388654
rect 135004 388334 135604 388418
rect 135004 388098 135186 388334
rect 135422 388098 135604 388334
rect 135004 352654 135604 388098
rect 135004 352418 135186 352654
rect 135422 352418 135604 352654
rect 135004 352334 135604 352418
rect 135004 352098 135186 352334
rect 135422 352098 135604 352334
rect 135004 316654 135604 352098
rect 135004 316418 135186 316654
rect 135422 316418 135604 316654
rect 135004 316334 135604 316418
rect 135004 316098 135186 316334
rect 135422 316098 135604 316334
rect 135004 280654 135604 316098
rect 135004 280418 135186 280654
rect 135422 280418 135604 280654
rect 135004 280334 135604 280418
rect 135004 280098 135186 280334
rect 135422 280098 135604 280334
rect 135004 244654 135604 280098
rect 135004 244418 135186 244654
rect 135422 244418 135604 244654
rect 135004 244334 135604 244418
rect 135004 244098 135186 244334
rect 135422 244098 135604 244334
rect 135004 208654 135604 244098
rect 135004 208418 135186 208654
rect 135422 208418 135604 208654
rect 135004 208334 135604 208418
rect 135004 208098 135186 208334
rect 135422 208098 135604 208334
rect 135004 172654 135604 208098
rect 135004 172418 135186 172654
rect 135422 172418 135604 172654
rect 135004 172334 135604 172418
rect 135004 172098 135186 172334
rect 135422 172098 135604 172334
rect 135004 136654 135604 172098
rect 135004 136418 135186 136654
rect 135422 136418 135604 136654
rect 135004 136334 135604 136418
rect 135004 136098 135186 136334
rect 135422 136098 135604 136334
rect 135004 100654 135604 136098
rect 135004 100418 135186 100654
rect 135422 100418 135604 100654
rect 135004 100334 135604 100418
rect 135004 100098 135186 100334
rect 135422 100098 135604 100334
rect 135004 64654 135604 100098
rect 135004 64418 135186 64654
rect 135422 64418 135604 64654
rect 135004 64334 135604 64418
rect 135004 64098 135186 64334
rect 135422 64098 135604 64334
rect 135004 28654 135604 64098
rect 135004 28418 135186 28654
rect 135422 28418 135604 28654
rect 135004 28334 135604 28418
rect 135004 28098 135186 28334
rect 135422 28098 135604 28334
rect 135004 -5046 135604 28098
rect 135004 -5282 135186 -5046
rect 135422 -5282 135604 -5046
rect 135004 -5366 135604 -5282
rect 135004 -5602 135186 -5366
rect 135422 -5602 135604 -5366
rect 135004 -5624 135604 -5602
rect 138604 680254 139204 710862
rect 156604 710478 157204 711440
rect 156604 710242 156786 710478
rect 157022 710242 157204 710478
rect 156604 710158 157204 710242
rect 156604 709922 156786 710158
rect 157022 709922 157204 710158
rect 153004 708598 153604 709560
rect 153004 708362 153186 708598
rect 153422 708362 153604 708598
rect 153004 708278 153604 708362
rect 153004 708042 153186 708278
rect 153422 708042 153604 708278
rect 149404 706718 150004 707680
rect 149404 706482 149586 706718
rect 149822 706482 150004 706718
rect 149404 706398 150004 706482
rect 149404 706162 149586 706398
rect 149822 706162 150004 706398
rect 138604 680018 138786 680254
rect 139022 680018 139204 680254
rect 138604 679934 139204 680018
rect 138604 679698 138786 679934
rect 139022 679698 139204 679934
rect 138604 644254 139204 679698
rect 138604 644018 138786 644254
rect 139022 644018 139204 644254
rect 138604 643934 139204 644018
rect 138604 643698 138786 643934
rect 139022 643698 139204 643934
rect 138604 608254 139204 643698
rect 138604 608018 138786 608254
rect 139022 608018 139204 608254
rect 138604 607934 139204 608018
rect 138604 607698 138786 607934
rect 139022 607698 139204 607934
rect 138604 572254 139204 607698
rect 138604 572018 138786 572254
rect 139022 572018 139204 572254
rect 138604 571934 139204 572018
rect 138604 571698 138786 571934
rect 139022 571698 139204 571934
rect 138604 536254 139204 571698
rect 138604 536018 138786 536254
rect 139022 536018 139204 536254
rect 138604 535934 139204 536018
rect 138604 535698 138786 535934
rect 139022 535698 139204 535934
rect 138604 500254 139204 535698
rect 138604 500018 138786 500254
rect 139022 500018 139204 500254
rect 138604 499934 139204 500018
rect 138604 499698 138786 499934
rect 139022 499698 139204 499934
rect 138604 464254 139204 499698
rect 138604 464018 138786 464254
rect 139022 464018 139204 464254
rect 138604 463934 139204 464018
rect 138604 463698 138786 463934
rect 139022 463698 139204 463934
rect 138604 428254 139204 463698
rect 138604 428018 138786 428254
rect 139022 428018 139204 428254
rect 138604 427934 139204 428018
rect 138604 427698 138786 427934
rect 139022 427698 139204 427934
rect 138604 392254 139204 427698
rect 138604 392018 138786 392254
rect 139022 392018 139204 392254
rect 138604 391934 139204 392018
rect 138604 391698 138786 391934
rect 139022 391698 139204 391934
rect 138604 356254 139204 391698
rect 138604 356018 138786 356254
rect 139022 356018 139204 356254
rect 138604 355934 139204 356018
rect 138604 355698 138786 355934
rect 139022 355698 139204 355934
rect 138604 320254 139204 355698
rect 138604 320018 138786 320254
rect 139022 320018 139204 320254
rect 138604 319934 139204 320018
rect 138604 319698 138786 319934
rect 139022 319698 139204 319934
rect 138604 284254 139204 319698
rect 138604 284018 138786 284254
rect 139022 284018 139204 284254
rect 138604 283934 139204 284018
rect 138604 283698 138786 283934
rect 139022 283698 139204 283934
rect 138604 248254 139204 283698
rect 138604 248018 138786 248254
rect 139022 248018 139204 248254
rect 138604 247934 139204 248018
rect 138604 247698 138786 247934
rect 139022 247698 139204 247934
rect 138604 212254 139204 247698
rect 138604 212018 138786 212254
rect 139022 212018 139204 212254
rect 138604 211934 139204 212018
rect 138604 211698 138786 211934
rect 139022 211698 139204 211934
rect 138604 176254 139204 211698
rect 138604 176018 138786 176254
rect 139022 176018 139204 176254
rect 138604 175934 139204 176018
rect 138604 175698 138786 175934
rect 139022 175698 139204 175934
rect 138604 140254 139204 175698
rect 138604 140018 138786 140254
rect 139022 140018 139204 140254
rect 138604 139934 139204 140018
rect 138604 139698 138786 139934
rect 139022 139698 139204 139934
rect 138604 104254 139204 139698
rect 138604 104018 138786 104254
rect 139022 104018 139204 104254
rect 138604 103934 139204 104018
rect 138604 103698 138786 103934
rect 139022 103698 139204 103934
rect 138604 68254 139204 103698
rect 138604 68018 138786 68254
rect 139022 68018 139204 68254
rect 138604 67934 139204 68018
rect 138604 67698 138786 67934
rect 139022 67698 139204 67934
rect 138604 32254 139204 67698
rect 138604 32018 138786 32254
rect 139022 32018 139204 32254
rect 138604 31934 139204 32018
rect 138604 31698 138786 31934
rect 139022 31698 139204 31934
rect 120604 -6222 120786 -5986
rect 121022 -6222 121204 -5986
rect 120604 -6306 121204 -6222
rect 120604 -6542 120786 -6306
rect 121022 -6542 121204 -6306
rect 120604 -7504 121204 -6542
rect 138604 -6926 139204 31698
rect 145804 704838 146404 705800
rect 145804 704602 145986 704838
rect 146222 704602 146404 704838
rect 145804 704518 146404 704602
rect 145804 704282 145986 704518
rect 146222 704282 146404 704518
rect 145804 687454 146404 704282
rect 145804 687218 145986 687454
rect 146222 687218 146404 687454
rect 145804 687134 146404 687218
rect 145804 686898 145986 687134
rect 146222 686898 146404 687134
rect 145804 651454 146404 686898
rect 145804 651218 145986 651454
rect 146222 651218 146404 651454
rect 145804 651134 146404 651218
rect 145804 650898 145986 651134
rect 146222 650898 146404 651134
rect 145804 615454 146404 650898
rect 145804 615218 145986 615454
rect 146222 615218 146404 615454
rect 145804 615134 146404 615218
rect 145804 614898 145986 615134
rect 146222 614898 146404 615134
rect 145804 579454 146404 614898
rect 145804 579218 145986 579454
rect 146222 579218 146404 579454
rect 145804 579134 146404 579218
rect 145804 578898 145986 579134
rect 146222 578898 146404 579134
rect 145804 543454 146404 578898
rect 145804 543218 145986 543454
rect 146222 543218 146404 543454
rect 145804 543134 146404 543218
rect 145804 542898 145986 543134
rect 146222 542898 146404 543134
rect 145804 507454 146404 542898
rect 145804 507218 145986 507454
rect 146222 507218 146404 507454
rect 145804 507134 146404 507218
rect 145804 506898 145986 507134
rect 146222 506898 146404 507134
rect 145804 471454 146404 506898
rect 145804 471218 145986 471454
rect 146222 471218 146404 471454
rect 145804 471134 146404 471218
rect 145804 470898 145986 471134
rect 146222 470898 146404 471134
rect 145804 435454 146404 470898
rect 145804 435218 145986 435454
rect 146222 435218 146404 435454
rect 145804 435134 146404 435218
rect 145804 434898 145986 435134
rect 146222 434898 146404 435134
rect 145804 399454 146404 434898
rect 145804 399218 145986 399454
rect 146222 399218 146404 399454
rect 145804 399134 146404 399218
rect 145804 398898 145986 399134
rect 146222 398898 146404 399134
rect 145804 363454 146404 398898
rect 145804 363218 145986 363454
rect 146222 363218 146404 363454
rect 145804 363134 146404 363218
rect 145804 362898 145986 363134
rect 146222 362898 146404 363134
rect 145804 327454 146404 362898
rect 145804 327218 145986 327454
rect 146222 327218 146404 327454
rect 145804 327134 146404 327218
rect 145804 326898 145986 327134
rect 146222 326898 146404 327134
rect 145804 291454 146404 326898
rect 145804 291218 145986 291454
rect 146222 291218 146404 291454
rect 145804 291134 146404 291218
rect 145804 290898 145986 291134
rect 146222 290898 146404 291134
rect 145804 255454 146404 290898
rect 145804 255218 145986 255454
rect 146222 255218 146404 255454
rect 145804 255134 146404 255218
rect 145804 254898 145986 255134
rect 146222 254898 146404 255134
rect 145804 219454 146404 254898
rect 145804 219218 145986 219454
rect 146222 219218 146404 219454
rect 145804 219134 146404 219218
rect 145804 218898 145986 219134
rect 146222 218898 146404 219134
rect 145804 183454 146404 218898
rect 145804 183218 145986 183454
rect 146222 183218 146404 183454
rect 145804 183134 146404 183218
rect 145804 182898 145986 183134
rect 146222 182898 146404 183134
rect 145804 147454 146404 182898
rect 145804 147218 145986 147454
rect 146222 147218 146404 147454
rect 145804 147134 146404 147218
rect 145804 146898 145986 147134
rect 146222 146898 146404 147134
rect 145804 111454 146404 146898
rect 145804 111218 145986 111454
rect 146222 111218 146404 111454
rect 145804 111134 146404 111218
rect 145804 110898 145986 111134
rect 146222 110898 146404 111134
rect 145804 75454 146404 110898
rect 145804 75218 145986 75454
rect 146222 75218 146404 75454
rect 145804 75134 146404 75218
rect 145804 74898 145986 75134
rect 146222 74898 146404 75134
rect 145804 39454 146404 74898
rect 145804 39218 145986 39454
rect 146222 39218 146404 39454
rect 145804 39134 146404 39218
rect 145804 38898 145986 39134
rect 146222 38898 146404 39134
rect 145804 3454 146404 38898
rect 145804 3218 145986 3454
rect 146222 3218 146404 3454
rect 145804 3134 146404 3218
rect 145804 2898 145986 3134
rect 146222 2898 146404 3134
rect 145804 -346 146404 2898
rect 145804 -582 145986 -346
rect 146222 -582 146404 -346
rect 145804 -666 146404 -582
rect 145804 -902 145986 -666
rect 146222 -902 146404 -666
rect 145804 -1864 146404 -902
rect 149404 691054 150004 706162
rect 149404 690818 149586 691054
rect 149822 690818 150004 691054
rect 149404 690734 150004 690818
rect 149404 690498 149586 690734
rect 149822 690498 150004 690734
rect 149404 655054 150004 690498
rect 149404 654818 149586 655054
rect 149822 654818 150004 655054
rect 149404 654734 150004 654818
rect 149404 654498 149586 654734
rect 149822 654498 150004 654734
rect 149404 619054 150004 654498
rect 149404 618818 149586 619054
rect 149822 618818 150004 619054
rect 149404 618734 150004 618818
rect 149404 618498 149586 618734
rect 149822 618498 150004 618734
rect 149404 583054 150004 618498
rect 149404 582818 149586 583054
rect 149822 582818 150004 583054
rect 149404 582734 150004 582818
rect 149404 582498 149586 582734
rect 149822 582498 150004 582734
rect 149404 547054 150004 582498
rect 149404 546818 149586 547054
rect 149822 546818 150004 547054
rect 149404 546734 150004 546818
rect 149404 546498 149586 546734
rect 149822 546498 150004 546734
rect 149404 511054 150004 546498
rect 149404 510818 149586 511054
rect 149822 510818 150004 511054
rect 149404 510734 150004 510818
rect 149404 510498 149586 510734
rect 149822 510498 150004 510734
rect 149404 475054 150004 510498
rect 149404 474818 149586 475054
rect 149822 474818 150004 475054
rect 149404 474734 150004 474818
rect 149404 474498 149586 474734
rect 149822 474498 150004 474734
rect 149404 439054 150004 474498
rect 149404 438818 149586 439054
rect 149822 438818 150004 439054
rect 149404 438734 150004 438818
rect 149404 438498 149586 438734
rect 149822 438498 150004 438734
rect 149404 403054 150004 438498
rect 149404 402818 149586 403054
rect 149822 402818 150004 403054
rect 149404 402734 150004 402818
rect 149404 402498 149586 402734
rect 149822 402498 150004 402734
rect 149404 367054 150004 402498
rect 149404 366818 149586 367054
rect 149822 366818 150004 367054
rect 149404 366734 150004 366818
rect 149404 366498 149586 366734
rect 149822 366498 150004 366734
rect 149404 331054 150004 366498
rect 149404 330818 149586 331054
rect 149822 330818 150004 331054
rect 149404 330734 150004 330818
rect 149404 330498 149586 330734
rect 149822 330498 150004 330734
rect 149404 295054 150004 330498
rect 149404 294818 149586 295054
rect 149822 294818 150004 295054
rect 149404 294734 150004 294818
rect 149404 294498 149586 294734
rect 149822 294498 150004 294734
rect 149404 259054 150004 294498
rect 149404 258818 149586 259054
rect 149822 258818 150004 259054
rect 149404 258734 150004 258818
rect 149404 258498 149586 258734
rect 149822 258498 150004 258734
rect 149404 223054 150004 258498
rect 149404 222818 149586 223054
rect 149822 222818 150004 223054
rect 149404 222734 150004 222818
rect 149404 222498 149586 222734
rect 149822 222498 150004 222734
rect 149404 187054 150004 222498
rect 149404 186818 149586 187054
rect 149822 186818 150004 187054
rect 149404 186734 150004 186818
rect 149404 186498 149586 186734
rect 149822 186498 150004 186734
rect 149404 151054 150004 186498
rect 149404 150818 149586 151054
rect 149822 150818 150004 151054
rect 149404 150734 150004 150818
rect 149404 150498 149586 150734
rect 149822 150498 150004 150734
rect 149404 115054 150004 150498
rect 149404 114818 149586 115054
rect 149822 114818 150004 115054
rect 149404 114734 150004 114818
rect 149404 114498 149586 114734
rect 149822 114498 150004 114734
rect 149404 79054 150004 114498
rect 149404 78818 149586 79054
rect 149822 78818 150004 79054
rect 149404 78734 150004 78818
rect 149404 78498 149586 78734
rect 149822 78498 150004 78734
rect 149404 43054 150004 78498
rect 149404 42818 149586 43054
rect 149822 42818 150004 43054
rect 149404 42734 150004 42818
rect 149404 42498 149586 42734
rect 149822 42498 150004 42734
rect 149404 7054 150004 42498
rect 149404 6818 149586 7054
rect 149822 6818 150004 7054
rect 149404 6734 150004 6818
rect 149404 6498 149586 6734
rect 149822 6498 150004 6734
rect 149404 -2226 150004 6498
rect 149404 -2462 149586 -2226
rect 149822 -2462 150004 -2226
rect 149404 -2546 150004 -2462
rect 149404 -2782 149586 -2546
rect 149822 -2782 150004 -2546
rect 149404 -3744 150004 -2782
rect 153004 694654 153604 708042
rect 153004 694418 153186 694654
rect 153422 694418 153604 694654
rect 153004 694334 153604 694418
rect 153004 694098 153186 694334
rect 153422 694098 153604 694334
rect 153004 658654 153604 694098
rect 153004 658418 153186 658654
rect 153422 658418 153604 658654
rect 153004 658334 153604 658418
rect 153004 658098 153186 658334
rect 153422 658098 153604 658334
rect 153004 622654 153604 658098
rect 153004 622418 153186 622654
rect 153422 622418 153604 622654
rect 153004 622334 153604 622418
rect 153004 622098 153186 622334
rect 153422 622098 153604 622334
rect 153004 586654 153604 622098
rect 153004 586418 153186 586654
rect 153422 586418 153604 586654
rect 153004 586334 153604 586418
rect 153004 586098 153186 586334
rect 153422 586098 153604 586334
rect 153004 550654 153604 586098
rect 153004 550418 153186 550654
rect 153422 550418 153604 550654
rect 153004 550334 153604 550418
rect 153004 550098 153186 550334
rect 153422 550098 153604 550334
rect 153004 514654 153604 550098
rect 153004 514418 153186 514654
rect 153422 514418 153604 514654
rect 153004 514334 153604 514418
rect 153004 514098 153186 514334
rect 153422 514098 153604 514334
rect 153004 478654 153604 514098
rect 156604 698254 157204 709922
rect 174604 711418 175204 711440
rect 174604 711182 174786 711418
rect 175022 711182 175204 711418
rect 174604 711098 175204 711182
rect 174604 710862 174786 711098
rect 175022 710862 175204 711098
rect 171004 709538 171604 709560
rect 171004 709302 171186 709538
rect 171422 709302 171604 709538
rect 171004 709218 171604 709302
rect 171004 708982 171186 709218
rect 171422 708982 171604 709218
rect 167404 707658 168004 707680
rect 167404 707422 167586 707658
rect 167822 707422 168004 707658
rect 167404 707338 168004 707422
rect 167404 707102 167586 707338
rect 167822 707102 168004 707338
rect 156604 698018 156786 698254
rect 157022 698018 157204 698254
rect 156604 697934 157204 698018
rect 156604 697698 156786 697934
rect 157022 697698 157204 697934
rect 156604 662254 157204 697698
rect 156604 662018 156786 662254
rect 157022 662018 157204 662254
rect 156604 661934 157204 662018
rect 156604 661698 156786 661934
rect 157022 661698 157204 661934
rect 156604 626254 157204 661698
rect 156604 626018 156786 626254
rect 157022 626018 157204 626254
rect 156604 625934 157204 626018
rect 156604 625698 156786 625934
rect 157022 625698 157204 625934
rect 156604 590254 157204 625698
rect 156604 590018 156786 590254
rect 157022 590018 157204 590254
rect 156604 589934 157204 590018
rect 156604 589698 156786 589934
rect 157022 589698 157204 589934
rect 156604 554254 157204 589698
rect 156604 554018 156786 554254
rect 157022 554018 157204 554254
rect 156604 553934 157204 554018
rect 156604 553698 156786 553934
rect 157022 553698 157204 553934
rect 156604 518254 157204 553698
rect 156604 518018 156786 518254
rect 157022 518018 157204 518254
rect 156604 517934 157204 518018
rect 156604 517698 156786 517934
rect 157022 517698 157204 517934
rect 156604 510000 157204 517698
rect 163804 705778 164404 705800
rect 163804 705542 163986 705778
rect 164222 705542 164404 705778
rect 163804 705458 164404 705542
rect 163804 705222 163986 705458
rect 164222 705222 164404 705458
rect 163804 669454 164404 705222
rect 163804 669218 163986 669454
rect 164222 669218 164404 669454
rect 163804 669134 164404 669218
rect 163804 668898 163986 669134
rect 164222 668898 164404 669134
rect 163804 633454 164404 668898
rect 163804 633218 163986 633454
rect 164222 633218 164404 633454
rect 163804 633134 164404 633218
rect 163804 632898 163986 633134
rect 164222 632898 164404 633134
rect 163804 597454 164404 632898
rect 163804 597218 163986 597454
rect 164222 597218 164404 597454
rect 163804 597134 164404 597218
rect 163804 596898 163986 597134
rect 164222 596898 164404 597134
rect 163804 561454 164404 596898
rect 163804 561218 163986 561454
rect 164222 561218 164404 561454
rect 163804 561134 164404 561218
rect 163804 560898 163986 561134
rect 164222 560898 164404 561134
rect 163804 525454 164404 560898
rect 163804 525218 163986 525454
rect 164222 525218 164404 525454
rect 163804 525134 164404 525218
rect 163804 524898 163986 525134
rect 164222 524898 164404 525134
rect 163804 510000 164404 524898
rect 167404 673054 168004 707102
rect 167404 672818 167586 673054
rect 167822 672818 168004 673054
rect 167404 672734 168004 672818
rect 167404 672498 167586 672734
rect 167822 672498 168004 672734
rect 167404 637054 168004 672498
rect 167404 636818 167586 637054
rect 167822 636818 168004 637054
rect 167404 636734 168004 636818
rect 167404 636498 167586 636734
rect 167822 636498 168004 636734
rect 167404 601054 168004 636498
rect 167404 600818 167586 601054
rect 167822 600818 168004 601054
rect 167404 600734 168004 600818
rect 167404 600498 167586 600734
rect 167822 600498 168004 600734
rect 167404 565054 168004 600498
rect 167404 564818 167586 565054
rect 167822 564818 168004 565054
rect 167404 564734 168004 564818
rect 167404 564498 167586 564734
rect 167822 564498 168004 564734
rect 167404 529054 168004 564498
rect 167404 528818 167586 529054
rect 167822 528818 168004 529054
rect 167404 528734 168004 528818
rect 167404 528498 167586 528734
rect 167822 528498 168004 528734
rect 167404 510000 168004 528498
rect 171004 676654 171604 708982
rect 171004 676418 171186 676654
rect 171422 676418 171604 676654
rect 171004 676334 171604 676418
rect 171004 676098 171186 676334
rect 171422 676098 171604 676334
rect 171004 640654 171604 676098
rect 171004 640418 171186 640654
rect 171422 640418 171604 640654
rect 171004 640334 171604 640418
rect 171004 640098 171186 640334
rect 171422 640098 171604 640334
rect 171004 604654 171604 640098
rect 171004 604418 171186 604654
rect 171422 604418 171604 604654
rect 171004 604334 171604 604418
rect 171004 604098 171186 604334
rect 171422 604098 171604 604334
rect 171004 568654 171604 604098
rect 171004 568418 171186 568654
rect 171422 568418 171604 568654
rect 171004 568334 171604 568418
rect 171004 568098 171186 568334
rect 171422 568098 171604 568334
rect 171004 532654 171604 568098
rect 171004 532418 171186 532654
rect 171422 532418 171604 532654
rect 171004 532334 171604 532418
rect 171004 532098 171186 532334
rect 171422 532098 171604 532334
rect 171004 510000 171604 532098
rect 174604 680254 175204 710862
rect 192604 710478 193204 711440
rect 192604 710242 192786 710478
rect 193022 710242 193204 710478
rect 192604 710158 193204 710242
rect 192604 709922 192786 710158
rect 193022 709922 193204 710158
rect 189004 708598 189604 709560
rect 189004 708362 189186 708598
rect 189422 708362 189604 708598
rect 189004 708278 189604 708362
rect 189004 708042 189186 708278
rect 189422 708042 189604 708278
rect 185404 706718 186004 707680
rect 185404 706482 185586 706718
rect 185822 706482 186004 706718
rect 185404 706398 186004 706482
rect 185404 706162 185586 706398
rect 185822 706162 186004 706398
rect 174604 680018 174786 680254
rect 175022 680018 175204 680254
rect 174604 679934 175204 680018
rect 174604 679698 174786 679934
rect 175022 679698 175204 679934
rect 174604 644254 175204 679698
rect 174604 644018 174786 644254
rect 175022 644018 175204 644254
rect 174604 643934 175204 644018
rect 174604 643698 174786 643934
rect 175022 643698 175204 643934
rect 174604 608254 175204 643698
rect 174604 608018 174786 608254
rect 175022 608018 175204 608254
rect 174604 607934 175204 608018
rect 174604 607698 174786 607934
rect 175022 607698 175204 607934
rect 174604 572254 175204 607698
rect 174604 572018 174786 572254
rect 175022 572018 175204 572254
rect 174604 571934 175204 572018
rect 174604 571698 174786 571934
rect 175022 571698 175204 571934
rect 174604 536254 175204 571698
rect 174604 536018 174786 536254
rect 175022 536018 175204 536254
rect 174604 535934 175204 536018
rect 174604 535698 174786 535934
rect 175022 535698 175204 535934
rect 174604 510000 175204 535698
rect 181804 704838 182404 705800
rect 181804 704602 181986 704838
rect 182222 704602 182404 704838
rect 181804 704518 182404 704602
rect 181804 704282 181986 704518
rect 182222 704282 182404 704518
rect 181804 687454 182404 704282
rect 181804 687218 181986 687454
rect 182222 687218 182404 687454
rect 181804 687134 182404 687218
rect 181804 686898 181986 687134
rect 182222 686898 182404 687134
rect 181804 651454 182404 686898
rect 181804 651218 181986 651454
rect 182222 651218 182404 651454
rect 181804 651134 182404 651218
rect 181804 650898 181986 651134
rect 182222 650898 182404 651134
rect 181804 615454 182404 650898
rect 181804 615218 181986 615454
rect 182222 615218 182404 615454
rect 181804 615134 182404 615218
rect 181804 614898 181986 615134
rect 182222 614898 182404 615134
rect 181804 579454 182404 614898
rect 181804 579218 181986 579454
rect 182222 579218 182404 579454
rect 181804 579134 182404 579218
rect 181804 578898 181986 579134
rect 182222 578898 182404 579134
rect 181804 543454 182404 578898
rect 181804 543218 181986 543454
rect 182222 543218 182404 543454
rect 181804 543134 182404 543218
rect 181804 542898 181986 543134
rect 182222 542898 182404 543134
rect 181804 510000 182404 542898
rect 185404 691054 186004 706162
rect 185404 690818 185586 691054
rect 185822 690818 186004 691054
rect 185404 690734 186004 690818
rect 185404 690498 185586 690734
rect 185822 690498 186004 690734
rect 185404 655054 186004 690498
rect 185404 654818 185586 655054
rect 185822 654818 186004 655054
rect 185404 654734 186004 654818
rect 185404 654498 185586 654734
rect 185822 654498 186004 654734
rect 185404 619054 186004 654498
rect 185404 618818 185586 619054
rect 185822 618818 186004 619054
rect 185404 618734 186004 618818
rect 185404 618498 185586 618734
rect 185822 618498 186004 618734
rect 185404 583054 186004 618498
rect 185404 582818 185586 583054
rect 185822 582818 186004 583054
rect 185404 582734 186004 582818
rect 185404 582498 185586 582734
rect 185822 582498 186004 582734
rect 185404 547054 186004 582498
rect 185404 546818 185586 547054
rect 185822 546818 186004 547054
rect 185404 546734 186004 546818
rect 185404 546498 185586 546734
rect 185822 546498 186004 546734
rect 185404 511054 186004 546498
rect 185404 510818 185586 511054
rect 185822 510818 186004 511054
rect 185404 510734 186004 510818
rect 185404 510498 185586 510734
rect 185822 510498 186004 510734
rect 185404 510000 186004 510498
rect 189004 694654 189604 708042
rect 189004 694418 189186 694654
rect 189422 694418 189604 694654
rect 189004 694334 189604 694418
rect 189004 694098 189186 694334
rect 189422 694098 189604 694334
rect 189004 658654 189604 694098
rect 189004 658418 189186 658654
rect 189422 658418 189604 658654
rect 189004 658334 189604 658418
rect 189004 658098 189186 658334
rect 189422 658098 189604 658334
rect 189004 622654 189604 658098
rect 189004 622418 189186 622654
rect 189422 622418 189604 622654
rect 189004 622334 189604 622418
rect 189004 622098 189186 622334
rect 189422 622098 189604 622334
rect 189004 586654 189604 622098
rect 189004 586418 189186 586654
rect 189422 586418 189604 586654
rect 189004 586334 189604 586418
rect 189004 586098 189186 586334
rect 189422 586098 189604 586334
rect 189004 550654 189604 586098
rect 189004 550418 189186 550654
rect 189422 550418 189604 550654
rect 189004 550334 189604 550418
rect 189004 550098 189186 550334
rect 189422 550098 189604 550334
rect 189004 514654 189604 550098
rect 189004 514418 189186 514654
rect 189422 514418 189604 514654
rect 189004 514334 189604 514418
rect 189004 514098 189186 514334
rect 189422 514098 189604 514334
rect 189004 510000 189604 514098
rect 192604 698254 193204 709922
rect 210604 711418 211204 711440
rect 210604 711182 210786 711418
rect 211022 711182 211204 711418
rect 210604 711098 211204 711182
rect 210604 710862 210786 711098
rect 211022 710862 211204 711098
rect 207004 709538 207604 709560
rect 207004 709302 207186 709538
rect 207422 709302 207604 709538
rect 207004 709218 207604 709302
rect 207004 708982 207186 709218
rect 207422 708982 207604 709218
rect 203404 707658 204004 707680
rect 203404 707422 203586 707658
rect 203822 707422 204004 707658
rect 203404 707338 204004 707422
rect 203404 707102 203586 707338
rect 203822 707102 204004 707338
rect 192604 698018 192786 698254
rect 193022 698018 193204 698254
rect 192604 697934 193204 698018
rect 192604 697698 192786 697934
rect 193022 697698 193204 697934
rect 192604 662254 193204 697698
rect 192604 662018 192786 662254
rect 193022 662018 193204 662254
rect 192604 661934 193204 662018
rect 192604 661698 192786 661934
rect 193022 661698 193204 661934
rect 192604 626254 193204 661698
rect 192604 626018 192786 626254
rect 193022 626018 193204 626254
rect 192604 625934 193204 626018
rect 192604 625698 192786 625934
rect 193022 625698 193204 625934
rect 192604 590254 193204 625698
rect 192604 590018 192786 590254
rect 193022 590018 193204 590254
rect 192604 589934 193204 590018
rect 192604 589698 192786 589934
rect 193022 589698 193204 589934
rect 192604 554254 193204 589698
rect 192604 554018 192786 554254
rect 193022 554018 193204 554254
rect 192604 553934 193204 554018
rect 192604 553698 192786 553934
rect 193022 553698 193204 553934
rect 192604 518254 193204 553698
rect 192604 518018 192786 518254
rect 193022 518018 193204 518254
rect 192604 517934 193204 518018
rect 192604 517698 192786 517934
rect 193022 517698 193204 517934
rect 192604 510000 193204 517698
rect 199804 705778 200404 705800
rect 199804 705542 199986 705778
rect 200222 705542 200404 705778
rect 199804 705458 200404 705542
rect 199804 705222 199986 705458
rect 200222 705222 200404 705458
rect 199804 669454 200404 705222
rect 199804 669218 199986 669454
rect 200222 669218 200404 669454
rect 199804 669134 200404 669218
rect 199804 668898 199986 669134
rect 200222 668898 200404 669134
rect 199804 633454 200404 668898
rect 199804 633218 199986 633454
rect 200222 633218 200404 633454
rect 199804 633134 200404 633218
rect 199804 632898 199986 633134
rect 200222 632898 200404 633134
rect 199804 597454 200404 632898
rect 199804 597218 199986 597454
rect 200222 597218 200404 597454
rect 199804 597134 200404 597218
rect 199804 596898 199986 597134
rect 200222 596898 200404 597134
rect 199804 561454 200404 596898
rect 199804 561218 199986 561454
rect 200222 561218 200404 561454
rect 199804 561134 200404 561218
rect 199804 560898 199986 561134
rect 200222 560898 200404 561134
rect 199804 525454 200404 560898
rect 199804 525218 199986 525454
rect 200222 525218 200404 525454
rect 199804 525134 200404 525218
rect 199804 524898 199986 525134
rect 200222 524898 200404 525134
rect 199804 510000 200404 524898
rect 203404 673054 204004 707102
rect 203404 672818 203586 673054
rect 203822 672818 204004 673054
rect 203404 672734 204004 672818
rect 203404 672498 203586 672734
rect 203822 672498 204004 672734
rect 203404 637054 204004 672498
rect 203404 636818 203586 637054
rect 203822 636818 204004 637054
rect 203404 636734 204004 636818
rect 203404 636498 203586 636734
rect 203822 636498 204004 636734
rect 203404 601054 204004 636498
rect 203404 600818 203586 601054
rect 203822 600818 204004 601054
rect 203404 600734 204004 600818
rect 203404 600498 203586 600734
rect 203822 600498 204004 600734
rect 203404 565054 204004 600498
rect 203404 564818 203586 565054
rect 203822 564818 204004 565054
rect 203404 564734 204004 564818
rect 203404 564498 203586 564734
rect 203822 564498 204004 564734
rect 203404 529054 204004 564498
rect 203404 528818 203586 529054
rect 203822 528818 204004 529054
rect 203404 528734 204004 528818
rect 203404 528498 203586 528734
rect 203822 528498 204004 528734
rect 203404 510000 204004 528498
rect 207004 676654 207604 708982
rect 207004 676418 207186 676654
rect 207422 676418 207604 676654
rect 207004 676334 207604 676418
rect 207004 676098 207186 676334
rect 207422 676098 207604 676334
rect 207004 640654 207604 676098
rect 207004 640418 207186 640654
rect 207422 640418 207604 640654
rect 207004 640334 207604 640418
rect 207004 640098 207186 640334
rect 207422 640098 207604 640334
rect 207004 604654 207604 640098
rect 207004 604418 207186 604654
rect 207422 604418 207604 604654
rect 207004 604334 207604 604418
rect 207004 604098 207186 604334
rect 207422 604098 207604 604334
rect 207004 568654 207604 604098
rect 207004 568418 207186 568654
rect 207422 568418 207604 568654
rect 207004 568334 207604 568418
rect 207004 568098 207186 568334
rect 207422 568098 207604 568334
rect 207004 532654 207604 568098
rect 207004 532418 207186 532654
rect 207422 532418 207604 532654
rect 207004 532334 207604 532418
rect 207004 532098 207186 532334
rect 207422 532098 207604 532334
rect 207004 510000 207604 532098
rect 210604 680254 211204 710862
rect 228604 710478 229204 711440
rect 228604 710242 228786 710478
rect 229022 710242 229204 710478
rect 228604 710158 229204 710242
rect 228604 709922 228786 710158
rect 229022 709922 229204 710158
rect 225004 708598 225604 709560
rect 225004 708362 225186 708598
rect 225422 708362 225604 708598
rect 225004 708278 225604 708362
rect 225004 708042 225186 708278
rect 225422 708042 225604 708278
rect 221404 706718 222004 707680
rect 221404 706482 221586 706718
rect 221822 706482 222004 706718
rect 221404 706398 222004 706482
rect 221404 706162 221586 706398
rect 221822 706162 222004 706398
rect 210604 680018 210786 680254
rect 211022 680018 211204 680254
rect 210604 679934 211204 680018
rect 210604 679698 210786 679934
rect 211022 679698 211204 679934
rect 210604 644254 211204 679698
rect 210604 644018 210786 644254
rect 211022 644018 211204 644254
rect 210604 643934 211204 644018
rect 210604 643698 210786 643934
rect 211022 643698 211204 643934
rect 210604 608254 211204 643698
rect 210604 608018 210786 608254
rect 211022 608018 211204 608254
rect 210604 607934 211204 608018
rect 210604 607698 210786 607934
rect 211022 607698 211204 607934
rect 210604 572254 211204 607698
rect 210604 572018 210786 572254
rect 211022 572018 211204 572254
rect 210604 571934 211204 572018
rect 210604 571698 210786 571934
rect 211022 571698 211204 571934
rect 210604 536254 211204 571698
rect 210604 536018 210786 536254
rect 211022 536018 211204 536254
rect 210604 535934 211204 536018
rect 210604 535698 210786 535934
rect 211022 535698 211204 535934
rect 210604 510000 211204 535698
rect 217804 704838 218404 705800
rect 217804 704602 217986 704838
rect 218222 704602 218404 704838
rect 217804 704518 218404 704602
rect 217804 704282 217986 704518
rect 218222 704282 218404 704518
rect 217804 687454 218404 704282
rect 217804 687218 217986 687454
rect 218222 687218 218404 687454
rect 217804 687134 218404 687218
rect 217804 686898 217986 687134
rect 218222 686898 218404 687134
rect 217804 651454 218404 686898
rect 217804 651218 217986 651454
rect 218222 651218 218404 651454
rect 217804 651134 218404 651218
rect 217804 650898 217986 651134
rect 218222 650898 218404 651134
rect 217804 615454 218404 650898
rect 217804 615218 217986 615454
rect 218222 615218 218404 615454
rect 217804 615134 218404 615218
rect 217804 614898 217986 615134
rect 218222 614898 218404 615134
rect 217804 579454 218404 614898
rect 217804 579218 217986 579454
rect 218222 579218 218404 579454
rect 217804 579134 218404 579218
rect 217804 578898 217986 579134
rect 218222 578898 218404 579134
rect 217804 543454 218404 578898
rect 217804 543218 217986 543454
rect 218222 543218 218404 543454
rect 217804 543134 218404 543218
rect 217804 542898 217986 543134
rect 218222 542898 218404 543134
rect 217804 510000 218404 542898
rect 221404 691054 222004 706162
rect 221404 690818 221586 691054
rect 221822 690818 222004 691054
rect 221404 690734 222004 690818
rect 221404 690498 221586 690734
rect 221822 690498 222004 690734
rect 221404 655054 222004 690498
rect 221404 654818 221586 655054
rect 221822 654818 222004 655054
rect 221404 654734 222004 654818
rect 221404 654498 221586 654734
rect 221822 654498 222004 654734
rect 221404 619054 222004 654498
rect 221404 618818 221586 619054
rect 221822 618818 222004 619054
rect 221404 618734 222004 618818
rect 221404 618498 221586 618734
rect 221822 618498 222004 618734
rect 221404 583054 222004 618498
rect 221404 582818 221586 583054
rect 221822 582818 222004 583054
rect 221404 582734 222004 582818
rect 221404 582498 221586 582734
rect 221822 582498 222004 582734
rect 221404 547054 222004 582498
rect 221404 546818 221586 547054
rect 221822 546818 222004 547054
rect 221404 546734 222004 546818
rect 221404 546498 221586 546734
rect 221822 546498 222004 546734
rect 221404 511054 222004 546498
rect 221404 510818 221586 511054
rect 221822 510818 222004 511054
rect 221404 510734 222004 510818
rect 221404 510498 221586 510734
rect 221822 510498 222004 510734
rect 221404 510000 222004 510498
rect 225004 694654 225604 708042
rect 225004 694418 225186 694654
rect 225422 694418 225604 694654
rect 225004 694334 225604 694418
rect 225004 694098 225186 694334
rect 225422 694098 225604 694334
rect 225004 658654 225604 694098
rect 225004 658418 225186 658654
rect 225422 658418 225604 658654
rect 225004 658334 225604 658418
rect 225004 658098 225186 658334
rect 225422 658098 225604 658334
rect 225004 622654 225604 658098
rect 225004 622418 225186 622654
rect 225422 622418 225604 622654
rect 225004 622334 225604 622418
rect 225004 622098 225186 622334
rect 225422 622098 225604 622334
rect 225004 586654 225604 622098
rect 225004 586418 225186 586654
rect 225422 586418 225604 586654
rect 225004 586334 225604 586418
rect 225004 586098 225186 586334
rect 225422 586098 225604 586334
rect 225004 550654 225604 586098
rect 225004 550418 225186 550654
rect 225422 550418 225604 550654
rect 225004 550334 225604 550418
rect 225004 550098 225186 550334
rect 225422 550098 225604 550334
rect 225004 514654 225604 550098
rect 225004 514418 225186 514654
rect 225422 514418 225604 514654
rect 225004 514334 225604 514418
rect 225004 514098 225186 514334
rect 225422 514098 225604 514334
rect 225004 510000 225604 514098
rect 228604 698254 229204 709922
rect 246604 711418 247204 711440
rect 246604 711182 246786 711418
rect 247022 711182 247204 711418
rect 246604 711098 247204 711182
rect 246604 710862 246786 711098
rect 247022 710862 247204 711098
rect 243004 709538 243604 709560
rect 243004 709302 243186 709538
rect 243422 709302 243604 709538
rect 243004 709218 243604 709302
rect 243004 708982 243186 709218
rect 243422 708982 243604 709218
rect 239404 707658 240004 707680
rect 239404 707422 239586 707658
rect 239822 707422 240004 707658
rect 239404 707338 240004 707422
rect 239404 707102 239586 707338
rect 239822 707102 240004 707338
rect 228604 698018 228786 698254
rect 229022 698018 229204 698254
rect 228604 697934 229204 698018
rect 228604 697698 228786 697934
rect 229022 697698 229204 697934
rect 228604 662254 229204 697698
rect 228604 662018 228786 662254
rect 229022 662018 229204 662254
rect 228604 661934 229204 662018
rect 228604 661698 228786 661934
rect 229022 661698 229204 661934
rect 228604 626254 229204 661698
rect 228604 626018 228786 626254
rect 229022 626018 229204 626254
rect 228604 625934 229204 626018
rect 228604 625698 228786 625934
rect 229022 625698 229204 625934
rect 228604 590254 229204 625698
rect 228604 590018 228786 590254
rect 229022 590018 229204 590254
rect 228604 589934 229204 590018
rect 228604 589698 228786 589934
rect 229022 589698 229204 589934
rect 228604 554254 229204 589698
rect 228604 554018 228786 554254
rect 229022 554018 229204 554254
rect 228604 553934 229204 554018
rect 228604 553698 228786 553934
rect 229022 553698 229204 553934
rect 228604 518254 229204 553698
rect 228604 518018 228786 518254
rect 229022 518018 229204 518254
rect 228604 517934 229204 518018
rect 228604 517698 228786 517934
rect 229022 517698 229204 517934
rect 228604 510000 229204 517698
rect 235804 705778 236404 705800
rect 235804 705542 235986 705778
rect 236222 705542 236404 705778
rect 235804 705458 236404 705542
rect 235804 705222 235986 705458
rect 236222 705222 236404 705458
rect 235804 669454 236404 705222
rect 235804 669218 235986 669454
rect 236222 669218 236404 669454
rect 235804 669134 236404 669218
rect 235804 668898 235986 669134
rect 236222 668898 236404 669134
rect 235804 633454 236404 668898
rect 235804 633218 235986 633454
rect 236222 633218 236404 633454
rect 235804 633134 236404 633218
rect 235804 632898 235986 633134
rect 236222 632898 236404 633134
rect 235804 597454 236404 632898
rect 235804 597218 235986 597454
rect 236222 597218 236404 597454
rect 235804 597134 236404 597218
rect 235804 596898 235986 597134
rect 236222 596898 236404 597134
rect 235804 561454 236404 596898
rect 235804 561218 235986 561454
rect 236222 561218 236404 561454
rect 235804 561134 236404 561218
rect 235804 560898 235986 561134
rect 236222 560898 236404 561134
rect 235804 525454 236404 560898
rect 235804 525218 235986 525454
rect 236222 525218 236404 525454
rect 235804 525134 236404 525218
rect 235804 524898 235986 525134
rect 236222 524898 236404 525134
rect 235804 510000 236404 524898
rect 239404 673054 240004 707102
rect 239404 672818 239586 673054
rect 239822 672818 240004 673054
rect 239404 672734 240004 672818
rect 239404 672498 239586 672734
rect 239822 672498 240004 672734
rect 239404 637054 240004 672498
rect 239404 636818 239586 637054
rect 239822 636818 240004 637054
rect 239404 636734 240004 636818
rect 239404 636498 239586 636734
rect 239822 636498 240004 636734
rect 239404 601054 240004 636498
rect 239404 600818 239586 601054
rect 239822 600818 240004 601054
rect 239404 600734 240004 600818
rect 239404 600498 239586 600734
rect 239822 600498 240004 600734
rect 239404 565054 240004 600498
rect 239404 564818 239586 565054
rect 239822 564818 240004 565054
rect 239404 564734 240004 564818
rect 239404 564498 239586 564734
rect 239822 564498 240004 564734
rect 239404 529054 240004 564498
rect 239404 528818 239586 529054
rect 239822 528818 240004 529054
rect 239404 528734 240004 528818
rect 239404 528498 239586 528734
rect 239822 528498 240004 528734
rect 239404 510000 240004 528498
rect 243004 676654 243604 708982
rect 243004 676418 243186 676654
rect 243422 676418 243604 676654
rect 243004 676334 243604 676418
rect 243004 676098 243186 676334
rect 243422 676098 243604 676334
rect 243004 640654 243604 676098
rect 243004 640418 243186 640654
rect 243422 640418 243604 640654
rect 243004 640334 243604 640418
rect 243004 640098 243186 640334
rect 243422 640098 243604 640334
rect 243004 604654 243604 640098
rect 243004 604418 243186 604654
rect 243422 604418 243604 604654
rect 243004 604334 243604 604418
rect 243004 604098 243186 604334
rect 243422 604098 243604 604334
rect 243004 568654 243604 604098
rect 243004 568418 243186 568654
rect 243422 568418 243604 568654
rect 243004 568334 243604 568418
rect 243004 568098 243186 568334
rect 243422 568098 243604 568334
rect 243004 532654 243604 568098
rect 243004 532418 243186 532654
rect 243422 532418 243604 532654
rect 243004 532334 243604 532418
rect 243004 532098 243186 532334
rect 243422 532098 243604 532334
rect 243004 510000 243604 532098
rect 246604 680254 247204 710862
rect 264604 710478 265204 711440
rect 264604 710242 264786 710478
rect 265022 710242 265204 710478
rect 264604 710158 265204 710242
rect 264604 709922 264786 710158
rect 265022 709922 265204 710158
rect 261004 708598 261604 709560
rect 261004 708362 261186 708598
rect 261422 708362 261604 708598
rect 261004 708278 261604 708362
rect 261004 708042 261186 708278
rect 261422 708042 261604 708278
rect 257404 706718 258004 707680
rect 257404 706482 257586 706718
rect 257822 706482 258004 706718
rect 257404 706398 258004 706482
rect 257404 706162 257586 706398
rect 257822 706162 258004 706398
rect 246604 680018 246786 680254
rect 247022 680018 247204 680254
rect 246604 679934 247204 680018
rect 246604 679698 246786 679934
rect 247022 679698 247204 679934
rect 246604 644254 247204 679698
rect 246604 644018 246786 644254
rect 247022 644018 247204 644254
rect 246604 643934 247204 644018
rect 246604 643698 246786 643934
rect 247022 643698 247204 643934
rect 246604 608254 247204 643698
rect 246604 608018 246786 608254
rect 247022 608018 247204 608254
rect 246604 607934 247204 608018
rect 246604 607698 246786 607934
rect 247022 607698 247204 607934
rect 246604 572254 247204 607698
rect 246604 572018 246786 572254
rect 247022 572018 247204 572254
rect 246604 571934 247204 572018
rect 246604 571698 246786 571934
rect 247022 571698 247204 571934
rect 246604 536254 247204 571698
rect 246604 536018 246786 536254
rect 247022 536018 247204 536254
rect 246604 535934 247204 536018
rect 246604 535698 246786 535934
rect 247022 535698 247204 535934
rect 246604 510000 247204 535698
rect 253804 704838 254404 705800
rect 253804 704602 253986 704838
rect 254222 704602 254404 704838
rect 253804 704518 254404 704602
rect 253804 704282 253986 704518
rect 254222 704282 254404 704518
rect 253804 687454 254404 704282
rect 253804 687218 253986 687454
rect 254222 687218 254404 687454
rect 253804 687134 254404 687218
rect 253804 686898 253986 687134
rect 254222 686898 254404 687134
rect 253804 651454 254404 686898
rect 253804 651218 253986 651454
rect 254222 651218 254404 651454
rect 253804 651134 254404 651218
rect 253804 650898 253986 651134
rect 254222 650898 254404 651134
rect 253804 615454 254404 650898
rect 253804 615218 253986 615454
rect 254222 615218 254404 615454
rect 253804 615134 254404 615218
rect 253804 614898 253986 615134
rect 254222 614898 254404 615134
rect 253804 579454 254404 614898
rect 253804 579218 253986 579454
rect 254222 579218 254404 579454
rect 253804 579134 254404 579218
rect 253804 578898 253986 579134
rect 254222 578898 254404 579134
rect 253804 543454 254404 578898
rect 253804 543218 253986 543454
rect 254222 543218 254404 543454
rect 253804 543134 254404 543218
rect 253804 542898 253986 543134
rect 254222 542898 254404 543134
rect 253804 510000 254404 542898
rect 257404 691054 258004 706162
rect 257404 690818 257586 691054
rect 257822 690818 258004 691054
rect 257404 690734 258004 690818
rect 257404 690498 257586 690734
rect 257822 690498 258004 690734
rect 257404 655054 258004 690498
rect 257404 654818 257586 655054
rect 257822 654818 258004 655054
rect 257404 654734 258004 654818
rect 257404 654498 257586 654734
rect 257822 654498 258004 654734
rect 257404 619054 258004 654498
rect 257404 618818 257586 619054
rect 257822 618818 258004 619054
rect 257404 618734 258004 618818
rect 257404 618498 257586 618734
rect 257822 618498 258004 618734
rect 257404 583054 258004 618498
rect 257404 582818 257586 583054
rect 257822 582818 258004 583054
rect 257404 582734 258004 582818
rect 257404 582498 257586 582734
rect 257822 582498 258004 582734
rect 257404 547054 258004 582498
rect 257404 546818 257586 547054
rect 257822 546818 258004 547054
rect 257404 546734 258004 546818
rect 257404 546498 257586 546734
rect 257822 546498 258004 546734
rect 257404 511054 258004 546498
rect 257404 510818 257586 511054
rect 257822 510818 258004 511054
rect 257404 510734 258004 510818
rect 257404 510498 257586 510734
rect 257822 510498 258004 510734
rect 257404 510000 258004 510498
rect 261004 694654 261604 708042
rect 261004 694418 261186 694654
rect 261422 694418 261604 694654
rect 261004 694334 261604 694418
rect 261004 694098 261186 694334
rect 261422 694098 261604 694334
rect 261004 658654 261604 694098
rect 261004 658418 261186 658654
rect 261422 658418 261604 658654
rect 261004 658334 261604 658418
rect 261004 658098 261186 658334
rect 261422 658098 261604 658334
rect 261004 622654 261604 658098
rect 261004 622418 261186 622654
rect 261422 622418 261604 622654
rect 261004 622334 261604 622418
rect 261004 622098 261186 622334
rect 261422 622098 261604 622334
rect 261004 586654 261604 622098
rect 261004 586418 261186 586654
rect 261422 586418 261604 586654
rect 261004 586334 261604 586418
rect 261004 586098 261186 586334
rect 261422 586098 261604 586334
rect 261004 550654 261604 586098
rect 261004 550418 261186 550654
rect 261422 550418 261604 550654
rect 261004 550334 261604 550418
rect 261004 550098 261186 550334
rect 261422 550098 261604 550334
rect 261004 514654 261604 550098
rect 261004 514418 261186 514654
rect 261422 514418 261604 514654
rect 261004 514334 261604 514418
rect 261004 514098 261186 514334
rect 261422 514098 261604 514334
rect 261004 510000 261604 514098
rect 264604 698254 265204 709922
rect 282604 711418 283204 711440
rect 282604 711182 282786 711418
rect 283022 711182 283204 711418
rect 282604 711098 283204 711182
rect 282604 710862 282786 711098
rect 283022 710862 283204 711098
rect 279004 709538 279604 709560
rect 279004 709302 279186 709538
rect 279422 709302 279604 709538
rect 279004 709218 279604 709302
rect 279004 708982 279186 709218
rect 279422 708982 279604 709218
rect 275404 707658 276004 707680
rect 275404 707422 275586 707658
rect 275822 707422 276004 707658
rect 275404 707338 276004 707422
rect 275404 707102 275586 707338
rect 275822 707102 276004 707338
rect 264604 698018 264786 698254
rect 265022 698018 265204 698254
rect 264604 697934 265204 698018
rect 264604 697698 264786 697934
rect 265022 697698 265204 697934
rect 264604 662254 265204 697698
rect 264604 662018 264786 662254
rect 265022 662018 265204 662254
rect 264604 661934 265204 662018
rect 264604 661698 264786 661934
rect 265022 661698 265204 661934
rect 264604 626254 265204 661698
rect 264604 626018 264786 626254
rect 265022 626018 265204 626254
rect 264604 625934 265204 626018
rect 264604 625698 264786 625934
rect 265022 625698 265204 625934
rect 264604 590254 265204 625698
rect 264604 590018 264786 590254
rect 265022 590018 265204 590254
rect 264604 589934 265204 590018
rect 264604 589698 264786 589934
rect 265022 589698 265204 589934
rect 264604 554254 265204 589698
rect 264604 554018 264786 554254
rect 265022 554018 265204 554254
rect 264604 553934 265204 554018
rect 264604 553698 264786 553934
rect 265022 553698 265204 553934
rect 264604 518254 265204 553698
rect 264604 518018 264786 518254
rect 265022 518018 265204 518254
rect 264604 517934 265204 518018
rect 264604 517698 264786 517934
rect 265022 517698 265204 517934
rect 264604 510000 265204 517698
rect 271804 705778 272404 705800
rect 271804 705542 271986 705778
rect 272222 705542 272404 705778
rect 271804 705458 272404 705542
rect 271804 705222 271986 705458
rect 272222 705222 272404 705458
rect 271804 669454 272404 705222
rect 271804 669218 271986 669454
rect 272222 669218 272404 669454
rect 271804 669134 272404 669218
rect 271804 668898 271986 669134
rect 272222 668898 272404 669134
rect 271804 633454 272404 668898
rect 271804 633218 271986 633454
rect 272222 633218 272404 633454
rect 271804 633134 272404 633218
rect 271804 632898 271986 633134
rect 272222 632898 272404 633134
rect 271804 597454 272404 632898
rect 271804 597218 271986 597454
rect 272222 597218 272404 597454
rect 271804 597134 272404 597218
rect 271804 596898 271986 597134
rect 272222 596898 272404 597134
rect 271804 561454 272404 596898
rect 271804 561218 271986 561454
rect 272222 561218 272404 561454
rect 271804 561134 272404 561218
rect 271804 560898 271986 561134
rect 272222 560898 272404 561134
rect 271804 525454 272404 560898
rect 271804 525218 271986 525454
rect 272222 525218 272404 525454
rect 271804 525134 272404 525218
rect 271804 524898 271986 525134
rect 272222 524898 272404 525134
rect 271804 510000 272404 524898
rect 275404 673054 276004 707102
rect 275404 672818 275586 673054
rect 275822 672818 276004 673054
rect 275404 672734 276004 672818
rect 275404 672498 275586 672734
rect 275822 672498 276004 672734
rect 275404 637054 276004 672498
rect 275404 636818 275586 637054
rect 275822 636818 276004 637054
rect 275404 636734 276004 636818
rect 275404 636498 275586 636734
rect 275822 636498 276004 636734
rect 275404 601054 276004 636498
rect 275404 600818 275586 601054
rect 275822 600818 276004 601054
rect 275404 600734 276004 600818
rect 275404 600498 275586 600734
rect 275822 600498 276004 600734
rect 275404 565054 276004 600498
rect 275404 564818 275586 565054
rect 275822 564818 276004 565054
rect 275404 564734 276004 564818
rect 275404 564498 275586 564734
rect 275822 564498 276004 564734
rect 275404 529054 276004 564498
rect 275404 528818 275586 529054
rect 275822 528818 276004 529054
rect 275404 528734 276004 528818
rect 275404 528498 275586 528734
rect 275822 528498 276004 528734
rect 275404 510000 276004 528498
rect 279004 676654 279604 708982
rect 279004 676418 279186 676654
rect 279422 676418 279604 676654
rect 279004 676334 279604 676418
rect 279004 676098 279186 676334
rect 279422 676098 279604 676334
rect 279004 640654 279604 676098
rect 279004 640418 279186 640654
rect 279422 640418 279604 640654
rect 279004 640334 279604 640418
rect 279004 640098 279186 640334
rect 279422 640098 279604 640334
rect 279004 604654 279604 640098
rect 279004 604418 279186 604654
rect 279422 604418 279604 604654
rect 279004 604334 279604 604418
rect 279004 604098 279186 604334
rect 279422 604098 279604 604334
rect 279004 568654 279604 604098
rect 279004 568418 279186 568654
rect 279422 568418 279604 568654
rect 279004 568334 279604 568418
rect 279004 568098 279186 568334
rect 279422 568098 279604 568334
rect 279004 532654 279604 568098
rect 279004 532418 279186 532654
rect 279422 532418 279604 532654
rect 279004 532334 279604 532418
rect 279004 532098 279186 532334
rect 279422 532098 279604 532334
rect 279004 510000 279604 532098
rect 282604 680254 283204 710862
rect 300604 710478 301204 711440
rect 300604 710242 300786 710478
rect 301022 710242 301204 710478
rect 300604 710158 301204 710242
rect 300604 709922 300786 710158
rect 301022 709922 301204 710158
rect 297004 708598 297604 709560
rect 297004 708362 297186 708598
rect 297422 708362 297604 708598
rect 297004 708278 297604 708362
rect 297004 708042 297186 708278
rect 297422 708042 297604 708278
rect 293404 706718 294004 707680
rect 293404 706482 293586 706718
rect 293822 706482 294004 706718
rect 293404 706398 294004 706482
rect 293404 706162 293586 706398
rect 293822 706162 294004 706398
rect 282604 680018 282786 680254
rect 283022 680018 283204 680254
rect 282604 679934 283204 680018
rect 282604 679698 282786 679934
rect 283022 679698 283204 679934
rect 282604 644254 283204 679698
rect 282604 644018 282786 644254
rect 283022 644018 283204 644254
rect 282604 643934 283204 644018
rect 282604 643698 282786 643934
rect 283022 643698 283204 643934
rect 282604 608254 283204 643698
rect 282604 608018 282786 608254
rect 283022 608018 283204 608254
rect 282604 607934 283204 608018
rect 282604 607698 282786 607934
rect 283022 607698 283204 607934
rect 282604 572254 283204 607698
rect 282604 572018 282786 572254
rect 283022 572018 283204 572254
rect 282604 571934 283204 572018
rect 282604 571698 282786 571934
rect 283022 571698 283204 571934
rect 282604 536254 283204 571698
rect 282604 536018 282786 536254
rect 283022 536018 283204 536254
rect 282604 535934 283204 536018
rect 282604 535698 282786 535934
rect 283022 535698 283204 535934
rect 282604 510000 283204 535698
rect 289804 704838 290404 705800
rect 289804 704602 289986 704838
rect 290222 704602 290404 704838
rect 289804 704518 290404 704602
rect 289804 704282 289986 704518
rect 290222 704282 290404 704518
rect 289804 687454 290404 704282
rect 289804 687218 289986 687454
rect 290222 687218 290404 687454
rect 289804 687134 290404 687218
rect 289804 686898 289986 687134
rect 290222 686898 290404 687134
rect 289804 651454 290404 686898
rect 289804 651218 289986 651454
rect 290222 651218 290404 651454
rect 289804 651134 290404 651218
rect 289804 650898 289986 651134
rect 290222 650898 290404 651134
rect 289804 615454 290404 650898
rect 289804 615218 289986 615454
rect 290222 615218 290404 615454
rect 289804 615134 290404 615218
rect 289804 614898 289986 615134
rect 290222 614898 290404 615134
rect 289804 579454 290404 614898
rect 289804 579218 289986 579454
rect 290222 579218 290404 579454
rect 289804 579134 290404 579218
rect 289804 578898 289986 579134
rect 290222 578898 290404 579134
rect 289804 543454 290404 578898
rect 289804 543218 289986 543454
rect 290222 543218 290404 543454
rect 289804 543134 290404 543218
rect 289804 542898 289986 543134
rect 290222 542898 290404 543134
rect 289804 510000 290404 542898
rect 293404 691054 294004 706162
rect 293404 690818 293586 691054
rect 293822 690818 294004 691054
rect 293404 690734 294004 690818
rect 293404 690498 293586 690734
rect 293822 690498 294004 690734
rect 293404 655054 294004 690498
rect 293404 654818 293586 655054
rect 293822 654818 294004 655054
rect 293404 654734 294004 654818
rect 293404 654498 293586 654734
rect 293822 654498 294004 654734
rect 293404 619054 294004 654498
rect 293404 618818 293586 619054
rect 293822 618818 294004 619054
rect 293404 618734 294004 618818
rect 293404 618498 293586 618734
rect 293822 618498 294004 618734
rect 293404 583054 294004 618498
rect 293404 582818 293586 583054
rect 293822 582818 294004 583054
rect 293404 582734 294004 582818
rect 293404 582498 293586 582734
rect 293822 582498 294004 582734
rect 293404 547054 294004 582498
rect 293404 546818 293586 547054
rect 293822 546818 294004 547054
rect 293404 546734 294004 546818
rect 293404 546498 293586 546734
rect 293822 546498 294004 546734
rect 293404 511054 294004 546498
rect 293404 510818 293586 511054
rect 293822 510818 294004 511054
rect 293404 510734 294004 510818
rect 293404 510498 293586 510734
rect 293822 510498 294004 510734
rect 293404 510000 294004 510498
rect 297004 694654 297604 708042
rect 297004 694418 297186 694654
rect 297422 694418 297604 694654
rect 297004 694334 297604 694418
rect 297004 694098 297186 694334
rect 297422 694098 297604 694334
rect 297004 658654 297604 694098
rect 297004 658418 297186 658654
rect 297422 658418 297604 658654
rect 297004 658334 297604 658418
rect 297004 658098 297186 658334
rect 297422 658098 297604 658334
rect 297004 622654 297604 658098
rect 297004 622418 297186 622654
rect 297422 622418 297604 622654
rect 297004 622334 297604 622418
rect 297004 622098 297186 622334
rect 297422 622098 297604 622334
rect 297004 586654 297604 622098
rect 297004 586418 297186 586654
rect 297422 586418 297604 586654
rect 297004 586334 297604 586418
rect 297004 586098 297186 586334
rect 297422 586098 297604 586334
rect 297004 550654 297604 586098
rect 297004 550418 297186 550654
rect 297422 550418 297604 550654
rect 297004 550334 297604 550418
rect 297004 550098 297186 550334
rect 297422 550098 297604 550334
rect 297004 514654 297604 550098
rect 297004 514418 297186 514654
rect 297422 514418 297604 514654
rect 297004 514334 297604 514418
rect 297004 514098 297186 514334
rect 297422 514098 297604 514334
rect 297004 510000 297604 514098
rect 300604 698254 301204 709922
rect 318604 711418 319204 711440
rect 318604 711182 318786 711418
rect 319022 711182 319204 711418
rect 318604 711098 319204 711182
rect 318604 710862 318786 711098
rect 319022 710862 319204 711098
rect 315004 709538 315604 709560
rect 315004 709302 315186 709538
rect 315422 709302 315604 709538
rect 315004 709218 315604 709302
rect 315004 708982 315186 709218
rect 315422 708982 315604 709218
rect 311404 707658 312004 707680
rect 311404 707422 311586 707658
rect 311822 707422 312004 707658
rect 311404 707338 312004 707422
rect 311404 707102 311586 707338
rect 311822 707102 312004 707338
rect 300604 698018 300786 698254
rect 301022 698018 301204 698254
rect 300604 697934 301204 698018
rect 300604 697698 300786 697934
rect 301022 697698 301204 697934
rect 300604 662254 301204 697698
rect 300604 662018 300786 662254
rect 301022 662018 301204 662254
rect 300604 661934 301204 662018
rect 300604 661698 300786 661934
rect 301022 661698 301204 661934
rect 300604 626254 301204 661698
rect 300604 626018 300786 626254
rect 301022 626018 301204 626254
rect 300604 625934 301204 626018
rect 300604 625698 300786 625934
rect 301022 625698 301204 625934
rect 300604 590254 301204 625698
rect 300604 590018 300786 590254
rect 301022 590018 301204 590254
rect 300604 589934 301204 590018
rect 300604 589698 300786 589934
rect 301022 589698 301204 589934
rect 300604 554254 301204 589698
rect 300604 554018 300786 554254
rect 301022 554018 301204 554254
rect 300604 553934 301204 554018
rect 300604 553698 300786 553934
rect 301022 553698 301204 553934
rect 300604 518254 301204 553698
rect 300604 518018 300786 518254
rect 301022 518018 301204 518254
rect 300604 517934 301204 518018
rect 300604 517698 300786 517934
rect 301022 517698 301204 517934
rect 300604 510000 301204 517698
rect 307804 705778 308404 705800
rect 307804 705542 307986 705778
rect 308222 705542 308404 705778
rect 307804 705458 308404 705542
rect 307804 705222 307986 705458
rect 308222 705222 308404 705458
rect 307804 669454 308404 705222
rect 307804 669218 307986 669454
rect 308222 669218 308404 669454
rect 307804 669134 308404 669218
rect 307804 668898 307986 669134
rect 308222 668898 308404 669134
rect 307804 633454 308404 668898
rect 307804 633218 307986 633454
rect 308222 633218 308404 633454
rect 307804 633134 308404 633218
rect 307804 632898 307986 633134
rect 308222 632898 308404 633134
rect 307804 597454 308404 632898
rect 307804 597218 307986 597454
rect 308222 597218 308404 597454
rect 307804 597134 308404 597218
rect 307804 596898 307986 597134
rect 308222 596898 308404 597134
rect 307804 561454 308404 596898
rect 307804 561218 307986 561454
rect 308222 561218 308404 561454
rect 307804 561134 308404 561218
rect 307804 560898 307986 561134
rect 308222 560898 308404 561134
rect 307804 525454 308404 560898
rect 307804 525218 307986 525454
rect 308222 525218 308404 525454
rect 307804 525134 308404 525218
rect 307804 524898 307986 525134
rect 308222 524898 308404 525134
rect 307804 510000 308404 524898
rect 311404 673054 312004 707102
rect 311404 672818 311586 673054
rect 311822 672818 312004 673054
rect 311404 672734 312004 672818
rect 311404 672498 311586 672734
rect 311822 672498 312004 672734
rect 311404 637054 312004 672498
rect 311404 636818 311586 637054
rect 311822 636818 312004 637054
rect 311404 636734 312004 636818
rect 311404 636498 311586 636734
rect 311822 636498 312004 636734
rect 311404 601054 312004 636498
rect 311404 600818 311586 601054
rect 311822 600818 312004 601054
rect 311404 600734 312004 600818
rect 311404 600498 311586 600734
rect 311822 600498 312004 600734
rect 311404 565054 312004 600498
rect 311404 564818 311586 565054
rect 311822 564818 312004 565054
rect 311404 564734 312004 564818
rect 311404 564498 311586 564734
rect 311822 564498 312004 564734
rect 311404 529054 312004 564498
rect 311404 528818 311586 529054
rect 311822 528818 312004 529054
rect 311404 528734 312004 528818
rect 311404 528498 311586 528734
rect 311822 528498 312004 528734
rect 311404 510000 312004 528498
rect 315004 676654 315604 708982
rect 315004 676418 315186 676654
rect 315422 676418 315604 676654
rect 315004 676334 315604 676418
rect 315004 676098 315186 676334
rect 315422 676098 315604 676334
rect 315004 640654 315604 676098
rect 315004 640418 315186 640654
rect 315422 640418 315604 640654
rect 315004 640334 315604 640418
rect 315004 640098 315186 640334
rect 315422 640098 315604 640334
rect 315004 604654 315604 640098
rect 315004 604418 315186 604654
rect 315422 604418 315604 604654
rect 315004 604334 315604 604418
rect 315004 604098 315186 604334
rect 315422 604098 315604 604334
rect 315004 568654 315604 604098
rect 315004 568418 315186 568654
rect 315422 568418 315604 568654
rect 315004 568334 315604 568418
rect 315004 568098 315186 568334
rect 315422 568098 315604 568334
rect 315004 532654 315604 568098
rect 315004 532418 315186 532654
rect 315422 532418 315604 532654
rect 315004 532334 315604 532418
rect 315004 532098 315186 532334
rect 315422 532098 315604 532334
rect 315004 510000 315604 532098
rect 318604 680254 319204 710862
rect 336604 710478 337204 711440
rect 336604 710242 336786 710478
rect 337022 710242 337204 710478
rect 336604 710158 337204 710242
rect 336604 709922 336786 710158
rect 337022 709922 337204 710158
rect 333004 708598 333604 709560
rect 333004 708362 333186 708598
rect 333422 708362 333604 708598
rect 333004 708278 333604 708362
rect 333004 708042 333186 708278
rect 333422 708042 333604 708278
rect 329404 706718 330004 707680
rect 329404 706482 329586 706718
rect 329822 706482 330004 706718
rect 329404 706398 330004 706482
rect 329404 706162 329586 706398
rect 329822 706162 330004 706398
rect 318604 680018 318786 680254
rect 319022 680018 319204 680254
rect 318604 679934 319204 680018
rect 318604 679698 318786 679934
rect 319022 679698 319204 679934
rect 318604 644254 319204 679698
rect 318604 644018 318786 644254
rect 319022 644018 319204 644254
rect 318604 643934 319204 644018
rect 318604 643698 318786 643934
rect 319022 643698 319204 643934
rect 318604 608254 319204 643698
rect 318604 608018 318786 608254
rect 319022 608018 319204 608254
rect 318604 607934 319204 608018
rect 318604 607698 318786 607934
rect 319022 607698 319204 607934
rect 318604 572254 319204 607698
rect 318604 572018 318786 572254
rect 319022 572018 319204 572254
rect 318604 571934 319204 572018
rect 318604 571698 318786 571934
rect 319022 571698 319204 571934
rect 318604 536254 319204 571698
rect 318604 536018 318786 536254
rect 319022 536018 319204 536254
rect 318604 535934 319204 536018
rect 318604 535698 318786 535934
rect 319022 535698 319204 535934
rect 318604 510000 319204 535698
rect 325804 704838 326404 705800
rect 325804 704602 325986 704838
rect 326222 704602 326404 704838
rect 325804 704518 326404 704602
rect 325804 704282 325986 704518
rect 326222 704282 326404 704518
rect 325804 687454 326404 704282
rect 325804 687218 325986 687454
rect 326222 687218 326404 687454
rect 325804 687134 326404 687218
rect 325804 686898 325986 687134
rect 326222 686898 326404 687134
rect 325804 651454 326404 686898
rect 325804 651218 325986 651454
rect 326222 651218 326404 651454
rect 325804 651134 326404 651218
rect 325804 650898 325986 651134
rect 326222 650898 326404 651134
rect 325804 615454 326404 650898
rect 325804 615218 325986 615454
rect 326222 615218 326404 615454
rect 325804 615134 326404 615218
rect 325804 614898 325986 615134
rect 326222 614898 326404 615134
rect 325804 579454 326404 614898
rect 325804 579218 325986 579454
rect 326222 579218 326404 579454
rect 325804 579134 326404 579218
rect 325804 578898 325986 579134
rect 326222 578898 326404 579134
rect 325804 543454 326404 578898
rect 325804 543218 325986 543454
rect 326222 543218 326404 543454
rect 325804 543134 326404 543218
rect 325804 542898 325986 543134
rect 326222 542898 326404 543134
rect 325804 510000 326404 542898
rect 329404 691054 330004 706162
rect 329404 690818 329586 691054
rect 329822 690818 330004 691054
rect 329404 690734 330004 690818
rect 329404 690498 329586 690734
rect 329822 690498 330004 690734
rect 329404 655054 330004 690498
rect 329404 654818 329586 655054
rect 329822 654818 330004 655054
rect 329404 654734 330004 654818
rect 329404 654498 329586 654734
rect 329822 654498 330004 654734
rect 329404 619054 330004 654498
rect 329404 618818 329586 619054
rect 329822 618818 330004 619054
rect 329404 618734 330004 618818
rect 329404 618498 329586 618734
rect 329822 618498 330004 618734
rect 329404 583054 330004 618498
rect 329404 582818 329586 583054
rect 329822 582818 330004 583054
rect 329404 582734 330004 582818
rect 329404 582498 329586 582734
rect 329822 582498 330004 582734
rect 329404 547054 330004 582498
rect 329404 546818 329586 547054
rect 329822 546818 330004 547054
rect 329404 546734 330004 546818
rect 329404 546498 329586 546734
rect 329822 546498 330004 546734
rect 329404 511054 330004 546498
rect 329404 510818 329586 511054
rect 329822 510818 330004 511054
rect 329404 510734 330004 510818
rect 329404 510498 329586 510734
rect 329822 510498 330004 510734
rect 329404 510000 330004 510498
rect 333004 694654 333604 708042
rect 333004 694418 333186 694654
rect 333422 694418 333604 694654
rect 333004 694334 333604 694418
rect 333004 694098 333186 694334
rect 333422 694098 333604 694334
rect 333004 658654 333604 694098
rect 333004 658418 333186 658654
rect 333422 658418 333604 658654
rect 333004 658334 333604 658418
rect 333004 658098 333186 658334
rect 333422 658098 333604 658334
rect 333004 622654 333604 658098
rect 333004 622418 333186 622654
rect 333422 622418 333604 622654
rect 333004 622334 333604 622418
rect 333004 622098 333186 622334
rect 333422 622098 333604 622334
rect 333004 586654 333604 622098
rect 333004 586418 333186 586654
rect 333422 586418 333604 586654
rect 333004 586334 333604 586418
rect 333004 586098 333186 586334
rect 333422 586098 333604 586334
rect 333004 550654 333604 586098
rect 333004 550418 333186 550654
rect 333422 550418 333604 550654
rect 333004 550334 333604 550418
rect 333004 550098 333186 550334
rect 333422 550098 333604 550334
rect 333004 514654 333604 550098
rect 333004 514418 333186 514654
rect 333422 514418 333604 514654
rect 333004 514334 333604 514418
rect 333004 514098 333186 514334
rect 333422 514098 333604 514334
rect 333004 510000 333604 514098
rect 336604 698254 337204 709922
rect 354604 711418 355204 711440
rect 354604 711182 354786 711418
rect 355022 711182 355204 711418
rect 354604 711098 355204 711182
rect 354604 710862 354786 711098
rect 355022 710862 355204 711098
rect 351004 709538 351604 709560
rect 351004 709302 351186 709538
rect 351422 709302 351604 709538
rect 351004 709218 351604 709302
rect 351004 708982 351186 709218
rect 351422 708982 351604 709218
rect 347404 707658 348004 707680
rect 347404 707422 347586 707658
rect 347822 707422 348004 707658
rect 347404 707338 348004 707422
rect 347404 707102 347586 707338
rect 347822 707102 348004 707338
rect 336604 698018 336786 698254
rect 337022 698018 337204 698254
rect 336604 697934 337204 698018
rect 336604 697698 336786 697934
rect 337022 697698 337204 697934
rect 336604 662254 337204 697698
rect 336604 662018 336786 662254
rect 337022 662018 337204 662254
rect 336604 661934 337204 662018
rect 336604 661698 336786 661934
rect 337022 661698 337204 661934
rect 336604 626254 337204 661698
rect 336604 626018 336786 626254
rect 337022 626018 337204 626254
rect 336604 625934 337204 626018
rect 336604 625698 336786 625934
rect 337022 625698 337204 625934
rect 336604 590254 337204 625698
rect 336604 590018 336786 590254
rect 337022 590018 337204 590254
rect 336604 589934 337204 590018
rect 336604 589698 336786 589934
rect 337022 589698 337204 589934
rect 336604 554254 337204 589698
rect 336604 554018 336786 554254
rect 337022 554018 337204 554254
rect 336604 553934 337204 554018
rect 336604 553698 336786 553934
rect 337022 553698 337204 553934
rect 336604 518254 337204 553698
rect 336604 518018 336786 518254
rect 337022 518018 337204 518254
rect 336604 517934 337204 518018
rect 336604 517698 336786 517934
rect 337022 517698 337204 517934
rect 336604 510000 337204 517698
rect 343804 705778 344404 705800
rect 343804 705542 343986 705778
rect 344222 705542 344404 705778
rect 343804 705458 344404 705542
rect 343804 705222 343986 705458
rect 344222 705222 344404 705458
rect 343804 669454 344404 705222
rect 343804 669218 343986 669454
rect 344222 669218 344404 669454
rect 343804 669134 344404 669218
rect 343804 668898 343986 669134
rect 344222 668898 344404 669134
rect 343804 633454 344404 668898
rect 343804 633218 343986 633454
rect 344222 633218 344404 633454
rect 343804 633134 344404 633218
rect 343804 632898 343986 633134
rect 344222 632898 344404 633134
rect 343804 597454 344404 632898
rect 343804 597218 343986 597454
rect 344222 597218 344404 597454
rect 343804 597134 344404 597218
rect 343804 596898 343986 597134
rect 344222 596898 344404 597134
rect 343804 561454 344404 596898
rect 343804 561218 343986 561454
rect 344222 561218 344404 561454
rect 343804 561134 344404 561218
rect 343804 560898 343986 561134
rect 344222 560898 344404 561134
rect 343804 525454 344404 560898
rect 343804 525218 343986 525454
rect 344222 525218 344404 525454
rect 343804 525134 344404 525218
rect 343804 524898 343986 525134
rect 344222 524898 344404 525134
rect 343804 510000 344404 524898
rect 347404 673054 348004 707102
rect 347404 672818 347586 673054
rect 347822 672818 348004 673054
rect 347404 672734 348004 672818
rect 347404 672498 347586 672734
rect 347822 672498 348004 672734
rect 347404 637054 348004 672498
rect 347404 636818 347586 637054
rect 347822 636818 348004 637054
rect 347404 636734 348004 636818
rect 347404 636498 347586 636734
rect 347822 636498 348004 636734
rect 347404 601054 348004 636498
rect 347404 600818 347586 601054
rect 347822 600818 348004 601054
rect 347404 600734 348004 600818
rect 347404 600498 347586 600734
rect 347822 600498 348004 600734
rect 347404 565054 348004 600498
rect 347404 564818 347586 565054
rect 347822 564818 348004 565054
rect 347404 564734 348004 564818
rect 347404 564498 347586 564734
rect 347822 564498 348004 564734
rect 347404 529054 348004 564498
rect 347404 528818 347586 529054
rect 347822 528818 348004 529054
rect 347404 528734 348004 528818
rect 347404 528498 347586 528734
rect 347822 528498 348004 528734
rect 347404 510000 348004 528498
rect 351004 676654 351604 708982
rect 351004 676418 351186 676654
rect 351422 676418 351604 676654
rect 351004 676334 351604 676418
rect 351004 676098 351186 676334
rect 351422 676098 351604 676334
rect 351004 640654 351604 676098
rect 351004 640418 351186 640654
rect 351422 640418 351604 640654
rect 351004 640334 351604 640418
rect 351004 640098 351186 640334
rect 351422 640098 351604 640334
rect 351004 604654 351604 640098
rect 351004 604418 351186 604654
rect 351422 604418 351604 604654
rect 351004 604334 351604 604418
rect 351004 604098 351186 604334
rect 351422 604098 351604 604334
rect 351004 568654 351604 604098
rect 351004 568418 351186 568654
rect 351422 568418 351604 568654
rect 351004 568334 351604 568418
rect 351004 568098 351186 568334
rect 351422 568098 351604 568334
rect 351004 532654 351604 568098
rect 351004 532418 351186 532654
rect 351422 532418 351604 532654
rect 351004 532334 351604 532418
rect 351004 532098 351186 532334
rect 351422 532098 351604 532334
rect 351004 510000 351604 532098
rect 354604 680254 355204 710862
rect 372604 710478 373204 711440
rect 372604 710242 372786 710478
rect 373022 710242 373204 710478
rect 372604 710158 373204 710242
rect 372604 709922 372786 710158
rect 373022 709922 373204 710158
rect 369004 708598 369604 709560
rect 369004 708362 369186 708598
rect 369422 708362 369604 708598
rect 369004 708278 369604 708362
rect 369004 708042 369186 708278
rect 369422 708042 369604 708278
rect 365404 706718 366004 707680
rect 365404 706482 365586 706718
rect 365822 706482 366004 706718
rect 365404 706398 366004 706482
rect 365404 706162 365586 706398
rect 365822 706162 366004 706398
rect 354604 680018 354786 680254
rect 355022 680018 355204 680254
rect 354604 679934 355204 680018
rect 354604 679698 354786 679934
rect 355022 679698 355204 679934
rect 354604 644254 355204 679698
rect 354604 644018 354786 644254
rect 355022 644018 355204 644254
rect 354604 643934 355204 644018
rect 354604 643698 354786 643934
rect 355022 643698 355204 643934
rect 354604 608254 355204 643698
rect 354604 608018 354786 608254
rect 355022 608018 355204 608254
rect 354604 607934 355204 608018
rect 354604 607698 354786 607934
rect 355022 607698 355204 607934
rect 354604 572254 355204 607698
rect 354604 572018 354786 572254
rect 355022 572018 355204 572254
rect 354604 571934 355204 572018
rect 354604 571698 354786 571934
rect 355022 571698 355204 571934
rect 354604 536254 355204 571698
rect 354604 536018 354786 536254
rect 355022 536018 355204 536254
rect 354604 535934 355204 536018
rect 354604 535698 354786 535934
rect 355022 535698 355204 535934
rect 354604 510000 355204 535698
rect 361804 704838 362404 705800
rect 361804 704602 361986 704838
rect 362222 704602 362404 704838
rect 361804 704518 362404 704602
rect 361804 704282 361986 704518
rect 362222 704282 362404 704518
rect 361804 687454 362404 704282
rect 361804 687218 361986 687454
rect 362222 687218 362404 687454
rect 361804 687134 362404 687218
rect 361804 686898 361986 687134
rect 362222 686898 362404 687134
rect 361804 651454 362404 686898
rect 361804 651218 361986 651454
rect 362222 651218 362404 651454
rect 361804 651134 362404 651218
rect 361804 650898 361986 651134
rect 362222 650898 362404 651134
rect 361804 615454 362404 650898
rect 361804 615218 361986 615454
rect 362222 615218 362404 615454
rect 361804 615134 362404 615218
rect 361804 614898 361986 615134
rect 362222 614898 362404 615134
rect 361804 579454 362404 614898
rect 361804 579218 361986 579454
rect 362222 579218 362404 579454
rect 361804 579134 362404 579218
rect 361804 578898 361986 579134
rect 362222 578898 362404 579134
rect 361804 543454 362404 578898
rect 361804 543218 361986 543454
rect 362222 543218 362404 543454
rect 361804 543134 362404 543218
rect 361804 542898 361986 543134
rect 362222 542898 362404 543134
rect 361804 510000 362404 542898
rect 365404 691054 366004 706162
rect 365404 690818 365586 691054
rect 365822 690818 366004 691054
rect 365404 690734 366004 690818
rect 365404 690498 365586 690734
rect 365822 690498 366004 690734
rect 365404 655054 366004 690498
rect 365404 654818 365586 655054
rect 365822 654818 366004 655054
rect 365404 654734 366004 654818
rect 365404 654498 365586 654734
rect 365822 654498 366004 654734
rect 365404 619054 366004 654498
rect 365404 618818 365586 619054
rect 365822 618818 366004 619054
rect 365404 618734 366004 618818
rect 365404 618498 365586 618734
rect 365822 618498 366004 618734
rect 365404 583054 366004 618498
rect 365404 582818 365586 583054
rect 365822 582818 366004 583054
rect 365404 582734 366004 582818
rect 365404 582498 365586 582734
rect 365822 582498 366004 582734
rect 365404 547054 366004 582498
rect 365404 546818 365586 547054
rect 365822 546818 366004 547054
rect 365404 546734 366004 546818
rect 365404 546498 365586 546734
rect 365822 546498 366004 546734
rect 365404 511054 366004 546498
rect 365404 510818 365586 511054
rect 365822 510818 366004 511054
rect 365404 510734 366004 510818
rect 365404 510498 365586 510734
rect 365822 510498 366004 510734
rect 365404 510000 366004 510498
rect 369004 694654 369604 708042
rect 369004 694418 369186 694654
rect 369422 694418 369604 694654
rect 369004 694334 369604 694418
rect 369004 694098 369186 694334
rect 369422 694098 369604 694334
rect 369004 658654 369604 694098
rect 369004 658418 369186 658654
rect 369422 658418 369604 658654
rect 369004 658334 369604 658418
rect 369004 658098 369186 658334
rect 369422 658098 369604 658334
rect 369004 622654 369604 658098
rect 369004 622418 369186 622654
rect 369422 622418 369604 622654
rect 369004 622334 369604 622418
rect 369004 622098 369186 622334
rect 369422 622098 369604 622334
rect 369004 586654 369604 622098
rect 369004 586418 369186 586654
rect 369422 586418 369604 586654
rect 369004 586334 369604 586418
rect 369004 586098 369186 586334
rect 369422 586098 369604 586334
rect 369004 550654 369604 586098
rect 369004 550418 369186 550654
rect 369422 550418 369604 550654
rect 369004 550334 369604 550418
rect 369004 550098 369186 550334
rect 369422 550098 369604 550334
rect 369004 514654 369604 550098
rect 369004 514418 369186 514654
rect 369422 514418 369604 514654
rect 369004 514334 369604 514418
rect 369004 514098 369186 514334
rect 369422 514098 369604 514334
rect 369004 510000 369604 514098
rect 372604 698254 373204 709922
rect 390604 711418 391204 711440
rect 390604 711182 390786 711418
rect 391022 711182 391204 711418
rect 390604 711098 391204 711182
rect 390604 710862 390786 711098
rect 391022 710862 391204 711098
rect 387004 709538 387604 709560
rect 387004 709302 387186 709538
rect 387422 709302 387604 709538
rect 387004 709218 387604 709302
rect 387004 708982 387186 709218
rect 387422 708982 387604 709218
rect 383404 707658 384004 707680
rect 383404 707422 383586 707658
rect 383822 707422 384004 707658
rect 383404 707338 384004 707422
rect 383404 707102 383586 707338
rect 383822 707102 384004 707338
rect 372604 698018 372786 698254
rect 373022 698018 373204 698254
rect 372604 697934 373204 698018
rect 372604 697698 372786 697934
rect 373022 697698 373204 697934
rect 372604 662254 373204 697698
rect 372604 662018 372786 662254
rect 373022 662018 373204 662254
rect 372604 661934 373204 662018
rect 372604 661698 372786 661934
rect 373022 661698 373204 661934
rect 372604 626254 373204 661698
rect 372604 626018 372786 626254
rect 373022 626018 373204 626254
rect 372604 625934 373204 626018
rect 372604 625698 372786 625934
rect 373022 625698 373204 625934
rect 372604 590254 373204 625698
rect 372604 590018 372786 590254
rect 373022 590018 373204 590254
rect 372604 589934 373204 590018
rect 372604 589698 372786 589934
rect 373022 589698 373204 589934
rect 372604 554254 373204 589698
rect 372604 554018 372786 554254
rect 373022 554018 373204 554254
rect 372604 553934 373204 554018
rect 372604 553698 372786 553934
rect 373022 553698 373204 553934
rect 372604 518254 373204 553698
rect 372604 518018 372786 518254
rect 373022 518018 373204 518254
rect 372604 517934 373204 518018
rect 372604 517698 372786 517934
rect 373022 517698 373204 517934
rect 372604 510000 373204 517698
rect 379804 705778 380404 705800
rect 379804 705542 379986 705778
rect 380222 705542 380404 705778
rect 379804 705458 380404 705542
rect 379804 705222 379986 705458
rect 380222 705222 380404 705458
rect 379804 669454 380404 705222
rect 379804 669218 379986 669454
rect 380222 669218 380404 669454
rect 379804 669134 380404 669218
rect 379804 668898 379986 669134
rect 380222 668898 380404 669134
rect 379804 633454 380404 668898
rect 379804 633218 379986 633454
rect 380222 633218 380404 633454
rect 379804 633134 380404 633218
rect 379804 632898 379986 633134
rect 380222 632898 380404 633134
rect 379804 597454 380404 632898
rect 379804 597218 379986 597454
rect 380222 597218 380404 597454
rect 379804 597134 380404 597218
rect 379804 596898 379986 597134
rect 380222 596898 380404 597134
rect 379804 561454 380404 596898
rect 379804 561218 379986 561454
rect 380222 561218 380404 561454
rect 379804 561134 380404 561218
rect 379804 560898 379986 561134
rect 380222 560898 380404 561134
rect 379804 525454 380404 560898
rect 379804 525218 379986 525454
rect 380222 525218 380404 525454
rect 379804 525134 380404 525218
rect 379804 524898 379986 525134
rect 380222 524898 380404 525134
rect 379804 510000 380404 524898
rect 383404 673054 384004 707102
rect 383404 672818 383586 673054
rect 383822 672818 384004 673054
rect 383404 672734 384004 672818
rect 383404 672498 383586 672734
rect 383822 672498 384004 672734
rect 383404 637054 384004 672498
rect 383404 636818 383586 637054
rect 383822 636818 384004 637054
rect 383404 636734 384004 636818
rect 383404 636498 383586 636734
rect 383822 636498 384004 636734
rect 383404 601054 384004 636498
rect 383404 600818 383586 601054
rect 383822 600818 384004 601054
rect 383404 600734 384004 600818
rect 383404 600498 383586 600734
rect 383822 600498 384004 600734
rect 383404 565054 384004 600498
rect 383404 564818 383586 565054
rect 383822 564818 384004 565054
rect 383404 564734 384004 564818
rect 383404 564498 383586 564734
rect 383822 564498 384004 564734
rect 383404 529054 384004 564498
rect 383404 528818 383586 529054
rect 383822 528818 384004 529054
rect 383404 528734 384004 528818
rect 383404 528498 383586 528734
rect 383822 528498 384004 528734
rect 383404 510000 384004 528498
rect 387004 676654 387604 708982
rect 387004 676418 387186 676654
rect 387422 676418 387604 676654
rect 387004 676334 387604 676418
rect 387004 676098 387186 676334
rect 387422 676098 387604 676334
rect 387004 640654 387604 676098
rect 387004 640418 387186 640654
rect 387422 640418 387604 640654
rect 387004 640334 387604 640418
rect 387004 640098 387186 640334
rect 387422 640098 387604 640334
rect 387004 604654 387604 640098
rect 387004 604418 387186 604654
rect 387422 604418 387604 604654
rect 387004 604334 387604 604418
rect 387004 604098 387186 604334
rect 387422 604098 387604 604334
rect 387004 568654 387604 604098
rect 387004 568418 387186 568654
rect 387422 568418 387604 568654
rect 387004 568334 387604 568418
rect 387004 568098 387186 568334
rect 387422 568098 387604 568334
rect 387004 532654 387604 568098
rect 387004 532418 387186 532654
rect 387422 532418 387604 532654
rect 387004 532334 387604 532418
rect 387004 532098 387186 532334
rect 387422 532098 387604 532334
rect 387004 510000 387604 532098
rect 390604 680254 391204 710862
rect 408604 710478 409204 711440
rect 408604 710242 408786 710478
rect 409022 710242 409204 710478
rect 408604 710158 409204 710242
rect 408604 709922 408786 710158
rect 409022 709922 409204 710158
rect 405004 708598 405604 709560
rect 405004 708362 405186 708598
rect 405422 708362 405604 708598
rect 405004 708278 405604 708362
rect 405004 708042 405186 708278
rect 405422 708042 405604 708278
rect 401404 706718 402004 707680
rect 401404 706482 401586 706718
rect 401822 706482 402004 706718
rect 401404 706398 402004 706482
rect 401404 706162 401586 706398
rect 401822 706162 402004 706398
rect 390604 680018 390786 680254
rect 391022 680018 391204 680254
rect 390604 679934 391204 680018
rect 390604 679698 390786 679934
rect 391022 679698 391204 679934
rect 390604 644254 391204 679698
rect 390604 644018 390786 644254
rect 391022 644018 391204 644254
rect 390604 643934 391204 644018
rect 390604 643698 390786 643934
rect 391022 643698 391204 643934
rect 390604 608254 391204 643698
rect 390604 608018 390786 608254
rect 391022 608018 391204 608254
rect 390604 607934 391204 608018
rect 390604 607698 390786 607934
rect 391022 607698 391204 607934
rect 390604 572254 391204 607698
rect 390604 572018 390786 572254
rect 391022 572018 391204 572254
rect 390604 571934 391204 572018
rect 390604 571698 390786 571934
rect 391022 571698 391204 571934
rect 390604 536254 391204 571698
rect 390604 536018 390786 536254
rect 391022 536018 391204 536254
rect 390604 535934 391204 536018
rect 390604 535698 390786 535934
rect 391022 535698 391204 535934
rect 390604 510000 391204 535698
rect 397804 704838 398404 705800
rect 397804 704602 397986 704838
rect 398222 704602 398404 704838
rect 397804 704518 398404 704602
rect 397804 704282 397986 704518
rect 398222 704282 398404 704518
rect 397804 687454 398404 704282
rect 397804 687218 397986 687454
rect 398222 687218 398404 687454
rect 397804 687134 398404 687218
rect 397804 686898 397986 687134
rect 398222 686898 398404 687134
rect 397804 651454 398404 686898
rect 397804 651218 397986 651454
rect 398222 651218 398404 651454
rect 397804 651134 398404 651218
rect 397804 650898 397986 651134
rect 398222 650898 398404 651134
rect 397804 615454 398404 650898
rect 397804 615218 397986 615454
rect 398222 615218 398404 615454
rect 397804 615134 398404 615218
rect 397804 614898 397986 615134
rect 398222 614898 398404 615134
rect 397804 579454 398404 614898
rect 397804 579218 397986 579454
rect 398222 579218 398404 579454
rect 397804 579134 398404 579218
rect 397804 578898 397986 579134
rect 398222 578898 398404 579134
rect 397804 543454 398404 578898
rect 397804 543218 397986 543454
rect 398222 543218 398404 543454
rect 397804 543134 398404 543218
rect 397804 542898 397986 543134
rect 398222 542898 398404 543134
rect 397804 510000 398404 542898
rect 401404 691054 402004 706162
rect 401404 690818 401586 691054
rect 401822 690818 402004 691054
rect 401404 690734 402004 690818
rect 401404 690498 401586 690734
rect 401822 690498 402004 690734
rect 401404 655054 402004 690498
rect 401404 654818 401586 655054
rect 401822 654818 402004 655054
rect 401404 654734 402004 654818
rect 401404 654498 401586 654734
rect 401822 654498 402004 654734
rect 401404 619054 402004 654498
rect 401404 618818 401586 619054
rect 401822 618818 402004 619054
rect 401404 618734 402004 618818
rect 401404 618498 401586 618734
rect 401822 618498 402004 618734
rect 401404 583054 402004 618498
rect 401404 582818 401586 583054
rect 401822 582818 402004 583054
rect 401404 582734 402004 582818
rect 401404 582498 401586 582734
rect 401822 582498 402004 582734
rect 401404 547054 402004 582498
rect 401404 546818 401586 547054
rect 401822 546818 402004 547054
rect 401404 546734 402004 546818
rect 401404 546498 401586 546734
rect 401822 546498 402004 546734
rect 401404 511054 402004 546498
rect 401404 510818 401586 511054
rect 401822 510818 402004 511054
rect 401404 510734 402004 510818
rect 401404 510498 401586 510734
rect 401822 510498 402004 510734
rect 401404 510000 402004 510498
rect 405004 694654 405604 708042
rect 405004 694418 405186 694654
rect 405422 694418 405604 694654
rect 405004 694334 405604 694418
rect 405004 694098 405186 694334
rect 405422 694098 405604 694334
rect 405004 658654 405604 694098
rect 405004 658418 405186 658654
rect 405422 658418 405604 658654
rect 405004 658334 405604 658418
rect 405004 658098 405186 658334
rect 405422 658098 405604 658334
rect 405004 622654 405604 658098
rect 405004 622418 405186 622654
rect 405422 622418 405604 622654
rect 405004 622334 405604 622418
rect 405004 622098 405186 622334
rect 405422 622098 405604 622334
rect 405004 586654 405604 622098
rect 405004 586418 405186 586654
rect 405422 586418 405604 586654
rect 405004 586334 405604 586418
rect 405004 586098 405186 586334
rect 405422 586098 405604 586334
rect 405004 550654 405604 586098
rect 405004 550418 405186 550654
rect 405422 550418 405604 550654
rect 405004 550334 405604 550418
rect 405004 550098 405186 550334
rect 405422 550098 405604 550334
rect 405004 514654 405604 550098
rect 405004 514418 405186 514654
rect 405422 514418 405604 514654
rect 405004 514334 405604 514418
rect 405004 514098 405186 514334
rect 405422 514098 405604 514334
rect 405004 510000 405604 514098
rect 408604 698254 409204 709922
rect 426604 711418 427204 711440
rect 426604 711182 426786 711418
rect 427022 711182 427204 711418
rect 426604 711098 427204 711182
rect 426604 710862 426786 711098
rect 427022 710862 427204 711098
rect 423004 709538 423604 709560
rect 423004 709302 423186 709538
rect 423422 709302 423604 709538
rect 423004 709218 423604 709302
rect 423004 708982 423186 709218
rect 423422 708982 423604 709218
rect 419404 707658 420004 707680
rect 419404 707422 419586 707658
rect 419822 707422 420004 707658
rect 419404 707338 420004 707422
rect 419404 707102 419586 707338
rect 419822 707102 420004 707338
rect 408604 698018 408786 698254
rect 409022 698018 409204 698254
rect 408604 697934 409204 698018
rect 408604 697698 408786 697934
rect 409022 697698 409204 697934
rect 408604 662254 409204 697698
rect 408604 662018 408786 662254
rect 409022 662018 409204 662254
rect 408604 661934 409204 662018
rect 408604 661698 408786 661934
rect 409022 661698 409204 661934
rect 408604 626254 409204 661698
rect 408604 626018 408786 626254
rect 409022 626018 409204 626254
rect 408604 625934 409204 626018
rect 408604 625698 408786 625934
rect 409022 625698 409204 625934
rect 408604 590254 409204 625698
rect 408604 590018 408786 590254
rect 409022 590018 409204 590254
rect 408604 589934 409204 590018
rect 408604 589698 408786 589934
rect 409022 589698 409204 589934
rect 408604 554254 409204 589698
rect 408604 554018 408786 554254
rect 409022 554018 409204 554254
rect 408604 553934 409204 554018
rect 408604 553698 408786 553934
rect 409022 553698 409204 553934
rect 408604 518254 409204 553698
rect 408604 518018 408786 518254
rect 409022 518018 409204 518254
rect 408604 517934 409204 518018
rect 408604 517698 408786 517934
rect 409022 517698 409204 517934
rect 408604 510000 409204 517698
rect 415804 705778 416404 705800
rect 415804 705542 415986 705778
rect 416222 705542 416404 705778
rect 415804 705458 416404 705542
rect 415804 705222 415986 705458
rect 416222 705222 416404 705458
rect 415804 669454 416404 705222
rect 415804 669218 415986 669454
rect 416222 669218 416404 669454
rect 415804 669134 416404 669218
rect 415804 668898 415986 669134
rect 416222 668898 416404 669134
rect 415804 633454 416404 668898
rect 415804 633218 415986 633454
rect 416222 633218 416404 633454
rect 415804 633134 416404 633218
rect 415804 632898 415986 633134
rect 416222 632898 416404 633134
rect 415804 597454 416404 632898
rect 415804 597218 415986 597454
rect 416222 597218 416404 597454
rect 415804 597134 416404 597218
rect 415804 596898 415986 597134
rect 416222 596898 416404 597134
rect 415804 561454 416404 596898
rect 415804 561218 415986 561454
rect 416222 561218 416404 561454
rect 415804 561134 416404 561218
rect 415804 560898 415986 561134
rect 416222 560898 416404 561134
rect 415804 525454 416404 560898
rect 415804 525218 415986 525454
rect 416222 525218 416404 525454
rect 415804 525134 416404 525218
rect 415804 524898 415986 525134
rect 416222 524898 416404 525134
rect 415804 510000 416404 524898
rect 419404 673054 420004 707102
rect 419404 672818 419586 673054
rect 419822 672818 420004 673054
rect 419404 672734 420004 672818
rect 419404 672498 419586 672734
rect 419822 672498 420004 672734
rect 419404 637054 420004 672498
rect 419404 636818 419586 637054
rect 419822 636818 420004 637054
rect 419404 636734 420004 636818
rect 419404 636498 419586 636734
rect 419822 636498 420004 636734
rect 419404 601054 420004 636498
rect 419404 600818 419586 601054
rect 419822 600818 420004 601054
rect 419404 600734 420004 600818
rect 419404 600498 419586 600734
rect 419822 600498 420004 600734
rect 419404 565054 420004 600498
rect 419404 564818 419586 565054
rect 419822 564818 420004 565054
rect 419404 564734 420004 564818
rect 419404 564498 419586 564734
rect 419822 564498 420004 564734
rect 419404 529054 420004 564498
rect 419404 528818 419586 529054
rect 419822 528818 420004 529054
rect 419404 528734 420004 528818
rect 419404 528498 419586 528734
rect 419822 528498 420004 528734
rect 419404 510000 420004 528498
rect 423004 676654 423604 708982
rect 423004 676418 423186 676654
rect 423422 676418 423604 676654
rect 423004 676334 423604 676418
rect 423004 676098 423186 676334
rect 423422 676098 423604 676334
rect 423004 640654 423604 676098
rect 423004 640418 423186 640654
rect 423422 640418 423604 640654
rect 423004 640334 423604 640418
rect 423004 640098 423186 640334
rect 423422 640098 423604 640334
rect 423004 604654 423604 640098
rect 423004 604418 423186 604654
rect 423422 604418 423604 604654
rect 423004 604334 423604 604418
rect 423004 604098 423186 604334
rect 423422 604098 423604 604334
rect 423004 568654 423604 604098
rect 423004 568418 423186 568654
rect 423422 568418 423604 568654
rect 423004 568334 423604 568418
rect 423004 568098 423186 568334
rect 423422 568098 423604 568334
rect 423004 532654 423604 568098
rect 423004 532418 423186 532654
rect 423422 532418 423604 532654
rect 423004 532334 423604 532418
rect 423004 532098 423186 532334
rect 423422 532098 423604 532334
rect 423004 510000 423604 532098
rect 426604 680254 427204 710862
rect 444604 710478 445204 711440
rect 444604 710242 444786 710478
rect 445022 710242 445204 710478
rect 444604 710158 445204 710242
rect 444604 709922 444786 710158
rect 445022 709922 445204 710158
rect 441004 708598 441604 709560
rect 441004 708362 441186 708598
rect 441422 708362 441604 708598
rect 441004 708278 441604 708362
rect 441004 708042 441186 708278
rect 441422 708042 441604 708278
rect 437404 706718 438004 707680
rect 437404 706482 437586 706718
rect 437822 706482 438004 706718
rect 437404 706398 438004 706482
rect 437404 706162 437586 706398
rect 437822 706162 438004 706398
rect 426604 680018 426786 680254
rect 427022 680018 427204 680254
rect 426604 679934 427204 680018
rect 426604 679698 426786 679934
rect 427022 679698 427204 679934
rect 426604 644254 427204 679698
rect 426604 644018 426786 644254
rect 427022 644018 427204 644254
rect 426604 643934 427204 644018
rect 426604 643698 426786 643934
rect 427022 643698 427204 643934
rect 426604 608254 427204 643698
rect 426604 608018 426786 608254
rect 427022 608018 427204 608254
rect 426604 607934 427204 608018
rect 426604 607698 426786 607934
rect 427022 607698 427204 607934
rect 426604 572254 427204 607698
rect 426604 572018 426786 572254
rect 427022 572018 427204 572254
rect 426604 571934 427204 572018
rect 426604 571698 426786 571934
rect 427022 571698 427204 571934
rect 426604 536254 427204 571698
rect 426604 536018 426786 536254
rect 427022 536018 427204 536254
rect 426604 535934 427204 536018
rect 426604 535698 426786 535934
rect 427022 535698 427204 535934
rect 426604 510000 427204 535698
rect 433804 704838 434404 705800
rect 433804 704602 433986 704838
rect 434222 704602 434404 704838
rect 433804 704518 434404 704602
rect 433804 704282 433986 704518
rect 434222 704282 434404 704518
rect 433804 687454 434404 704282
rect 433804 687218 433986 687454
rect 434222 687218 434404 687454
rect 433804 687134 434404 687218
rect 433804 686898 433986 687134
rect 434222 686898 434404 687134
rect 433804 651454 434404 686898
rect 433804 651218 433986 651454
rect 434222 651218 434404 651454
rect 433804 651134 434404 651218
rect 433804 650898 433986 651134
rect 434222 650898 434404 651134
rect 433804 615454 434404 650898
rect 433804 615218 433986 615454
rect 434222 615218 434404 615454
rect 433804 615134 434404 615218
rect 433804 614898 433986 615134
rect 434222 614898 434404 615134
rect 433804 579454 434404 614898
rect 433804 579218 433986 579454
rect 434222 579218 434404 579454
rect 433804 579134 434404 579218
rect 433804 578898 433986 579134
rect 434222 578898 434404 579134
rect 433804 543454 434404 578898
rect 433804 543218 433986 543454
rect 434222 543218 434404 543454
rect 433804 543134 434404 543218
rect 433804 542898 433986 543134
rect 434222 542898 434404 543134
rect 433804 510000 434404 542898
rect 437404 691054 438004 706162
rect 437404 690818 437586 691054
rect 437822 690818 438004 691054
rect 437404 690734 438004 690818
rect 437404 690498 437586 690734
rect 437822 690498 438004 690734
rect 437404 655054 438004 690498
rect 437404 654818 437586 655054
rect 437822 654818 438004 655054
rect 437404 654734 438004 654818
rect 437404 654498 437586 654734
rect 437822 654498 438004 654734
rect 437404 619054 438004 654498
rect 437404 618818 437586 619054
rect 437822 618818 438004 619054
rect 437404 618734 438004 618818
rect 437404 618498 437586 618734
rect 437822 618498 438004 618734
rect 437404 583054 438004 618498
rect 437404 582818 437586 583054
rect 437822 582818 438004 583054
rect 437404 582734 438004 582818
rect 437404 582498 437586 582734
rect 437822 582498 438004 582734
rect 437404 547054 438004 582498
rect 437404 546818 437586 547054
rect 437822 546818 438004 547054
rect 437404 546734 438004 546818
rect 437404 546498 437586 546734
rect 437822 546498 438004 546734
rect 437404 511054 438004 546498
rect 437404 510818 437586 511054
rect 437822 510818 438004 511054
rect 437404 510734 438004 510818
rect 437404 510498 437586 510734
rect 437822 510498 438004 510734
rect 437404 510000 438004 510498
rect 441004 694654 441604 708042
rect 441004 694418 441186 694654
rect 441422 694418 441604 694654
rect 441004 694334 441604 694418
rect 441004 694098 441186 694334
rect 441422 694098 441604 694334
rect 441004 658654 441604 694098
rect 441004 658418 441186 658654
rect 441422 658418 441604 658654
rect 441004 658334 441604 658418
rect 441004 658098 441186 658334
rect 441422 658098 441604 658334
rect 441004 622654 441604 658098
rect 441004 622418 441186 622654
rect 441422 622418 441604 622654
rect 441004 622334 441604 622418
rect 441004 622098 441186 622334
rect 441422 622098 441604 622334
rect 441004 586654 441604 622098
rect 441004 586418 441186 586654
rect 441422 586418 441604 586654
rect 441004 586334 441604 586418
rect 441004 586098 441186 586334
rect 441422 586098 441604 586334
rect 441004 550654 441604 586098
rect 441004 550418 441186 550654
rect 441422 550418 441604 550654
rect 441004 550334 441604 550418
rect 441004 550098 441186 550334
rect 441422 550098 441604 550334
rect 441004 514654 441604 550098
rect 441004 514418 441186 514654
rect 441422 514418 441604 514654
rect 441004 514334 441604 514418
rect 441004 514098 441186 514334
rect 441422 514098 441604 514334
rect 153004 478418 153186 478654
rect 153422 478418 153604 478654
rect 153004 478334 153604 478418
rect 153004 478098 153186 478334
rect 153422 478098 153604 478334
rect 153004 442654 153604 478098
rect 153004 442418 153186 442654
rect 153422 442418 153604 442654
rect 153004 442334 153604 442418
rect 153004 442098 153186 442334
rect 153422 442098 153604 442334
rect 153004 406654 153604 442098
rect 153004 406418 153186 406654
rect 153422 406418 153604 406654
rect 153004 406334 153604 406418
rect 153004 406098 153186 406334
rect 153422 406098 153604 406334
rect 153004 370654 153604 406098
rect 153004 370418 153186 370654
rect 153422 370418 153604 370654
rect 153004 370334 153604 370418
rect 153004 370098 153186 370334
rect 153422 370098 153604 370334
rect 153004 334654 153604 370098
rect 441004 478654 441604 514098
rect 441004 478418 441186 478654
rect 441422 478418 441604 478654
rect 441004 478334 441604 478418
rect 441004 478098 441186 478334
rect 441422 478098 441604 478334
rect 441004 442654 441604 478098
rect 441004 442418 441186 442654
rect 441422 442418 441604 442654
rect 441004 442334 441604 442418
rect 441004 442098 441186 442334
rect 441422 442098 441604 442334
rect 441004 406654 441604 442098
rect 441004 406418 441186 406654
rect 441422 406418 441604 406654
rect 441004 406334 441604 406418
rect 441004 406098 441186 406334
rect 441422 406098 441604 406334
rect 441004 370654 441604 406098
rect 441004 370418 441186 370654
rect 441422 370418 441604 370654
rect 441004 370334 441604 370418
rect 441004 370098 441186 370334
rect 441422 370098 441604 370334
rect 429699 342548 429765 342549
rect 429699 342484 429700 342548
rect 429764 342484 429765 342548
rect 429699 342483 429765 342484
rect 153004 334418 153186 334654
rect 153422 334418 153604 334654
rect 153004 334334 153604 334418
rect 153004 334098 153186 334334
rect 153422 334098 153604 334334
rect 153004 298654 153604 334098
rect 153004 298418 153186 298654
rect 153422 298418 153604 298654
rect 153004 298334 153604 298418
rect 153004 298098 153186 298334
rect 153422 298098 153604 298334
rect 153004 262654 153604 298098
rect 153004 262418 153186 262654
rect 153422 262418 153604 262654
rect 153004 262334 153604 262418
rect 153004 262098 153186 262334
rect 153422 262098 153604 262334
rect 153004 226654 153604 262098
rect 153004 226418 153186 226654
rect 153422 226418 153604 226654
rect 153004 226334 153604 226418
rect 153004 226098 153186 226334
rect 153422 226098 153604 226334
rect 153004 190654 153604 226098
rect 153004 190418 153186 190654
rect 153422 190418 153604 190654
rect 153004 190334 153604 190418
rect 153004 190098 153186 190334
rect 153422 190098 153604 190334
rect 153004 154654 153604 190098
rect 153004 154418 153186 154654
rect 153422 154418 153604 154654
rect 153004 154334 153604 154418
rect 153004 154098 153186 154334
rect 153422 154098 153604 154334
rect 153004 118654 153604 154098
rect 153004 118418 153186 118654
rect 153422 118418 153604 118654
rect 153004 118334 153604 118418
rect 153004 118098 153186 118334
rect 153422 118098 153604 118334
rect 153004 82654 153604 118098
rect 153004 82418 153186 82654
rect 153422 82418 153604 82654
rect 153004 82334 153604 82418
rect 153004 82098 153186 82334
rect 153422 82098 153604 82334
rect 153004 46654 153604 82098
rect 153004 46418 153186 46654
rect 153422 46418 153604 46654
rect 153004 46334 153604 46418
rect 153004 46098 153186 46334
rect 153422 46098 153604 46334
rect 153004 10654 153604 46098
rect 153004 10418 153186 10654
rect 153422 10418 153604 10654
rect 153004 10334 153604 10418
rect 153004 10098 153186 10334
rect 153422 10098 153604 10334
rect 153004 -4106 153604 10098
rect 153004 -4342 153186 -4106
rect 153422 -4342 153604 -4106
rect 153004 -4426 153604 -4342
rect 153004 -4662 153186 -4426
rect 153422 -4662 153604 -4426
rect 153004 -5624 153604 -4662
rect 156604 302254 157204 326000
rect 156604 302018 156786 302254
rect 157022 302018 157204 302254
rect 156604 301934 157204 302018
rect 156604 301698 156786 301934
rect 157022 301698 157204 301934
rect 156604 266254 157204 301698
rect 156604 266018 156786 266254
rect 157022 266018 157204 266254
rect 156604 265934 157204 266018
rect 156604 265698 156786 265934
rect 157022 265698 157204 265934
rect 156604 230254 157204 265698
rect 156604 230018 156786 230254
rect 157022 230018 157204 230254
rect 156604 229934 157204 230018
rect 156604 229698 156786 229934
rect 157022 229698 157204 229934
rect 156604 194254 157204 229698
rect 156604 194018 156786 194254
rect 157022 194018 157204 194254
rect 156604 193934 157204 194018
rect 156604 193698 156786 193934
rect 157022 193698 157204 193934
rect 156604 158254 157204 193698
rect 156604 158018 156786 158254
rect 157022 158018 157204 158254
rect 156604 157934 157204 158018
rect 156604 157698 156786 157934
rect 157022 157698 157204 157934
rect 156604 122254 157204 157698
rect 156604 122018 156786 122254
rect 157022 122018 157204 122254
rect 156604 121934 157204 122018
rect 156604 121698 156786 121934
rect 157022 121698 157204 121934
rect 156604 86254 157204 121698
rect 156604 86018 156786 86254
rect 157022 86018 157204 86254
rect 156604 85934 157204 86018
rect 156604 85698 156786 85934
rect 157022 85698 157204 85934
rect 156604 50254 157204 85698
rect 156604 50018 156786 50254
rect 157022 50018 157204 50254
rect 156604 49934 157204 50018
rect 156604 49698 156786 49934
rect 157022 49698 157204 49934
rect 156604 14254 157204 49698
rect 156604 14018 156786 14254
rect 157022 14018 157204 14254
rect 156604 13934 157204 14018
rect 156604 13698 156786 13934
rect 157022 13698 157204 13934
rect 138604 -7162 138786 -6926
rect 139022 -7162 139204 -6926
rect 138604 -7246 139204 -7162
rect 138604 -7482 138786 -7246
rect 139022 -7482 139204 -7246
rect 138604 -7504 139204 -7482
rect 156604 -5986 157204 13698
rect 163804 309454 164404 326000
rect 163804 309218 163986 309454
rect 164222 309218 164404 309454
rect 163804 309134 164404 309218
rect 163804 308898 163986 309134
rect 164222 308898 164404 309134
rect 163804 273454 164404 308898
rect 163804 273218 163986 273454
rect 164222 273218 164404 273454
rect 163804 273134 164404 273218
rect 163804 272898 163986 273134
rect 164222 272898 164404 273134
rect 163804 237454 164404 272898
rect 163804 237218 163986 237454
rect 164222 237218 164404 237454
rect 163804 237134 164404 237218
rect 163804 236898 163986 237134
rect 164222 236898 164404 237134
rect 163804 201454 164404 236898
rect 163804 201218 163986 201454
rect 164222 201218 164404 201454
rect 163804 201134 164404 201218
rect 163804 200898 163986 201134
rect 164222 200898 164404 201134
rect 163804 165454 164404 200898
rect 163804 165218 163986 165454
rect 164222 165218 164404 165454
rect 163804 165134 164404 165218
rect 163804 164898 163986 165134
rect 164222 164898 164404 165134
rect 163804 129454 164404 164898
rect 163804 129218 163986 129454
rect 164222 129218 164404 129454
rect 163804 129134 164404 129218
rect 163804 128898 163986 129134
rect 164222 128898 164404 129134
rect 163804 93454 164404 128898
rect 163804 93218 163986 93454
rect 164222 93218 164404 93454
rect 163804 93134 164404 93218
rect 163804 92898 163986 93134
rect 164222 92898 164404 93134
rect 163804 57454 164404 92898
rect 163804 57218 163986 57454
rect 164222 57218 164404 57454
rect 163804 57134 164404 57218
rect 163804 56898 163986 57134
rect 164222 56898 164404 57134
rect 163804 21454 164404 56898
rect 163804 21218 163986 21454
rect 164222 21218 164404 21454
rect 163804 21134 164404 21218
rect 163804 20898 163986 21134
rect 164222 20898 164404 21134
rect 163804 -1286 164404 20898
rect 163804 -1522 163986 -1286
rect 164222 -1522 164404 -1286
rect 163804 -1606 164404 -1522
rect 163804 -1842 163986 -1606
rect 164222 -1842 164404 -1606
rect 163804 -1864 164404 -1842
rect 167404 313054 168004 326000
rect 167404 312818 167586 313054
rect 167822 312818 168004 313054
rect 167404 312734 168004 312818
rect 167404 312498 167586 312734
rect 167822 312498 168004 312734
rect 167404 277054 168004 312498
rect 167404 276818 167586 277054
rect 167822 276818 168004 277054
rect 167404 276734 168004 276818
rect 167404 276498 167586 276734
rect 167822 276498 168004 276734
rect 167404 241054 168004 276498
rect 167404 240818 167586 241054
rect 167822 240818 168004 241054
rect 167404 240734 168004 240818
rect 167404 240498 167586 240734
rect 167822 240498 168004 240734
rect 167404 205054 168004 240498
rect 167404 204818 167586 205054
rect 167822 204818 168004 205054
rect 167404 204734 168004 204818
rect 167404 204498 167586 204734
rect 167822 204498 168004 204734
rect 167404 169054 168004 204498
rect 167404 168818 167586 169054
rect 167822 168818 168004 169054
rect 167404 168734 168004 168818
rect 167404 168498 167586 168734
rect 167822 168498 168004 168734
rect 167404 133054 168004 168498
rect 167404 132818 167586 133054
rect 167822 132818 168004 133054
rect 167404 132734 168004 132818
rect 167404 132498 167586 132734
rect 167822 132498 168004 132734
rect 167404 97054 168004 132498
rect 167404 96818 167586 97054
rect 167822 96818 168004 97054
rect 167404 96734 168004 96818
rect 167404 96498 167586 96734
rect 167822 96498 168004 96734
rect 167404 61054 168004 96498
rect 167404 60818 167586 61054
rect 167822 60818 168004 61054
rect 167404 60734 168004 60818
rect 167404 60498 167586 60734
rect 167822 60498 168004 60734
rect 167404 25054 168004 60498
rect 167404 24818 167586 25054
rect 167822 24818 168004 25054
rect 167404 24734 168004 24818
rect 167404 24498 167586 24734
rect 167822 24498 168004 24734
rect 167404 -3166 168004 24498
rect 167404 -3402 167586 -3166
rect 167822 -3402 168004 -3166
rect 167404 -3486 168004 -3402
rect 167404 -3722 167586 -3486
rect 167822 -3722 168004 -3486
rect 167404 -3744 168004 -3722
rect 171004 316654 171604 326000
rect 171004 316418 171186 316654
rect 171422 316418 171604 316654
rect 171004 316334 171604 316418
rect 171004 316098 171186 316334
rect 171422 316098 171604 316334
rect 171004 280654 171604 316098
rect 171004 280418 171186 280654
rect 171422 280418 171604 280654
rect 171004 280334 171604 280418
rect 171004 280098 171186 280334
rect 171422 280098 171604 280334
rect 171004 244654 171604 280098
rect 171004 244418 171186 244654
rect 171422 244418 171604 244654
rect 171004 244334 171604 244418
rect 171004 244098 171186 244334
rect 171422 244098 171604 244334
rect 171004 208654 171604 244098
rect 171004 208418 171186 208654
rect 171422 208418 171604 208654
rect 171004 208334 171604 208418
rect 171004 208098 171186 208334
rect 171422 208098 171604 208334
rect 171004 172654 171604 208098
rect 171004 172418 171186 172654
rect 171422 172418 171604 172654
rect 171004 172334 171604 172418
rect 171004 172098 171186 172334
rect 171422 172098 171604 172334
rect 171004 136654 171604 172098
rect 171004 136418 171186 136654
rect 171422 136418 171604 136654
rect 171004 136334 171604 136418
rect 171004 136098 171186 136334
rect 171422 136098 171604 136334
rect 171004 100654 171604 136098
rect 171004 100418 171186 100654
rect 171422 100418 171604 100654
rect 171004 100334 171604 100418
rect 171004 100098 171186 100334
rect 171422 100098 171604 100334
rect 171004 64654 171604 100098
rect 171004 64418 171186 64654
rect 171422 64418 171604 64654
rect 171004 64334 171604 64418
rect 171004 64098 171186 64334
rect 171422 64098 171604 64334
rect 171004 28654 171604 64098
rect 171004 28418 171186 28654
rect 171422 28418 171604 28654
rect 171004 28334 171604 28418
rect 171004 28098 171186 28334
rect 171422 28098 171604 28334
rect 171004 -5046 171604 28098
rect 171004 -5282 171186 -5046
rect 171422 -5282 171604 -5046
rect 171004 -5366 171604 -5282
rect 171004 -5602 171186 -5366
rect 171422 -5602 171604 -5366
rect 171004 -5624 171604 -5602
rect 174604 320254 175204 326000
rect 174604 320018 174786 320254
rect 175022 320018 175204 320254
rect 174604 319934 175204 320018
rect 174604 319698 174786 319934
rect 175022 319698 175204 319934
rect 174604 284254 175204 319698
rect 174604 284018 174786 284254
rect 175022 284018 175204 284254
rect 174604 283934 175204 284018
rect 174604 283698 174786 283934
rect 175022 283698 175204 283934
rect 174604 248254 175204 283698
rect 174604 248018 174786 248254
rect 175022 248018 175204 248254
rect 174604 247934 175204 248018
rect 174604 247698 174786 247934
rect 175022 247698 175204 247934
rect 174604 212254 175204 247698
rect 174604 212018 174786 212254
rect 175022 212018 175204 212254
rect 174604 211934 175204 212018
rect 174604 211698 174786 211934
rect 175022 211698 175204 211934
rect 174604 176254 175204 211698
rect 174604 176018 174786 176254
rect 175022 176018 175204 176254
rect 174604 175934 175204 176018
rect 174604 175698 174786 175934
rect 175022 175698 175204 175934
rect 174604 140254 175204 175698
rect 174604 140018 174786 140254
rect 175022 140018 175204 140254
rect 174604 139934 175204 140018
rect 174604 139698 174786 139934
rect 175022 139698 175204 139934
rect 174604 104254 175204 139698
rect 174604 104018 174786 104254
rect 175022 104018 175204 104254
rect 174604 103934 175204 104018
rect 174604 103698 174786 103934
rect 175022 103698 175204 103934
rect 174604 68254 175204 103698
rect 174604 68018 174786 68254
rect 175022 68018 175204 68254
rect 174604 67934 175204 68018
rect 174604 67698 174786 67934
rect 175022 67698 175204 67934
rect 174604 32254 175204 67698
rect 174604 32018 174786 32254
rect 175022 32018 175204 32254
rect 174604 31934 175204 32018
rect 174604 31698 174786 31934
rect 175022 31698 175204 31934
rect 156604 -6222 156786 -5986
rect 157022 -6222 157204 -5986
rect 156604 -6306 157204 -6222
rect 156604 -6542 156786 -6306
rect 157022 -6542 157204 -6306
rect 156604 -7504 157204 -6542
rect 174604 -6926 175204 31698
rect 181804 291454 182404 326000
rect 181804 291218 181986 291454
rect 182222 291218 182404 291454
rect 181804 291134 182404 291218
rect 181804 290898 181986 291134
rect 182222 290898 182404 291134
rect 181804 255454 182404 290898
rect 181804 255218 181986 255454
rect 182222 255218 182404 255454
rect 181804 255134 182404 255218
rect 181804 254898 181986 255134
rect 182222 254898 182404 255134
rect 181804 219454 182404 254898
rect 181804 219218 181986 219454
rect 182222 219218 182404 219454
rect 181804 219134 182404 219218
rect 181804 218898 181986 219134
rect 182222 218898 182404 219134
rect 181804 183454 182404 218898
rect 181804 183218 181986 183454
rect 182222 183218 182404 183454
rect 181804 183134 182404 183218
rect 181804 182898 181986 183134
rect 182222 182898 182404 183134
rect 181804 147454 182404 182898
rect 181804 147218 181986 147454
rect 182222 147218 182404 147454
rect 181804 147134 182404 147218
rect 181804 146898 181986 147134
rect 182222 146898 182404 147134
rect 181804 111454 182404 146898
rect 181804 111218 181986 111454
rect 182222 111218 182404 111454
rect 181804 111134 182404 111218
rect 181804 110898 181986 111134
rect 182222 110898 182404 111134
rect 181804 75454 182404 110898
rect 181804 75218 181986 75454
rect 182222 75218 182404 75454
rect 181804 75134 182404 75218
rect 181804 74898 181986 75134
rect 182222 74898 182404 75134
rect 181804 39454 182404 74898
rect 181804 39218 181986 39454
rect 182222 39218 182404 39454
rect 181804 39134 182404 39218
rect 181804 38898 181986 39134
rect 182222 38898 182404 39134
rect 181804 3454 182404 38898
rect 181804 3218 181986 3454
rect 182222 3218 182404 3454
rect 181804 3134 182404 3218
rect 181804 2898 181986 3134
rect 182222 2898 182404 3134
rect 181804 -346 182404 2898
rect 181804 -582 181986 -346
rect 182222 -582 182404 -346
rect 181804 -666 182404 -582
rect 181804 -902 181986 -666
rect 182222 -902 182404 -666
rect 181804 -1864 182404 -902
rect 185404 295054 186004 326000
rect 185404 294818 185586 295054
rect 185822 294818 186004 295054
rect 185404 294734 186004 294818
rect 185404 294498 185586 294734
rect 185822 294498 186004 294734
rect 185404 259054 186004 294498
rect 185404 258818 185586 259054
rect 185822 258818 186004 259054
rect 185404 258734 186004 258818
rect 185404 258498 185586 258734
rect 185822 258498 186004 258734
rect 185404 223054 186004 258498
rect 185404 222818 185586 223054
rect 185822 222818 186004 223054
rect 185404 222734 186004 222818
rect 185404 222498 185586 222734
rect 185822 222498 186004 222734
rect 185404 187054 186004 222498
rect 185404 186818 185586 187054
rect 185822 186818 186004 187054
rect 185404 186734 186004 186818
rect 185404 186498 185586 186734
rect 185822 186498 186004 186734
rect 185404 151054 186004 186498
rect 185404 150818 185586 151054
rect 185822 150818 186004 151054
rect 185404 150734 186004 150818
rect 185404 150498 185586 150734
rect 185822 150498 186004 150734
rect 185404 115054 186004 150498
rect 185404 114818 185586 115054
rect 185822 114818 186004 115054
rect 185404 114734 186004 114818
rect 185404 114498 185586 114734
rect 185822 114498 186004 114734
rect 185404 79054 186004 114498
rect 185404 78818 185586 79054
rect 185822 78818 186004 79054
rect 185404 78734 186004 78818
rect 185404 78498 185586 78734
rect 185822 78498 186004 78734
rect 185404 43054 186004 78498
rect 185404 42818 185586 43054
rect 185822 42818 186004 43054
rect 185404 42734 186004 42818
rect 185404 42498 185586 42734
rect 185822 42498 186004 42734
rect 185404 7054 186004 42498
rect 185404 6818 185586 7054
rect 185822 6818 186004 7054
rect 185404 6734 186004 6818
rect 185404 6498 185586 6734
rect 185822 6498 186004 6734
rect 185404 -2226 186004 6498
rect 185404 -2462 185586 -2226
rect 185822 -2462 186004 -2226
rect 185404 -2546 186004 -2462
rect 185404 -2782 185586 -2546
rect 185822 -2782 186004 -2546
rect 185404 -3744 186004 -2782
rect 189004 298654 189604 326000
rect 189004 298418 189186 298654
rect 189422 298418 189604 298654
rect 189004 298334 189604 298418
rect 189004 298098 189186 298334
rect 189422 298098 189604 298334
rect 189004 262654 189604 298098
rect 189004 262418 189186 262654
rect 189422 262418 189604 262654
rect 189004 262334 189604 262418
rect 189004 262098 189186 262334
rect 189422 262098 189604 262334
rect 189004 226654 189604 262098
rect 189004 226418 189186 226654
rect 189422 226418 189604 226654
rect 189004 226334 189604 226418
rect 189004 226098 189186 226334
rect 189422 226098 189604 226334
rect 189004 190654 189604 226098
rect 189004 190418 189186 190654
rect 189422 190418 189604 190654
rect 189004 190334 189604 190418
rect 189004 190098 189186 190334
rect 189422 190098 189604 190334
rect 189004 154654 189604 190098
rect 189004 154418 189186 154654
rect 189422 154418 189604 154654
rect 189004 154334 189604 154418
rect 189004 154098 189186 154334
rect 189422 154098 189604 154334
rect 189004 118654 189604 154098
rect 189004 118418 189186 118654
rect 189422 118418 189604 118654
rect 189004 118334 189604 118418
rect 189004 118098 189186 118334
rect 189422 118098 189604 118334
rect 189004 82654 189604 118098
rect 189004 82418 189186 82654
rect 189422 82418 189604 82654
rect 189004 82334 189604 82418
rect 189004 82098 189186 82334
rect 189422 82098 189604 82334
rect 189004 46654 189604 82098
rect 189004 46418 189186 46654
rect 189422 46418 189604 46654
rect 189004 46334 189604 46418
rect 189004 46098 189186 46334
rect 189422 46098 189604 46334
rect 189004 10654 189604 46098
rect 189004 10418 189186 10654
rect 189422 10418 189604 10654
rect 189004 10334 189604 10418
rect 189004 10098 189186 10334
rect 189422 10098 189604 10334
rect 189004 -4106 189604 10098
rect 189004 -4342 189186 -4106
rect 189422 -4342 189604 -4106
rect 189004 -4426 189604 -4342
rect 189004 -4662 189186 -4426
rect 189422 -4662 189604 -4426
rect 189004 -5624 189604 -4662
rect 192604 302254 193204 326000
rect 192604 302018 192786 302254
rect 193022 302018 193204 302254
rect 192604 301934 193204 302018
rect 192604 301698 192786 301934
rect 193022 301698 193204 301934
rect 192604 266254 193204 301698
rect 192604 266018 192786 266254
rect 193022 266018 193204 266254
rect 192604 265934 193204 266018
rect 192604 265698 192786 265934
rect 193022 265698 193204 265934
rect 192604 230254 193204 265698
rect 192604 230018 192786 230254
rect 193022 230018 193204 230254
rect 192604 229934 193204 230018
rect 192604 229698 192786 229934
rect 193022 229698 193204 229934
rect 192604 194254 193204 229698
rect 192604 194018 192786 194254
rect 193022 194018 193204 194254
rect 192604 193934 193204 194018
rect 192604 193698 192786 193934
rect 193022 193698 193204 193934
rect 192604 158254 193204 193698
rect 192604 158018 192786 158254
rect 193022 158018 193204 158254
rect 192604 157934 193204 158018
rect 192604 157698 192786 157934
rect 193022 157698 193204 157934
rect 192604 122254 193204 157698
rect 192604 122018 192786 122254
rect 193022 122018 193204 122254
rect 192604 121934 193204 122018
rect 192604 121698 192786 121934
rect 193022 121698 193204 121934
rect 192604 86254 193204 121698
rect 192604 86018 192786 86254
rect 193022 86018 193204 86254
rect 192604 85934 193204 86018
rect 192604 85698 192786 85934
rect 193022 85698 193204 85934
rect 192604 50254 193204 85698
rect 192604 50018 192786 50254
rect 193022 50018 193204 50254
rect 192604 49934 193204 50018
rect 192604 49698 192786 49934
rect 193022 49698 193204 49934
rect 192604 14254 193204 49698
rect 192604 14018 192786 14254
rect 193022 14018 193204 14254
rect 192604 13934 193204 14018
rect 192604 13698 192786 13934
rect 193022 13698 193204 13934
rect 174604 -7162 174786 -6926
rect 175022 -7162 175204 -6926
rect 174604 -7246 175204 -7162
rect 174604 -7482 174786 -7246
rect 175022 -7482 175204 -7246
rect 174604 -7504 175204 -7482
rect 192604 -5986 193204 13698
rect 199804 309454 200404 326000
rect 199804 309218 199986 309454
rect 200222 309218 200404 309454
rect 199804 309134 200404 309218
rect 199804 308898 199986 309134
rect 200222 308898 200404 309134
rect 199804 273454 200404 308898
rect 199804 273218 199986 273454
rect 200222 273218 200404 273454
rect 199804 273134 200404 273218
rect 199804 272898 199986 273134
rect 200222 272898 200404 273134
rect 199804 237454 200404 272898
rect 199804 237218 199986 237454
rect 200222 237218 200404 237454
rect 199804 237134 200404 237218
rect 199804 236898 199986 237134
rect 200222 236898 200404 237134
rect 199804 201454 200404 236898
rect 199804 201218 199986 201454
rect 200222 201218 200404 201454
rect 199804 201134 200404 201218
rect 199804 200898 199986 201134
rect 200222 200898 200404 201134
rect 199804 165454 200404 200898
rect 199804 165218 199986 165454
rect 200222 165218 200404 165454
rect 199804 165134 200404 165218
rect 199804 164898 199986 165134
rect 200222 164898 200404 165134
rect 199804 129454 200404 164898
rect 199804 129218 199986 129454
rect 200222 129218 200404 129454
rect 199804 129134 200404 129218
rect 199804 128898 199986 129134
rect 200222 128898 200404 129134
rect 199804 93454 200404 128898
rect 199804 93218 199986 93454
rect 200222 93218 200404 93454
rect 199804 93134 200404 93218
rect 199804 92898 199986 93134
rect 200222 92898 200404 93134
rect 199804 57454 200404 92898
rect 199804 57218 199986 57454
rect 200222 57218 200404 57454
rect 199804 57134 200404 57218
rect 199804 56898 199986 57134
rect 200222 56898 200404 57134
rect 199804 21454 200404 56898
rect 199804 21218 199986 21454
rect 200222 21218 200404 21454
rect 199804 21134 200404 21218
rect 199804 20898 199986 21134
rect 200222 20898 200404 21134
rect 199804 -1286 200404 20898
rect 199804 -1522 199986 -1286
rect 200222 -1522 200404 -1286
rect 199804 -1606 200404 -1522
rect 199804 -1842 199986 -1606
rect 200222 -1842 200404 -1606
rect 199804 -1864 200404 -1842
rect 203404 313054 204004 326000
rect 203404 312818 203586 313054
rect 203822 312818 204004 313054
rect 203404 312734 204004 312818
rect 203404 312498 203586 312734
rect 203822 312498 204004 312734
rect 203404 277054 204004 312498
rect 203404 276818 203586 277054
rect 203822 276818 204004 277054
rect 203404 276734 204004 276818
rect 203404 276498 203586 276734
rect 203822 276498 204004 276734
rect 203404 241054 204004 276498
rect 203404 240818 203586 241054
rect 203822 240818 204004 241054
rect 203404 240734 204004 240818
rect 203404 240498 203586 240734
rect 203822 240498 204004 240734
rect 203404 205054 204004 240498
rect 203404 204818 203586 205054
rect 203822 204818 204004 205054
rect 203404 204734 204004 204818
rect 203404 204498 203586 204734
rect 203822 204498 204004 204734
rect 203404 169054 204004 204498
rect 203404 168818 203586 169054
rect 203822 168818 204004 169054
rect 203404 168734 204004 168818
rect 203404 168498 203586 168734
rect 203822 168498 204004 168734
rect 203404 133054 204004 168498
rect 203404 132818 203586 133054
rect 203822 132818 204004 133054
rect 203404 132734 204004 132818
rect 203404 132498 203586 132734
rect 203822 132498 204004 132734
rect 203404 97054 204004 132498
rect 203404 96818 203586 97054
rect 203822 96818 204004 97054
rect 203404 96734 204004 96818
rect 203404 96498 203586 96734
rect 203822 96498 204004 96734
rect 203404 61054 204004 96498
rect 203404 60818 203586 61054
rect 203822 60818 204004 61054
rect 203404 60734 204004 60818
rect 203404 60498 203586 60734
rect 203822 60498 204004 60734
rect 203404 25054 204004 60498
rect 203404 24818 203586 25054
rect 203822 24818 204004 25054
rect 203404 24734 204004 24818
rect 203404 24498 203586 24734
rect 203822 24498 204004 24734
rect 203404 -3166 204004 24498
rect 203404 -3402 203586 -3166
rect 203822 -3402 204004 -3166
rect 203404 -3486 204004 -3402
rect 203404 -3722 203586 -3486
rect 203822 -3722 204004 -3486
rect 203404 -3744 204004 -3722
rect 207004 316654 207604 326000
rect 207004 316418 207186 316654
rect 207422 316418 207604 316654
rect 207004 316334 207604 316418
rect 207004 316098 207186 316334
rect 207422 316098 207604 316334
rect 207004 280654 207604 316098
rect 207004 280418 207186 280654
rect 207422 280418 207604 280654
rect 207004 280334 207604 280418
rect 207004 280098 207186 280334
rect 207422 280098 207604 280334
rect 207004 244654 207604 280098
rect 207004 244418 207186 244654
rect 207422 244418 207604 244654
rect 207004 244334 207604 244418
rect 207004 244098 207186 244334
rect 207422 244098 207604 244334
rect 207004 208654 207604 244098
rect 207004 208418 207186 208654
rect 207422 208418 207604 208654
rect 207004 208334 207604 208418
rect 207004 208098 207186 208334
rect 207422 208098 207604 208334
rect 207004 172654 207604 208098
rect 207004 172418 207186 172654
rect 207422 172418 207604 172654
rect 207004 172334 207604 172418
rect 207004 172098 207186 172334
rect 207422 172098 207604 172334
rect 207004 136654 207604 172098
rect 207004 136418 207186 136654
rect 207422 136418 207604 136654
rect 207004 136334 207604 136418
rect 207004 136098 207186 136334
rect 207422 136098 207604 136334
rect 207004 100654 207604 136098
rect 207004 100418 207186 100654
rect 207422 100418 207604 100654
rect 207004 100334 207604 100418
rect 207004 100098 207186 100334
rect 207422 100098 207604 100334
rect 207004 64654 207604 100098
rect 207004 64418 207186 64654
rect 207422 64418 207604 64654
rect 207004 64334 207604 64418
rect 207004 64098 207186 64334
rect 207422 64098 207604 64334
rect 207004 28654 207604 64098
rect 207004 28418 207186 28654
rect 207422 28418 207604 28654
rect 207004 28334 207604 28418
rect 207004 28098 207186 28334
rect 207422 28098 207604 28334
rect 207004 -5046 207604 28098
rect 207004 -5282 207186 -5046
rect 207422 -5282 207604 -5046
rect 207004 -5366 207604 -5282
rect 207004 -5602 207186 -5366
rect 207422 -5602 207604 -5366
rect 207004 -5624 207604 -5602
rect 210604 320254 211204 326000
rect 210604 320018 210786 320254
rect 211022 320018 211204 320254
rect 210604 319934 211204 320018
rect 210604 319698 210786 319934
rect 211022 319698 211204 319934
rect 210604 284254 211204 319698
rect 210604 284018 210786 284254
rect 211022 284018 211204 284254
rect 210604 283934 211204 284018
rect 210604 283698 210786 283934
rect 211022 283698 211204 283934
rect 210604 248254 211204 283698
rect 210604 248018 210786 248254
rect 211022 248018 211204 248254
rect 210604 247934 211204 248018
rect 210604 247698 210786 247934
rect 211022 247698 211204 247934
rect 210604 212254 211204 247698
rect 210604 212018 210786 212254
rect 211022 212018 211204 212254
rect 210604 211934 211204 212018
rect 210604 211698 210786 211934
rect 211022 211698 211204 211934
rect 210604 176254 211204 211698
rect 210604 176018 210786 176254
rect 211022 176018 211204 176254
rect 210604 175934 211204 176018
rect 210604 175698 210786 175934
rect 211022 175698 211204 175934
rect 210604 140254 211204 175698
rect 210604 140018 210786 140254
rect 211022 140018 211204 140254
rect 210604 139934 211204 140018
rect 210604 139698 210786 139934
rect 211022 139698 211204 139934
rect 210604 104254 211204 139698
rect 210604 104018 210786 104254
rect 211022 104018 211204 104254
rect 210604 103934 211204 104018
rect 210604 103698 210786 103934
rect 211022 103698 211204 103934
rect 210604 68254 211204 103698
rect 210604 68018 210786 68254
rect 211022 68018 211204 68254
rect 210604 67934 211204 68018
rect 210604 67698 210786 67934
rect 211022 67698 211204 67934
rect 210604 32254 211204 67698
rect 210604 32018 210786 32254
rect 211022 32018 211204 32254
rect 210604 31934 211204 32018
rect 210604 31698 210786 31934
rect 211022 31698 211204 31934
rect 192604 -6222 192786 -5986
rect 193022 -6222 193204 -5986
rect 192604 -6306 193204 -6222
rect 192604 -6542 192786 -6306
rect 193022 -6542 193204 -6306
rect 192604 -7504 193204 -6542
rect 210604 -6926 211204 31698
rect 217804 291454 218404 326000
rect 217804 291218 217986 291454
rect 218222 291218 218404 291454
rect 217804 291134 218404 291218
rect 217804 290898 217986 291134
rect 218222 290898 218404 291134
rect 217804 255454 218404 290898
rect 217804 255218 217986 255454
rect 218222 255218 218404 255454
rect 217804 255134 218404 255218
rect 217804 254898 217986 255134
rect 218222 254898 218404 255134
rect 217804 219454 218404 254898
rect 217804 219218 217986 219454
rect 218222 219218 218404 219454
rect 217804 219134 218404 219218
rect 217804 218898 217986 219134
rect 218222 218898 218404 219134
rect 217804 183454 218404 218898
rect 217804 183218 217986 183454
rect 218222 183218 218404 183454
rect 217804 183134 218404 183218
rect 217804 182898 217986 183134
rect 218222 182898 218404 183134
rect 217804 147454 218404 182898
rect 217804 147218 217986 147454
rect 218222 147218 218404 147454
rect 217804 147134 218404 147218
rect 217804 146898 217986 147134
rect 218222 146898 218404 147134
rect 217804 111454 218404 146898
rect 217804 111218 217986 111454
rect 218222 111218 218404 111454
rect 217804 111134 218404 111218
rect 217804 110898 217986 111134
rect 218222 110898 218404 111134
rect 217804 75454 218404 110898
rect 217804 75218 217986 75454
rect 218222 75218 218404 75454
rect 217804 75134 218404 75218
rect 217804 74898 217986 75134
rect 218222 74898 218404 75134
rect 217804 39454 218404 74898
rect 217804 39218 217986 39454
rect 218222 39218 218404 39454
rect 217804 39134 218404 39218
rect 217804 38898 217986 39134
rect 218222 38898 218404 39134
rect 217804 3454 218404 38898
rect 217804 3218 217986 3454
rect 218222 3218 218404 3454
rect 217804 3134 218404 3218
rect 217804 2898 217986 3134
rect 218222 2898 218404 3134
rect 217804 -346 218404 2898
rect 217804 -582 217986 -346
rect 218222 -582 218404 -346
rect 217804 -666 218404 -582
rect 217804 -902 217986 -666
rect 218222 -902 218404 -666
rect 217804 -1864 218404 -902
rect 221404 295054 222004 326000
rect 221404 294818 221586 295054
rect 221822 294818 222004 295054
rect 221404 294734 222004 294818
rect 221404 294498 221586 294734
rect 221822 294498 222004 294734
rect 221404 259054 222004 294498
rect 221404 258818 221586 259054
rect 221822 258818 222004 259054
rect 221404 258734 222004 258818
rect 221404 258498 221586 258734
rect 221822 258498 222004 258734
rect 221404 223054 222004 258498
rect 221404 222818 221586 223054
rect 221822 222818 222004 223054
rect 221404 222734 222004 222818
rect 221404 222498 221586 222734
rect 221822 222498 222004 222734
rect 221404 187054 222004 222498
rect 221404 186818 221586 187054
rect 221822 186818 222004 187054
rect 221404 186734 222004 186818
rect 221404 186498 221586 186734
rect 221822 186498 222004 186734
rect 221404 151054 222004 186498
rect 221404 150818 221586 151054
rect 221822 150818 222004 151054
rect 221404 150734 222004 150818
rect 221404 150498 221586 150734
rect 221822 150498 222004 150734
rect 221404 115054 222004 150498
rect 221404 114818 221586 115054
rect 221822 114818 222004 115054
rect 221404 114734 222004 114818
rect 221404 114498 221586 114734
rect 221822 114498 222004 114734
rect 221404 79054 222004 114498
rect 221404 78818 221586 79054
rect 221822 78818 222004 79054
rect 221404 78734 222004 78818
rect 221404 78498 221586 78734
rect 221822 78498 222004 78734
rect 221404 43054 222004 78498
rect 221404 42818 221586 43054
rect 221822 42818 222004 43054
rect 221404 42734 222004 42818
rect 221404 42498 221586 42734
rect 221822 42498 222004 42734
rect 221404 7054 222004 42498
rect 221404 6818 221586 7054
rect 221822 6818 222004 7054
rect 221404 6734 222004 6818
rect 221404 6498 221586 6734
rect 221822 6498 222004 6734
rect 221404 -2226 222004 6498
rect 221404 -2462 221586 -2226
rect 221822 -2462 222004 -2226
rect 221404 -2546 222004 -2462
rect 221404 -2782 221586 -2546
rect 221822 -2782 222004 -2546
rect 221404 -3744 222004 -2782
rect 225004 298654 225604 326000
rect 225004 298418 225186 298654
rect 225422 298418 225604 298654
rect 225004 298334 225604 298418
rect 225004 298098 225186 298334
rect 225422 298098 225604 298334
rect 225004 262654 225604 298098
rect 225004 262418 225186 262654
rect 225422 262418 225604 262654
rect 225004 262334 225604 262418
rect 225004 262098 225186 262334
rect 225422 262098 225604 262334
rect 225004 226654 225604 262098
rect 225004 226418 225186 226654
rect 225422 226418 225604 226654
rect 225004 226334 225604 226418
rect 225004 226098 225186 226334
rect 225422 226098 225604 226334
rect 225004 190654 225604 226098
rect 225004 190418 225186 190654
rect 225422 190418 225604 190654
rect 225004 190334 225604 190418
rect 225004 190098 225186 190334
rect 225422 190098 225604 190334
rect 225004 154654 225604 190098
rect 225004 154418 225186 154654
rect 225422 154418 225604 154654
rect 225004 154334 225604 154418
rect 225004 154098 225186 154334
rect 225422 154098 225604 154334
rect 225004 118654 225604 154098
rect 225004 118418 225186 118654
rect 225422 118418 225604 118654
rect 225004 118334 225604 118418
rect 225004 118098 225186 118334
rect 225422 118098 225604 118334
rect 225004 82654 225604 118098
rect 225004 82418 225186 82654
rect 225422 82418 225604 82654
rect 225004 82334 225604 82418
rect 225004 82098 225186 82334
rect 225422 82098 225604 82334
rect 225004 46654 225604 82098
rect 225004 46418 225186 46654
rect 225422 46418 225604 46654
rect 225004 46334 225604 46418
rect 225004 46098 225186 46334
rect 225422 46098 225604 46334
rect 225004 10654 225604 46098
rect 225004 10418 225186 10654
rect 225422 10418 225604 10654
rect 225004 10334 225604 10418
rect 225004 10098 225186 10334
rect 225422 10098 225604 10334
rect 225004 -4106 225604 10098
rect 225004 -4342 225186 -4106
rect 225422 -4342 225604 -4106
rect 225004 -4426 225604 -4342
rect 225004 -4662 225186 -4426
rect 225422 -4662 225604 -4426
rect 225004 -5624 225604 -4662
rect 228604 302254 229204 326000
rect 228604 302018 228786 302254
rect 229022 302018 229204 302254
rect 228604 301934 229204 302018
rect 228604 301698 228786 301934
rect 229022 301698 229204 301934
rect 228604 266254 229204 301698
rect 228604 266018 228786 266254
rect 229022 266018 229204 266254
rect 228604 265934 229204 266018
rect 228604 265698 228786 265934
rect 229022 265698 229204 265934
rect 228604 230254 229204 265698
rect 228604 230018 228786 230254
rect 229022 230018 229204 230254
rect 228604 229934 229204 230018
rect 228604 229698 228786 229934
rect 229022 229698 229204 229934
rect 228604 194254 229204 229698
rect 228604 194018 228786 194254
rect 229022 194018 229204 194254
rect 228604 193934 229204 194018
rect 228604 193698 228786 193934
rect 229022 193698 229204 193934
rect 228604 158254 229204 193698
rect 228604 158018 228786 158254
rect 229022 158018 229204 158254
rect 228604 157934 229204 158018
rect 228604 157698 228786 157934
rect 229022 157698 229204 157934
rect 228604 122254 229204 157698
rect 228604 122018 228786 122254
rect 229022 122018 229204 122254
rect 228604 121934 229204 122018
rect 228604 121698 228786 121934
rect 229022 121698 229204 121934
rect 228604 86254 229204 121698
rect 228604 86018 228786 86254
rect 229022 86018 229204 86254
rect 228604 85934 229204 86018
rect 228604 85698 228786 85934
rect 229022 85698 229204 85934
rect 228604 50254 229204 85698
rect 228604 50018 228786 50254
rect 229022 50018 229204 50254
rect 228604 49934 229204 50018
rect 228604 49698 228786 49934
rect 229022 49698 229204 49934
rect 228604 14254 229204 49698
rect 228604 14018 228786 14254
rect 229022 14018 229204 14254
rect 228604 13934 229204 14018
rect 228604 13698 228786 13934
rect 229022 13698 229204 13934
rect 210604 -7162 210786 -6926
rect 211022 -7162 211204 -6926
rect 210604 -7246 211204 -7162
rect 210604 -7482 210786 -7246
rect 211022 -7482 211204 -7246
rect 210604 -7504 211204 -7482
rect 228604 -5986 229204 13698
rect 235804 309454 236404 326000
rect 235804 309218 235986 309454
rect 236222 309218 236404 309454
rect 235804 309134 236404 309218
rect 235804 308898 235986 309134
rect 236222 308898 236404 309134
rect 235804 273454 236404 308898
rect 235804 273218 235986 273454
rect 236222 273218 236404 273454
rect 235804 273134 236404 273218
rect 235804 272898 235986 273134
rect 236222 272898 236404 273134
rect 235804 237454 236404 272898
rect 235804 237218 235986 237454
rect 236222 237218 236404 237454
rect 235804 237134 236404 237218
rect 235804 236898 235986 237134
rect 236222 236898 236404 237134
rect 235804 201454 236404 236898
rect 235804 201218 235986 201454
rect 236222 201218 236404 201454
rect 235804 201134 236404 201218
rect 235804 200898 235986 201134
rect 236222 200898 236404 201134
rect 235804 165454 236404 200898
rect 235804 165218 235986 165454
rect 236222 165218 236404 165454
rect 235804 165134 236404 165218
rect 235804 164898 235986 165134
rect 236222 164898 236404 165134
rect 235804 129454 236404 164898
rect 235804 129218 235986 129454
rect 236222 129218 236404 129454
rect 235804 129134 236404 129218
rect 235804 128898 235986 129134
rect 236222 128898 236404 129134
rect 235804 93454 236404 128898
rect 235804 93218 235986 93454
rect 236222 93218 236404 93454
rect 235804 93134 236404 93218
rect 235804 92898 235986 93134
rect 236222 92898 236404 93134
rect 235804 57454 236404 92898
rect 235804 57218 235986 57454
rect 236222 57218 236404 57454
rect 235804 57134 236404 57218
rect 235804 56898 235986 57134
rect 236222 56898 236404 57134
rect 235804 21454 236404 56898
rect 235804 21218 235986 21454
rect 236222 21218 236404 21454
rect 235804 21134 236404 21218
rect 235804 20898 235986 21134
rect 236222 20898 236404 21134
rect 235804 -1286 236404 20898
rect 235804 -1522 235986 -1286
rect 236222 -1522 236404 -1286
rect 235804 -1606 236404 -1522
rect 235804 -1842 235986 -1606
rect 236222 -1842 236404 -1606
rect 235804 -1864 236404 -1842
rect 239404 313054 240004 326000
rect 239404 312818 239586 313054
rect 239822 312818 240004 313054
rect 239404 312734 240004 312818
rect 239404 312498 239586 312734
rect 239822 312498 240004 312734
rect 239404 277054 240004 312498
rect 239404 276818 239586 277054
rect 239822 276818 240004 277054
rect 239404 276734 240004 276818
rect 239404 276498 239586 276734
rect 239822 276498 240004 276734
rect 239404 241054 240004 276498
rect 239404 240818 239586 241054
rect 239822 240818 240004 241054
rect 239404 240734 240004 240818
rect 239404 240498 239586 240734
rect 239822 240498 240004 240734
rect 239404 205054 240004 240498
rect 239404 204818 239586 205054
rect 239822 204818 240004 205054
rect 239404 204734 240004 204818
rect 239404 204498 239586 204734
rect 239822 204498 240004 204734
rect 239404 169054 240004 204498
rect 239404 168818 239586 169054
rect 239822 168818 240004 169054
rect 239404 168734 240004 168818
rect 239404 168498 239586 168734
rect 239822 168498 240004 168734
rect 239404 133054 240004 168498
rect 239404 132818 239586 133054
rect 239822 132818 240004 133054
rect 239404 132734 240004 132818
rect 239404 132498 239586 132734
rect 239822 132498 240004 132734
rect 239404 97054 240004 132498
rect 239404 96818 239586 97054
rect 239822 96818 240004 97054
rect 239404 96734 240004 96818
rect 239404 96498 239586 96734
rect 239822 96498 240004 96734
rect 239404 61054 240004 96498
rect 239404 60818 239586 61054
rect 239822 60818 240004 61054
rect 239404 60734 240004 60818
rect 239404 60498 239586 60734
rect 239822 60498 240004 60734
rect 239404 25054 240004 60498
rect 239404 24818 239586 25054
rect 239822 24818 240004 25054
rect 239404 24734 240004 24818
rect 239404 24498 239586 24734
rect 239822 24498 240004 24734
rect 239404 -3166 240004 24498
rect 239404 -3402 239586 -3166
rect 239822 -3402 240004 -3166
rect 239404 -3486 240004 -3402
rect 239404 -3722 239586 -3486
rect 239822 -3722 240004 -3486
rect 239404 -3744 240004 -3722
rect 243004 316654 243604 326000
rect 243004 316418 243186 316654
rect 243422 316418 243604 316654
rect 243004 316334 243604 316418
rect 243004 316098 243186 316334
rect 243422 316098 243604 316334
rect 243004 280654 243604 316098
rect 243004 280418 243186 280654
rect 243422 280418 243604 280654
rect 243004 280334 243604 280418
rect 243004 280098 243186 280334
rect 243422 280098 243604 280334
rect 243004 244654 243604 280098
rect 243004 244418 243186 244654
rect 243422 244418 243604 244654
rect 243004 244334 243604 244418
rect 243004 244098 243186 244334
rect 243422 244098 243604 244334
rect 243004 208654 243604 244098
rect 243004 208418 243186 208654
rect 243422 208418 243604 208654
rect 243004 208334 243604 208418
rect 243004 208098 243186 208334
rect 243422 208098 243604 208334
rect 243004 172654 243604 208098
rect 243004 172418 243186 172654
rect 243422 172418 243604 172654
rect 243004 172334 243604 172418
rect 243004 172098 243186 172334
rect 243422 172098 243604 172334
rect 243004 136654 243604 172098
rect 243004 136418 243186 136654
rect 243422 136418 243604 136654
rect 243004 136334 243604 136418
rect 243004 136098 243186 136334
rect 243422 136098 243604 136334
rect 243004 100654 243604 136098
rect 243004 100418 243186 100654
rect 243422 100418 243604 100654
rect 243004 100334 243604 100418
rect 243004 100098 243186 100334
rect 243422 100098 243604 100334
rect 243004 64654 243604 100098
rect 243004 64418 243186 64654
rect 243422 64418 243604 64654
rect 243004 64334 243604 64418
rect 243004 64098 243186 64334
rect 243422 64098 243604 64334
rect 243004 28654 243604 64098
rect 243004 28418 243186 28654
rect 243422 28418 243604 28654
rect 243004 28334 243604 28418
rect 243004 28098 243186 28334
rect 243422 28098 243604 28334
rect 243004 -5046 243604 28098
rect 243004 -5282 243186 -5046
rect 243422 -5282 243604 -5046
rect 243004 -5366 243604 -5282
rect 243004 -5602 243186 -5366
rect 243422 -5602 243604 -5366
rect 243004 -5624 243604 -5602
rect 246604 320254 247204 326000
rect 246604 320018 246786 320254
rect 247022 320018 247204 320254
rect 246604 319934 247204 320018
rect 246604 319698 246786 319934
rect 247022 319698 247204 319934
rect 246604 284254 247204 319698
rect 246604 284018 246786 284254
rect 247022 284018 247204 284254
rect 246604 283934 247204 284018
rect 246604 283698 246786 283934
rect 247022 283698 247204 283934
rect 246604 248254 247204 283698
rect 246604 248018 246786 248254
rect 247022 248018 247204 248254
rect 246604 247934 247204 248018
rect 246604 247698 246786 247934
rect 247022 247698 247204 247934
rect 246604 212254 247204 247698
rect 246604 212018 246786 212254
rect 247022 212018 247204 212254
rect 246604 211934 247204 212018
rect 246604 211698 246786 211934
rect 247022 211698 247204 211934
rect 246604 176254 247204 211698
rect 246604 176018 246786 176254
rect 247022 176018 247204 176254
rect 246604 175934 247204 176018
rect 246604 175698 246786 175934
rect 247022 175698 247204 175934
rect 246604 140254 247204 175698
rect 246604 140018 246786 140254
rect 247022 140018 247204 140254
rect 246604 139934 247204 140018
rect 246604 139698 246786 139934
rect 247022 139698 247204 139934
rect 246604 104254 247204 139698
rect 246604 104018 246786 104254
rect 247022 104018 247204 104254
rect 246604 103934 247204 104018
rect 246604 103698 246786 103934
rect 247022 103698 247204 103934
rect 246604 68254 247204 103698
rect 246604 68018 246786 68254
rect 247022 68018 247204 68254
rect 246604 67934 247204 68018
rect 246604 67698 246786 67934
rect 247022 67698 247204 67934
rect 246604 32254 247204 67698
rect 246604 32018 246786 32254
rect 247022 32018 247204 32254
rect 246604 31934 247204 32018
rect 246604 31698 246786 31934
rect 247022 31698 247204 31934
rect 228604 -6222 228786 -5986
rect 229022 -6222 229204 -5986
rect 228604 -6306 229204 -6222
rect 228604 -6542 228786 -6306
rect 229022 -6542 229204 -6306
rect 228604 -7504 229204 -6542
rect 246604 -6926 247204 31698
rect 253804 291454 254404 326000
rect 253804 291218 253986 291454
rect 254222 291218 254404 291454
rect 253804 291134 254404 291218
rect 253804 290898 253986 291134
rect 254222 290898 254404 291134
rect 253804 255454 254404 290898
rect 253804 255218 253986 255454
rect 254222 255218 254404 255454
rect 253804 255134 254404 255218
rect 253804 254898 253986 255134
rect 254222 254898 254404 255134
rect 253804 219454 254404 254898
rect 253804 219218 253986 219454
rect 254222 219218 254404 219454
rect 253804 219134 254404 219218
rect 253804 218898 253986 219134
rect 254222 218898 254404 219134
rect 253804 183454 254404 218898
rect 253804 183218 253986 183454
rect 254222 183218 254404 183454
rect 253804 183134 254404 183218
rect 253804 182898 253986 183134
rect 254222 182898 254404 183134
rect 253804 147454 254404 182898
rect 253804 147218 253986 147454
rect 254222 147218 254404 147454
rect 253804 147134 254404 147218
rect 253804 146898 253986 147134
rect 254222 146898 254404 147134
rect 253804 111454 254404 146898
rect 253804 111218 253986 111454
rect 254222 111218 254404 111454
rect 253804 111134 254404 111218
rect 253804 110898 253986 111134
rect 254222 110898 254404 111134
rect 253804 75454 254404 110898
rect 253804 75218 253986 75454
rect 254222 75218 254404 75454
rect 253804 75134 254404 75218
rect 253804 74898 253986 75134
rect 254222 74898 254404 75134
rect 253804 39454 254404 74898
rect 253804 39218 253986 39454
rect 254222 39218 254404 39454
rect 253804 39134 254404 39218
rect 253804 38898 253986 39134
rect 254222 38898 254404 39134
rect 253804 3454 254404 38898
rect 253804 3218 253986 3454
rect 254222 3218 254404 3454
rect 253804 3134 254404 3218
rect 253804 2898 253986 3134
rect 254222 2898 254404 3134
rect 253804 -346 254404 2898
rect 253804 -582 253986 -346
rect 254222 -582 254404 -346
rect 253804 -666 254404 -582
rect 253804 -902 253986 -666
rect 254222 -902 254404 -666
rect 253804 -1864 254404 -902
rect 257404 295054 258004 326000
rect 257404 294818 257586 295054
rect 257822 294818 258004 295054
rect 257404 294734 258004 294818
rect 257404 294498 257586 294734
rect 257822 294498 258004 294734
rect 257404 259054 258004 294498
rect 257404 258818 257586 259054
rect 257822 258818 258004 259054
rect 257404 258734 258004 258818
rect 257404 258498 257586 258734
rect 257822 258498 258004 258734
rect 257404 223054 258004 258498
rect 257404 222818 257586 223054
rect 257822 222818 258004 223054
rect 257404 222734 258004 222818
rect 257404 222498 257586 222734
rect 257822 222498 258004 222734
rect 257404 187054 258004 222498
rect 257404 186818 257586 187054
rect 257822 186818 258004 187054
rect 257404 186734 258004 186818
rect 257404 186498 257586 186734
rect 257822 186498 258004 186734
rect 257404 151054 258004 186498
rect 257404 150818 257586 151054
rect 257822 150818 258004 151054
rect 257404 150734 258004 150818
rect 257404 150498 257586 150734
rect 257822 150498 258004 150734
rect 257404 115054 258004 150498
rect 257404 114818 257586 115054
rect 257822 114818 258004 115054
rect 257404 114734 258004 114818
rect 257404 114498 257586 114734
rect 257822 114498 258004 114734
rect 257404 79054 258004 114498
rect 257404 78818 257586 79054
rect 257822 78818 258004 79054
rect 257404 78734 258004 78818
rect 257404 78498 257586 78734
rect 257822 78498 258004 78734
rect 257404 43054 258004 78498
rect 257404 42818 257586 43054
rect 257822 42818 258004 43054
rect 257404 42734 258004 42818
rect 257404 42498 257586 42734
rect 257822 42498 258004 42734
rect 257404 7054 258004 42498
rect 257404 6818 257586 7054
rect 257822 6818 258004 7054
rect 257404 6734 258004 6818
rect 257404 6498 257586 6734
rect 257822 6498 258004 6734
rect 257404 -2226 258004 6498
rect 257404 -2462 257586 -2226
rect 257822 -2462 258004 -2226
rect 257404 -2546 258004 -2462
rect 257404 -2782 257586 -2546
rect 257822 -2782 258004 -2546
rect 257404 -3744 258004 -2782
rect 261004 298654 261604 326000
rect 261004 298418 261186 298654
rect 261422 298418 261604 298654
rect 261004 298334 261604 298418
rect 261004 298098 261186 298334
rect 261422 298098 261604 298334
rect 261004 262654 261604 298098
rect 261004 262418 261186 262654
rect 261422 262418 261604 262654
rect 261004 262334 261604 262418
rect 261004 262098 261186 262334
rect 261422 262098 261604 262334
rect 261004 226654 261604 262098
rect 261004 226418 261186 226654
rect 261422 226418 261604 226654
rect 261004 226334 261604 226418
rect 261004 226098 261186 226334
rect 261422 226098 261604 226334
rect 261004 190654 261604 226098
rect 261004 190418 261186 190654
rect 261422 190418 261604 190654
rect 261004 190334 261604 190418
rect 261004 190098 261186 190334
rect 261422 190098 261604 190334
rect 261004 154654 261604 190098
rect 261004 154418 261186 154654
rect 261422 154418 261604 154654
rect 261004 154334 261604 154418
rect 261004 154098 261186 154334
rect 261422 154098 261604 154334
rect 261004 118654 261604 154098
rect 261004 118418 261186 118654
rect 261422 118418 261604 118654
rect 261004 118334 261604 118418
rect 261004 118098 261186 118334
rect 261422 118098 261604 118334
rect 261004 82654 261604 118098
rect 261004 82418 261186 82654
rect 261422 82418 261604 82654
rect 261004 82334 261604 82418
rect 261004 82098 261186 82334
rect 261422 82098 261604 82334
rect 261004 46654 261604 82098
rect 261004 46418 261186 46654
rect 261422 46418 261604 46654
rect 261004 46334 261604 46418
rect 261004 46098 261186 46334
rect 261422 46098 261604 46334
rect 261004 10654 261604 46098
rect 261004 10418 261186 10654
rect 261422 10418 261604 10654
rect 261004 10334 261604 10418
rect 261004 10098 261186 10334
rect 261422 10098 261604 10334
rect 261004 -4106 261604 10098
rect 261004 -4342 261186 -4106
rect 261422 -4342 261604 -4106
rect 261004 -4426 261604 -4342
rect 261004 -4662 261186 -4426
rect 261422 -4662 261604 -4426
rect 261004 -5624 261604 -4662
rect 264604 302254 265204 326000
rect 264604 302018 264786 302254
rect 265022 302018 265204 302254
rect 264604 301934 265204 302018
rect 264604 301698 264786 301934
rect 265022 301698 265204 301934
rect 264604 266254 265204 301698
rect 264604 266018 264786 266254
rect 265022 266018 265204 266254
rect 264604 265934 265204 266018
rect 264604 265698 264786 265934
rect 265022 265698 265204 265934
rect 264604 230254 265204 265698
rect 264604 230018 264786 230254
rect 265022 230018 265204 230254
rect 264604 229934 265204 230018
rect 264604 229698 264786 229934
rect 265022 229698 265204 229934
rect 264604 194254 265204 229698
rect 264604 194018 264786 194254
rect 265022 194018 265204 194254
rect 264604 193934 265204 194018
rect 264604 193698 264786 193934
rect 265022 193698 265204 193934
rect 264604 158254 265204 193698
rect 264604 158018 264786 158254
rect 265022 158018 265204 158254
rect 264604 157934 265204 158018
rect 264604 157698 264786 157934
rect 265022 157698 265204 157934
rect 264604 122254 265204 157698
rect 264604 122018 264786 122254
rect 265022 122018 265204 122254
rect 264604 121934 265204 122018
rect 264604 121698 264786 121934
rect 265022 121698 265204 121934
rect 264604 86254 265204 121698
rect 264604 86018 264786 86254
rect 265022 86018 265204 86254
rect 264604 85934 265204 86018
rect 264604 85698 264786 85934
rect 265022 85698 265204 85934
rect 264604 50254 265204 85698
rect 264604 50018 264786 50254
rect 265022 50018 265204 50254
rect 264604 49934 265204 50018
rect 264604 49698 264786 49934
rect 265022 49698 265204 49934
rect 264604 14254 265204 49698
rect 264604 14018 264786 14254
rect 265022 14018 265204 14254
rect 264604 13934 265204 14018
rect 264604 13698 264786 13934
rect 265022 13698 265204 13934
rect 246604 -7162 246786 -6926
rect 247022 -7162 247204 -6926
rect 246604 -7246 247204 -7162
rect 246604 -7482 246786 -7246
rect 247022 -7482 247204 -7246
rect 246604 -7504 247204 -7482
rect 264604 -5986 265204 13698
rect 271804 309454 272404 326000
rect 271804 309218 271986 309454
rect 272222 309218 272404 309454
rect 271804 309134 272404 309218
rect 271804 308898 271986 309134
rect 272222 308898 272404 309134
rect 271804 273454 272404 308898
rect 271804 273218 271986 273454
rect 272222 273218 272404 273454
rect 271804 273134 272404 273218
rect 271804 272898 271986 273134
rect 272222 272898 272404 273134
rect 271804 237454 272404 272898
rect 271804 237218 271986 237454
rect 272222 237218 272404 237454
rect 271804 237134 272404 237218
rect 271804 236898 271986 237134
rect 272222 236898 272404 237134
rect 271804 201454 272404 236898
rect 271804 201218 271986 201454
rect 272222 201218 272404 201454
rect 271804 201134 272404 201218
rect 271804 200898 271986 201134
rect 272222 200898 272404 201134
rect 271804 165454 272404 200898
rect 271804 165218 271986 165454
rect 272222 165218 272404 165454
rect 271804 165134 272404 165218
rect 271804 164898 271986 165134
rect 272222 164898 272404 165134
rect 271804 129454 272404 164898
rect 271804 129218 271986 129454
rect 272222 129218 272404 129454
rect 271804 129134 272404 129218
rect 271804 128898 271986 129134
rect 272222 128898 272404 129134
rect 271804 93454 272404 128898
rect 271804 93218 271986 93454
rect 272222 93218 272404 93454
rect 271804 93134 272404 93218
rect 271804 92898 271986 93134
rect 272222 92898 272404 93134
rect 271804 57454 272404 92898
rect 271804 57218 271986 57454
rect 272222 57218 272404 57454
rect 271804 57134 272404 57218
rect 271804 56898 271986 57134
rect 272222 56898 272404 57134
rect 271804 21454 272404 56898
rect 271804 21218 271986 21454
rect 272222 21218 272404 21454
rect 271804 21134 272404 21218
rect 271804 20898 271986 21134
rect 272222 20898 272404 21134
rect 271804 -1286 272404 20898
rect 271804 -1522 271986 -1286
rect 272222 -1522 272404 -1286
rect 271804 -1606 272404 -1522
rect 271804 -1842 271986 -1606
rect 272222 -1842 272404 -1606
rect 271804 -1864 272404 -1842
rect 275404 313054 276004 326000
rect 275404 312818 275586 313054
rect 275822 312818 276004 313054
rect 275404 312734 276004 312818
rect 275404 312498 275586 312734
rect 275822 312498 276004 312734
rect 275404 277054 276004 312498
rect 275404 276818 275586 277054
rect 275822 276818 276004 277054
rect 275404 276734 276004 276818
rect 275404 276498 275586 276734
rect 275822 276498 276004 276734
rect 275404 241054 276004 276498
rect 275404 240818 275586 241054
rect 275822 240818 276004 241054
rect 275404 240734 276004 240818
rect 275404 240498 275586 240734
rect 275822 240498 276004 240734
rect 275404 205054 276004 240498
rect 275404 204818 275586 205054
rect 275822 204818 276004 205054
rect 275404 204734 276004 204818
rect 275404 204498 275586 204734
rect 275822 204498 276004 204734
rect 275404 169054 276004 204498
rect 275404 168818 275586 169054
rect 275822 168818 276004 169054
rect 275404 168734 276004 168818
rect 275404 168498 275586 168734
rect 275822 168498 276004 168734
rect 275404 133054 276004 168498
rect 275404 132818 275586 133054
rect 275822 132818 276004 133054
rect 275404 132734 276004 132818
rect 275404 132498 275586 132734
rect 275822 132498 276004 132734
rect 275404 97054 276004 132498
rect 275404 96818 275586 97054
rect 275822 96818 276004 97054
rect 275404 96734 276004 96818
rect 275404 96498 275586 96734
rect 275822 96498 276004 96734
rect 275404 61054 276004 96498
rect 275404 60818 275586 61054
rect 275822 60818 276004 61054
rect 275404 60734 276004 60818
rect 275404 60498 275586 60734
rect 275822 60498 276004 60734
rect 275404 25054 276004 60498
rect 275404 24818 275586 25054
rect 275822 24818 276004 25054
rect 275404 24734 276004 24818
rect 275404 24498 275586 24734
rect 275822 24498 276004 24734
rect 275404 -3166 276004 24498
rect 275404 -3402 275586 -3166
rect 275822 -3402 276004 -3166
rect 275404 -3486 276004 -3402
rect 275404 -3722 275586 -3486
rect 275822 -3722 276004 -3486
rect 275404 -3744 276004 -3722
rect 279004 316654 279604 326000
rect 279004 316418 279186 316654
rect 279422 316418 279604 316654
rect 279004 316334 279604 316418
rect 279004 316098 279186 316334
rect 279422 316098 279604 316334
rect 279004 280654 279604 316098
rect 279004 280418 279186 280654
rect 279422 280418 279604 280654
rect 279004 280334 279604 280418
rect 279004 280098 279186 280334
rect 279422 280098 279604 280334
rect 279004 244654 279604 280098
rect 279004 244418 279186 244654
rect 279422 244418 279604 244654
rect 279004 244334 279604 244418
rect 279004 244098 279186 244334
rect 279422 244098 279604 244334
rect 279004 208654 279604 244098
rect 279004 208418 279186 208654
rect 279422 208418 279604 208654
rect 279004 208334 279604 208418
rect 279004 208098 279186 208334
rect 279422 208098 279604 208334
rect 279004 172654 279604 208098
rect 279004 172418 279186 172654
rect 279422 172418 279604 172654
rect 279004 172334 279604 172418
rect 279004 172098 279186 172334
rect 279422 172098 279604 172334
rect 279004 136654 279604 172098
rect 279004 136418 279186 136654
rect 279422 136418 279604 136654
rect 279004 136334 279604 136418
rect 279004 136098 279186 136334
rect 279422 136098 279604 136334
rect 279004 100654 279604 136098
rect 279004 100418 279186 100654
rect 279422 100418 279604 100654
rect 279004 100334 279604 100418
rect 279004 100098 279186 100334
rect 279422 100098 279604 100334
rect 279004 64654 279604 100098
rect 279004 64418 279186 64654
rect 279422 64418 279604 64654
rect 279004 64334 279604 64418
rect 279004 64098 279186 64334
rect 279422 64098 279604 64334
rect 279004 28654 279604 64098
rect 279004 28418 279186 28654
rect 279422 28418 279604 28654
rect 279004 28334 279604 28418
rect 279004 28098 279186 28334
rect 279422 28098 279604 28334
rect 279004 -5046 279604 28098
rect 279004 -5282 279186 -5046
rect 279422 -5282 279604 -5046
rect 279004 -5366 279604 -5282
rect 279004 -5602 279186 -5366
rect 279422 -5602 279604 -5366
rect 279004 -5624 279604 -5602
rect 282604 320254 283204 326000
rect 282604 320018 282786 320254
rect 283022 320018 283204 320254
rect 282604 319934 283204 320018
rect 282604 319698 282786 319934
rect 283022 319698 283204 319934
rect 282604 284254 283204 319698
rect 282604 284018 282786 284254
rect 283022 284018 283204 284254
rect 282604 283934 283204 284018
rect 282604 283698 282786 283934
rect 283022 283698 283204 283934
rect 282604 248254 283204 283698
rect 282604 248018 282786 248254
rect 283022 248018 283204 248254
rect 282604 247934 283204 248018
rect 282604 247698 282786 247934
rect 283022 247698 283204 247934
rect 282604 212254 283204 247698
rect 282604 212018 282786 212254
rect 283022 212018 283204 212254
rect 282604 211934 283204 212018
rect 282604 211698 282786 211934
rect 283022 211698 283204 211934
rect 282604 176254 283204 211698
rect 282604 176018 282786 176254
rect 283022 176018 283204 176254
rect 282604 175934 283204 176018
rect 282604 175698 282786 175934
rect 283022 175698 283204 175934
rect 282604 140254 283204 175698
rect 282604 140018 282786 140254
rect 283022 140018 283204 140254
rect 282604 139934 283204 140018
rect 282604 139698 282786 139934
rect 283022 139698 283204 139934
rect 282604 104254 283204 139698
rect 282604 104018 282786 104254
rect 283022 104018 283204 104254
rect 282604 103934 283204 104018
rect 282604 103698 282786 103934
rect 283022 103698 283204 103934
rect 282604 68254 283204 103698
rect 282604 68018 282786 68254
rect 283022 68018 283204 68254
rect 282604 67934 283204 68018
rect 282604 67698 282786 67934
rect 283022 67698 283204 67934
rect 282604 32254 283204 67698
rect 282604 32018 282786 32254
rect 283022 32018 283204 32254
rect 282604 31934 283204 32018
rect 282604 31698 282786 31934
rect 283022 31698 283204 31934
rect 264604 -6222 264786 -5986
rect 265022 -6222 265204 -5986
rect 264604 -6306 265204 -6222
rect 264604 -6542 264786 -6306
rect 265022 -6542 265204 -6306
rect 264604 -7504 265204 -6542
rect 282604 -6926 283204 31698
rect 289804 291454 290404 326000
rect 289804 291218 289986 291454
rect 290222 291218 290404 291454
rect 289804 291134 290404 291218
rect 289804 290898 289986 291134
rect 290222 290898 290404 291134
rect 289804 255454 290404 290898
rect 289804 255218 289986 255454
rect 290222 255218 290404 255454
rect 289804 255134 290404 255218
rect 289804 254898 289986 255134
rect 290222 254898 290404 255134
rect 289804 219454 290404 254898
rect 289804 219218 289986 219454
rect 290222 219218 290404 219454
rect 289804 219134 290404 219218
rect 289804 218898 289986 219134
rect 290222 218898 290404 219134
rect 289804 183454 290404 218898
rect 289804 183218 289986 183454
rect 290222 183218 290404 183454
rect 289804 183134 290404 183218
rect 289804 182898 289986 183134
rect 290222 182898 290404 183134
rect 289804 147454 290404 182898
rect 289804 147218 289986 147454
rect 290222 147218 290404 147454
rect 289804 147134 290404 147218
rect 289804 146898 289986 147134
rect 290222 146898 290404 147134
rect 289804 111454 290404 146898
rect 289804 111218 289986 111454
rect 290222 111218 290404 111454
rect 289804 111134 290404 111218
rect 289804 110898 289986 111134
rect 290222 110898 290404 111134
rect 289804 75454 290404 110898
rect 289804 75218 289986 75454
rect 290222 75218 290404 75454
rect 289804 75134 290404 75218
rect 289804 74898 289986 75134
rect 290222 74898 290404 75134
rect 289804 39454 290404 74898
rect 289804 39218 289986 39454
rect 290222 39218 290404 39454
rect 289804 39134 290404 39218
rect 289804 38898 289986 39134
rect 290222 38898 290404 39134
rect 289804 3454 290404 38898
rect 289804 3218 289986 3454
rect 290222 3218 290404 3454
rect 289804 3134 290404 3218
rect 289804 2898 289986 3134
rect 290222 2898 290404 3134
rect 289804 -346 290404 2898
rect 289804 -582 289986 -346
rect 290222 -582 290404 -346
rect 289804 -666 290404 -582
rect 289804 -902 289986 -666
rect 290222 -902 290404 -666
rect 289804 -1864 290404 -902
rect 293404 295054 294004 326000
rect 293404 294818 293586 295054
rect 293822 294818 294004 295054
rect 293404 294734 294004 294818
rect 293404 294498 293586 294734
rect 293822 294498 294004 294734
rect 293404 259054 294004 294498
rect 293404 258818 293586 259054
rect 293822 258818 294004 259054
rect 293404 258734 294004 258818
rect 293404 258498 293586 258734
rect 293822 258498 294004 258734
rect 293404 223054 294004 258498
rect 293404 222818 293586 223054
rect 293822 222818 294004 223054
rect 293404 222734 294004 222818
rect 293404 222498 293586 222734
rect 293822 222498 294004 222734
rect 293404 187054 294004 222498
rect 293404 186818 293586 187054
rect 293822 186818 294004 187054
rect 293404 186734 294004 186818
rect 293404 186498 293586 186734
rect 293822 186498 294004 186734
rect 293404 151054 294004 186498
rect 293404 150818 293586 151054
rect 293822 150818 294004 151054
rect 293404 150734 294004 150818
rect 293404 150498 293586 150734
rect 293822 150498 294004 150734
rect 293404 115054 294004 150498
rect 293404 114818 293586 115054
rect 293822 114818 294004 115054
rect 293404 114734 294004 114818
rect 293404 114498 293586 114734
rect 293822 114498 294004 114734
rect 293404 79054 294004 114498
rect 293404 78818 293586 79054
rect 293822 78818 294004 79054
rect 293404 78734 294004 78818
rect 293404 78498 293586 78734
rect 293822 78498 294004 78734
rect 293404 43054 294004 78498
rect 293404 42818 293586 43054
rect 293822 42818 294004 43054
rect 293404 42734 294004 42818
rect 293404 42498 293586 42734
rect 293822 42498 294004 42734
rect 293404 7054 294004 42498
rect 293404 6818 293586 7054
rect 293822 6818 294004 7054
rect 293404 6734 294004 6818
rect 293404 6498 293586 6734
rect 293822 6498 294004 6734
rect 293404 -2226 294004 6498
rect 293404 -2462 293586 -2226
rect 293822 -2462 294004 -2226
rect 293404 -2546 294004 -2462
rect 293404 -2782 293586 -2546
rect 293822 -2782 294004 -2546
rect 293404 -3744 294004 -2782
rect 297004 298654 297604 326000
rect 297004 298418 297186 298654
rect 297422 298418 297604 298654
rect 297004 298334 297604 298418
rect 297004 298098 297186 298334
rect 297422 298098 297604 298334
rect 297004 262654 297604 298098
rect 297004 262418 297186 262654
rect 297422 262418 297604 262654
rect 297004 262334 297604 262418
rect 297004 262098 297186 262334
rect 297422 262098 297604 262334
rect 297004 226654 297604 262098
rect 297004 226418 297186 226654
rect 297422 226418 297604 226654
rect 297004 226334 297604 226418
rect 297004 226098 297186 226334
rect 297422 226098 297604 226334
rect 297004 190654 297604 226098
rect 297004 190418 297186 190654
rect 297422 190418 297604 190654
rect 297004 190334 297604 190418
rect 297004 190098 297186 190334
rect 297422 190098 297604 190334
rect 297004 154654 297604 190098
rect 297004 154418 297186 154654
rect 297422 154418 297604 154654
rect 297004 154334 297604 154418
rect 297004 154098 297186 154334
rect 297422 154098 297604 154334
rect 297004 118654 297604 154098
rect 297004 118418 297186 118654
rect 297422 118418 297604 118654
rect 297004 118334 297604 118418
rect 297004 118098 297186 118334
rect 297422 118098 297604 118334
rect 297004 82654 297604 118098
rect 297004 82418 297186 82654
rect 297422 82418 297604 82654
rect 297004 82334 297604 82418
rect 297004 82098 297186 82334
rect 297422 82098 297604 82334
rect 297004 46654 297604 82098
rect 297004 46418 297186 46654
rect 297422 46418 297604 46654
rect 297004 46334 297604 46418
rect 297004 46098 297186 46334
rect 297422 46098 297604 46334
rect 297004 10654 297604 46098
rect 297004 10418 297186 10654
rect 297422 10418 297604 10654
rect 297004 10334 297604 10418
rect 297004 10098 297186 10334
rect 297422 10098 297604 10334
rect 297004 -4106 297604 10098
rect 297004 -4342 297186 -4106
rect 297422 -4342 297604 -4106
rect 297004 -4426 297604 -4342
rect 297004 -4662 297186 -4426
rect 297422 -4662 297604 -4426
rect 297004 -5624 297604 -4662
rect 300604 302254 301204 326000
rect 300604 302018 300786 302254
rect 301022 302018 301204 302254
rect 300604 301934 301204 302018
rect 300604 301698 300786 301934
rect 301022 301698 301204 301934
rect 300604 266254 301204 301698
rect 300604 266018 300786 266254
rect 301022 266018 301204 266254
rect 300604 265934 301204 266018
rect 300604 265698 300786 265934
rect 301022 265698 301204 265934
rect 300604 230254 301204 265698
rect 300604 230018 300786 230254
rect 301022 230018 301204 230254
rect 300604 229934 301204 230018
rect 300604 229698 300786 229934
rect 301022 229698 301204 229934
rect 300604 194254 301204 229698
rect 300604 194018 300786 194254
rect 301022 194018 301204 194254
rect 300604 193934 301204 194018
rect 300604 193698 300786 193934
rect 301022 193698 301204 193934
rect 300604 158254 301204 193698
rect 300604 158018 300786 158254
rect 301022 158018 301204 158254
rect 300604 157934 301204 158018
rect 300604 157698 300786 157934
rect 301022 157698 301204 157934
rect 300604 122254 301204 157698
rect 300604 122018 300786 122254
rect 301022 122018 301204 122254
rect 300604 121934 301204 122018
rect 300604 121698 300786 121934
rect 301022 121698 301204 121934
rect 300604 86254 301204 121698
rect 300604 86018 300786 86254
rect 301022 86018 301204 86254
rect 300604 85934 301204 86018
rect 300604 85698 300786 85934
rect 301022 85698 301204 85934
rect 300604 50254 301204 85698
rect 300604 50018 300786 50254
rect 301022 50018 301204 50254
rect 300604 49934 301204 50018
rect 300604 49698 300786 49934
rect 301022 49698 301204 49934
rect 300604 14254 301204 49698
rect 300604 14018 300786 14254
rect 301022 14018 301204 14254
rect 300604 13934 301204 14018
rect 300604 13698 300786 13934
rect 301022 13698 301204 13934
rect 282604 -7162 282786 -6926
rect 283022 -7162 283204 -6926
rect 282604 -7246 283204 -7162
rect 282604 -7482 282786 -7246
rect 283022 -7482 283204 -7246
rect 282604 -7504 283204 -7482
rect 300604 -5986 301204 13698
rect 307804 309454 308404 326000
rect 307804 309218 307986 309454
rect 308222 309218 308404 309454
rect 307804 309134 308404 309218
rect 307804 308898 307986 309134
rect 308222 308898 308404 309134
rect 307804 273454 308404 308898
rect 307804 273218 307986 273454
rect 308222 273218 308404 273454
rect 307804 273134 308404 273218
rect 307804 272898 307986 273134
rect 308222 272898 308404 273134
rect 307804 237454 308404 272898
rect 307804 237218 307986 237454
rect 308222 237218 308404 237454
rect 307804 237134 308404 237218
rect 307804 236898 307986 237134
rect 308222 236898 308404 237134
rect 307804 201454 308404 236898
rect 307804 201218 307986 201454
rect 308222 201218 308404 201454
rect 307804 201134 308404 201218
rect 307804 200898 307986 201134
rect 308222 200898 308404 201134
rect 307804 165454 308404 200898
rect 307804 165218 307986 165454
rect 308222 165218 308404 165454
rect 307804 165134 308404 165218
rect 307804 164898 307986 165134
rect 308222 164898 308404 165134
rect 307804 129454 308404 164898
rect 307804 129218 307986 129454
rect 308222 129218 308404 129454
rect 307804 129134 308404 129218
rect 307804 128898 307986 129134
rect 308222 128898 308404 129134
rect 307804 93454 308404 128898
rect 307804 93218 307986 93454
rect 308222 93218 308404 93454
rect 307804 93134 308404 93218
rect 307804 92898 307986 93134
rect 308222 92898 308404 93134
rect 307804 57454 308404 92898
rect 307804 57218 307986 57454
rect 308222 57218 308404 57454
rect 307804 57134 308404 57218
rect 307804 56898 307986 57134
rect 308222 56898 308404 57134
rect 307804 21454 308404 56898
rect 307804 21218 307986 21454
rect 308222 21218 308404 21454
rect 307804 21134 308404 21218
rect 307804 20898 307986 21134
rect 308222 20898 308404 21134
rect 307804 -1286 308404 20898
rect 307804 -1522 307986 -1286
rect 308222 -1522 308404 -1286
rect 307804 -1606 308404 -1522
rect 307804 -1842 307986 -1606
rect 308222 -1842 308404 -1606
rect 307804 -1864 308404 -1842
rect 311404 313054 312004 326000
rect 311404 312818 311586 313054
rect 311822 312818 312004 313054
rect 311404 312734 312004 312818
rect 311404 312498 311586 312734
rect 311822 312498 312004 312734
rect 311404 277054 312004 312498
rect 311404 276818 311586 277054
rect 311822 276818 312004 277054
rect 311404 276734 312004 276818
rect 311404 276498 311586 276734
rect 311822 276498 312004 276734
rect 311404 241054 312004 276498
rect 311404 240818 311586 241054
rect 311822 240818 312004 241054
rect 311404 240734 312004 240818
rect 311404 240498 311586 240734
rect 311822 240498 312004 240734
rect 311404 205054 312004 240498
rect 311404 204818 311586 205054
rect 311822 204818 312004 205054
rect 311404 204734 312004 204818
rect 311404 204498 311586 204734
rect 311822 204498 312004 204734
rect 311404 169054 312004 204498
rect 311404 168818 311586 169054
rect 311822 168818 312004 169054
rect 311404 168734 312004 168818
rect 311404 168498 311586 168734
rect 311822 168498 312004 168734
rect 311404 133054 312004 168498
rect 311404 132818 311586 133054
rect 311822 132818 312004 133054
rect 311404 132734 312004 132818
rect 311404 132498 311586 132734
rect 311822 132498 312004 132734
rect 311404 97054 312004 132498
rect 311404 96818 311586 97054
rect 311822 96818 312004 97054
rect 311404 96734 312004 96818
rect 311404 96498 311586 96734
rect 311822 96498 312004 96734
rect 311404 61054 312004 96498
rect 311404 60818 311586 61054
rect 311822 60818 312004 61054
rect 311404 60734 312004 60818
rect 311404 60498 311586 60734
rect 311822 60498 312004 60734
rect 311404 25054 312004 60498
rect 311404 24818 311586 25054
rect 311822 24818 312004 25054
rect 311404 24734 312004 24818
rect 311404 24498 311586 24734
rect 311822 24498 312004 24734
rect 311404 -3166 312004 24498
rect 311404 -3402 311586 -3166
rect 311822 -3402 312004 -3166
rect 311404 -3486 312004 -3402
rect 311404 -3722 311586 -3486
rect 311822 -3722 312004 -3486
rect 311404 -3744 312004 -3722
rect 315004 316654 315604 326000
rect 315004 316418 315186 316654
rect 315422 316418 315604 316654
rect 315004 316334 315604 316418
rect 315004 316098 315186 316334
rect 315422 316098 315604 316334
rect 315004 280654 315604 316098
rect 315004 280418 315186 280654
rect 315422 280418 315604 280654
rect 315004 280334 315604 280418
rect 315004 280098 315186 280334
rect 315422 280098 315604 280334
rect 315004 244654 315604 280098
rect 315004 244418 315186 244654
rect 315422 244418 315604 244654
rect 315004 244334 315604 244418
rect 315004 244098 315186 244334
rect 315422 244098 315604 244334
rect 315004 208654 315604 244098
rect 315004 208418 315186 208654
rect 315422 208418 315604 208654
rect 315004 208334 315604 208418
rect 315004 208098 315186 208334
rect 315422 208098 315604 208334
rect 315004 172654 315604 208098
rect 315004 172418 315186 172654
rect 315422 172418 315604 172654
rect 315004 172334 315604 172418
rect 315004 172098 315186 172334
rect 315422 172098 315604 172334
rect 315004 136654 315604 172098
rect 315004 136418 315186 136654
rect 315422 136418 315604 136654
rect 315004 136334 315604 136418
rect 315004 136098 315186 136334
rect 315422 136098 315604 136334
rect 315004 100654 315604 136098
rect 315004 100418 315186 100654
rect 315422 100418 315604 100654
rect 315004 100334 315604 100418
rect 315004 100098 315186 100334
rect 315422 100098 315604 100334
rect 315004 64654 315604 100098
rect 315004 64418 315186 64654
rect 315422 64418 315604 64654
rect 315004 64334 315604 64418
rect 315004 64098 315186 64334
rect 315422 64098 315604 64334
rect 315004 28654 315604 64098
rect 315004 28418 315186 28654
rect 315422 28418 315604 28654
rect 315004 28334 315604 28418
rect 315004 28098 315186 28334
rect 315422 28098 315604 28334
rect 315004 -5046 315604 28098
rect 315004 -5282 315186 -5046
rect 315422 -5282 315604 -5046
rect 315004 -5366 315604 -5282
rect 315004 -5602 315186 -5366
rect 315422 -5602 315604 -5366
rect 315004 -5624 315604 -5602
rect 318604 320254 319204 326000
rect 318604 320018 318786 320254
rect 319022 320018 319204 320254
rect 318604 319934 319204 320018
rect 318604 319698 318786 319934
rect 319022 319698 319204 319934
rect 318604 284254 319204 319698
rect 318604 284018 318786 284254
rect 319022 284018 319204 284254
rect 318604 283934 319204 284018
rect 318604 283698 318786 283934
rect 319022 283698 319204 283934
rect 318604 248254 319204 283698
rect 318604 248018 318786 248254
rect 319022 248018 319204 248254
rect 318604 247934 319204 248018
rect 318604 247698 318786 247934
rect 319022 247698 319204 247934
rect 318604 212254 319204 247698
rect 318604 212018 318786 212254
rect 319022 212018 319204 212254
rect 318604 211934 319204 212018
rect 318604 211698 318786 211934
rect 319022 211698 319204 211934
rect 318604 176254 319204 211698
rect 318604 176018 318786 176254
rect 319022 176018 319204 176254
rect 318604 175934 319204 176018
rect 318604 175698 318786 175934
rect 319022 175698 319204 175934
rect 318604 140254 319204 175698
rect 318604 140018 318786 140254
rect 319022 140018 319204 140254
rect 318604 139934 319204 140018
rect 318604 139698 318786 139934
rect 319022 139698 319204 139934
rect 318604 104254 319204 139698
rect 318604 104018 318786 104254
rect 319022 104018 319204 104254
rect 318604 103934 319204 104018
rect 318604 103698 318786 103934
rect 319022 103698 319204 103934
rect 318604 68254 319204 103698
rect 318604 68018 318786 68254
rect 319022 68018 319204 68254
rect 318604 67934 319204 68018
rect 318604 67698 318786 67934
rect 319022 67698 319204 67934
rect 318604 32254 319204 67698
rect 318604 32018 318786 32254
rect 319022 32018 319204 32254
rect 318604 31934 319204 32018
rect 318604 31698 318786 31934
rect 319022 31698 319204 31934
rect 300604 -6222 300786 -5986
rect 301022 -6222 301204 -5986
rect 300604 -6306 301204 -6222
rect 300604 -6542 300786 -6306
rect 301022 -6542 301204 -6306
rect 300604 -7504 301204 -6542
rect 318604 -6926 319204 31698
rect 325804 291454 326404 326000
rect 325804 291218 325986 291454
rect 326222 291218 326404 291454
rect 325804 291134 326404 291218
rect 325804 290898 325986 291134
rect 326222 290898 326404 291134
rect 325804 255454 326404 290898
rect 325804 255218 325986 255454
rect 326222 255218 326404 255454
rect 325804 255134 326404 255218
rect 325804 254898 325986 255134
rect 326222 254898 326404 255134
rect 325804 219454 326404 254898
rect 325804 219218 325986 219454
rect 326222 219218 326404 219454
rect 325804 219134 326404 219218
rect 325804 218898 325986 219134
rect 326222 218898 326404 219134
rect 325804 183454 326404 218898
rect 325804 183218 325986 183454
rect 326222 183218 326404 183454
rect 325804 183134 326404 183218
rect 325804 182898 325986 183134
rect 326222 182898 326404 183134
rect 325804 147454 326404 182898
rect 325804 147218 325986 147454
rect 326222 147218 326404 147454
rect 325804 147134 326404 147218
rect 325804 146898 325986 147134
rect 326222 146898 326404 147134
rect 325804 111454 326404 146898
rect 325804 111218 325986 111454
rect 326222 111218 326404 111454
rect 325804 111134 326404 111218
rect 325804 110898 325986 111134
rect 326222 110898 326404 111134
rect 325804 75454 326404 110898
rect 325804 75218 325986 75454
rect 326222 75218 326404 75454
rect 325804 75134 326404 75218
rect 325804 74898 325986 75134
rect 326222 74898 326404 75134
rect 325804 39454 326404 74898
rect 325804 39218 325986 39454
rect 326222 39218 326404 39454
rect 325804 39134 326404 39218
rect 325804 38898 325986 39134
rect 326222 38898 326404 39134
rect 325804 3454 326404 38898
rect 325804 3218 325986 3454
rect 326222 3218 326404 3454
rect 325804 3134 326404 3218
rect 325804 2898 325986 3134
rect 326222 2898 326404 3134
rect 325804 -346 326404 2898
rect 325804 -582 325986 -346
rect 326222 -582 326404 -346
rect 325804 -666 326404 -582
rect 325804 -902 325986 -666
rect 326222 -902 326404 -666
rect 325804 -1864 326404 -902
rect 329404 295054 330004 326000
rect 329404 294818 329586 295054
rect 329822 294818 330004 295054
rect 329404 294734 330004 294818
rect 329404 294498 329586 294734
rect 329822 294498 330004 294734
rect 329404 259054 330004 294498
rect 329404 258818 329586 259054
rect 329822 258818 330004 259054
rect 329404 258734 330004 258818
rect 329404 258498 329586 258734
rect 329822 258498 330004 258734
rect 329404 223054 330004 258498
rect 329404 222818 329586 223054
rect 329822 222818 330004 223054
rect 329404 222734 330004 222818
rect 329404 222498 329586 222734
rect 329822 222498 330004 222734
rect 329404 187054 330004 222498
rect 329404 186818 329586 187054
rect 329822 186818 330004 187054
rect 329404 186734 330004 186818
rect 329404 186498 329586 186734
rect 329822 186498 330004 186734
rect 329404 151054 330004 186498
rect 329404 150818 329586 151054
rect 329822 150818 330004 151054
rect 329404 150734 330004 150818
rect 329404 150498 329586 150734
rect 329822 150498 330004 150734
rect 329404 115054 330004 150498
rect 329404 114818 329586 115054
rect 329822 114818 330004 115054
rect 329404 114734 330004 114818
rect 329404 114498 329586 114734
rect 329822 114498 330004 114734
rect 329404 79054 330004 114498
rect 329404 78818 329586 79054
rect 329822 78818 330004 79054
rect 329404 78734 330004 78818
rect 329404 78498 329586 78734
rect 329822 78498 330004 78734
rect 329404 43054 330004 78498
rect 329404 42818 329586 43054
rect 329822 42818 330004 43054
rect 329404 42734 330004 42818
rect 329404 42498 329586 42734
rect 329822 42498 330004 42734
rect 329404 7054 330004 42498
rect 329404 6818 329586 7054
rect 329822 6818 330004 7054
rect 329404 6734 330004 6818
rect 329404 6498 329586 6734
rect 329822 6498 330004 6734
rect 329404 -2226 330004 6498
rect 329404 -2462 329586 -2226
rect 329822 -2462 330004 -2226
rect 329404 -2546 330004 -2462
rect 329404 -2782 329586 -2546
rect 329822 -2782 330004 -2546
rect 329404 -3744 330004 -2782
rect 333004 298654 333604 326000
rect 333004 298418 333186 298654
rect 333422 298418 333604 298654
rect 333004 298334 333604 298418
rect 333004 298098 333186 298334
rect 333422 298098 333604 298334
rect 333004 262654 333604 298098
rect 333004 262418 333186 262654
rect 333422 262418 333604 262654
rect 333004 262334 333604 262418
rect 333004 262098 333186 262334
rect 333422 262098 333604 262334
rect 333004 226654 333604 262098
rect 333004 226418 333186 226654
rect 333422 226418 333604 226654
rect 333004 226334 333604 226418
rect 333004 226098 333186 226334
rect 333422 226098 333604 226334
rect 333004 190654 333604 226098
rect 333004 190418 333186 190654
rect 333422 190418 333604 190654
rect 333004 190334 333604 190418
rect 333004 190098 333186 190334
rect 333422 190098 333604 190334
rect 333004 154654 333604 190098
rect 333004 154418 333186 154654
rect 333422 154418 333604 154654
rect 333004 154334 333604 154418
rect 333004 154098 333186 154334
rect 333422 154098 333604 154334
rect 333004 118654 333604 154098
rect 333004 118418 333186 118654
rect 333422 118418 333604 118654
rect 333004 118334 333604 118418
rect 333004 118098 333186 118334
rect 333422 118098 333604 118334
rect 333004 82654 333604 118098
rect 333004 82418 333186 82654
rect 333422 82418 333604 82654
rect 333004 82334 333604 82418
rect 333004 82098 333186 82334
rect 333422 82098 333604 82334
rect 333004 46654 333604 82098
rect 333004 46418 333186 46654
rect 333422 46418 333604 46654
rect 333004 46334 333604 46418
rect 333004 46098 333186 46334
rect 333422 46098 333604 46334
rect 333004 10654 333604 46098
rect 333004 10418 333186 10654
rect 333422 10418 333604 10654
rect 333004 10334 333604 10418
rect 333004 10098 333186 10334
rect 333422 10098 333604 10334
rect 333004 -4106 333604 10098
rect 333004 -4342 333186 -4106
rect 333422 -4342 333604 -4106
rect 333004 -4426 333604 -4342
rect 333004 -4662 333186 -4426
rect 333422 -4662 333604 -4426
rect 333004 -5624 333604 -4662
rect 336604 302254 337204 326000
rect 336604 302018 336786 302254
rect 337022 302018 337204 302254
rect 336604 301934 337204 302018
rect 336604 301698 336786 301934
rect 337022 301698 337204 301934
rect 336604 266254 337204 301698
rect 336604 266018 336786 266254
rect 337022 266018 337204 266254
rect 336604 265934 337204 266018
rect 336604 265698 336786 265934
rect 337022 265698 337204 265934
rect 336604 230254 337204 265698
rect 336604 230018 336786 230254
rect 337022 230018 337204 230254
rect 336604 229934 337204 230018
rect 336604 229698 336786 229934
rect 337022 229698 337204 229934
rect 336604 194254 337204 229698
rect 336604 194018 336786 194254
rect 337022 194018 337204 194254
rect 336604 193934 337204 194018
rect 336604 193698 336786 193934
rect 337022 193698 337204 193934
rect 336604 158254 337204 193698
rect 336604 158018 336786 158254
rect 337022 158018 337204 158254
rect 336604 157934 337204 158018
rect 336604 157698 336786 157934
rect 337022 157698 337204 157934
rect 336604 122254 337204 157698
rect 336604 122018 336786 122254
rect 337022 122018 337204 122254
rect 336604 121934 337204 122018
rect 336604 121698 336786 121934
rect 337022 121698 337204 121934
rect 336604 86254 337204 121698
rect 336604 86018 336786 86254
rect 337022 86018 337204 86254
rect 336604 85934 337204 86018
rect 336604 85698 336786 85934
rect 337022 85698 337204 85934
rect 336604 50254 337204 85698
rect 336604 50018 336786 50254
rect 337022 50018 337204 50254
rect 336604 49934 337204 50018
rect 336604 49698 336786 49934
rect 337022 49698 337204 49934
rect 336604 14254 337204 49698
rect 336604 14018 336786 14254
rect 337022 14018 337204 14254
rect 336604 13934 337204 14018
rect 336604 13698 336786 13934
rect 337022 13698 337204 13934
rect 318604 -7162 318786 -6926
rect 319022 -7162 319204 -6926
rect 318604 -7246 319204 -7162
rect 318604 -7482 318786 -7246
rect 319022 -7482 319204 -7246
rect 318604 -7504 319204 -7482
rect 336604 -5986 337204 13698
rect 343804 309454 344404 326000
rect 343804 309218 343986 309454
rect 344222 309218 344404 309454
rect 343804 309134 344404 309218
rect 343804 308898 343986 309134
rect 344222 308898 344404 309134
rect 343804 273454 344404 308898
rect 343804 273218 343986 273454
rect 344222 273218 344404 273454
rect 343804 273134 344404 273218
rect 343804 272898 343986 273134
rect 344222 272898 344404 273134
rect 343804 237454 344404 272898
rect 343804 237218 343986 237454
rect 344222 237218 344404 237454
rect 343804 237134 344404 237218
rect 343804 236898 343986 237134
rect 344222 236898 344404 237134
rect 343804 201454 344404 236898
rect 343804 201218 343986 201454
rect 344222 201218 344404 201454
rect 343804 201134 344404 201218
rect 343804 200898 343986 201134
rect 344222 200898 344404 201134
rect 343804 165454 344404 200898
rect 343804 165218 343986 165454
rect 344222 165218 344404 165454
rect 343804 165134 344404 165218
rect 343804 164898 343986 165134
rect 344222 164898 344404 165134
rect 343804 129454 344404 164898
rect 343804 129218 343986 129454
rect 344222 129218 344404 129454
rect 343804 129134 344404 129218
rect 343804 128898 343986 129134
rect 344222 128898 344404 129134
rect 343804 93454 344404 128898
rect 343804 93218 343986 93454
rect 344222 93218 344404 93454
rect 343804 93134 344404 93218
rect 343804 92898 343986 93134
rect 344222 92898 344404 93134
rect 343804 57454 344404 92898
rect 343804 57218 343986 57454
rect 344222 57218 344404 57454
rect 343804 57134 344404 57218
rect 343804 56898 343986 57134
rect 344222 56898 344404 57134
rect 343804 21454 344404 56898
rect 343804 21218 343986 21454
rect 344222 21218 344404 21454
rect 343804 21134 344404 21218
rect 343804 20898 343986 21134
rect 344222 20898 344404 21134
rect 343804 -1286 344404 20898
rect 343804 -1522 343986 -1286
rect 344222 -1522 344404 -1286
rect 343804 -1606 344404 -1522
rect 343804 -1842 343986 -1606
rect 344222 -1842 344404 -1606
rect 343804 -1864 344404 -1842
rect 347404 313054 348004 326000
rect 347404 312818 347586 313054
rect 347822 312818 348004 313054
rect 347404 312734 348004 312818
rect 347404 312498 347586 312734
rect 347822 312498 348004 312734
rect 347404 277054 348004 312498
rect 347404 276818 347586 277054
rect 347822 276818 348004 277054
rect 347404 276734 348004 276818
rect 347404 276498 347586 276734
rect 347822 276498 348004 276734
rect 347404 241054 348004 276498
rect 347404 240818 347586 241054
rect 347822 240818 348004 241054
rect 347404 240734 348004 240818
rect 347404 240498 347586 240734
rect 347822 240498 348004 240734
rect 347404 205054 348004 240498
rect 347404 204818 347586 205054
rect 347822 204818 348004 205054
rect 347404 204734 348004 204818
rect 347404 204498 347586 204734
rect 347822 204498 348004 204734
rect 347404 169054 348004 204498
rect 347404 168818 347586 169054
rect 347822 168818 348004 169054
rect 347404 168734 348004 168818
rect 347404 168498 347586 168734
rect 347822 168498 348004 168734
rect 347404 133054 348004 168498
rect 347404 132818 347586 133054
rect 347822 132818 348004 133054
rect 347404 132734 348004 132818
rect 347404 132498 347586 132734
rect 347822 132498 348004 132734
rect 347404 97054 348004 132498
rect 347404 96818 347586 97054
rect 347822 96818 348004 97054
rect 347404 96734 348004 96818
rect 347404 96498 347586 96734
rect 347822 96498 348004 96734
rect 347404 61054 348004 96498
rect 347404 60818 347586 61054
rect 347822 60818 348004 61054
rect 347404 60734 348004 60818
rect 347404 60498 347586 60734
rect 347822 60498 348004 60734
rect 347404 25054 348004 60498
rect 347404 24818 347586 25054
rect 347822 24818 348004 25054
rect 347404 24734 348004 24818
rect 347404 24498 347586 24734
rect 347822 24498 348004 24734
rect 347404 -3166 348004 24498
rect 347404 -3402 347586 -3166
rect 347822 -3402 348004 -3166
rect 347404 -3486 348004 -3402
rect 347404 -3722 347586 -3486
rect 347822 -3722 348004 -3486
rect 347404 -3744 348004 -3722
rect 351004 316654 351604 326000
rect 351004 316418 351186 316654
rect 351422 316418 351604 316654
rect 351004 316334 351604 316418
rect 351004 316098 351186 316334
rect 351422 316098 351604 316334
rect 351004 280654 351604 316098
rect 351004 280418 351186 280654
rect 351422 280418 351604 280654
rect 351004 280334 351604 280418
rect 351004 280098 351186 280334
rect 351422 280098 351604 280334
rect 351004 244654 351604 280098
rect 351004 244418 351186 244654
rect 351422 244418 351604 244654
rect 351004 244334 351604 244418
rect 351004 244098 351186 244334
rect 351422 244098 351604 244334
rect 351004 208654 351604 244098
rect 351004 208418 351186 208654
rect 351422 208418 351604 208654
rect 351004 208334 351604 208418
rect 351004 208098 351186 208334
rect 351422 208098 351604 208334
rect 351004 172654 351604 208098
rect 351004 172418 351186 172654
rect 351422 172418 351604 172654
rect 351004 172334 351604 172418
rect 351004 172098 351186 172334
rect 351422 172098 351604 172334
rect 351004 136654 351604 172098
rect 351004 136418 351186 136654
rect 351422 136418 351604 136654
rect 351004 136334 351604 136418
rect 351004 136098 351186 136334
rect 351422 136098 351604 136334
rect 351004 100654 351604 136098
rect 351004 100418 351186 100654
rect 351422 100418 351604 100654
rect 351004 100334 351604 100418
rect 351004 100098 351186 100334
rect 351422 100098 351604 100334
rect 351004 64654 351604 100098
rect 351004 64418 351186 64654
rect 351422 64418 351604 64654
rect 351004 64334 351604 64418
rect 351004 64098 351186 64334
rect 351422 64098 351604 64334
rect 351004 28654 351604 64098
rect 351004 28418 351186 28654
rect 351422 28418 351604 28654
rect 351004 28334 351604 28418
rect 351004 28098 351186 28334
rect 351422 28098 351604 28334
rect 351004 -5046 351604 28098
rect 351004 -5282 351186 -5046
rect 351422 -5282 351604 -5046
rect 351004 -5366 351604 -5282
rect 351004 -5602 351186 -5366
rect 351422 -5602 351604 -5366
rect 351004 -5624 351604 -5602
rect 354604 320254 355204 326000
rect 354604 320018 354786 320254
rect 355022 320018 355204 320254
rect 354604 319934 355204 320018
rect 354604 319698 354786 319934
rect 355022 319698 355204 319934
rect 354604 284254 355204 319698
rect 354604 284018 354786 284254
rect 355022 284018 355204 284254
rect 354604 283934 355204 284018
rect 354604 283698 354786 283934
rect 355022 283698 355204 283934
rect 354604 248254 355204 283698
rect 354604 248018 354786 248254
rect 355022 248018 355204 248254
rect 354604 247934 355204 248018
rect 354604 247698 354786 247934
rect 355022 247698 355204 247934
rect 354604 212254 355204 247698
rect 354604 212018 354786 212254
rect 355022 212018 355204 212254
rect 354604 211934 355204 212018
rect 354604 211698 354786 211934
rect 355022 211698 355204 211934
rect 354604 176254 355204 211698
rect 354604 176018 354786 176254
rect 355022 176018 355204 176254
rect 354604 175934 355204 176018
rect 354604 175698 354786 175934
rect 355022 175698 355204 175934
rect 354604 140254 355204 175698
rect 354604 140018 354786 140254
rect 355022 140018 355204 140254
rect 354604 139934 355204 140018
rect 354604 139698 354786 139934
rect 355022 139698 355204 139934
rect 354604 104254 355204 139698
rect 354604 104018 354786 104254
rect 355022 104018 355204 104254
rect 354604 103934 355204 104018
rect 354604 103698 354786 103934
rect 355022 103698 355204 103934
rect 354604 68254 355204 103698
rect 354604 68018 354786 68254
rect 355022 68018 355204 68254
rect 354604 67934 355204 68018
rect 354604 67698 354786 67934
rect 355022 67698 355204 67934
rect 354604 32254 355204 67698
rect 354604 32018 354786 32254
rect 355022 32018 355204 32254
rect 354604 31934 355204 32018
rect 354604 31698 354786 31934
rect 355022 31698 355204 31934
rect 336604 -6222 336786 -5986
rect 337022 -6222 337204 -5986
rect 336604 -6306 337204 -6222
rect 336604 -6542 336786 -6306
rect 337022 -6542 337204 -6306
rect 336604 -7504 337204 -6542
rect 354604 -6926 355204 31698
rect 361804 291454 362404 326000
rect 361804 291218 361986 291454
rect 362222 291218 362404 291454
rect 361804 291134 362404 291218
rect 361804 290898 361986 291134
rect 362222 290898 362404 291134
rect 361804 255454 362404 290898
rect 361804 255218 361986 255454
rect 362222 255218 362404 255454
rect 361804 255134 362404 255218
rect 361804 254898 361986 255134
rect 362222 254898 362404 255134
rect 361804 219454 362404 254898
rect 361804 219218 361986 219454
rect 362222 219218 362404 219454
rect 361804 219134 362404 219218
rect 361804 218898 361986 219134
rect 362222 218898 362404 219134
rect 361804 183454 362404 218898
rect 361804 183218 361986 183454
rect 362222 183218 362404 183454
rect 361804 183134 362404 183218
rect 361804 182898 361986 183134
rect 362222 182898 362404 183134
rect 361804 147454 362404 182898
rect 361804 147218 361986 147454
rect 362222 147218 362404 147454
rect 361804 147134 362404 147218
rect 361804 146898 361986 147134
rect 362222 146898 362404 147134
rect 361804 111454 362404 146898
rect 361804 111218 361986 111454
rect 362222 111218 362404 111454
rect 361804 111134 362404 111218
rect 361804 110898 361986 111134
rect 362222 110898 362404 111134
rect 361804 75454 362404 110898
rect 361804 75218 361986 75454
rect 362222 75218 362404 75454
rect 361804 75134 362404 75218
rect 361804 74898 361986 75134
rect 362222 74898 362404 75134
rect 361804 39454 362404 74898
rect 361804 39218 361986 39454
rect 362222 39218 362404 39454
rect 361804 39134 362404 39218
rect 361804 38898 361986 39134
rect 362222 38898 362404 39134
rect 361804 3454 362404 38898
rect 361804 3218 361986 3454
rect 362222 3218 362404 3454
rect 361804 3134 362404 3218
rect 361804 2898 361986 3134
rect 362222 2898 362404 3134
rect 361804 -346 362404 2898
rect 361804 -582 361986 -346
rect 362222 -582 362404 -346
rect 361804 -666 362404 -582
rect 361804 -902 361986 -666
rect 362222 -902 362404 -666
rect 361804 -1864 362404 -902
rect 365404 295054 366004 326000
rect 365404 294818 365586 295054
rect 365822 294818 366004 295054
rect 365404 294734 366004 294818
rect 365404 294498 365586 294734
rect 365822 294498 366004 294734
rect 365404 259054 366004 294498
rect 365404 258818 365586 259054
rect 365822 258818 366004 259054
rect 365404 258734 366004 258818
rect 365404 258498 365586 258734
rect 365822 258498 366004 258734
rect 365404 223054 366004 258498
rect 365404 222818 365586 223054
rect 365822 222818 366004 223054
rect 365404 222734 366004 222818
rect 365404 222498 365586 222734
rect 365822 222498 366004 222734
rect 365404 187054 366004 222498
rect 365404 186818 365586 187054
rect 365822 186818 366004 187054
rect 365404 186734 366004 186818
rect 365404 186498 365586 186734
rect 365822 186498 366004 186734
rect 365404 151054 366004 186498
rect 365404 150818 365586 151054
rect 365822 150818 366004 151054
rect 365404 150734 366004 150818
rect 365404 150498 365586 150734
rect 365822 150498 366004 150734
rect 365404 115054 366004 150498
rect 365404 114818 365586 115054
rect 365822 114818 366004 115054
rect 365404 114734 366004 114818
rect 365404 114498 365586 114734
rect 365822 114498 366004 114734
rect 365404 79054 366004 114498
rect 365404 78818 365586 79054
rect 365822 78818 366004 79054
rect 365404 78734 366004 78818
rect 365404 78498 365586 78734
rect 365822 78498 366004 78734
rect 365404 43054 366004 78498
rect 365404 42818 365586 43054
rect 365822 42818 366004 43054
rect 365404 42734 366004 42818
rect 365404 42498 365586 42734
rect 365822 42498 366004 42734
rect 365404 7054 366004 42498
rect 365404 6818 365586 7054
rect 365822 6818 366004 7054
rect 365404 6734 366004 6818
rect 365404 6498 365586 6734
rect 365822 6498 366004 6734
rect 365404 -2226 366004 6498
rect 365404 -2462 365586 -2226
rect 365822 -2462 366004 -2226
rect 365404 -2546 366004 -2462
rect 365404 -2782 365586 -2546
rect 365822 -2782 366004 -2546
rect 365404 -3744 366004 -2782
rect 369004 298654 369604 326000
rect 369004 298418 369186 298654
rect 369422 298418 369604 298654
rect 369004 298334 369604 298418
rect 369004 298098 369186 298334
rect 369422 298098 369604 298334
rect 369004 262654 369604 298098
rect 369004 262418 369186 262654
rect 369422 262418 369604 262654
rect 369004 262334 369604 262418
rect 369004 262098 369186 262334
rect 369422 262098 369604 262334
rect 369004 226654 369604 262098
rect 369004 226418 369186 226654
rect 369422 226418 369604 226654
rect 369004 226334 369604 226418
rect 369004 226098 369186 226334
rect 369422 226098 369604 226334
rect 369004 190654 369604 226098
rect 369004 190418 369186 190654
rect 369422 190418 369604 190654
rect 369004 190334 369604 190418
rect 369004 190098 369186 190334
rect 369422 190098 369604 190334
rect 369004 154654 369604 190098
rect 369004 154418 369186 154654
rect 369422 154418 369604 154654
rect 369004 154334 369604 154418
rect 369004 154098 369186 154334
rect 369422 154098 369604 154334
rect 369004 118654 369604 154098
rect 369004 118418 369186 118654
rect 369422 118418 369604 118654
rect 369004 118334 369604 118418
rect 369004 118098 369186 118334
rect 369422 118098 369604 118334
rect 369004 82654 369604 118098
rect 369004 82418 369186 82654
rect 369422 82418 369604 82654
rect 369004 82334 369604 82418
rect 369004 82098 369186 82334
rect 369422 82098 369604 82334
rect 369004 46654 369604 82098
rect 369004 46418 369186 46654
rect 369422 46418 369604 46654
rect 369004 46334 369604 46418
rect 369004 46098 369186 46334
rect 369422 46098 369604 46334
rect 369004 10654 369604 46098
rect 369004 10418 369186 10654
rect 369422 10418 369604 10654
rect 369004 10334 369604 10418
rect 369004 10098 369186 10334
rect 369422 10098 369604 10334
rect 369004 -4106 369604 10098
rect 369004 -4342 369186 -4106
rect 369422 -4342 369604 -4106
rect 369004 -4426 369604 -4342
rect 369004 -4662 369186 -4426
rect 369422 -4662 369604 -4426
rect 369004 -5624 369604 -4662
rect 372604 302254 373204 326000
rect 372604 302018 372786 302254
rect 373022 302018 373204 302254
rect 372604 301934 373204 302018
rect 372604 301698 372786 301934
rect 373022 301698 373204 301934
rect 372604 266254 373204 301698
rect 372604 266018 372786 266254
rect 373022 266018 373204 266254
rect 372604 265934 373204 266018
rect 372604 265698 372786 265934
rect 373022 265698 373204 265934
rect 372604 230254 373204 265698
rect 372604 230018 372786 230254
rect 373022 230018 373204 230254
rect 372604 229934 373204 230018
rect 372604 229698 372786 229934
rect 373022 229698 373204 229934
rect 372604 194254 373204 229698
rect 372604 194018 372786 194254
rect 373022 194018 373204 194254
rect 372604 193934 373204 194018
rect 372604 193698 372786 193934
rect 373022 193698 373204 193934
rect 372604 158254 373204 193698
rect 372604 158018 372786 158254
rect 373022 158018 373204 158254
rect 372604 157934 373204 158018
rect 372604 157698 372786 157934
rect 373022 157698 373204 157934
rect 372604 122254 373204 157698
rect 372604 122018 372786 122254
rect 373022 122018 373204 122254
rect 372604 121934 373204 122018
rect 372604 121698 372786 121934
rect 373022 121698 373204 121934
rect 372604 86254 373204 121698
rect 372604 86018 372786 86254
rect 373022 86018 373204 86254
rect 372604 85934 373204 86018
rect 372604 85698 372786 85934
rect 373022 85698 373204 85934
rect 372604 50254 373204 85698
rect 372604 50018 372786 50254
rect 373022 50018 373204 50254
rect 372604 49934 373204 50018
rect 372604 49698 372786 49934
rect 373022 49698 373204 49934
rect 372604 14254 373204 49698
rect 372604 14018 372786 14254
rect 373022 14018 373204 14254
rect 372604 13934 373204 14018
rect 372604 13698 372786 13934
rect 373022 13698 373204 13934
rect 354604 -7162 354786 -6926
rect 355022 -7162 355204 -6926
rect 354604 -7246 355204 -7162
rect 354604 -7482 354786 -7246
rect 355022 -7482 355204 -7246
rect 354604 -7504 355204 -7482
rect 372604 -5986 373204 13698
rect 379804 309454 380404 326000
rect 379804 309218 379986 309454
rect 380222 309218 380404 309454
rect 379804 309134 380404 309218
rect 379804 308898 379986 309134
rect 380222 308898 380404 309134
rect 379804 273454 380404 308898
rect 379804 273218 379986 273454
rect 380222 273218 380404 273454
rect 379804 273134 380404 273218
rect 379804 272898 379986 273134
rect 380222 272898 380404 273134
rect 379804 237454 380404 272898
rect 379804 237218 379986 237454
rect 380222 237218 380404 237454
rect 379804 237134 380404 237218
rect 379804 236898 379986 237134
rect 380222 236898 380404 237134
rect 379804 201454 380404 236898
rect 379804 201218 379986 201454
rect 380222 201218 380404 201454
rect 379804 201134 380404 201218
rect 379804 200898 379986 201134
rect 380222 200898 380404 201134
rect 379804 165454 380404 200898
rect 379804 165218 379986 165454
rect 380222 165218 380404 165454
rect 379804 165134 380404 165218
rect 379804 164898 379986 165134
rect 380222 164898 380404 165134
rect 379804 129454 380404 164898
rect 379804 129218 379986 129454
rect 380222 129218 380404 129454
rect 379804 129134 380404 129218
rect 379804 128898 379986 129134
rect 380222 128898 380404 129134
rect 379804 93454 380404 128898
rect 379804 93218 379986 93454
rect 380222 93218 380404 93454
rect 379804 93134 380404 93218
rect 379804 92898 379986 93134
rect 380222 92898 380404 93134
rect 379804 57454 380404 92898
rect 379804 57218 379986 57454
rect 380222 57218 380404 57454
rect 379804 57134 380404 57218
rect 379804 56898 379986 57134
rect 380222 56898 380404 57134
rect 379804 21454 380404 56898
rect 379804 21218 379986 21454
rect 380222 21218 380404 21454
rect 379804 21134 380404 21218
rect 379804 20898 379986 21134
rect 380222 20898 380404 21134
rect 379804 -1286 380404 20898
rect 379804 -1522 379986 -1286
rect 380222 -1522 380404 -1286
rect 379804 -1606 380404 -1522
rect 379804 -1842 379986 -1606
rect 380222 -1842 380404 -1606
rect 379804 -1864 380404 -1842
rect 383404 313054 384004 326000
rect 383404 312818 383586 313054
rect 383822 312818 384004 313054
rect 383404 312734 384004 312818
rect 383404 312498 383586 312734
rect 383822 312498 384004 312734
rect 383404 277054 384004 312498
rect 383404 276818 383586 277054
rect 383822 276818 384004 277054
rect 383404 276734 384004 276818
rect 383404 276498 383586 276734
rect 383822 276498 384004 276734
rect 383404 241054 384004 276498
rect 383404 240818 383586 241054
rect 383822 240818 384004 241054
rect 383404 240734 384004 240818
rect 383404 240498 383586 240734
rect 383822 240498 384004 240734
rect 383404 205054 384004 240498
rect 383404 204818 383586 205054
rect 383822 204818 384004 205054
rect 383404 204734 384004 204818
rect 383404 204498 383586 204734
rect 383822 204498 384004 204734
rect 383404 169054 384004 204498
rect 383404 168818 383586 169054
rect 383822 168818 384004 169054
rect 383404 168734 384004 168818
rect 383404 168498 383586 168734
rect 383822 168498 384004 168734
rect 383404 133054 384004 168498
rect 383404 132818 383586 133054
rect 383822 132818 384004 133054
rect 383404 132734 384004 132818
rect 383404 132498 383586 132734
rect 383822 132498 384004 132734
rect 383404 97054 384004 132498
rect 383404 96818 383586 97054
rect 383822 96818 384004 97054
rect 383404 96734 384004 96818
rect 383404 96498 383586 96734
rect 383822 96498 384004 96734
rect 383404 61054 384004 96498
rect 383404 60818 383586 61054
rect 383822 60818 384004 61054
rect 383404 60734 384004 60818
rect 383404 60498 383586 60734
rect 383822 60498 384004 60734
rect 383404 25054 384004 60498
rect 383404 24818 383586 25054
rect 383822 24818 384004 25054
rect 383404 24734 384004 24818
rect 383404 24498 383586 24734
rect 383822 24498 384004 24734
rect 383404 -3166 384004 24498
rect 383404 -3402 383586 -3166
rect 383822 -3402 384004 -3166
rect 383404 -3486 384004 -3402
rect 383404 -3722 383586 -3486
rect 383822 -3722 384004 -3486
rect 383404 -3744 384004 -3722
rect 387004 316654 387604 326000
rect 387004 316418 387186 316654
rect 387422 316418 387604 316654
rect 387004 316334 387604 316418
rect 387004 316098 387186 316334
rect 387422 316098 387604 316334
rect 387004 280654 387604 316098
rect 387004 280418 387186 280654
rect 387422 280418 387604 280654
rect 387004 280334 387604 280418
rect 387004 280098 387186 280334
rect 387422 280098 387604 280334
rect 387004 244654 387604 280098
rect 387004 244418 387186 244654
rect 387422 244418 387604 244654
rect 387004 244334 387604 244418
rect 387004 244098 387186 244334
rect 387422 244098 387604 244334
rect 387004 208654 387604 244098
rect 387004 208418 387186 208654
rect 387422 208418 387604 208654
rect 387004 208334 387604 208418
rect 387004 208098 387186 208334
rect 387422 208098 387604 208334
rect 387004 172654 387604 208098
rect 387004 172418 387186 172654
rect 387422 172418 387604 172654
rect 387004 172334 387604 172418
rect 387004 172098 387186 172334
rect 387422 172098 387604 172334
rect 387004 136654 387604 172098
rect 387004 136418 387186 136654
rect 387422 136418 387604 136654
rect 387004 136334 387604 136418
rect 387004 136098 387186 136334
rect 387422 136098 387604 136334
rect 387004 100654 387604 136098
rect 387004 100418 387186 100654
rect 387422 100418 387604 100654
rect 387004 100334 387604 100418
rect 387004 100098 387186 100334
rect 387422 100098 387604 100334
rect 387004 64654 387604 100098
rect 387004 64418 387186 64654
rect 387422 64418 387604 64654
rect 387004 64334 387604 64418
rect 387004 64098 387186 64334
rect 387422 64098 387604 64334
rect 387004 28654 387604 64098
rect 387004 28418 387186 28654
rect 387422 28418 387604 28654
rect 387004 28334 387604 28418
rect 387004 28098 387186 28334
rect 387422 28098 387604 28334
rect 387004 -5046 387604 28098
rect 387004 -5282 387186 -5046
rect 387422 -5282 387604 -5046
rect 387004 -5366 387604 -5282
rect 387004 -5602 387186 -5366
rect 387422 -5602 387604 -5366
rect 387004 -5624 387604 -5602
rect 390604 320254 391204 326000
rect 390604 320018 390786 320254
rect 391022 320018 391204 320254
rect 390604 319934 391204 320018
rect 390604 319698 390786 319934
rect 391022 319698 391204 319934
rect 390604 284254 391204 319698
rect 390604 284018 390786 284254
rect 391022 284018 391204 284254
rect 390604 283934 391204 284018
rect 390604 283698 390786 283934
rect 391022 283698 391204 283934
rect 390604 248254 391204 283698
rect 390604 248018 390786 248254
rect 391022 248018 391204 248254
rect 390604 247934 391204 248018
rect 390604 247698 390786 247934
rect 391022 247698 391204 247934
rect 390604 212254 391204 247698
rect 390604 212018 390786 212254
rect 391022 212018 391204 212254
rect 390604 211934 391204 212018
rect 390604 211698 390786 211934
rect 391022 211698 391204 211934
rect 390604 176254 391204 211698
rect 390604 176018 390786 176254
rect 391022 176018 391204 176254
rect 390604 175934 391204 176018
rect 390604 175698 390786 175934
rect 391022 175698 391204 175934
rect 390604 140254 391204 175698
rect 390604 140018 390786 140254
rect 391022 140018 391204 140254
rect 390604 139934 391204 140018
rect 390604 139698 390786 139934
rect 391022 139698 391204 139934
rect 390604 104254 391204 139698
rect 390604 104018 390786 104254
rect 391022 104018 391204 104254
rect 390604 103934 391204 104018
rect 390604 103698 390786 103934
rect 391022 103698 391204 103934
rect 390604 68254 391204 103698
rect 390604 68018 390786 68254
rect 391022 68018 391204 68254
rect 390604 67934 391204 68018
rect 390604 67698 390786 67934
rect 391022 67698 391204 67934
rect 390604 32254 391204 67698
rect 390604 32018 390786 32254
rect 391022 32018 391204 32254
rect 390604 31934 391204 32018
rect 390604 31698 390786 31934
rect 391022 31698 391204 31934
rect 372604 -6222 372786 -5986
rect 373022 -6222 373204 -5986
rect 372604 -6306 373204 -6222
rect 372604 -6542 372786 -6306
rect 373022 -6542 373204 -6306
rect 372604 -7504 373204 -6542
rect 390604 -6926 391204 31698
rect 397804 291454 398404 326000
rect 397804 291218 397986 291454
rect 398222 291218 398404 291454
rect 397804 291134 398404 291218
rect 397804 290898 397986 291134
rect 398222 290898 398404 291134
rect 397804 255454 398404 290898
rect 397804 255218 397986 255454
rect 398222 255218 398404 255454
rect 397804 255134 398404 255218
rect 397804 254898 397986 255134
rect 398222 254898 398404 255134
rect 397804 219454 398404 254898
rect 397804 219218 397986 219454
rect 398222 219218 398404 219454
rect 397804 219134 398404 219218
rect 397804 218898 397986 219134
rect 398222 218898 398404 219134
rect 397804 183454 398404 218898
rect 397804 183218 397986 183454
rect 398222 183218 398404 183454
rect 397804 183134 398404 183218
rect 397804 182898 397986 183134
rect 398222 182898 398404 183134
rect 397804 147454 398404 182898
rect 397804 147218 397986 147454
rect 398222 147218 398404 147454
rect 397804 147134 398404 147218
rect 397804 146898 397986 147134
rect 398222 146898 398404 147134
rect 397804 111454 398404 146898
rect 397804 111218 397986 111454
rect 398222 111218 398404 111454
rect 397804 111134 398404 111218
rect 397804 110898 397986 111134
rect 398222 110898 398404 111134
rect 397804 75454 398404 110898
rect 397804 75218 397986 75454
rect 398222 75218 398404 75454
rect 397804 75134 398404 75218
rect 397804 74898 397986 75134
rect 398222 74898 398404 75134
rect 397804 39454 398404 74898
rect 397804 39218 397986 39454
rect 398222 39218 398404 39454
rect 397804 39134 398404 39218
rect 397804 38898 397986 39134
rect 398222 38898 398404 39134
rect 397804 3454 398404 38898
rect 397804 3218 397986 3454
rect 398222 3218 398404 3454
rect 397804 3134 398404 3218
rect 397804 2898 397986 3134
rect 398222 2898 398404 3134
rect 397804 -346 398404 2898
rect 397804 -582 397986 -346
rect 398222 -582 398404 -346
rect 397804 -666 398404 -582
rect 397804 -902 397986 -666
rect 398222 -902 398404 -666
rect 397804 -1864 398404 -902
rect 401404 295054 402004 326000
rect 401404 294818 401586 295054
rect 401822 294818 402004 295054
rect 401404 294734 402004 294818
rect 401404 294498 401586 294734
rect 401822 294498 402004 294734
rect 401404 259054 402004 294498
rect 401404 258818 401586 259054
rect 401822 258818 402004 259054
rect 401404 258734 402004 258818
rect 401404 258498 401586 258734
rect 401822 258498 402004 258734
rect 401404 223054 402004 258498
rect 401404 222818 401586 223054
rect 401822 222818 402004 223054
rect 401404 222734 402004 222818
rect 401404 222498 401586 222734
rect 401822 222498 402004 222734
rect 401404 187054 402004 222498
rect 401404 186818 401586 187054
rect 401822 186818 402004 187054
rect 401404 186734 402004 186818
rect 401404 186498 401586 186734
rect 401822 186498 402004 186734
rect 401404 151054 402004 186498
rect 401404 150818 401586 151054
rect 401822 150818 402004 151054
rect 401404 150734 402004 150818
rect 401404 150498 401586 150734
rect 401822 150498 402004 150734
rect 401404 115054 402004 150498
rect 401404 114818 401586 115054
rect 401822 114818 402004 115054
rect 401404 114734 402004 114818
rect 401404 114498 401586 114734
rect 401822 114498 402004 114734
rect 401404 79054 402004 114498
rect 401404 78818 401586 79054
rect 401822 78818 402004 79054
rect 401404 78734 402004 78818
rect 401404 78498 401586 78734
rect 401822 78498 402004 78734
rect 401404 43054 402004 78498
rect 401404 42818 401586 43054
rect 401822 42818 402004 43054
rect 401404 42734 402004 42818
rect 401404 42498 401586 42734
rect 401822 42498 402004 42734
rect 401404 7054 402004 42498
rect 401404 6818 401586 7054
rect 401822 6818 402004 7054
rect 401404 6734 402004 6818
rect 401404 6498 401586 6734
rect 401822 6498 402004 6734
rect 401404 -2226 402004 6498
rect 401404 -2462 401586 -2226
rect 401822 -2462 402004 -2226
rect 401404 -2546 402004 -2462
rect 401404 -2782 401586 -2546
rect 401822 -2782 402004 -2546
rect 401404 -3744 402004 -2782
rect 405004 298654 405604 326000
rect 405004 298418 405186 298654
rect 405422 298418 405604 298654
rect 405004 298334 405604 298418
rect 405004 298098 405186 298334
rect 405422 298098 405604 298334
rect 405004 262654 405604 298098
rect 405004 262418 405186 262654
rect 405422 262418 405604 262654
rect 405004 262334 405604 262418
rect 405004 262098 405186 262334
rect 405422 262098 405604 262334
rect 405004 226654 405604 262098
rect 405004 226418 405186 226654
rect 405422 226418 405604 226654
rect 405004 226334 405604 226418
rect 405004 226098 405186 226334
rect 405422 226098 405604 226334
rect 405004 190654 405604 226098
rect 405004 190418 405186 190654
rect 405422 190418 405604 190654
rect 405004 190334 405604 190418
rect 405004 190098 405186 190334
rect 405422 190098 405604 190334
rect 405004 154654 405604 190098
rect 405004 154418 405186 154654
rect 405422 154418 405604 154654
rect 405004 154334 405604 154418
rect 405004 154098 405186 154334
rect 405422 154098 405604 154334
rect 405004 118654 405604 154098
rect 405004 118418 405186 118654
rect 405422 118418 405604 118654
rect 405004 118334 405604 118418
rect 405004 118098 405186 118334
rect 405422 118098 405604 118334
rect 405004 82654 405604 118098
rect 405004 82418 405186 82654
rect 405422 82418 405604 82654
rect 405004 82334 405604 82418
rect 405004 82098 405186 82334
rect 405422 82098 405604 82334
rect 405004 46654 405604 82098
rect 405004 46418 405186 46654
rect 405422 46418 405604 46654
rect 405004 46334 405604 46418
rect 405004 46098 405186 46334
rect 405422 46098 405604 46334
rect 405004 10654 405604 46098
rect 405004 10418 405186 10654
rect 405422 10418 405604 10654
rect 405004 10334 405604 10418
rect 405004 10098 405186 10334
rect 405422 10098 405604 10334
rect 405004 -4106 405604 10098
rect 405004 -4342 405186 -4106
rect 405422 -4342 405604 -4106
rect 405004 -4426 405604 -4342
rect 405004 -4662 405186 -4426
rect 405422 -4662 405604 -4426
rect 405004 -5624 405604 -4662
rect 408604 302254 409204 326000
rect 408604 302018 408786 302254
rect 409022 302018 409204 302254
rect 408604 301934 409204 302018
rect 408604 301698 408786 301934
rect 409022 301698 409204 301934
rect 408604 266254 409204 301698
rect 408604 266018 408786 266254
rect 409022 266018 409204 266254
rect 408604 265934 409204 266018
rect 408604 265698 408786 265934
rect 409022 265698 409204 265934
rect 408604 230254 409204 265698
rect 408604 230018 408786 230254
rect 409022 230018 409204 230254
rect 408604 229934 409204 230018
rect 408604 229698 408786 229934
rect 409022 229698 409204 229934
rect 408604 194254 409204 229698
rect 408604 194018 408786 194254
rect 409022 194018 409204 194254
rect 408604 193934 409204 194018
rect 408604 193698 408786 193934
rect 409022 193698 409204 193934
rect 408604 158254 409204 193698
rect 408604 158018 408786 158254
rect 409022 158018 409204 158254
rect 408604 157934 409204 158018
rect 408604 157698 408786 157934
rect 409022 157698 409204 157934
rect 408604 122254 409204 157698
rect 408604 122018 408786 122254
rect 409022 122018 409204 122254
rect 408604 121934 409204 122018
rect 408604 121698 408786 121934
rect 409022 121698 409204 121934
rect 408604 86254 409204 121698
rect 408604 86018 408786 86254
rect 409022 86018 409204 86254
rect 408604 85934 409204 86018
rect 408604 85698 408786 85934
rect 409022 85698 409204 85934
rect 408604 50254 409204 85698
rect 408604 50018 408786 50254
rect 409022 50018 409204 50254
rect 408604 49934 409204 50018
rect 408604 49698 408786 49934
rect 409022 49698 409204 49934
rect 408604 14254 409204 49698
rect 408604 14018 408786 14254
rect 409022 14018 409204 14254
rect 408604 13934 409204 14018
rect 408604 13698 408786 13934
rect 409022 13698 409204 13934
rect 390604 -7162 390786 -6926
rect 391022 -7162 391204 -6926
rect 390604 -7246 391204 -7162
rect 390604 -7482 390786 -7246
rect 391022 -7482 391204 -7246
rect 390604 -7504 391204 -7482
rect 408604 -5986 409204 13698
rect 415804 309454 416404 326000
rect 415804 309218 415986 309454
rect 416222 309218 416404 309454
rect 415804 309134 416404 309218
rect 415804 308898 415986 309134
rect 416222 308898 416404 309134
rect 415804 273454 416404 308898
rect 415804 273218 415986 273454
rect 416222 273218 416404 273454
rect 415804 273134 416404 273218
rect 415804 272898 415986 273134
rect 416222 272898 416404 273134
rect 415804 237454 416404 272898
rect 415804 237218 415986 237454
rect 416222 237218 416404 237454
rect 415804 237134 416404 237218
rect 415804 236898 415986 237134
rect 416222 236898 416404 237134
rect 415804 201454 416404 236898
rect 415804 201218 415986 201454
rect 416222 201218 416404 201454
rect 415804 201134 416404 201218
rect 415804 200898 415986 201134
rect 416222 200898 416404 201134
rect 415804 165454 416404 200898
rect 415804 165218 415986 165454
rect 416222 165218 416404 165454
rect 415804 165134 416404 165218
rect 415804 164898 415986 165134
rect 416222 164898 416404 165134
rect 415804 129454 416404 164898
rect 415804 129218 415986 129454
rect 416222 129218 416404 129454
rect 415804 129134 416404 129218
rect 415804 128898 415986 129134
rect 416222 128898 416404 129134
rect 415804 93454 416404 128898
rect 415804 93218 415986 93454
rect 416222 93218 416404 93454
rect 415804 93134 416404 93218
rect 415804 92898 415986 93134
rect 416222 92898 416404 93134
rect 415804 57454 416404 92898
rect 415804 57218 415986 57454
rect 416222 57218 416404 57454
rect 415804 57134 416404 57218
rect 415804 56898 415986 57134
rect 416222 56898 416404 57134
rect 415804 21454 416404 56898
rect 415804 21218 415986 21454
rect 416222 21218 416404 21454
rect 415804 21134 416404 21218
rect 415804 20898 415986 21134
rect 416222 20898 416404 21134
rect 415804 -1286 416404 20898
rect 415804 -1522 415986 -1286
rect 416222 -1522 416404 -1286
rect 415804 -1606 416404 -1522
rect 415804 -1842 415986 -1606
rect 416222 -1842 416404 -1606
rect 415804 -1864 416404 -1842
rect 419404 313054 420004 326000
rect 419404 312818 419586 313054
rect 419822 312818 420004 313054
rect 419404 312734 420004 312818
rect 419404 312498 419586 312734
rect 419822 312498 420004 312734
rect 419404 277054 420004 312498
rect 419404 276818 419586 277054
rect 419822 276818 420004 277054
rect 419404 276734 420004 276818
rect 419404 276498 419586 276734
rect 419822 276498 420004 276734
rect 419404 241054 420004 276498
rect 419404 240818 419586 241054
rect 419822 240818 420004 241054
rect 419404 240734 420004 240818
rect 419404 240498 419586 240734
rect 419822 240498 420004 240734
rect 419404 205054 420004 240498
rect 419404 204818 419586 205054
rect 419822 204818 420004 205054
rect 419404 204734 420004 204818
rect 419404 204498 419586 204734
rect 419822 204498 420004 204734
rect 419404 169054 420004 204498
rect 419404 168818 419586 169054
rect 419822 168818 420004 169054
rect 419404 168734 420004 168818
rect 419404 168498 419586 168734
rect 419822 168498 420004 168734
rect 419404 133054 420004 168498
rect 419404 132818 419586 133054
rect 419822 132818 420004 133054
rect 419404 132734 420004 132818
rect 419404 132498 419586 132734
rect 419822 132498 420004 132734
rect 419404 97054 420004 132498
rect 419404 96818 419586 97054
rect 419822 96818 420004 97054
rect 419404 96734 420004 96818
rect 419404 96498 419586 96734
rect 419822 96498 420004 96734
rect 419404 61054 420004 96498
rect 419404 60818 419586 61054
rect 419822 60818 420004 61054
rect 419404 60734 420004 60818
rect 419404 60498 419586 60734
rect 419822 60498 420004 60734
rect 419404 25054 420004 60498
rect 419404 24818 419586 25054
rect 419822 24818 420004 25054
rect 419404 24734 420004 24818
rect 419404 24498 419586 24734
rect 419822 24498 420004 24734
rect 419404 -3166 420004 24498
rect 419404 -3402 419586 -3166
rect 419822 -3402 420004 -3166
rect 419404 -3486 420004 -3402
rect 419404 -3722 419586 -3486
rect 419822 -3722 420004 -3486
rect 419404 -3744 420004 -3722
rect 423004 316654 423604 326000
rect 423004 316418 423186 316654
rect 423422 316418 423604 316654
rect 423004 316334 423604 316418
rect 423004 316098 423186 316334
rect 423422 316098 423604 316334
rect 423004 280654 423604 316098
rect 423004 280418 423186 280654
rect 423422 280418 423604 280654
rect 423004 280334 423604 280418
rect 423004 280098 423186 280334
rect 423422 280098 423604 280334
rect 423004 244654 423604 280098
rect 423004 244418 423186 244654
rect 423422 244418 423604 244654
rect 423004 244334 423604 244418
rect 423004 244098 423186 244334
rect 423422 244098 423604 244334
rect 423004 208654 423604 244098
rect 423004 208418 423186 208654
rect 423422 208418 423604 208654
rect 423004 208334 423604 208418
rect 423004 208098 423186 208334
rect 423422 208098 423604 208334
rect 423004 172654 423604 208098
rect 423004 172418 423186 172654
rect 423422 172418 423604 172654
rect 423004 172334 423604 172418
rect 423004 172098 423186 172334
rect 423422 172098 423604 172334
rect 423004 136654 423604 172098
rect 423004 136418 423186 136654
rect 423422 136418 423604 136654
rect 423004 136334 423604 136418
rect 423004 136098 423186 136334
rect 423422 136098 423604 136334
rect 423004 100654 423604 136098
rect 423004 100418 423186 100654
rect 423422 100418 423604 100654
rect 423004 100334 423604 100418
rect 423004 100098 423186 100334
rect 423422 100098 423604 100334
rect 423004 64654 423604 100098
rect 423004 64418 423186 64654
rect 423422 64418 423604 64654
rect 423004 64334 423604 64418
rect 423004 64098 423186 64334
rect 423422 64098 423604 64334
rect 423004 28654 423604 64098
rect 423004 28418 423186 28654
rect 423422 28418 423604 28654
rect 423004 28334 423604 28418
rect 423004 28098 423186 28334
rect 423422 28098 423604 28334
rect 423004 -5046 423604 28098
rect 423004 -5282 423186 -5046
rect 423422 -5282 423604 -5046
rect 423004 -5366 423604 -5282
rect 423004 -5602 423186 -5366
rect 423422 -5602 423604 -5366
rect 423004 -5624 423604 -5602
rect 426604 320254 427204 326000
rect 426604 320018 426786 320254
rect 427022 320018 427204 320254
rect 426604 319934 427204 320018
rect 426604 319698 426786 319934
rect 427022 319698 427204 319934
rect 426604 284254 427204 319698
rect 426604 284018 426786 284254
rect 427022 284018 427204 284254
rect 426604 283934 427204 284018
rect 426604 283698 426786 283934
rect 427022 283698 427204 283934
rect 426604 248254 427204 283698
rect 426604 248018 426786 248254
rect 427022 248018 427204 248254
rect 426604 247934 427204 248018
rect 426604 247698 426786 247934
rect 427022 247698 427204 247934
rect 426604 212254 427204 247698
rect 426604 212018 426786 212254
rect 427022 212018 427204 212254
rect 426604 211934 427204 212018
rect 426604 211698 426786 211934
rect 427022 211698 427204 211934
rect 426604 176254 427204 211698
rect 426604 176018 426786 176254
rect 427022 176018 427204 176254
rect 426604 175934 427204 176018
rect 426604 175698 426786 175934
rect 427022 175698 427204 175934
rect 426604 140254 427204 175698
rect 426604 140018 426786 140254
rect 427022 140018 427204 140254
rect 426604 139934 427204 140018
rect 426604 139698 426786 139934
rect 427022 139698 427204 139934
rect 426604 104254 427204 139698
rect 426604 104018 426786 104254
rect 427022 104018 427204 104254
rect 426604 103934 427204 104018
rect 426604 103698 426786 103934
rect 427022 103698 427204 103934
rect 426604 68254 427204 103698
rect 426604 68018 426786 68254
rect 427022 68018 427204 68254
rect 426604 67934 427204 68018
rect 426604 67698 426786 67934
rect 427022 67698 427204 67934
rect 426604 32254 427204 67698
rect 426604 32018 426786 32254
rect 427022 32018 427204 32254
rect 426604 31934 427204 32018
rect 426604 31698 426786 31934
rect 427022 31698 427204 31934
rect 408604 -6222 408786 -5986
rect 409022 -6222 409204 -5986
rect 408604 -6306 409204 -6222
rect 408604 -6542 408786 -6306
rect 409022 -6542 409204 -6306
rect 408604 -7504 409204 -6542
rect 426604 -6926 427204 31698
rect 429702 19413 429762 342483
rect 441004 334654 441604 370098
rect 441004 334418 441186 334654
rect 441422 334418 441604 334654
rect 441004 334334 441604 334418
rect 441004 334098 441186 334334
rect 441422 334098 441604 334334
rect 433804 291454 434404 326000
rect 433804 291218 433986 291454
rect 434222 291218 434404 291454
rect 433804 291134 434404 291218
rect 433804 290898 433986 291134
rect 434222 290898 434404 291134
rect 433804 255454 434404 290898
rect 433804 255218 433986 255454
rect 434222 255218 434404 255454
rect 433804 255134 434404 255218
rect 433804 254898 433986 255134
rect 434222 254898 434404 255134
rect 433804 219454 434404 254898
rect 433804 219218 433986 219454
rect 434222 219218 434404 219454
rect 433804 219134 434404 219218
rect 433804 218898 433986 219134
rect 434222 218898 434404 219134
rect 433804 183454 434404 218898
rect 433804 183218 433986 183454
rect 434222 183218 434404 183454
rect 433804 183134 434404 183218
rect 433804 182898 433986 183134
rect 434222 182898 434404 183134
rect 433804 147454 434404 182898
rect 433804 147218 433986 147454
rect 434222 147218 434404 147454
rect 433804 147134 434404 147218
rect 433804 146898 433986 147134
rect 434222 146898 434404 147134
rect 433804 111454 434404 146898
rect 433804 111218 433986 111454
rect 434222 111218 434404 111454
rect 433804 111134 434404 111218
rect 433804 110898 433986 111134
rect 434222 110898 434404 111134
rect 433804 75454 434404 110898
rect 433804 75218 433986 75454
rect 434222 75218 434404 75454
rect 433804 75134 434404 75218
rect 433804 74898 433986 75134
rect 434222 74898 434404 75134
rect 433804 39454 434404 74898
rect 433804 39218 433986 39454
rect 434222 39218 434404 39454
rect 433804 39134 434404 39218
rect 433804 38898 433986 39134
rect 434222 38898 434404 39134
rect 429699 19412 429765 19413
rect 429699 19348 429700 19412
rect 429764 19348 429765 19412
rect 429699 19347 429765 19348
rect 433804 3454 434404 38898
rect 433804 3218 433986 3454
rect 434222 3218 434404 3454
rect 433804 3134 434404 3218
rect 433804 2898 433986 3134
rect 434222 2898 434404 3134
rect 433804 -346 434404 2898
rect 433804 -582 433986 -346
rect 434222 -582 434404 -346
rect 433804 -666 434404 -582
rect 433804 -902 433986 -666
rect 434222 -902 434404 -666
rect 433804 -1864 434404 -902
rect 437404 295054 438004 326000
rect 437404 294818 437586 295054
rect 437822 294818 438004 295054
rect 437404 294734 438004 294818
rect 437404 294498 437586 294734
rect 437822 294498 438004 294734
rect 437404 259054 438004 294498
rect 437404 258818 437586 259054
rect 437822 258818 438004 259054
rect 437404 258734 438004 258818
rect 437404 258498 437586 258734
rect 437822 258498 438004 258734
rect 437404 223054 438004 258498
rect 437404 222818 437586 223054
rect 437822 222818 438004 223054
rect 437404 222734 438004 222818
rect 437404 222498 437586 222734
rect 437822 222498 438004 222734
rect 437404 187054 438004 222498
rect 437404 186818 437586 187054
rect 437822 186818 438004 187054
rect 437404 186734 438004 186818
rect 437404 186498 437586 186734
rect 437822 186498 438004 186734
rect 437404 151054 438004 186498
rect 437404 150818 437586 151054
rect 437822 150818 438004 151054
rect 437404 150734 438004 150818
rect 437404 150498 437586 150734
rect 437822 150498 438004 150734
rect 437404 115054 438004 150498
rect 437404 114818 437586 115054
rect 437822 114818 438004 115054
rect 437404 114734 438004 114818
rect 437404 114498 437586 114734
rect 437822 114498 438004 114734
rect 437404 79054 438004 114498
rect 437404 78818 437586 79054
rect 437822 78818 438004 79054
rect 437404 78734 438004 78818
rect 437404 78498 437586 78734
rect 437822 78498 438004 78734
rect 437404 43054 438004 78498
rect 437404 42818 437586 43054
rect 437822 42818 438004 43054
rect 437404 42734 438004 42818
rect 437404 42498 437586 42734
rect 437822 42498 438004 42734
rect 437404 7054 438004 42498
rect 437404 6818 437586 7054
rect 437822 6818 438004 7054
rect 437404 6734 438004 6818
rect 437404 6498 437586 6734
rect 437822 6498 438004 6734
rect 437404 -2226 438004 6498
rect 437404 -2462 437586 -2226
rect 437822 -2462 438004 -2226
rect 437404 -2546 438004 -2462
rect 437404 -2782 437586 -2546
rect 437822 -2782 438004 -2546
rect 437404 -3744 438004 -2782
rect 441004 298654 441604 334098
rect 441004 298418 441186 298654
rect 441422 298418 441604 298654
rect 441004 298334 441604 298418
rect 441004 298098 441186 298334
rect 441422 298098 441604 298334
rect 441004 262654 441604 298098
rect 441004 262418 441186 262654
rect 441422 262418 441604 262654
rect 441004 262334 441604 262418
rect 441004 262098 441186 262334
rect 441422 262098 441604 262334
rect 441004 226654 441604 262098
rect 441004 226418 441186 226654
rect 441422 226418 441604 226654
rect 441004 226334 441604 226418
rect 441004 226098 441186 226334
rect 441422 226098 441604 226334
rect 441004 190654 441604 226098
rect 441004 190418 441186 190654
rect 441422 190418 441604 190654
rect 441004 190334 441604 190418
rect 441004 190098 441186 190334
rect 441422 190098 441604 190334
rect 441004 154654 441604 190098
rect 441004 154418 441186 154654
rect 441422 154418 441604 154654
rect 441004 154334 441604 154418
rect 441004 154098 441186 154334
rect 441422 154098 441604 154334
rect 441004 118654 441604 154098
rect 441004 118418 441186 118654
rect 441422 118418 441604 118654
rect 441004 118334 441604 118418
rect 441004 118098 441186 118334
rect 441422 118098 441604 118334
rect 441004 82654 441604 118098
rect 441004 82418 441186 82654
rect 441422 82418 441604 82654
rect 441004 82334 441604 82418
rect 441004 82098 441186 82334
rect 441422 82098 441604 82334
rect 441004 46654 441604 82098
rect 441004 46418 441186 46654
rect 441422 46418 441604 46654
rect 441004 46334 441604 46418
rect 441004 46098 441186 46334
rect 441422 46098 441604 46334
rect 441004 10654 441604 46098
rect 441004 10418 441186 10654
rect 441422 10418 441604 10654
rect 441004 10334 441604 10418
rect 441004 10098 441186 10334
rect 441422 10098 441604 10334
rect 441004 -4106 441604 10098
rect 441004 -4342 441186 -4106
rect 441422 -4342 441604 -4106
rect 441004 -4426 441604 -4342
rect 441004 -4662 441186 -4426
rect 441422 -4662 441604 -4426
rect 441004 -5624 441604 -4662
rect 444604 698254 445204 709922
rect 462604 711418 463204 711440
rect 462604 711182 462786 711418
rect 463022 711182 463204 711418
rect 462604 711098 463204 711182
rect 462604 710862 462786 711098
rect 463022 710862 463204 711098
rect 459004 709538 459604 709560
rect 459004 709302 459186 709538
rect 459422 709302 459604 709538
rect 459004 709218 459604 709302
rect 459004 708982 459186 709218
rect 459422 708982 459604 709218
rect 455404 707658 456004 707680
rect 455404 707422 455586 707658
rect 455822 707422 456004 707658
rect 455404 707338 456004 707422
rect 455404 707102 455586 707338
rect 455822 707102 456004 707338
rect 444604 698018 444786 698254
rect 445022 698018 445204 698254
rect 444604 697934 445204 698018
rect 444604 697698 444786 697934
rect 445022 697698 445204 697934
rect 444604 662254 445204 697698
rect 444604 662018 444786 662254
rect 445022 662018 445204 662254
rect 444604 661934 445204 662018
rect 444604 661698 444786 661934
rect 445022 661698 445204 661934
rect 444604 626254 445204 661698
rect 444604 626018 444786 626254
rect 445022 626018 445204 626254
rect 444604 625934 445204 626018
rect 444604 625698 444786 625934
rect 445022 625698 445204 625934
rect 444604 590254 445204 625698
rect 444604 590018 444786 590254
rect 445022 590018 445204 590254
rect 444604 589934 445204 590018
rect 444604 589698 444786 589934
rect 445022 589698 445204 589934
rect 444604 554254 445204 589698
rect 444604 554018 444786 554254
rect 445022 554018 445204 554254
rect 444604 553934 445204 554018
rect 444604 553698 444786 553934
rect 445022 553698 445204 553934
rect 444604 518254 445204 553698
rect 444604 518018 444786 518254
rect 445022 518018 445204 518254
rect 444604 517934 445204 518018
rect 444604 517698 444786 517934
rect 445022 517698 445204 517934
rect 444604 482254 445204 517698
rect 444604 482018 444786 482254
rect 445022 482018 445204 482254
rect 444604 481934 445204 482018
rect 444604 481698 444786 481934
rect 445022 481698 445204 481934
rect 444604 446254 445204 481698
rect 444604 446018 444786 446254
rect 445022 446018 445204 446254
rect 444604 445934 445204 446018
rect 444604 445698 444786 445934
rect 445022 445698 445204 445934
rect 444604 410254 445204 445698
rect 444604 410018 444786 410254
rect 445022 410018 445204 410254
rect 444604 409934 445204 410018
rect 444604 409698 444786 409934
rect 445022 409698 445204 409934
rect 444604 374254 445204 409698
rect 444604 374018 444786 374254
rect 445022 374018 445204 374254
rect 444604 373934 445204 374018
rect 444604 373698 444786 373934
rect 445022 373698 445204 373934
rect 444604 338254 445204 373698
rect 444604 338018 444786 338254
rect 445022 338018 445204 338254
rect 444604 337934 445204 338018
rect 444604 337698 444786 337934
rect 445022 337698 445204 337934
rect 444604 302254 445204 337698
rect 444604 302018 444786 302254
rect 445022 302018 445204 302254
rect 444604 301934 445204 302018
rect 444604 301698 444786 301934
rect 445022 301698 445204 301934
rect 444604 266254 445204 301698
rect 444604 266018 444786 266254
rect 445022 266018 445204 266254
rect 444604 265934 445204 266018
rect 444604 265698 444786 265934
rect 445022 265698 445204 265934
rect 444604 230254 445204 265698
rect 444604 230018 444786 230254
rect 445022 230018 445204 230254
rect 444604 229934 445204 230018
rect 444604 229698 444786 229934
rect 445022 229698 445204 229934
rect 444604 194254 445204 229698
rect 444604 194018 444786 194254
rect 445022 194018 445204 194254
rect 444604 193934 445204 194018
rect 444604 193698 444786 193934
rect 445022 193698 445204 193934
rect 444604 158254 445204 193698
rect 444604 158018 444786 158254
rect 445022 158018 445204 158254
rect 444604 157934 445204 158018
rect 444604 157698 444786 157934
rect 445022 157698 445204 157934
rect 444604 122254 445204 157698
rect 444604 122018 444786 122254
rect 445022 122018 445204 122254
rect 444604 121934 445204 122018
rect 444604 121698 444786 121934
rect 445022 121698 445204 121934
rect 444604 86254 445204 121698
rect 444604 86018 444786 86254
rect 445022 86018 445204 86254
rect 444604 85934 445204 86018
rect 444604 85698 444786 85934
rect 445022 85698 445204 85934
rect 444604 50254 445204 85698
rect 444604 50018 444786 50254
rect 445022 50018 445204 50254
rect 444604 49934 445204 50018
rect 444604 49698 444786 49934
rect 445022 49698 445204 49934
rect 444604 14254 445204 49698
rect 444604 14018 444786 14254
rect 445022 14018 445204 14254
rect 444604 13934 445204 14018
rect 444604 13698 444786 13934
rect 445022 13698 445204 13934
rect 426604 -7162 426786 -6926
rect 427022 -7162 427204 -6926
rect 426604 -7246 427204 -7162
rect 426604 -7482 426786 -7246
rect 427022 -7482 427204 -7246
rect 426604 -7504 427204 -7482
rect 444604 -5986 445204 13698
rect 451804 705778 452404 705800
rect 451804 705542 451986 705778
rect 452222 705542 452404 705778
rect 451804 705458 452404 705542
rect 451804 705222 451986 705458
rect 452222 705222 452404 705458
rect 451804 669454 452404 705222
rect 451804 669218 451986 669454
rect 452222 669218 452404 669454
rect 451804 669134 452404 669218
rect 451804 668898 451986 669134
rect 452222 668898 452404 669134
rect 451804 633454 452404 668898
rect 451804 633218 451986 633454
rect 452222 633218 452404 633454
rect 451804 633134 452404 633218
rect 451804 632898 451986 633134
rect 452222 632898 452404 633134
rect 451804 597454 452404 632898
rect 451804 597218 451986 597454
rect 452222 597218 452404 597454
rect 451804 597134 452404 597218
rect 451804 596898 451986 597134
rect 452222 596898 452404 597134
rect 451804 561454 452404 596898
rect 451804 561218 451986 561454
rect 452222 561218 452404 561454
rect 451804 561134 452404 561218
rect 451804 560898 451986 561134
rect 452222 560898 452404 561134
rect 451804 525454 452404 560898
rect 451804 525218 451986 525454
rect 452222 525218 452404 525454
rect 451804 525134 452404 525218
rect 451804 524898 451986 525134
rect 452222 524898 452404 525134
rect 451804 489454 452404 524898
rect 451804 489218 451986 489454
rect 452222 489218 452404 489454
rect 451804 489134 452404 489218
rect 451804 488898 451986 489134
rect 452222 488898 452404 489134
rect 451804 453454 452404 488898
rect 451804 453218 451986 453454
rect 452222 453218 452404 453454
rect 451804 453134 452404 453218
rect 451804 452898 451986 453134
rect 452222 452898 452404 453134
rect 451804 417454 452404 452898
rect 451804 417218 451986 417454
rect 452222 417218 452404 417454
rect 451804 417134 452404 417218
rect 451804 416898 451986 417134
rect 452222 416898 452404 417134
rect 451804 381454 452404 416898
rect 451804 381218 451986 381454
rect 452222 381218 452404 381454
rect 451804 381134 452404 381218
rect 451804 380898 451986 381134
rect 452222 380898 452404 381134
rect 451804 345454 452404 380898
rect 451804 345218 451986 345454
rect 452222 345218 452404 345454
rect 451804 345134 452404 345218
rect 451804 344898 451986 345134
rect 452222 344898 452404 345134
rect 451804 309454 452404 344898
rect 451804 309218 451986 309454
rect 452222 309218 452404 309454
rect 451804 309134 452404 309218
rect 451804 308898 451986 309134
rect 452222 308898 452404 309134
rect 451804 273454 452404 308898
rect 451804 273218 451986 273454
rect 452222 273218 452404 273454
rect 451804 273134 452404 273218
rect 451804 272898 451986 273134
rect 452222 272898 452404 273134
rect 451804 237454 452404 272898
rect 451804 237218 451986 237454
rect 452222 237218 452404 237454
rect 451804 237134 452404 237218
rect 451804 236898 451986 237134
rect 452222 236898 452404 237134
rect 451804 201454 452404 236898
rect 451804 201218 451986 201454
rect 452222 201218 452404 201454
rect 451804 201134 452404 201218
rect 451804 200898 451986 201134
rect 452222 200898 452404 201134
rect 451804 165454 452404 200898
rect 451804 165218 451986 165454
rect 452222 165218 452404 165454
rect 451804 165134 452404 165218
rect 451804 164898 451986 165134
rect 452222 164898 452404 165134
rect 451804 129454 452404 164898
rect 451804 129218 451986 129454
rect 452222 129218 452404 129454
rect 451804 129134 452404 129218
rect 451804 128898 451986 129134
rect 452222 128898 452404 129134
rect 451804 93454 452404 128898
rect 451804 93218 451986 93454
rect 452222 93218 452404 93454
rect 451804 93134 452404 93218
rect 451804 92898 451986 93134
rect 452222 92898 452404 93134
rect 451804 57454 452404 92898
rect 451804 57218 451986 57454
rect 452222 57218 452404 57454
rect 451804 57134 452404 57218
rect 451804 56898 451986 57134
rect 452222 56898 452404 57134
rect 451804 21454 452404 56898
rect 451804 21218 451986 21454
rect 452222 21218 452404 21454
rect 451804 21134 452404 21218
rect 451804 20898 451986 21134
rect 452222 20898 452404 21134
rect 451804 -1286 452404 20898
rect 451804 -1522 451986 -1286
rect 452222 -1522 452404 -1286
rect 451804 -1606 452404 -1522
rect 451804 -1842 451986 -1606
rect 452222 -1842 452404 -1606
rect 451804 -1864 452404 -1842
rect 455404 673054 456004 707102
rect 455404 672818 455586 673054
rect 455822 672818 456004 673054
rect 455404 672734 456004 672818
rect 455404 672498 455586 672734
rect 455822 672498 456004 672734
rect 455404 637054 456004 672498
rect 455404 636818 455586 637054
rect 455822 636818 456004 637054
rect 455404 636734 456004 636818
rect 455404 636498 455586 636734
rect 455822 636498 456004 636734
rect 455404 601054 456004 636498
rect 455404 600818 455586 601054
rect 455822 600818 456004 601054
rect 455404 600734 456004 600818
rect 455404 600498 455586 600734
rect 455822 600498 456004 600734
rect 455404 565054 456004 600498
rect 455404 564818 455586 565054
rect 455822 564818 456004 565054
rect 455404 564734 456004 564818
rect 455404 564498 455586 564734
rect 455822 564498 456004 564734
rect 455404 529054 456004 564498
rect 455404 528818 455586 529054
rect 455822 528818 456004 529054
rect 455404 528734 456004 528818
rect 455404 528498 455586 528734
rect 455822 528498 456004 528734
rect 455404 493054 456004 528498
rect 455404 492818 455586 493054
rect 455822 492818 456004 493054
rect 455404 492734 456004 492818
rect 455404 492498 455586 492734
rect 455822 492498 456004 492734
rect 455404 457054 456004 492498
rect 455404 456818 455586 457054
rect 455822 456818 456004 457054
rect 455404 456734 456004 456818
rect 455404 456498 455586 456734
rect 455822 456498 456004 456734
rect 455404 421054 456004 456498
rect 455404 420818 455586 421054
rect 455822 420818 456004 421054
rect 455404 420734 456004 420818
rect 455404 420498 455586 420734
rect 455822 420498 456004 420734
rect 455404 385054 456004 420498
rect 455404 384818 455586 385054
rect 455822 384818 456004 385054
rect 455404 384734 456004 384818
rect 455404 384498 455586 384734
rect 455822 384498 456004 384734
rect 455404 349054 456004 384498
rect 455404 348818 455586 349054
rect 455822 348818 456004 349054
rect 455404 348734 456004 348818
rect 455404 348498 455586 348734
rect 455822 348498 456004 348734
rect 455404 313054 456004 348498
rect 455404 312818 455586 313054
rect 455822 312818 456004 313054
rect 455404 312734 456004 312818
rect 455404 312498 455586 312734
rect 455822 312498 456004 312734
rect 455404 277054 456004 312498
rect 455404 276818 455586 277054
rect 455822 276818 456004 277054
rect 455404 276734 456004 276818
rect 455404 276498 455586 276734
rect 455822 276498 456004 276734
rect 455404 241054 456004 276498
rect 455404 240818 455586 241054
rect 455822 240818 456004 241054
rect 455404 240734 456004 240818
rect 455404 240498 455586 240734
rect 455822 240498 456004 240734
rect 455404 205054 456004 240498
rect 455404 204818 455586 205054
rect 455822 204818 456004 205054
rect 455404 204734 456004 204818
rect 455404 204498 455586 204734
rect 455822 204498 456004 204734
rect 455404 169054 456004 204498
rect 455404 168818 455586 169054
rect 455822 168818 456004 169054
rect 455404 168734 456004 168818
rect 455404 168498 455586 168734
rect 455822 168498 456004 168734
rect 455404 133054 456004 168498
rect 455404 132818 455586 133054
rect 455822 132818 456004 133054
rect 455404 132734 456004 132818
rect 455404 132498 455586 132734
rect 455822 132498 456004 132734
rect 455404 97054 456004 132498
rect 455404 96818 455586 97054
rect 455822 96818 456004 97054
rect 455404 96734 456004 96818
rect 455404 96498 455586 96734
rect 455822 96498 456004 96734
rect 455404 61054 456004 96498
rect 455404 60818 455586 61054
rect 455822 60818 456004 61054
rect 455404 60734 456004 60818
rect 455404 60498 455586 60734
rect 455822 60498 456004 60734
rect 455404 25054 456004 60498
rect 455404 24818 455586 25054
rect 455822 24818 456004 25054
rect 455404 24734 456004 24818
rect 455404 24498 455586 24734
rect 455822 24498 456004 24734
rect 455404 -3166 456004 24498
rect 455404 -3402 455586 -3166
rect 455822 -3402 456004 -3166
rect 455404 -3486 456004 -3402
rect 455404 -3722 455586 -3486
rect 455822 -3722 456004 -3486
rect 455404 -3744 456004 -3722
rect 459004 676654 459604 708982
rect 459004 676418 459186 676654
rect 459422 676418 459604 676654
rect 459004 676334 459604 676418
rect 459004 676098 459186 676334
rect 459422 676098 459604 676334
rect 459004 640654 459604 676098
rect 459004 640418 459186 640654
rect 459422 640418 459604 640654
rect 459004 640334 459604 640418
rect 459004 640098 459186 640334
rect 459422 640098 459604 640334
rect 459004 604654 459604 640098
rect 459004 604418 459186 604654
rect 459422 604418 459604 604654
rect 459004 604334 459604 604418
rect 459004 604098 459186 604334
rect 459422 604098 459604 604334
rect 459004 568654 459604 604098
rect 459004 568418 459186 568654
rect 459422 568418 459604 568654
rect 459004 568334 459604 568418
rect 459004 568098 459186 568334
rect 459422 568098 459604 568334
rect 459004 532654 459604 568098
rect 459004 532418 459186 532654
rect 459422 532418 459604 532654
rect 459004 532334 459604 532418
rect 459004 532098 459186 532334
rect 459422 532098 459604 532334
rect 459004 496654 459604 532098
rect 459004 496418 459186 496654
rect 459422 496418 459604 496654
rect 459004 496334 459604 496418
rect 459004 496098 459186 496334
rect 459422 496098 459604 496334
rect 459004 460654 459604 496098
rect 459004 460418 459186 460654
rect 459422 460418 459604 460654
rect 459004 460334 459604 460418
rect 459004 460098 459186 460334
rect 459422 460098 459604 460334
rect 459004 424654 459604 460098
rect 459004 424418 459186 424654
rect 459422 424418 459604 424654
rect 459004 424334 459604 424418
rect 459004 424098 459186 424334
rect 459422 424098 459604 424334
rect 459004 388654 459604 424098
rect 459004 388418 459186 388654
rect 459422 388418 459604 388654
rect 459004 388334 459604 388418
rect 459004 388098 459186 388334
rect 459422 388098 459604 388334
rect 459004 352654 459604 388098
rect 459004 352418 459186 352654
rect 459422 352418 459604 352654
rect 459004 352334 459604 352418
rect 459004 352098 459186 352334
rect 459422 352098 459604 352334
rect 459004 316654 459604 352098
rect 459004 316418 459186 316654
rect 459422 316418 459604 316654
rect 459004 316334 459604 316418
rect 459004 316098 459186 316334
rect 459422 316098 459604 316334
rect 459004 280654 459604 316098
rect 459004 280418 459186 280654
rect 459422 280418 459604 280654
rect 459004 280334 459604 280418
rect 459004 280098 459186 280334
rect 459422 280098 459604 280334
rect 459004 244654 459604 280098
rect 459004 244418 459186 244654
rect 459422 244418 459604 244654
rect 459004 244334 459604 244418
rect 459004 244098 459186 244334
rect 459422 244098 459604 244334
rect 459004 208654 459604 244098
rect 459004 208418 459186 208654
rect 459422 208418 459604 208654
rect 459004 208334 459604 208418
rect 459004 208098 459186 208334
rect 459422 208098 459604 208334
rect 459004 172654 459604 208098
rect 459004 172418 459186 172654
rect 459422 172418 459604 172654
rect 459004 172334 459604 172418
rect 459004 172098 459186 172334
rect 459422 172098 459604 172334
rect 459004 136654 459604 172098
rect 459004 136418 459186 136654
rect 459422 136418 459604 136654
rect 459004 136334 459604 136418
rect 459004 136098 459186 136334
rect 459422 136098 459604 136334
rect 459004 100654 459604 136098
rect 459004 100418 459186 100654
rect 459422 100418 459604 100654
rect 459004 100334 459604 100418
rect 459004 100098 459186 100334
rect 459422 100098 459604 100334
rect 459004 64654 459604 100098
rect 459004 64418 459186 64654
rect 459422 64418 459604 64654
rect 459004 64334 459604 64418
rect 459004 64098 459186 64334
rect 459422 64098 459604 64334
rect 459004 28654 459604 64098
rect 459004 28418 459186 28654
rect 459422 28418 459604 28654
rect 459004 28334 459604 28418
rect 459004 28098 459186 28334
rect 459422 28098 459604 28334
rect 459004 -5046 459604 28098
rect 459004 -5282 459186 -5046
rect 459422 -5282 459604 -5046
rect 459004 -5366 459604 -5282
rect 459004 -5602 459186 -5366
rect 459422 -5602 459604 -5366
rect 459004 -5624 459604 -5602
rect 462604 680254 463204 710862
rect 480604 710478 481204 711440
rect 480604 710242 480786 710478
rect 481022 710242 481204 710478
rect 480604 710158 481204 710242
rect 480604 709922 480786 710158
rect 481022 709922 481204 710158
rect 477004 708598 477604 709560
rect 477004 708362 477186 708598
rect 477422 708362 477604 708598
rect 477004 708278 477604 708362
rect 477004 708042 477186 708278
rect 477422 708042 477604 708278
rect 473404 706718 474004 707680
rect 473404 706482 473586 706718
rect 473822 706482 474004 706718
rect 473404 706398 474004 706482
rect 473404 706162 473586 706398
rect 473822 706162 474004 706398
rect 462604 680018 462786 680254
rect 463022 680018 463204 680254
rect 462604 679934 463204 680018
rect 462604 679698 462786 679934
rect 463022 679698 463204 679934
rect 462604 644254 463204 679698
rect 462604 644018 462786 644254
rect 463022 644018 463204 644254
rect 462604 643934 463204 644018
rect 462604 643698 462786 643934
rect 463022 643698 463204 643934
rect 462604 608254 463204 643698
rect 462604 608018 462786 608254
rect 463022 608018 463204 608254
rect 462604 607934 463204 608018
rect 462604 607698 462786 607934
rect 463022 607698 463204 607934
rect 462604 572254 463204 607698
rect 462604 572018 462786 572254
rect 463022 572018 463204 572254
rect 462604 571934 463204 572018
rect 462604 571698 462786 571934
rect 463022 571698 463204 571934
rect 462604 536254 463204 571698
rect 462604 536018 462786 536254
rect 463022 536018 463204 536254
rect 462604 535934 463204 536018
rect 462604 535698 462786 535934
rect 463022 535698 463204 535934
rect 462604 500254 463204 535698
rect 462604 500018 462786 500254
rect 463022 500018 463204 500254
rect 462604 499934 463204 500018
rect 462604 499698 462786 499934
rect 463022 499698 463204 499934
rect 462604 464254 463204 499698
rect 462604 464018 462786 464254
rect 463022 464018 463204 464254
rect 462604 463934 463204 464018
rect 462604 463698 462786 463934
rect 463022 463698 463204 463934
rect 462604 428254 463204 463698
rect 462604 428018 462786 428254
rect 463022 428018 463204 428254
rect 462604 427934 463204 428018
rect 462604 427698 462786 427934
rect 463022 427698 463204 427934
rect 462604 392254 463204 427698
rect 462604 392018 462786 392254
rect 463022 392018 463204 392254
rect 462604 391934 463204 392018
rect 462604 391698 462786 391934
rect 463022 391698 463204 391934
rect 462604 356254 463204 391698
rect 462604 356018 462786 356254
rect 463022 356018 463204 356254
rect 462604 355934 463204 356018
rect 462604 355698 462786 355934
rect 463022 355698 463204 355934
rect 462604 320254 463204 355698
rect 462604 320018 462786 320254
rect 463022 320018 463204 320254
rect 462604 319934 463204 320018
rect 462604 319698 462786 319934
rect 463022 319698 463204 319934
rect 462604 284254 463204 319698
rect 462604 284018 462786 284254
rect 463022 284018 463204 284254
rect 462604 283934 463204 284018
rect 462604 283698 462786 283934
rect 463022 283698 463204 283934
rect 462604 248254 463204 283698
rect 462604 248018 462786 248254
rect 463022 248018 463204 248254
rect 462604 247934 463204 248018
rect 462604 247698 462786 247934
rect 463022 247698 463204 247934
rect 462604 212254 463204 247698
rect 462604 212018 462786 212254
rect 463022 212018 463204 212254
rect 462604 211934 463204 212018
rect 462604 211698 462786 211934
rect 463022 211698 463204 211934
rect 462604 176254 463204 211698
rect 462604 176018 462786 176254
rect 463022 176018 463204 176254
rect 462604 175934 463204 176018
rect 462604 175698 462786 175934
rect 463022 175698 463204 175934
rect 462604 140254 463204 175698
rect 462604 140018 462786 140254
rect 463022 140018 463204 140254
rect 462604 139934 463204 140018
rect 462604 139698 462786 139934
rect 463022 139698 463204 139934
rect 462604 104254 463204 139698
rect 462604 104018 462786 104254
rect 463022 104018 463204 104254
rect 462604 103934 463204 104018
rect 462604 103698 462786 103934
rect 463022 103698 463204 103934
rect 462604 68254 463204 103698
rect 462604 68018 462786 68254
rect 463022 68018 463204 68254
rect 462604 67934 463204 68018
rect 462604 67698 462786 67934
rect 463022 67698 463204 67934
rect 462604 32254 463204 67698
rect 462604 32018 462786 32254
rect 463022 32018 463204 32254
rect 462604 31934 463204 32018
rect 462604 31698 462786 31934
rect 463022 31698 463204 31934
rect 444604 -6222 444786 -5986
rect 445022 -6222 445204 -5986
rect 444604 -6306 445204 -6222
rect 444604 -6542 444786 -6306
rect 445022 -6542 445204 -6306
rect 444604 -7504 445204 -6542
rect 462604 -6926 463204 31698
rect 469804 704838 470404 705800
rect 469804 704602 469986 704838
rect 470222 704602 470404 704838
rect 469804 704518 470404 704602
rect 469804 704282 469986 704518
rect 470222 704282 470404 704518
rect 469804 687454 470404 704282
rect 469804 687218 469986 687454
rect 470222 687218 470404 687454
rect 469804 687134 470404 687218
rect 469804 686898 469986 687134
rect 470222 686898 470404 687134
rect 469804 651454 470404 686898
rect 469804 651218 469986 651454
rect 470222 651218 470404 651454
rect 469804 651134 470404 651218
rect 469804 650898 469986 651134
rect 470222 650898 470404 651134
rect 469804 615454 470404 650898
rect 469804 615218 469986 615454
rect 470222 615218 470404 615454
rect 469804 615134 470404 615218
rect 469804 614898 469986 615134
rect 470222 614898 470404 615134
rect 469804 579454 470404 614898
rect 469804 579218 469986 579454
rect 470222 579218 470404 579454
rect 469804 579134 470404 579218
rect 469804 578898 469986 579134
rect 470222 578898 470404 579134
rect 469804 543454 470404 578898
rect 469804 543218 469986 543454
rect 470222 543218 470404 543454
rect 469804 543134 470404 543218
rect 469804 542898 469986 543134
rect 470222 542898 470404 543134
rect 469804 507454 470404 542898
rect 469804 507218 469986 507454
rect 470222 507218 470404 507454
rect 469804 507134 470404 507218
rect 469804 506898 469986 507134
rect 470222 506898 470404 507134
rect 469804 471454 470404 506898
rect 469804 471218 469986 471454
rect 470222 471218 470404 471454
rect 469804 471134 470404 471218
rect 469804 470898 469986 471134
rect 470222 470898 470404 471134
rect 469804 435454 470404 470898
rect 469804 435218 469986 435454
rect 470222 435218 470404 435454
rect 469804 435134 470404 435218
rect 469804 434898 469986 435134
rect 470222 434898 470404 435134
rect 469804 399454 470404 434898
rect 469804 399218 469986 399454
rect 470222 399218 470404 399454
rect 469804 399134 470404 399218
rect 469804 398898 469986 399134
rect 470222 398898 470404 399134
rect 469804 363454 470404 398898
rect 469804 363218 469986 363454
rect 470222 363218 470404 363454
rect 469804 363134 470404 363218
rect 469804 362898 469986 363134
rect 470222 362898 470404 363134
rect 469804 327454 470404 362898
rect 469804 327218 469986 327454
rect 470222 327218 470404 327454
rect 469804 327134 470404 327218
rect 469804 326898 469986 327134
rect 470222 326898 470404 327134
rect 469804 291454 470404 326898
rect 469804 291218 469986 291454
rect 470222 291218 470404 291454
rect 469804 291134 470404 291218
rect 469804 290898 469986 291134
rect 470222 290898 470404 291134
rect 469804 255454 470404 290898
rect 469804 255218 469986 255454
rect 470222 255218 470404 255454
rect 469804 255134 470404 255218
rect 469804 254898 469986 255134
rect 470222 254898 470404 255134
rect 469804 219454 470404 254898
rect 469804 219218 469986 219454
rect 470222 219218 470404 219454
rect 469804 219134 470404 219218
rect 469804 218898 469986 219134
rect 470222 218898 470404 219134
rect 469804 183454 470404 218898
rect 469804 183218 469986 183454
rect 470222 183218 470404 183454
rect 469804 183134 470404 183218
rect 469804 182898 469986 183134
rect 470222 182898 470404 183134
rect 469804 147454 470404 182898
rect 469804 147218 469986 147454
rect 470222 147218 470404 147454
rect 469804 147134 470404 147218
rect 469804 146898 469986 147134
rect 470222 146898 470404 147134
rect 469804 111454 470404 146898
rect 469804 111218 469986 111454
rect 470222 111218 470404 111454
rect 469804 111134 470404 111218
rect 469804 110898 469986 111134
rect 470222 110898 470404 111134
rect 469804 75454 470404 110898
rect 469804 75218 469986 75454
rect 470222 75218 470404 75454
rect 469804 75134 470404 75218
rect 469804 74898 469986 75134
rect 470222 74898 470404 75134
rect 469804 39454 470404 74898
rect 469804 39218 469986 39454
rect 470222 39218 470404 39454
rect 469804 39134 470404 39218
rect 469804 38898 469986 39134
rect 470222 38898 470404 39134
rect 469804 3454 470404 38898
rect 469804 3218 469986 3454
rect 470222 3218 470404 3454
rect 469804 3134 470404 3218
rect 469804 2898 469986 3134
rect 470222 2898 470404 3134
rect 469804 -346 470404 2898
rect 469804 -582 469986 -346
rect 470222 -582 470404 -346
rect 469804 -666 470404 -582
rect 469804 -902 469986 -666
rect 470222 -902 470404 -666
rect 469804 -1864 470404 -902
rect 473404 691054 474004 706162
rect 473404 690818 473586 691054
rect 473822 690818 474004 691054
rect 473404 690734 474004 690818
rect 473404 690498 473586 690734
rect 473822 690498 474004 690734
rect 473404 655054 474004 690498
rect 473404 654818 473586 655054
rect 473822 654818 474004 655054
rect 473404 654734 474004 654818
rect 473404 654498 473586 654734
rect 473822 654498 474004 654734
rect 473404 619054 474004 654498
rect 473404 618818 473586 619054
rect 473822 618818 474004 619054
rect 473404 618734 474004 618818
rect 473404 618498 473586 618734
rect 473822 618498 474004 618734
rect 473404 583054 474004 618498
rect 473404 582818 473586 583054
rect 473822 582818 474004 583054
rect 473404 582734 474004 582818
rect 473404 582498 473586 582734
rect 473822 582498 474004 582734
rect 473404 547054 474004 582498
rect 473404 546818 473586 547054
rect 473822 546818 474004 547054
rect 473404 546734 474004 546818
rect 473404 546498 473586 546734
rect 473822 546498 474004 546734
rect 473404 511054 474004 546498
rect 473404 510818 473586 511054
rect 473822 510818 474004 511054
rect 473404 510734 474004 510818
rect 473404 510498 473586 510734
rect 473822 510498 474004 510734
rect 473404 475054 474004 510498
rect 473404 474818 473586 475054
rect 473822 474818 474004 475054
rect 473404 474734 474004 474818
rect 473404 474498 473586 474734
rect 473822 474498 474004 474734
rect 473404 439054 474004 474498
rect 473404 438818 473586 439054
rect 473822 438818 474004 439054
rect 473404 438734 474004 438818
rect 473404 438498 473586 438734
rect 473822 438498 474004 438734
rect 473404 403054 474004 438498
rect 473404 402818 473586 403054
rect 473822 402818 474004 403054
rect 473404 402734 474004 402818
rect 473404 402498 473586 402734
rect 473822 402498 474004 402734
rect 473404 367054 474004 402498
rect 473404 366818 473586 367054
rect 473822 366818 474004 367054
rect 473404 366734 474004 366818
rect 473404 366498 473586 366734
rect 473822 366498 474004 366734
rect 473404 331054 474004 366498
rect 473404 330818 473586 331054
rect 473822 330818 474004 331054
rect 473404 330734 474004 330818
rect 473404 330498 473586 330734
rect 473822 330498 474004 330734
rect 473404 295054 474004 330498
rect 473404 294818 473586 295054
rect 473822 294818 474004 295054
rect 473404 294734 474004 294818
rect 473404 294498 473586 294734
rect 473822 294498 474004 294734
rect 473404 259054 474004 294498
rect 473404 258818 473586 259054
rect 473822 258818 474004 259054
rect 473404 258734 474004 258818
rect 473404 258498 473586 258734
rect 473822 258498 474004 258734
rect 473404 223054 474004 258498
rect 473404 222818 473586 223054
rect 473822 222818 474004 223054
rect 473404 222734 474004 222818
rect 473404 222498 473586 222734
rect 473822 222498 474004 222734
rect 473404 187054 474004 222498
rect 473404 186818 473586 187054
rect 473822 186818 474004 187054
rect 473404 186734 474004 186818
rect 473404 186498 473586 186734
rect 473822 186498 474004 186734
rect 473404 151054 474004 186498
rect 473404 150818 473586 151054
rect 473822 150818 474004 151054
rect 473404 150734 474004 150818
rect 473404 150498 473586 150734
rect 473822 150498 474004 150734
rect 473404 115054 474004 150498
rect 473404 114818 473586 115054
rect 473822 114818 474004 115054
rect 473404 114734 474004 114818
rect 473404 114498 473586 114734
rect 473822 114498 474004 114734
rect 473404 79054 474004 114498
rect 473404 78818 473586 79054
rect 473822 78818 474004 79054
rect 473404 78734 474004 78818
rect 473404 78498 473586 78734
rect 473822 78498 474004 78734
rect 473404 43054 474004 78498
rect 473404 42818 473586 43054
rect 473822 42818 474004 43054
rect 473404 42734 474004 42818
rect 473404 42498 473586 42734
rect 473822 42498 474004 42734
rect 473404 7054 474004 42498
rect 473404 6818 473586 7054
rect 473822 6818 474004 7054
rect 473404 6734 474004 6818
rect 473404 6498 473586 6734
rect 473822 6498 474004 6734
rect 473404 -2226 474004 6498
rect 473404 -2462 473586 -2226
rect 473822 -2462 474004 -2226
rect 473404 -2546 474004 -2462
rect 473404 -2782 473586 -2546
rect 473822 -2782 474004 -2546
rect 473404 -3744 474004 -2782
rect 477004 694654 477604 708042
rect 477004 694418 477186 694654
rect 477422 694418 477604 694654
rect 477004 694334 477604 694418
rect 477004 694098 477186 694334
rect 477422 694098 477604 694334
rect 477004 658654 477604 694098
rect 477004 658418 477186 658654
rect 477422 658418 477604 658654
rect 477004 658334 477604 658418
rect 477004 658098 477186 658334
rect 477422 658098 477604 658334
rect 477004 622654 477604 658098
rect 477004 622418 477186 622654
rect 477422 622418 477604 622654
rect 477004 622334 477604 622418
rect 477004 622098 477186 622334
rect 477422 622098 477604 622334
rect 477004 586654 477604 622098
rect 477004 586418 477186 586654
rect 477422 586418 477604 586654
rect 477004 586334 477604 586418
rect 477004 586098 477186 586334
rect 477422 586098 477604 586334
rect 477004 550654 477604 586098
rect 477004 550418 477186 550654
rect 477422 550418 477604 550654
rect 477004 550334 477604 550418
rect 477004 550098 477186 550334
rect 477422 550098 477604 550334
rect 477004 514654 477604 550098
rect 477004 514418 477186 514654
rect 477422 514418 477604 514654
rect 477004 514334 477604 514418
rect 477004 514098 477186 514334
rect 477422 514098 477604 514334
rect 477004 478654 477604 514098
rect 477004 478418 477186 478654
rect 477422 478418 477604 478654
rect 477004 478334 477604 478418
rect 477004 478098 477186 478334
rect 477422 478098 477604 478334
rect 477004 442654 477604 478098
rect 477004 442418 477186 442654
rect 477422 442418 477604 442654
rect 477004 442334 477604 442418
rect 477004 442098 477186 442334
rect 477422 442098 477604 442334
rect 477004 406654 477604 442098
rect 477004 406418 477186 406654
rect 477422 406418 477604 406654
rect 477004 406334 477604 406418
rect 477004 406098 477186 406334
rect 477422 406098 477604 406334
rect 477004 370654 477604 406098
rect 477004 370418 477186 370654
rect 477422 370418 477604 370654
rect 477004 370334 477604 370418
rect 477004 370098 477186 370334
rect 477422 370098 477604 370334
rect 477004 334654 477604 370098
rect 477004 334418 477186 334654
rect 477422 334418 477604 334654
rect 477004 334334 477604 334418
rect 477004 334098 477186 334334
rect 477422 334098 477604 334334
rect 477004 298654 477604 334098
rect 477004 298418 477186 298654
rect 477422 298418 477604 298654
rect 477004 298334 477604 298418
rect 477004 298098 477186 298334
rect 477422 298098 477604 298334
rect 477004 262654 477604 298098
rect 477004 262418 477186 262654
rect 477422 262418 477604 262654
rect 477004 262334 477604 262418
rect 477004 262098 477186 262334
rect 477422 262098 477604 262334
rect 477004 226654 477604 262098
rect 477004 226418 477186 226654
rect 477422 226418 477604 226654
rect 477004 226334 477604 226418
rect 477004 226098 477186 226334
rect 477422 226098 477604 226334
rect 477004 190654 477604 226098
rect 477004 190418 477186 190654
rect 477422 190418 477604 190654
rect 477004 190334 477604 190418
rect 477004 190098 477186 190334
rect 477422 190098 477604 190334
rect 477004 154654 477604 190098
rect 477004 154418 477186 154654
rect 477422 154418 477604 154654
rect 477004 154334 477604 154418
rect 477004 154098 477186 154334
rect 477422 154098 477604 154334
rect 477004 118654 477604 154098
rect 477004 118418 477186 118654
rect 477422 118418 477604 118654
rect 477004 118334 477604 118418
rect 477004 118098 477186 118334
rect 477422 118098 477604 118334
rect 477004 82654 477604 118098
rect 477004 82418 477186 82654
rect 477422 82418 477604 82654
rect 477004 82334 477604 82418
rect 477004 82098 477186 82334
rect 477422 82098 477604 82334
rect 477004 46654 477604 82098
rect 477004 46418 477186 46654
rect 477422 46418 477604 46654
rect 477004 46334 477604 46418
rect 477004 46098 477186 46334
rect 477422 46098 477604 46334
rect 477004 10654 477604 46098
rect 477004 10418 477186 10654
rect 477422 10418 477604 10654
rect 477004 10334 477604 10418
rect 477004 10098 477186 10334
rect 477422 10098 477604 10334
rect 477004 -4106 477604 10098
rect 477004 -4342 477186 -4106
rect 477422 -4342 477604 -4106
rect 477004 -4426 477604 -4342
rect 477004 -4662 477186 -4426
rect 477422 -4662 477604 -4426
rect 477004 -5624 477604 -4662
rect 480604 698254 481204 709922
rect 498604 711418 499204 711440
rect 498604 711182 498786 711418
rect 499022 711182 499204 711418
rect 498604 711098 499204 711182
rect 498604 710862 498786 711098
rect 499022 710862 499204 711098
rect 495004 709538 495604 709560
rect 495004 709302 495186 709538
rect 495422 709302 495604 709538
rect 495004 709218 495604 709302
rect 495004 708982 495186 709218
rect 495422 708982 495604 709218
rect 491404 707658 492004 707680
rect 491404 707422 491586 707658
rect 491822 707422 492004 707658
rect 491404 707338 492004 707422
rect 491404 707102 491586 707338
rect 491822 707102 492004 707338
rect 480604 698018 480786 698254
rect 481022 698018 481204 698254
rect 480604 697934 481204 698018
rect 480604 697698 480786 697934
rect 481022 697698 481204 697934
rect 480604 662254 481204 697698
rect 480604 662018 480786 662254
rect 481022 662018 481204 662254
rect 480604 661934 481204 662018
rect 480604 661698 480786 661934
rect 481022 661698 481204 661934
rect 480604 626254 481204 661698
rect 480604 626018 480786 626254
rect 481022 626018 481204 626254
rect 480604 625934 481204 626018
rect 480604 625698 480786 625934
rect 481022 625698 481204 625934
rect 480604 590254 481204 625698
rect 480604 590018 480786 590254
rect 481022 590018 481204 590254
rect 480604 589934 481204 590018
rect 480604 589698 480786 589934
rect 481022 589698 481204 589934
rect 480604 554254 481204 589698
rect 480604 554018 480786 554254
rect 481022 554018 481204 554254
rect 480604 553934 481204 554018
rect 480604 553698 480786 553934
rect 481022 553698 481204 553934
rect 480604 518254 481204 553698
rect 480604 518018 480786 518254
rect 481022 518018 481204 518254
rect 480604 517934 481204 518018
rect 480604 517698 480786 517934
rect 481022 517698 481204 517934
rect 480604 482254 481204 517698
rect 480604 482018 480786 482254
rect 481022 482018 481204 482254
rect 480604 481934 481204 482018
rect 480604 481698 480786 481934
rect 481022 481698 481204 481934
rect 480604 446254 481204 481698
rect 480604 446018 480786 446254
rect 481022 446018 481204 446254
rect 480604 445934 481204 446018
rect 480604 445698 480786 445934
rect 481022 445698 481204 445934
rect 480604 410254 481204 445698
rect 480604 410018 480786 410254
rect 481022 410018 481204 410254
rect 480604 409934 481204 410018
rect 480604 409698 480786 409934
rect 481022 409698 481204 409934
rect 480604 374254 481204 409698
rect 480604 374018 480786 374254
rect 481022 374018 481204 374254
rect 480604 373934 481204 374018
rect 480604 373698 480786 373934
rect 481022 373698 481204 373934
rect 480604 338254 481204 373698
rect 480604 338018 480786 338254
rect 481022 338018 481204 338254
rect 480604 337934 481204 338018
rect 480604 337698 480786 337934
rect 481022 337698 481204 337934
rect 480604 302254 481204 337698
rect 480604 302018 480786 302254
rect 481022 302018 481204 302254
rect 480604 301934 481204 302018
rect 480604 301698 480786 301934
rect 481022 301698 481204 301934
rect 480604 266254 481204 301698
rect 480604 266018 480786 266254
rect 481022 266018 481204 266254
rect 480604 265934 481204 266018
rect 480604 265698 480786 265934
rect 481022 265698 481204 265934
rect 480604 230254 481204 265698
rect 480604 230018 480786 230254
rect 481022 230018 481204 230254
rect 480604 229934 481204 230018
rect 480604 229698 480786 229934
rect 481022 229698 481204 229934
rect 480604 194254 481204 229698
rect 480604 194018 480786 194254
rect 481022 194018 481204 194254
rect 480604 193934 481204 194018
rect 480604 193698 480786 193934
rect 481022 193698 481204 193934
rect 480604 158254 481204 193698
rect 480604 158018 480786 158254
rect 481022 158018 481204 158254
rect 480604 157934 481204 158018
rect 480604 157698 480786 157934
rect 481022 157698 481204 157934
rect 480604 122254 481204 157698
rect 480604 122018 480786 122254
rect 481022 122018 481204 122254
rect 480604 121934 481204 122018
rect 480604 121698 480786 121934
rect 481022 121698 481204 121934
rect 480604 86254 481204 121698
rect 480604 86018 480786 86254
rect 481022 86018 481204 86254
rect 480604 85934 481204 86018
rect 480604 85698 480786 85934
rect 481022 85698 481204 85934
rect 480604 50254 481204 85698
rect 480604 50018 480786 50254
rect 481022 50018 481204 50254
rect 480604 49934 481204 50018
rect 480604 49698 480786 49934
rect 481022 49698 481204 49934
rect 480604 14254 481204 49698
rect 480604 14018 480786 14254
rect 481022 14018 481204 14254
rect 480604 13934 481204 14018
rect 480604 13698 480786 13934
rect 481022 13698 481204 13934
rect 462604 -7162 462786 -6926
rect 463022 -7162 463204 -6926
rect 462604 -7246 463204 -7162
rect 462604 -7482 462786 -7246
rect 463022 -7482 463204 -7246
rect 462604 -7504 463204 -7482
rect 480604 -5986 481204 13698
rect 487804 705778 488404 705800
rect 487804 705542 487986 705778
rect 488222 705542 488404 705778
rect 487804 705458 488404 705542
rect 487804 705222 487986 705458
rect 488222 705222 488404 705458
rect 487804 669454 488404 705222
rect 487804 669218 487986 669454
rect 488222 669218 488404 669454
rect 487804 669134 488404 669218
rect 487804 668898 487986 669134
rect 488222 668898 488404 669134
rect 487804 633454 488404 668898
rect 487804 633218 487986 633454
rect 488222 633218 488404 633454
rect 487804 633134 488404 633218
rect 487804 632898 487986 633134
rect 488222 632898 488404 633134
rect 487804 597454 488404 632898
rect 487804 597218 487986 597454
rect 488222 597218 488404 597454
rect 487804 597134 488404 597218
rect 487804 596898 487986 597134
rect 488222 596898 488404 597134
rect 487804 561454 488404 596898
rect 487804 561218 487986 561454
rect 488222 561218 488404 561454
rect 487804 561134 488404 561218
rect 487804 560898 487986 561134
rect 488222 560898 488404 561134
rect 487804 525454 488404 560898
rect 487804 525218 487986 525454
rect 488222 525218 488404 525454
rect 487804 525134 488404 525218
rect 487804 524898 487986 525134
rect 488222 524898 488404 525134
rect 487804 489454 488404 524898
rect 487804 489218 487986 489454
rect 488222 489218 488404 489454
rect 487804 489134 488404 489218
rect 487804 488898 487986 489134
rect 488222 488898 488404 489134
rect 487804 453454 488404 488898
rect 487804 453218 487986 453454
rect 488222 453218 488404 453454
rect 487804 453134 488404 453218
rect 487804 452898 487986 453134
rect 488222 452898 488404 453134
rect 487804 417454 488404 452898
rect 487804 417218 487986 417454
rect 488222 417218 488404 417454
rect 487804 417134 488404 417218
rect 487804 416898 487986 417134
rect 488222 416898 488404 417134
rect 487804 381454 488404 416898
rect 487804 381218 487986 381454
rect 488222 381218 488404 381454
rect 487804 381134 488404 381218
rect 487804 380898 487986 381134
rect 488222 380898 488404 381134
rect 487804 345454 488404 380898
rect 487804 345218 487986 345454
rect 488222 345218 488404 345454
rect 487804 345134 488404 345218
rect 487804 344898 487986 345134
rect 488222 344898 488404 345134
rect 487804 309454 488404 344898
rect 487804 309218 487986 309454
rect 488222 309218 488404 309454
rect 487804 309134 488404 309218
rect 487804 308898 487986 309134
rect 488222 308898 488404 309134
rect 487804 273454 488404 308898
rect 487804 273218 487986 273454
rect 488222 273218 488404 273454
rect 487804 273134 488404 273218
rect 487804 272898 487986 273134
rect 488222 272898 488404 273134
rect 487804 237454 488404 272898
rect 487804 237218 487986 237454
rect 488222 237218 488404 237454
rect 487804 237134 488404 237218
rect 487804 236898 487986 237134
rect 488222 236898 488404 237134
rect 487804 201454 488404 236898
rect 487804 201218 487986 201454
rect 488222 201218 488404 201454
rect 487804 201134 488404 201218
rect 487804 200898 487986 201134
rect 488222 200898 488404 201134
rect 487804 165454 488404 200898
rect 487804 165218 487986 165454
rect 488222 165218 488404 165454
rect 487804 165134 488404 165218
rect 487804 164898 487986 165134
rect 488222 164898 488404 165134
rect 487804 129454 488404 164898
rect 487804 129218 487986 129454
rect 488222 129218 488404 129454
rect 487804 129134 488404 129218
rect 487804 128898 487986 129134
rect 488222 128898 488404 129134
rect 487804 93454 488404 128898
rect 487804 93218 487986 93454
rect 488222 93218 488404 93454
rect 487804 93134 488404 93218
rect 487804 92898 487986 93134
rect 488222 92898 488404 93134
rect 487804 57454 488404 92898
rect 487804 57218 487986 57454
rect 488222 57218 488404 57454
rect 487804 57134 488404 57218
rect 487804 56898 487986 57134
rect 488222 56898 488404 57134
rect 487804 21454 488404 56898
rect 487804 21218 487986 21454
rect 488222 21218 488404 21454
rect 487804 21134 488404 21218
rect 487804 20898 487986 21134
rect 488222 20898 488404 21134
rect 487804 -1286 488404 20898
rect 487804 -1522 487986 -1286
rect 488222 -1522 488404 -1286
rect 487804 -1606 488404 -1522
rect 487804 -1842 487986 -1606
rect 488222 -1842 488404 -1606
rect 487804 -1864 488404 -1842
rect 491404 673054 492004 707102
rect 491404 672818 491586 673054
rect 491822 672818 492004 673054
rect 491404 672734 492004 672818
rect 491404 672498 491586 672734
rect 491822 672498 492004 672734
rect 491404 637054 492004 672498
rect 491404 636818 491586 637054
rect 491822 636818 492004 637054
rect 491404 636734 492004 636818
rect 491404 636498 491586 636734
rect 491822 636498 492004 636734
rect 491404 601054 492004 636498
rect 491404 600818 491586 601054
rect 491822 600818 492004 601054
rect 491404 600734 492004 600818
rect 491404 600498 491586 600734
rect 491822 600498 492004 600734
rect 491404 565054 492004 600498
rect 491404 564818 491586 565054
rect 491822 564818 492004 565054
rect 491404 564734 492004 564818
rect 491404 564498 491586 564734
rect 491822 564498 492004 564734
rect 491404 529054 492004 564498
rect 491404 528818 491586 529054
rect 491822 528818 492004 529054
rect 491404 528734 492004 528818
rect 491404 528498 491586 528734
rect 491822 528498 492004 528734
rect 491404 493054 492004 528498
rect 491404 492818 491586 493054
rect 491822 492818 492004 493054
rect 491404 492734 492004 492818
rect 491404 492498 491586 492734
rect 491822 492498 492004 492734
rect 491404 457054 492004 492498
rect 491404 456818 491586 457054
rect 491822 456818 492004 457054
rect 491404 456734 492004 456818
rect 491404 456498 491586 456734
rect 491822 456498 492004 456734
rect 491404 421054 492004 456498
rect 491404 420818 491586 421054
rect 491822 420818 492004 421054
rect 491404 420734 492004 420818
rect 491404 420498 491586 420734
rect 491822 420498 492004 420734
rect 491404 385054 492004 420498
rect 491404 384818 491586 385054
rect 491822 384818 492004 385054
rect 491404 384734 492004 384818
rect 491404 384498 491586 384734
rect 491822 384498 492004 384734
rect 491404 349054 492004 384498
rect 491404 348818 491586 349054
rect 491822 348818 492004 349054
rect 491404 348734 492004 348818
rect 491404 348498 491586 348734
rect 491822 348498 492004 348734
rect 491404 313054 492004 348498
rect 491404 312818 491586 313054
rect 491822 312818 492004 313054
rect 491404 312734 492004 312818
rect 491404 312498 491586 312734
rect 491822 312498 492004 312734
rect 491404 277054 492004 312498
rect 491404 276818 491586 277054
rect 491822 276818 492004 277054
rect 491404 276734 492004 276818
rect 491404 276498 491586 276734
rect 491822 276498 492004 276734
rect 491404 241054 492004 276498
rect 491404 240818 491586 241054
rect 491822 240818 492004 241054
rect 491404 240734 492004 240818
rect 491404 240498 491586 240734
rect 491822 240498 492004 240734
rect 491404 205054 492004 240498
rect 491404 204818 491586 205054
rect 491822 204818 492004 205054
rect 491404 204734 492004 204818
rect 491404 204498 491586 204734
rect 491822 204498 492004 204734
rect 491404 169054 492004 204498
rect 491404 168818 491586 169054
rect 491822 168818 492004 169054
rect 491404 168734 492004 168818
rect 491404 168498 491586 168734
rect 491822 168498 492004 168734
rect 491404 133054 492004 168498
rect 491404 132818 491586 133054
rect 491822 132818 492004 133054
rect 491404 132734 492004 132818
rect 491404 132498 491586 132734
rect 491822 132498 492004 132734
rect 491404 97054 492004 132498
rect 491404 96818 491586 97054
rect 491822 96818 492004 97054
rect 491404 96734 492004 96818
rect 491404 96498 491586 96734
rect 491822 96498 492004 96734
rect 491404 61054 492004 96498
rect 491404 60818 491586 61054
rect 491822 60818 492004 61054
rect 491404 60734 492004 60818
rect 491404 60498 491586 60734
rect 491822 60498 492004 60734
rect 491404 25054 492004 60498
rect 491404 24818 491586 25054
rect 491822 24818 492004 25054
rect 491404 24734 492004 24818
rect 491404 24498 491586 24734
rect 491822 24498 492004 24734
rect 491404 -3166 492004 24498
rect 491404 -3402 491586 -3166
rect 491822 -3402 492004 -3166
rect 491404 -3486 492004 -3402
rect 491404 -3722 491586 -3486
rect 491822 -3722 492004 -3486
rect 491404 -3744 492004 -3722
rect 495004 676654 495604 708982
rect 495004 676418 495186 676654
rect 495422 676418 495604 676654
rect 495004 676334 495604 676418
rect 495004 676098 495186 676334
rect 495422 676098 495604 676334
rect 495004 640654 495604 676098
rect 495004 640418 495186 640654
rect 495422 640418 495604 640654
rect 495004 640334 495604 640418
rect 495004 640098 495186 640334
rect 495422 640098 495604 640334
rect 495004 604654 495604 640098
rect 495004 604418 495186 604654
rect 495422 604418 495604 604654
rect 495004 604334 495604 604418
rect 495004 604098 495186 604334
rect 495422 604098 495604 604334
rect 495004 568654 495604 604098
rect 495004 568418 495186 568654
rect 495422 568418 495604 568654
rect 495004 568334 495604 568418
rect 495004 568098 495186 568334
rect 495422 568098 495604 568334
rect 495004 532654 495604 568098
rect 495004 532418 495186 532654
rect 495422 532418 495604 532654
rect 495004 532334 495604 532418
rect 495004 532098 495186 532334
rect 495422 532098 495604 532334
rect 495004 496654 495604 532098
rect 495004 496418 495186 496654
rect 495422 496418 495604 496654
rect 495004 496334 495604 496418
rect 495004 496098 495186 496334
rect 495422 496098 495604 496334
rect 495004 460654 495604 496098
rect 495004 460418 495186 460654
rect 495422 460418 495604 460654
rect 495004 460334 495604 460418
rect 495004 460098 495186 460334
rect 495422 460098 495604 460334
rect 495004 424654 495604 460098
rect 495004 424418 495186 424654
rect 495422 424418 495604 424654
rect 495004 424334 495604 424418
rect 495004 424098 495186 424334
rect 495422 424098 495604 424334
rect 495004 388654 495604 424098
rect 495004 388418 495186 388654
rect 495422 388418 495604 388654
rect 495004 388334 495604 388418
rect 495004 388098 495186 388334
rect 495422 388098 495604 388334
rect 495004 352654 495604 388098
rect 495004 352418 495186 352654
rect 495422 352418 495604 352654
rect 495004 352334 495604 352418
rect 495004 352098 495186 352334
rect 495422 352098 495604 352334
rect 495004 316654 495604 352098
rect 495004 316418 495186 316654
rect 495422 316418 495604 316654
rect 495004 316334 495604 316418
rect 495004 316098 495186 316334
rect 495422 316098 495604 316334
rect 495004 280654 495604 316098
rect 495004 280418 495186 280654
rect 495422 280418 495604 280654
rect 495004 280334 495604 280418
rect 495004 280098 495186 280334
rect 495422 280098 495604 280334
rect 495004 244654 495604 280098
rect 495004 244418 495186 244654
rect 495422 244418 495604 244654
rect 495004 244334 495604 244418
rect 495004 244098 495186 244334
rect 495422 244098 495604 244334
rect 495004 208654 495604 244098
rect 495004 208418 495186 208654
rect 495422 208418 495604 208654
rect 495004 208334 495604 208418
rect 495004 208098 495186 208334
rect 495422 208098 495604 208334
rect 495004 172654 495604 208098
rect 495004 172418 495186 172654
rect 495422 172418 495604 172654
rect 495004 172334 495604 172418
rect 495004 172098 495186 172334
rect 495422 172098 495604 172334
rect 495004 136654 495604 172098
rect 495004 136418 495186 136654
rect 495422 136418 495604 136654
rect 495004 136334 495604 136418
rect 495004 136098 495186 136334
rect 495422 136098 495604 136334
rect 495004 100654 495604 136098
rect 495004 100418 495186 100654
rect 495422 100418 495604 100654
rect 495004 100334 495604 100418
rect 495004 100098 495186 100334
rect 495422 100098 495604 100334
rect 495004 64654 495604 100098
rect 495004 64418 495186 64654
rect 495422 64418 495604 64654
rect 495004 64334 495604 64418
rect 495004 64098 495186 64334
rect 495422 64098 495604 64334
rect 495004 28654 495604 64098
rect 495004 28418 495186 28654
rect 495422 28418 495604 28654
rect 495004 28334 495604 28418
rect 495004 28098 495186 28334
rect 495422 28098 495604 28334
rect 495004 -5046 495604 28098
rect 495004 -5282 495186 -5046
rect 495422 -5282 495604 -5046
rect 495004 -5366 495604 -5282
rect 495004 -5602 495186 -5366
rect 495422 -5602 495604 -5366
rect 495004 -5624 495604 -5602
rect 498604 680254 499204 710862
rect 516604 710478 517204 711440
rect 516604 710242 516786 710478
rect 517022 710242 517204 710478
rect 516604 710158 517204 710242
rect 516604 709922 516786 710158
rect 517022 709922 517204 710158
rect 513004 708598 513604 709560
rect 513004 708362 513186 708598
rect 513422 708362 513604 708598
rect 513004 708278 513604 708362
rect 513004 708042 513186 708278
rect 513422 708042 513604 708278
rect 509404 706718 510004 707680
rect 509404 706482 509586 706718
rect 509822 706482 510004 706718
rect 509404 706398 510004 706482
rect 509404 706162 509586 706398
rect 509822 706162 510004 706398
rect 498604 680018 498786 680254
rect 499022 680018 499204 680254
rect 498604 679934 499204 680018
rect 498604 679698 498786 679934
rect 499022 679698 499204 679934
rect 498604 644254 499204 679698
rect 498604 644018 498786 644254
rect 499022 644018 499204 644254
rect 498604 643934 499204 644018
rect 498604 643698 498786 643934
rect 499022 643698 499204 643934
rect 498604 608254 499204 643698
rect 498604 608018 498786 608254
rect 499022 608018 499204 608254
rect 498604 607934 499204 608018
rect 498604 607698 498786 607934
rect 499022 607698 499204 607934
rect 498604 572254 499204 607698
rect 498604 572018 498786 572254
rect 499022 572018 499204 572254
rect 498604 571934 499204 572018
rect 498604 571698 498786 571934
rect 499022 571698 499204 571934
rect 498604 536254 499204 571698
rect 498604 536018 498786 536254
rect 499022 536018 499204 536254
rect 498604 535934 499204 536018
rect 498604 535698 498786 535934
rect 499022 535698 499204 535934
rect 498604 500254 499204 535698
rect 498604 500018 498786 500254
rect 499022 500018 499204 500254
rect 498604 499934 499204 500018
rect 498604 499698 498786 499934
rect 499022 499698 499204 499934
rect 498604 464254 499204 499698
rect 498604 464018 498786 464254
rect 499022 464018 499204 464254
rect 498604 463934 499204 464018
rect 498604 463698 498786 463934
rect 499022 463698 499204 463934
rect 498604 428254 499204 463698
rect 498604 428018 498786 428254
rect 499022 428018 499204 428254
rect 498604 427934 499204 428018
rect 498604 427698 498786 427934
rect 499022 427698 499204 427934
rect 498604 392254 499204 427698
rect 498604 392018 498786 392254
rect 499022 392018 499204 392254
rect 498604 391934 499204 392018
rect 498604 391698 498786 391934
rect 499022 391698 499204 391934
rect 498604 356254 499204 391698
rect 498604 356018 498786 356254
rect 499022 356018 499204 356254
rect 498604 355934 499204 356018
rect 498604 355698 498786 355934
rect 499022 355698 499204 355934
rect 498604 320254 499204 355698
rect 498604 320018 498786 320254
rect 499022 320018 499204 320254
rect 498604 319934 499204 320018
rect 498604 319698 498786 319934
rect 499022 319698 499204 319934
rect 498604 284254 499204 319698
rect 498604 284018 498786 284254
rect 499022 284018 499204 284254
rect 498604 283934 499204 284018
rect 498604 283698 498786 283934
rect 499022 283698 499204 283934
rect 498604 248254 499204 283698
rect 498604 248018 498786 248254
rect 499022 248018 499204 248254
rect 498604 247934 499204 248018
rect 498604 247698 498786 247934
rect 499022 247698 499204 247934
rect 498604 212254 499204 247698
rect 498604 212018 498786 212254
rect 499022 212018 499204 212254
rect 498604 211934 499204 212018
rect 498604 211698 498786 211934
rect 499022 211698 499204 211934
rect 498604 176254 499204 211698
rect 498604 176018 498786 176254
rect 499022 176018 499204 176254
rect 498604 175934 499204 176018
rect 498604 175698 498786 175934
rect 499022 175698 499204 175934
rect 498604 140254 499204 175698
rect 498604 140018 498786 140254
rect 499022 140018 499204 140254
rect 498604 139934 499204 140018
rect 498604 139698 498786 139934
rect 499022 139698 499204 139934
rect 498604 104254 499204 139698
rect 498604 104018 498786 104254
rect 499022 104018 499204 104254
rect 498604 103934 499204 104018
rect 498604 103698 498786 103934
rect 499022 103698 499204 103934
rect 498604 68254 499204 103698
rect 498604 68018 498786 68254
rect 499022 68018 499204 68254
rect 498604 67934 499204 68018
rect 498604 67698 498786 67934
rect 499022 67698 499204 67934
rect 498604 32254 499204 67698
rect 498604 32018 498786 32254
rect 499022 32018 499204 32254
rect 498604 31934 499204 32018
rect 498604 31698 498786 31934
rect 499022 31698 499204 31934
rect 480604 -6222 480786 -5986
rect 481022 -6222 481204 -5986
rect 480604 -6306 481204 -6222
rect 480604 -6542 480786 -6306
rect 481022 -6542 481204 -6306
rect 480604 -7504 481204 -6542
rect 498604 -6926 499204 31698
rect 505804 704838 506404 705800
rect 505804 704602 505986 704838
rect 506222 704602 506404 704838
rect 505804 704518 506404 704602
rect 505804 704282 505986 704518
rect 506222 704282 506404 704518
rect 505804 687454 506404 704282
rect 505804 687218 505986 687454
rect 506222 687218 506404 687454
rect 505804 687134 506404 687218
rect 505804 686898 505986 687134
rect 506222 686898 506404 687134
rect 505804 651454 506404 686898
rect 505804 651218 505986 651454
rect 506222 651218 506404 651454
rect 505804 651134 506404 651218
rect 505804 650898 505986 651134
rect 506222 650898 506404 651134
rect 505804 615454 506404 650898
rect 505804 615218 505986 615454
rect 506222 615218 506404 615454
rect 505804 615134 506404 615218
rect 505804 614898 505986 615134
rect 506222 614898 506404 615134
rect 505804 579454 506404 614898
rect 505804 579218 505986 579454
rect 506222 579218 506404 579454
rect 505804 579134 506404 579218
rect 505804 578898 505986 579134
rect 506222 578898 506404 579134
rect 505804 543454 506404 578898
rect 505804 543218 505986 543454
rect 506222 543218 506404 543454
rect 505804 543134 506404 543218
rect 505804 542898 505986 543134
rect 506222 542898 506404 543134
rect 505804 507454 506404 542898
rect 505804 507218 505986 507454
rect 506222 507218 506404 507454
rect 505804 507134 506404 507218
rect 505804 506898 505986 507134
rect 506222 506898 506404 507134
rect 505804 471454 506404 506898
rect 505804 471218 505986 471454
rect 506222 471218 506404 471454
rect 505804 471134 506404 471218
rect 505804 470898 505986 471134
rect 506222 470898 506404 471134
rect 505804 435454 506404 470898
rect 505804 435218 505986 435454
rect 506222 435218 506404 435454
rect 505804 435134 506404 435218
rect 505804 434898 505986 435134
rect 506222 434898 506404 435134
rect 505804 399454 506404 434898
rect 505804 399218 505986 399454
rect 506222 399218 506404 399454
rect 505804 399134 506404 399218
rect 505804 398898 505986 399134
rect 506222 398898 506404 399134
rect 505804 363454 506404 398898
rect 505804 363218 505986 363454
rect 506222 363218 506404 363454
rect 505804 363134 506404 363218
rect 505804 362898 505986 363134
rect 506222 362898 506404 363134
rect 505804 327454 506404 362898
rect 505804 327218 505986 327454
rect 506222 327218 506404 327454
rect 505804 327134 506404 327218
rect 505804 326898 505986 327134
rect 506222 326898 506404 327134
rect 505804 291454 506404 326898
rect 505804 291218 505986 291454
rect 506222 291218 506404 291454
rect 505804 291134 506404 291218
rect 505804 290898 505986 291134
rect 506222 290898 506404 291134
rect 505804 255454 506404 290898
rect 505804 255218 505986 255454
rect 506222 255218 506404 255454
rect 505804 255134 506404 255218
rect 505804 254898 505986 255134
rect 506222 254898 506404 255134
rect 505804 219454 506404 254898
rect 505804 219218 505986 219454
rect 506222 219218 506404 219454
rect 505804 219134 506404 219218
rect 505804 218898 505986 219134
rect 506222 218898 506404 219134
rect 505804 183454 506404 218898
rect 505804 183218 505986 183454
rect 506222 183218 506404 183454
rect 505804 183134 506404 183218
rect 505804 182898 505986 183134
rect 506222 182898 506404 183134
rect 505804 147454 506404 182898
rect 505804 147218 505986 147454
rect 506222 147218 506404 147454
rect 505804 147134 506404 147218
rect 505804 146898 505986 147134
rect 506222 146898 506404 147134
rect 505804 111454 506404 146898
rect 505804 111218 505986 111454
rect 506222 111218 506404 111454
rect 505804 111134 506404 111218
rect 505804 110898 505986 111134
rect 506222 110898 506404 111134
rect 505804 75454 506404 110898
rect 505804 75218 505986 75454
rect 506222 75218 506404 75454
rect 505804 75134 506404 75218
rect 505804 74898 505986 75134
rect 506222 74898 506404 75134
rect 505804 39454 506404 74898
rect 505804 39218 505986 39454
rect 506222 39218 506404 39454
rect 505804 39134 506404 39218
rect 505804 38898 505986 39134
rect 506222 38898 506404 39134
rect 505804 3454 506404 38898
rect 505804 3218 505986 3454
rect 506222 3218 506404 3454
rect 505804 3134 506404 3218
rect 505804 2898 505986 3134
rect 506222 2898 506404 3134
rect 505804 -346 506404 2898
rect 505804 -582 505986 -346
rect 506222 -582 506404 -346
rect 505804 -666 506404 -582
rect 505804 -902 505986 -666
rect 506222 -902 506404 -666
rect 505804 -1864 506404 -902
rect 509404 691054 510004 706162
rect 509404 690818 509586 691054
rect 509822 690818 510004 691054
rect 509404 690734 510004 690818
rect 509404 690498 509586 690734
rect 509822 690498 510004 690734
rect 509404 655054 510004 690498
rect 509404 654818 509586 655054
rect 509822 654818 510004 655054
rect 509404 654734 510004 654818
rect 509404 654498 509586 654734
rect 509822 654498 510004 654734
rect 509404 619054 510004 654498
rect 509404 618818 509586 619054
rect 509822 618818 510004 619054
rect 509404 618734 510004 618818
rect 509404 618498 509586 618734
rect 509822 618498 510004 618734
rect 509404 583054 510004 618498
rect 509404 582818 509586 583054
rect 509822 582818 510004 583054
rect 509404 582734 510004 582818
rect 509404 582498 509586 582734
rect 509822 582498 510004 582734
rect 509404 547054 510004 582498
rect 509404 546818 509586 547054
rect 509822 546818 510004 547054
rect 509404 546734 510004 546818
rect 509404 546498 509586 546734
rect 509822 546498 510004 546734
rect 509404 511054 510004 546498
rect 509404 510818 509586 511054
rect 509822 510818 510004 511054
rect 509404 510734 510004 510818
rect 509404 510498 509586 510734
rect 509822 510498 510004 510734
rect 509404 475054 510004 510498
rect 509404 474818 509586 475054
rect 509822 474818 510004 475054
rect 509404 474734 510004 474818
rect 509404 474498 509586 474734
rect 509822 474498 510004 474734
rect 509404 439054 510004 474498
rect 509404 438818 509586 439054
rect 509822 438818 510004 439054
rect 509404 438734 510004 438818
rect 509404 438498 509586 438734
rect 509822 438498 510004 438734
rect 509404 403054 510004 438498
rect 509404 402818 509586 403054
rect 509822 402818 510004 403054
rect 509404 402734 510004 402818
rect 509404 402498 509586 402734
rect 509822 402498 510004 402734
rect 509404 367054 510004 402498
rect 509404 366818 509586 367054
rect 509822 366818 510004 367054
rect 509404 366734 510004 366818
rect 509404 366498 509586 366734
rect 509822 366498 510004 366734
rect 509404 331054 510004 366498
rect 509404 330818 509586 331054
rect 509822 330818 510004 331054
rect 509404 330734 510004 330818
rect 509404 330498 509586 330734
rect 509822 330498 510004 330734
rect 509404 295054 510004 330498
rect 509404 294818 509586 295054
rect 509822 294818 510004 295054
rect 509404 294734 510004 294818
rect 509404 294498 509586 294734
rect 509822 294498 510004 294734
rect 509404 259054 510004 294498
rect 509404 258818 509586 259054
rect 509822 258818 510004 259054
rect 509404 258734 510004 258818
rect 509404 258498 509586 258734
rect 509822 258498 510004 258734
rect 509404 223054 510004 258498
rect 509404 222818 509586 223054
rect 509822 222818 510004 223054
rect 509404 222734 510004 222818
rect 509404 222498 509586 222734
rect 509822 222498 510004 222734
rect 509404 187054 510004 222498
rect 509404 186818 509586 187054
rect 509822 186818 510004 187054
rect 509404 186734 510004 186818
rect 509404 186498 509586 186734
rect 509822 186498 510004 186734
rect 509404 151054 510004 186498
rect 509404 150818 509586 151054
rect 509822 150818 510004 151054
rect 509404 150734 510004 150818
rect 509404 150498 509586 150734
rect 509822 150498 510004 150734
rect 509404 115054 510004 150498
rect 509404 114818 509586 115054
rect 509822 114818 510004 115054
rect 509404 114734 510004 114818
rect 509404 114498 509586 114734
rect 509822 114498 510004 114734
rect 509404 79054 510004 114498
rect 509404 78818 509586 79054
rect 509822 78818 510004 79054
rect 509404 78734 510004 78818
rect 509404 78498 509586 78734
rect 509822 78498 510004 78734
rect 509404 43054 510004 78498
rect 509404 42818 509586 43054
rect 509822 42818 510004 43054
rect 509404 42734 510004 42818
rect 509404 42498 509586 42734
rect 509822 42498 510004 42734
rect 509404 7054 510004 42498
rect 509404 6818 509586 7054
rect 509822 6818 510004 7054
rect 509404 6734 510004 6818
rect 509404 6498 509586 6734
rect 509822 6498 510004 6734
rect 509404 -2226 510004 6498
rect 509404 -2462 509586 -2226
rect 509822 -2462 510004 -2226
rect 509404 -2546 510004 -2462
rect 509404 -2782 509586 -2546
rect 509822 -2782 510004 -2546
rect 509404 -3744 510004 -2782
rect 513004 694654 513604 708042
rect 513004 694418 513186 694654
rect 513422 694418 513604 694654
rect 513004 694334 513604 694418
rect 513004 694098 513186 694334
rect 513422 694098 513604 694334
rect 513004 658654 513604 694098
rect 513004 658418 513186 658654
rect 513422 658418 513604 658654
rect 513004 658334 513604 658418
rect 513004 658098 513186 658334
rect 513422 658098 513604 658334
rect 513004 622654 513604 658098
rect 513004 622418 513186 622654
rect 513422 622418 513604 622654
rect 513004 622334 513604 622418
rect 513004 622098 513186 622334
rect 513422 622098 513604 622334
rect 513004 586654 513604 622098
rect 513004 586418 513186 586654
rect 513422 586418 513604 586654
rect 513004 586334 513604 586418
rect 513004 586098 513186 586334
rect 513422 586098 513604 586334
rect 513004 550654 513604 586098
rect 513004 550418 513186 550654
rect 513422 550418 513604 550654
rect 513004 550334 513604 550418
rect 513004 550098 513186 550334
rect 513422 550098 513604 550334
rect 513004 514654 513604 550098
rect 513004 514418 513186 514654
rect 513422 514418 513604 514654
rect 513004 514334 513604 514418
rect 513004 514098 513186 514334
rect 513422 514098 513604 514334
rect 513004 478654 513604 514098
rect 513004 478418 513186 478654
rect 513422 478418 513604 478654
rect 513004 478334 513604 478418
rect 513004 478098 513186 478334
rect 513422 478098 513604 478334
rect 513004 442654 513604 478098
rect 513004 442418 513186 442654
rect 513422 442418 513604 442654
rect 513004 442334 513604 442418
rect 513004 442098 513186 442334
rect 513422 442098 513604 442334
rect 513004 406654 513604 442098
rect 513004 406418 513186 406654
rect 513422 406418 513604 406654
rect 513004 406334 513604 406418
rect 513004 406098 513186 406334
rect 513422 406098 513604 406334
rect 513004 370654 513604 406098
rect 513004 370418 513186 370654
rect 513422 370418 513604 370654
rect 513004 370334 513604 370418
rect 513004 370098 513186 370334
rect 513422 370098 513604 370334
rect 513004 334654 513604 370098
rect 513004 334418 513186 334654
rect 513422 334418 513604 334654
rect 513004 334334 513604 334418
rect 513004 334098 513186 334334
rect 513422 334098 513604 334334
rect 513004 298654 513604 334098
rect 513004 298418 513186 298654
rect 513422 298418 513604 298654
rect 513004 298334 513604 298418
rect 513004 298098 513186 298334
rect 513422 298098 513604 298334
rect 513004 262654 513604 298098
rect 513004 262418 513186 262654
rect 513422 262418 513604 262654
rect 513004 262334 513604 262418
rect 513004 262098 513186 262334
rect 513422 262098 513604 262334
rect 513004 226654 513604 262098
rect 513004 226418 513186 226654
rect 513422 226418 513604 226654
rect 513004 226334 513604 226418
rect 513004 226098 513186 226334
rect 513422 226098 513604 226334
rect 513004 190654 513604 226098
rect 513004 190418 513186 190654
rect 513422 190418 513604 190654
rect 513004 190334 513604 190418
rect 513004 190098 513186 190334
rect 513422 190098 513604 190334
rect 513004 154654 513604 190098
rect 513004 154418 513186 154654
rect 513422 154418 513604 154654
rect 513004 154334 513604 154418
rect 513004 154098 513186 154334
rect 513422 154098 513604 154334
rect 513004 118654 513604 154098
rect 513004 118418 513186 118654
rect 513422 118418 513604 118654
rect 513004 118334 513604 118418
rect 513004 118098 513186 118334
rect 513422 118098 513604 118334
rect 513004 82654 513604 118098
rect 513004 82418 513186 82654
rect 513422 82418 513604 82654
rect 513004 82334 513604 82418
rect 513004 82098 513186 82334
rect 513422 82098 513604 82334
rect 513004 46654 513604 82098
rect 513004 46418 513186 46654
rect 513422 46418 513604 46654
rect 513004 46334 513604 46418
rect 513004 46098 513186 46334
rect 513422 46098 513604 46334
rect 513004 10654 513604 46098
rect 513004 10418 513186 10654
rect 513422 10418 513604 10654
rect 513004 10334 513604 10418
rect 513004 10098 513186 10334
rect 513422 10098 513604 10334
rect 513004 -4106 513604 10098
rect 513004 -4342 513186 -4106
rect 513422 -4342 513604 -4106
rect 513004 -4426 513604 -4342
rect 513004 -4662 513186 -4426
rect 513422 -4662 513604 -4426
rect 513004 -5624 513604 -4662
rect 516604 698254 517204 709922
rect 534604 711418 535204 711440
rect 534604 711182 534786 711418
rect 535022 711182 535204 711418
rect 534604 711098 535204 711182
rect 534604 710862 534786 711098
rect 535022 710862 535204 711098
rect 531004 709538 531604 709560
rect 531004 709302 531186 709538
rect 531422 709302 531604 709538
rect 531004 709218 531604 709302
rect 531004 708982 531186 709218
rect 531422 708982 531604 709218
rect 527404 707658 528004 707680
rect 527404 707422 527586 707658
rect 527822 707422 528004 707658
rect 527404 707338 528004 707422
rect 527404 707102 527586 707338
rect 527822 707102 528004 707338
rect 516604 698018 516786 698254
rect 517022 698018 517204 698254
rect 516604 697934 517204 698018
rect 516604 697698 516786 697934
rect 517022 697698 517204 697934
rect 516604 662254 517204 697698
rect 516604 662018 516786 662254
rect 517022 662018 517204 662254
rect 516604 661934 517204 662018
rect 516604 661698 516786 661934
rect 517022 661698 517204 661934
rect 516604 626254 517204 661698
rect 516604 626018 516786 626254
rect 517022 626018 517204 626254
rect 516604 625934 517204 626018
rect 516604 625698 516786 625934
rect 517022 625698 517204 625934
rect 516604 590254 517204 625698
rect 516604 590018 516786 590254
rect 517022 590018 517204 590254
rect 516604 589934 517204 590018
rect 516604 589698 516786 589934
rect 517022 589698 517204 589934
rect 516604 554254 517204 589698
rect 516604 554018 516786 554254
rect 517022 554018 517204 554254
rect 516604 553934 517204 554018
rect 516604 553698 516786 553934
rect 517022 553698 517204 553934
rect 516604 518254 517204 553698
rect 516604 518018 516786 518254
rect 517022 518018 517204 518254
rect 516604 517934 517204 518018
rect 516604 517698 516786 517934
rect 517022 517698 517204 517934
rect 516604 482254 517204 517698
rect 516604 482018 516786 482254
rect 517022 482018 517204 482254
rect 516604 481934 517204 482018
rect 516604 481698 516786 481934
rect 517022 481698 517204 481934
rect 516604 446254 517204 481698
rect 516604 446018 516786 446254
rect 517022 446018 517204 446254
rect 516604 445934 517204 446018
rect 516604 445698 516786 445934
rect 517022 445698 517204 445934
rect 516604 410254 517204 445698
rect 516604 410018 516786 410254
rect 517022 410018 517204 410254
rect 516604 409934 517204 410018
rect 516604 409698 516786 409934
rect 517022 409698 517204 409934
rect 516604 374254 517204 409698
rect 516604 374018 516786 374254
rect 517022 374018 517204 374254
rect 516604 373934 517204 374018
rect 516604 373698 516786 373934
rect 517022 373698 517204 373934
rect 516604 338254 517204 373698
rect 516604 338018 516786 338254
rect 517022 338018 517204 338254
rect 516604 337934 517204 338018
rect 516604 337698 516786 337934
rect 517022 337698 517204 337934
rect 516604 302254 517204 337698
rect 516604 302018 516786 302254
rect 517022 302018 517204 302254
rect 516604 301934 517204 302018
rect 516604 301698 516786 301934
rect 517022 301698 517204 301934
rect 516604 266254 517204 301698
rect 516604 266018 516786 266254
rect 517022 266018 517204 266254
rect 516604 265934 517204 266018
rect 516604 265698 516786 265934
rect 517022 265698 517204 265934
rect 516604 230254 517204 265698
rect 516604 230018 516786 230254
rect 517022 230018 517204 230254
rect 516604 229934 517204 230018
rect 516604 229698 516786 229934
rect 517022 229698 517204 229934
rect 516604 194254 517204 229698
rect 516604 194018 516786 194254
rect 517022 194018 517204 194254
rect 516604 193934 517204 194018
rect 516604 193698 516786 193934
rect 517022 193698 517204 193934
rect 516604 158254 517204 193698
rect 516604 158018 516786 158254
rect 517022 158018 517204 158254
rect 516604 157934 517204 158018
rect 516604 157698 516786 157934
rect 517022 157698 517204 157934
rect 516604 122254 517204 157698
rect 516604 122018 516786 122254
rect 517022 122018 517204 122254
rect 516604 121934 517204 122018
rect 516604 121698 516786 121934
rect 517022 121698 517204 121934
rect 516604 86254 517204 121698
rect 516604 86018 516786 86254
rect 517022 86018 517204 86254
rect 516604 85934 517204 86018
rect 516604 85698 516786 85934
rect 517022 85698 517204 85934
rect 516604 50254 517204 85698
rect 516604 50018 516786 50254
rect 517022 50018 517204 50254
rect 516604 49934 517204 50018
rect 516604 49698 516786 49934
rect 517022 49698 517204 49934
rect 516604 14254 517204 49698
rect 516604 14018 516786 14254
rect 517022 14018 517204 14254
rect 516604 13934 517204 14018
rect 516604 13698 516786 13934
rect 517022 13698 517204 13934
rect 498604 -7162 498786 -6926
rect 499022 -7162 499204 -6926
rect 498604 -7246 499204 -7162
rect 498604 -7482 498786 -7246
rect 499022 -7482 499204 -7246
rect 498604 -7504 499204 -7482
rect 516604 -5986 517204 13698
rect 523804 705778 524404 705800
rect 523804 705542 523986 705778
rect 524222 705542 524404 705778
rect 523804 705458 524404 705542
rect 523804 705222 523986 705458
rect 524222 705222 524404 705458
rect 523804 669454 524404 705222
rect 523804 669218 523986 669454
rect 524222 669218 524404 669454
rect 523804 669134 524404 669218
rect 523804 668898 523986 669134
rect 524222 668898 524404 669134
rect 523804 633454 524404 668898
rect 523804 633218 523986 633454
rect 524222 633218 524404 633454
rect 523804 633134 524404 633218
rect 523804 632898 523986 633134
rect 524222 632898 524404 633134
rect 523804 597454 524404 632898
rect 523804 597218 523986 597454
rect 524222 597218 524404 597454
rect 523804 597134 524404 597218
rect 523804 596898 523986 597134
rect 524222 596898 524404 597134
rect 523804 561454 524404 596898
rect 523804 561218 523986 561454
rect 524222 561218 524404 561454
rect 523804 561134 524404 561218
rect 523804 560898 523986 561134
rect 524222 560898 524404 561134
rect 523804 525454 524404 560898
rect 523804 525218 523986 525454
rect 524222 525218 524404 525454
rect 523804 525134 524404 525218
rect 523804 524898 523986 525134
rect 524222 524898 524404 525134
rect 523804 489454 524404 524898
rect 523804 489218 523986 489454
rect 524222 489218 524404 489454
rect 523804 489134 524404 489218
rect 523804 488898 523986 489134
rect 524222 488898 524404 489134
rect 523804 453454 524404 488898
rect 523804 453218 523986 453454
rect 524222 453218 524404 453454
rect 523804 453134 524404 453218
rect 523804 452898 523986 453134
rect 524222 452898 524404 453134
rect 523804 417454 524404 452898
rect 523804 417218 523986 417454
rect 524222 417218 524404 417454
rect 523804 417134 524404 417218
rect 523804 416898 523986 417134
rect 524222 416898 524404 417134
rect 523804 381454 524404 416898
rect 523804 381218 523986 381454
rect 524222 381218 524404 381454
rect 523804 381134 524404 381218
rect 523804 380898 523986 381134
rect 524222 380898 524404 381134
rect 523804 345454 524404 380898
rect 523804 345218 523986 345454
rect 524222 345218 524404 345454
rect 523804 345134 524404 345218
rect 523804 344898 523986 345134
rect 524222 344898 524404 345134
rect 523804 309454 524404 344898
rect 523804 309218 523986 309454
rect 524222 309218 524404 309454
rect 523804 309134 524404 309218
rect 523804 308898 523986 309134
rect 524222 308898 524404 309134
rect 523804 273454 524404 308898
rect 523804 273218 523986 273454
rect 524222 273218 524404 273454
rect 523804 273134 524404 273218
rect 523804 272898 523986 273134
rect 524222 272898 524404 273134
rect 523804 237454 524404 272898
rect 523804 237218 523986 237454
rect 524222 237218 524404 237454
rect 523804 237134 524404 237218
rect 523804 236898 523986 237134
rect 524222 236898 524404 237134
rect 523804 201454 524404 236898
rect 523804 201218 523986 201454
rect 524222 201218 524404 201454
rect 523804 201134 524404 201218
rect 523804 200898 523986 201134
rect 524222 200898 524404 201134
rect 523804 165454 524404 200898
rect 523804 165218 523986 165454
rect 524222 165218 524404 165454
rect 523804 165134 524404 165218
rect 523804 164898 523986 165134
rect 524222 164898 524404 165134
rect 523804 129454 524404 164898
rect 523804 129218 523986 129454
rect 524222 129218 524404 129454
rect 523804 129134 524404 129218
rect 523804 128898 523986 129134
rect 524222 128898 524404 129134
rect 523804 93454 524404 128898
rect 523804 93218 523986 93454
rect 524222 93218 524404 93454
rect 523804 93134 524404 93218
rect 523804 92898 523986 93134
rect 524222 92898 524404 93134
rect 523804 57454 524404 92898
rect 523804 57218 523986 57454
rect 524222 57218 524404 57454
rect 523804 57134 524404 57218
rect 523804 56898 523986 57134
rect 524222 56898 524404 57134
rect 523804 21454 524404 56898
rect 523804 21218 523986 21454
rect 524222 21218 524404 21454
rect 523804 21134 524404 21218
rect 523804 20898 523986 21134
rect 524222 20898 524404 21134
rect 523804 -1286 524404 20898
rect 523804 -1522 523986 -1286
rect 524222 -1522 524404 -1286
rect 523804 -1606 524404 -1522
rect 523804 -1842 523986 -1606
rect 524222 -1842 524404 -1606
rect 523804 -1864 524404 -1842
rect 527404 673054 528004 707102
rect 527404 672818 527586 673054
rect 527822 672818 528004 673054
rect 527404 672734 528004 672818
rect 527404 672498 527586 672734
rect 527822 672498 528004 672734
rect 527404 637054 528004 672498
rect 527404 636818 527586 637054
rect 527822 636818 528004 637054
rect 527404 636734 528004 636818
rect 527404 636498 527586 636734
rect 527822 636498 528004 636734
rect 527404 601054 528004 636498
rect 527404 600818 527586 601054
rect 527822 600818 528004 601054
rect 527404 600734 528004 600818
rect 527404 600498 527586 600734
rect 527822 600498 528004 600734
rect 527404 565054 528004 600498
rect 527404 564818 527586 565054
rect 527822 564818 528004 565054
rect 527404 564734 528004 564818
rect 527404 564498 527586 564734
rect 527822 564498 528004 564734
rect 527404 529054 528004 564498
rect 527404 528818 527586 529054
rect 527822 528818 528004 529054
rect 527404 528734 528004 528818
rect 527404 528498 527586 528734
rect 527822 528498 528004 528734
rect 527404 493054 528004 528498
rect 527404 492818 527586 493054
rect 527822 492818 528004 493054
rect 527404 492734 528004 492818
rect 527404 492498 527586 492734
rect 527822 492498 528004 492734
rect 527404 457054 528004 492498
rect 527404 456818 527586 457054
rect 527822 456818 528004 457054
rect 527404 456734 528004 456818
rect 527404 456498 527586 456734
rect 527822 456498 528004 456734
rect 527404 421054 528004 456498
rect 527404 420818 527586 421054
rect 527822 420818 528004 421054
rect 527404 420734 528004 420818
rect 527404 420498 527586 420734
rect 527822 420498 528004 420734
rect 527404 385054 528004 420498
rect 527404 384818 527586 385054
rect 527822 384818 528004 385054
rect 527404 384734 528004 384818
rect 527404 384498 527586 384734
rect 527822 384498 528004 384734
rect 527404 349054 528004 384498
rect 527404 348818 527586 349054
rect 527822 348818 528004 349054
rect 527404 348734 528004 348818
rect 527404 348498 527586 348734
rect 527822 348498 528004 348734
rect 527404 313054 528004 348498
rect 527404 312818 527586 313054
rect 527822 312818 528004 313054
rect 527404 312734 528004 312818
rect 527404 312498 527586 312734
rect 527822 312498 528004 312734
rect 527404 277054 528004 312498
rect 527404 276818 527586 277054
rect 527822 276818 528004 277054
rect 527404 276734 528004 276818
rect 527404 276498 527586 276734
rect 527822 276498 528004 276734
rect 527404 241054 528004 276498
rect 527404 240818 527586 241054
rect 527822 240818 528004 241054
rect 527404 240734 528004 240818
rect 527404 240498 527586 240734
rect 527822 240498 528004 240734
rect 527404 205054 528004 240498
rect 527404 204818 527586 205054
rect 527822 204818 528004 205054
rect 527404 204734 528004 204818
rect 527404 204498 527586 204734
rect 527822 204498 528004 204734
rect 527404 169054 528004 204498
rect 527404 168818 527586 169054
rect 527822 168818 528004 169054
rect 527404 168734 528004 168818
rect 527404 168498 527586 168734
rect 527822 168498 528004 168734
rect 527404 133054 528004 168498
rect 527404 132818 527586 133054
rect 527822 132818 528004 133054
rect 527404 132734 528004 132818
rect 527404 132498 527586 132734
rect 527822 132498 528004 132734
rect 527404 97054 528004 132498
rect 527404 96818 527586 97054
rect 527822 96818 528004 97054
rect 527404 96734 528004 96818
rect 527404 96498 527586 96734
rect 527822 96498 528004 96734
rect 527404 61054 528004 96498
rect 527404 60818 527586 61054
rect 527822 60818 528004 61054
rect 527404 60734 528004 60818
rect 527404 60498 527586 60734
rect 527822 60498 528004 60734
rect 527404 25054 528004 60498
rect 527404 24818 527586 25054
rect 527822 24818 528004 25054
rect 527404 24734 528004 24818
rect 527404 24498 527586 24734
rect 527822 24498 528004 24734
rect 527404 -3166 528004 24498
rect 527404 -3402 527586 -3166
rect 527822 -3402 528004 -3166
rect 527404 -3486 528004 -3402
rect 527404 -3722 527586 -3486
rect 527822 -3722 528004 -3486
rect 527404 -3744 528004 -3722
rect 531004 676654 531604 708982
rect 531004 676418 531186 676654
rect 531422 676418 531604 676654
rect 531004 676334 531604 676418
rect 531004 676098 531186 676334
rect 531422 676098 531604 676334
rect 531004 640654 531604 676098
rect 531004 640418 531186 640654
rect 531422 640418 531604 640654
rect 531004 640334 531604 640418
rect 531004 640098 531186 640334
rect 531422 640098 531604 640334
rect 531004 604654 531604 640098
rect 531004 604418 531186 604654
rect 531422 604418 531604 604654
rect 531004 604334 531604 604418
rect 531004 604098 531186 604334
rect 531422 604098 531604 604334
rect 531004 568654 531604 604098
rect 531004 568418 531186 568654
rect 531422 568418 531604 568654
rect 531004 568334 531604 568418
rect 531004 568098 531186 568334
rect 531422 568098 531604 568334
rect 531004 532654 531604 568098
rect 531004 532418 531186 532654
rect 531422 532418 531604 532654
rect 531004 532334 531604 532418
rect 531004 532098 531186 532334
rect 531422 532098 531604 532334
rect 531004 496654 531604 532098
rect 531004 496418 531186 496654
rect 531422 496418 531604 496654
rect 531004 496334 531604 496418
rect 531004 496098 531186 496334
rect 531422 496098 531604 496334
rect 531004 460654 531604 496098
rect 531004 460418 531186 460654
rect 531422 460418 531604 460654
rect 531004 460334 531604 460418
rect 531004 460098 531186 460334
rect 531422 460098 531604 460334
rect 531004 424654 531604 460098
rect 531004 424418 531186 424654
rect 531422 424418 531604 424654
rect 531004 424334 531604 424418
rect 531004 424098 531186 424334
rect 531422 424098 531604 424334
rect 531004 388654 531604 424098
rect 531004 388418 531186 388654
rect 531422 388418 531604 388654
rect 531004 388334 531604 388418
rect 531004 388098 531186 388334
rect 531422 388098 531604 388334
rect 531004 352654 531604 388098
rect 531004 352418 531186 352654
rect 531422 352418 531604 352654
rect 531004 352334 531604 352418
rect 531004 352098 531186 352334
rect 531422 352098 531604 352334
rect 531004 316654 531604 352098
rect 531004 316418 531186 316654
rect 531422 316418 531604 316654
rect 531004 316334 531604 316418
rect 531004 316098 531186 316334
rect 531422 316098 531604 316334
rect 531004 280654 531604 316098
rect 531004 280418 531186 280654
rect 531422 280418 531604 280654
rect 531004 280334 531604 280418
rect 531004 280098 531186 280334
rect 531422 280098 531604 280334
rect 531004 244654 531604 280098
rect 531004 244418 531186 244654
rect 531422 244418 531604 244654
rect 531004 244334 531604 244418
rect 531004 244098 531186 244334
rect 531422 244098 531604 244334
rect 531004 208654 531604 244098
rect 531004 208418 531186 208654
rect 531422 208418 531604 208654
rect 531004 208334 531604 208418
rect 531004 208098 531186 208334
rect 531422 208098 531604 208334
rect 531004 172654 531604 208098
rect 531004 172418 531186 172654
rect 531422 172418 531604 172654
rect 531004 172334 531604 172418
rect 531004 172098 531186 172334
rect 531422 172098 531604 172334
rect 531004 136654 531604 172098
rect 531004 136418 531186 136654
rect 531422 136418 531604 136654
rect 531004 136334 531604 136418
rect 531004 136098 531186 136334
rect 531422 136098 531604 136334
rect 531004 100654 531604 136098
rect 531004 100418 531186 100654
rect 531422 100418 531604 100654
rect 531004 100334 531604 100418
rect 531004 100098 531186 100334
rect 531422 100098 531604 100334
rect 531004 64654 531604 100098
rect 531004 64418 531186 64654
rect 531422 64418 531604 64654
rect 531004 64334 531604 64418
rect 531004 64098 531186 64334
rect 531422 64098 531604 64334
rect 531004 28654 531604 64098
rect 531004 28418 531186 28654
rect 531422 28418 531604 28654
rect 531004 28334 531604 28418
rect 531004 28098 531186 28334
rect 531422 28098 531604 28334
rect 531004 -5046 531604 28098
rect 531004 -5282 531186 -5046
rect 531422 -5282 531604 -5046
rect 531004 -5366 531604 -5282
rect 531004 -5602 531186 -5366
rect 531422 -5602 531604 -5366
rect 531004 -5624 531604 -5602
rect 534604 680254 535204 710862
rect 552604 710478 553204 711440
rect 552604 710242 552786 710478
rect 553022 710242 553204 710478
rect 552604 710158 553204 710242
rect 552604 709922 552786 710158
rect 553022 709922 553204 710158
rect 549004 708598 549604 709560
rect 549004 708362 549186 708598
rect 549422 708362 549604 708598
rect 549004 708278 549604 708362
rect 549004 708042 549186 708278
rect 549422 708042 549604 708278
rect 545404 706718 546004 707680
rect 545404 706482 545586 706718
rect 545822 706482 546004 706718
rect 545404 706398 546004 706482
rect 545404 706162 545586 706398
rect 545822 706162 546004 706398
rect 534604 680018 534786 680254
rect 535022 680018 535204 680254
rect 534604 679934 535204 680018
rect 534604 679698 534786 679934
rect 535022 679698 535204 679934
rect 534604 644254 535204 679698
rect 534604 644018 534786 644254
rect 535022 644018 535204 644254
rect 534604 643934 535204 644018
rect 534604 643698 534786 643934
rect 535022 643698 535204 643934
rect 534604 608254 535204 643698
rect 534604 608018 534786 608254
rect 535022 608018 535204 608254
rect 534604 607934 535204 608018
rect 534604 607698 534786 607934
rect 535022 607698 535204 607934
rect 534604 572254 535204 607698
rect 534604 572018 534786 572254
rect 535022 572018 535204 572254
rect 534604 571934 535204 572018
rect 534604 571698 534786 571934
rect 535022 571698 535204 571934
rect 534604 536254 535204 571698
rect 534604 536018 534786 536254
rect 535022 536018 535204 536254
rect 534604 535934 535204 536018
rect 534604 535698 534786 535934
rect 535022 535698 535204 535934
rect 534604 500254 535204 535698
rect 534604 500018 534786 500254
rect 535022 500018 535204 500254
rect 534604 499934 535204 500018
rect 534604 499698 534786 499934
rect 535022 499698 535204 499934
rect 534604 464254 535204 499698
rect 534604 464018 534786 464254
rect 535022 464018 535204 464254
rect 534604 463934 535204 464018
rect 534604 463698 534786 463934
rect 535022 463698 535204 463934
rect 534604 428254 535204 463698
rect 534604 428018 534786 428254
rect 535022 428018 535204 428254
rect 534604 427934 535204 428018
rect 534604 427698 534786 427934
rect 535022 427698 535204 427934
rect 534604 392254 535204 427698
rect 534604 392018 534786 392254
rect 535022 392018 535204 392254
rect 534604 391934 535204 392018
rect 534604 391698 534786 391934
rect 535022 391698 535204 391934
rect 534604 356254 535204 391698
rect 534604 356018 534786 356254
rect 535022 356018 535204 356254
rect 534604 355934 535204 356018
rect 534604 355698 534786 355934
rect 535022 355698 535204 355934
rect 534604 320254 535204 355698
rect 534604 320018 534786 320254
rect 535022 320018 535204 320254
rect 534604 319934 535204 320018
rect 534604 319698 534786 319934
rect 535022 319698 535204 319934
rect 534604 284254 535204 319698
rect 534604 284018 534786 284254
rect 535022 284018 535204 284254
rect 534604 283934 535204 284018
rect 534604 283698 534786 283934
rect 535022 283698 535204 283934
rect 534604 248254 535204 283698
rect 534604 248018 534786 248254
rect 535022 248018 535204 248254
rect 534604 247934 535204 248018
rect 534604 247698 534786 247934
rect 535022 247698 535204 247934
rect 534604 212254 535204 247698
rect 534604 212018 534786 212254
rect 535022 212018 535204 212254
rect 534604 211934 535204 212018
rect 534604 211698 534786 211934
rect 535022 211698 535204 211934
rect 534604 176254 535204 211698
rect 534604 176018 534786 176254
rect 535022 176018 535204 176254
rect 534604 175934 535204 176018
rect 534604 175698 534786 175934
rect 535022 175698 535204 175934
rect 534604 140254 535204 175698
rect 534604 140018 534786 140254
rect 535022 140018 535204 140254
rect 534604 139934 535204 140018
rect 534604 139698 534786 139934
rect 535022 139698 535204 139934
rect 534604 104254 535204 139698
rect 534604 104018 534786 104254
rect 535022 104018 535204 104254
rect 534604 103934 535204 104018
rect 534604 103698 534786 103934
rect 535022 103698 535204 103934
rect 534604 68254 535204 103698
rect 534604 68018 534786 68254
rect 535022 68018 535204 68254
rect 534604 67934 535204 68018
rect 534604 67698 534786 67934
rect 535022 67698 535204 67934
rect 534604 32254 535204 67698
rect 534604 32018 534786 32254
rect 535022 32018 535204 32254
rect 534604 31934 535204 32018
rect 534604 31698 534786 31934
rect 535022 31698 535204 31934
rect 516604 -6222 516786 -5986
rect 517022 -6222 517204 -5986
rect 516604 -6306 517204 -6222
rect 516604 -6542 516786 -6306
rect 517022 -6542 517204 -6306
rect 516604 -7504 517204 -6542
rect 534604 -6926 535204 31698
rect 541804 704838 542404 705800
rect 541804 704602 541986 704838
rect 542222 704602 542404 704838
rect 541804 704518 542404 704602
rect 541804 704282 541986 704518
rect 542222 704282 542404 704518
rect 541804 687454 542404 704282
rect 541804 687218 541986 687454
rect 542222 687218 542404 687454
rect 541804 687134 542404 687218
rect 541804 686898 541986 687134
rect 542222 686898 542404 687134
rect 541804 651454 542404 686898
rect 541804 651218 541986 651454
rect 542222 651218 542404 651454
rect 541804 651134 542404 651218
rect 541804 650898 541986 651134
rect 542222 650898 542404 651134
rect 541804 615454 542404 650898
rect 541804 615218 541986 615454
rect 542222 615218 542404 615454
rect 541804 615134 542404 615218
rect 541804 614898 541986 615134
rect 542222 614898 542404 615134
rect 541804 579454 542404 614898
rect 541804 579218 541986 579454
rect 542222 579218 542404 579454
rect 541804 579134 542404 579218
rect 541804 578898 541986 579134
rect 542222 578898 542404 579134
rect 541804 543454 542404 578898
rect 541804 543218 541986 543454
rect 542222 543218 542404 543454
rect 541804 543134 542404 543218
rect 541804 542898 541986 543134
rect 542222 542898 542404 543134
rect 541804 507454 542404 542898
rect 541804 507218 541986 507454
rect 542222 507218 542404 507454
rect 541804 507134 542404 507218
rect 541804 506898 541986 507134
rect 542222 506898 542404 507134
rect 541804 471454 542404 506898
rect 541804 471218 541986 471454
rect 542222 471218 542404 471454
rect 541804 471134 542404 471218
rect 541804 470898 541986 471134
rect 542222 470898 542404 471134
rect 541804 435454 542404 470898
rect 541804 435218 541986 435454
rect 542222 435218 542404 435454
rect 541804 435134 542404 435218
rect 541804 434898 541986 435134
rect 542222 434898 542404 435134
rect 541804 399454 542404 434898
rect 541804 399218 541986 399454
rect 542222 399218 542404 399454
rect 541804 399134 542404 399218
rect 541804 398898 541986 399134
rect 542222 398898 542404 399134
rect 541804 363454 542404 398898
rect 541804 363218 541986 363454
rect 542222 363218 542404 363454
rect 541804 363134 542404 363218
rect 541804 362898 541986 363134
rect 542222 362898 542404 363134
rect 541804 327454 542404 362898
rect 541804 327218 541986 327454
rect 542222 327218 542404 327454
rect 541804 327134 542404 327218
rect 541804 326898 541986 327134
rect 542222 326898 542404 327134
rect 541804 291454 542404 326898
rect 541804 291218 541986 291454
rect 542222 291218 542404 291454
rect 541804 291134 542404 291218
rect 541804 290898 541986 291134
rect 542222 290898 542404 291134
rect 541804 255454 542404 290898
rect 541804 255218 541986 255454
rect 542222 255218 542404 255454
rect 541804 255134 542404 255218
rect 541804 254898 541986 255134
rect 542222 254898 542404 255134
rect 541804 219454 542404 254898
rect 541804 219218 541986 219454
rect 542222 219218 542404 219454
rect 541804 219134 542404 219218
rect 541804 218898 541986 219134
rect 542222 218898 542404 219134
rect 541804 183454 542404 218898
rect 541804 183218 541986 183454
rect 542222 183218 542404 183454
rect 541804 183134 542404 183218
rect 541804 182898 541986 183134
rect 542222 182898 542404 183134
rect 541804 147454 542404 182898
rect 541804 147218 541986 147454
rect 542222 147218 542404 147454
rect 541804 147134 542404 147218
rect 541804 146898 541986 147134
rect 542222 146898 542404 147134
rect 541804 111454 542404 146898
rect 541804 111218 541986 111454
rect 542222 111218 542404 111454
rect 541804 111134 542404 111218
rect 541804 110898 541986 111134
rect 542222 110898 542404 111134
rect 541804 75454 542404 110898
rect 541804 75218 541986 75454
rect 542222 75218 542404 75454
rect 541804 75134 542404 75218
rect 541804 74898 541986 75134
rect 542222 74898 542404 75134
rect 541804 39454 542404 74898
rect 541804 39218 541986 39454
rect 542222 39218 542404 39454
rect 541804 39134 542404 39218
rect 541804 38898 541986 39134
rect 542222 38898 542404 39134
rect 541804 3454 542404 38898
rect 541804 3218 541986 3454
rect 542222 3218 542404 3454
rect 541804 3134 542404 3218
rect 541804 2898 541986 3134
rect 542222 2898 542404 3134
rect 541804 -346 542404 2898
rect 541804 -582 541986 -346
rect 542222 -582 542404 -346
rect 541804 -666 542404 -582
rect 541804 -902 541986 -666
rect 542222 -902 542404 -666
rect 541804 -1864 542404 -902
rect 545404 691054 546004 706162
rect 545404 690818 545586 691054
rect 545822 690818 546004 691054
rect 545404 690734 546004 690818
rect 545404 690498 545586 690734
rect 545822 690498 546004 690734
rect 545404 655054 546004 690498
rect 545404 654818 545586 655054
rect 545822 654818 546004 655054
rect 545404 654734 546004 654818
rect 545404 654498 545586 654734
rect 545822 654498 546004 654734
rect 545404 619054 546004 654498
rect 545404 618818 545586 619054
rect 545822 618818 546004 619054
rect 545404 618734 546004 618818
rect 545404 618498 545586 618734
rect 545822 618498 546004 618734
rect 545404 583054 546004 618498
rect 545404 582818 545586 583054
rect 545822 582818 546004 583054
rect 545404 582734 546004 582818
rect 545404 582498 545586 582734
rect 545822 582498 546004 582734
rect 545404 547054 546004 582498
rect 545404 546818 545586 547054
rect 545822 546818 546004 547054
rect 545404 546734 546004 546818
rect 545404 546498 545586 546734
rect 545822 546498 546004 546734
rect 545404 511054 546004 546498
rect 545404 510818 545586 511054
rect 545822 510818 546004 511054
rect 545404 510734 546004 510818
rect 545404 510498 545586 510734
rect 545822 510498 546004 510734
rect 545404 475054 546004 510498
rect 545404 474818 545586 475054
rect 545822 474818 546004 475054
rect 545404 474734 546004 474818
rect 545404 474498 545586 474734
rect 545822 474498 546004 474734
rect 545404 439054 546004 474498
rect 545404 438818 545586 439054
rect 545822 438818 546004 439054
rect 545404 438734 546004 438818
rect 545404 438498 545586 438734
rect 545822 438498 546004 438734
rect 545404 403054 546004 438498
rect 545404 402818 545586 403054
rect 545822 402818 546004 403054
rect 545404 402734 546004 402818
rect 545404 402498 545586 402734
rect 545822 402498 546004 402734
rect 545404 367054 546004 402498
rect 545404 366818 545586 367054
rect 545822 366818 546004 367054
rect 545404 366734 546004 366818
rect 545404 366498 545586 366734
rect 545822 366498 546004 366734
rect 545404 331054 546004 366498
rect 545404 330818 545586 331054
rect 545822 330818 546004 331054
rect 545404 330734 546004 330818
rect 545404 330498 545586 330734
rect 545822 330498 546004 330734
rect 545404 295054 546004 330498
rect 545404 294818 545586 295054
rect 545822 294818 546004 295054
rect 545404 294734 546004 294818
rect 545404 294498 545586 294734
rect 545822 294498 546004 294734
rect 545404 259054 546004 294498
rect 545404 258818 545586 259054
rect 545822 258818 546004 259054
rect 545404 258734 546004 258818
rect 545404 258498 545586 258734
rect 545822 258498 546004 258734
rect 545404 223054 546004 258498
rect 545404 222818 545586 223054
rect 545822 222818 546004 223054
rect 545404 222734 546004 222818
rect 545404 222498 545586 222734
rect 545822 222498 546004 222734
rect 545404 187054 546004 222498
rect 545404 186818 545586 187054
rect 545822 186818 546004 187054
rect 545404 186734 546004 186818
rect 545404 186498 545586 186734
rect 545822 186498 546004 186734
rect 545404 151054 546004 186498
rect 545404 150818 545586 151054
rect 545822 150818 546004 151054
rect 545404 150734 546004 150818
rect 545404 150498 545586 150734
rect 545822 150498 546004 150734
rect 545404 115054 546004 150498
rect 545404 114818 545586 115054
rect 545822 114818 546004 115054
rect 545404 114734 546004 114818
rect 545404 114498 545586 114734
rect 545822 114498 546004 114734
rect 545404 79054 546004 114498
rect 545404 78818 545586 79054
rect 545822 78818 546004 79054
rect 545404 78734 546004 78818
rect 545404 78498 545586 78734
rect 545822 78498 546004 78734
rect 545404 43054 546004 78498
rect 545404 42818 545586 43054
rect 545822 42818 546004 43054
rect 545404 42734 546004 42818
rect 545404 42498 545586 42734
rect 545822 42498 546004 42734
rect 545404 7054 546004 42498
rect 545404 6818 545586 7054
rect 545822 6818 546004 7054
rect 545404 6734 546004 6818
rect 545404 6498 545586 6734
rect 545822 6498 546004 6734
rect 545404 -2226 546004 6498
rect 545404 -2462 545586 -2226
rect 545822 -2462 546004 -2226
rect 545404 -2546 546004 -2462
rect 545404 -2782 545586 -2546
rect 545822 -2782 546004 -2546
rect 545404 -3744 546004 -2782
rect 549004 694654 549604 708042
rect 549004 694418 549186 694654
rect 549422 694418 549604 694654
rect 549004 694334 549604 694418
rect 549004 694098 549186 694334
rect 549422 694098 549604 694334
rect 549004 658654 549604 694098
rect 549004 658418 549186 658654
rect 549422 658418 549604 658654
rect 549004 658334 549604 658418
rect 549004 658098 549186 658334
rect 549422 658098 549604 658334
rect 549004 622654 549604 658098
rect 549004 622418 549186 622654
rect 549422 622418 549604 622654
rect 549004 622334 549604 622418
rect 549004 622098 549186 622334
rect 549422 622098 549604 622334
rect 549004 586654 549604 622098
rect 549004 586418 549186 586654
rect 549422 586418 549604 586654
rect 549004 586334 549604 586418
rect 549004 586098 549186 586334
rect 549422 586098 549604 586334
rect 549004 550654 549604 586098
rect 549004 550418 549186 550654
rect 549422 550418 549604 550654
rect 549004 550334 549604 550418
rect 549004 550098 549186 550334
rect 549422 550098 549604 550334
rect 549004 514654 549604 550098
rect 549004 514418 549186 514654
rect 549422 514418 549604 514654
rect 549004 514334 549604 514418
rect 549004 514098 549186 514334
rect 549422 514098 549604 514334
rect 549004 478654 549604 514098
rect 549004 478418 549186 478654
rect 549422 478418 549604 478654
rect 549004 478334 549604 478418
rect 549004 478098 549186 478334
rect 549422 478098 549604 478334
rect 549004 442654 549604 478098
rect 549004 442418 549186 442654
rect 549422 442418 549604 442654
rect 549004 442334 549604 442418
rect 549004 442098 549186 442334
rect 549422 442098 549604 442334
rect 549004 406654 549604 442098
rect 549004 406418 549186 406654
rect 549422 406418 549604 406654
rect 549004 406334 549604 406418
rect 549004 406098 549186 406334
rect 549422 406098 549604 406334
rect 549004 370654 549604 406098
rect 549004 370418 549186 370654
rect 549422 370418 549604 370654
rect 549004 370334 549604 370418
rect 549004 370098 549186 370334
rect 549422 370098 549604 370334
rect 549004 334654 549604 370098
rect 549004 334418 549186 334654
rect 549422 334418 549604 334654
rect 549004 334334 549604 334418
rect 549004 334098 549186 334334
rect 549422 334098 549604 334334
rect 549004 298654 549604 334098
rect 549004 298418 549186 298654
rect 549422 298418 549604 298654
rect 549004 298334 549604 298418
rect 549004 298098 549186 298334
rect 549422 298098 549604 298334
rect 549004 262654 549604 298098
rect 549004 262418 549186 262654
rect 549422 262418 549604 262654
rect 549004 262334 549604 262418
rect 549004 262098 549186 262334
rect 549422 262098 549604 262334
rect 549004 226654 549604 262098
rect 549004 226418 549186 226654
rect 549422 226418 549604 226654
rect 549004 226334 549604 226418
rect 549004 226098 549186 226334
rect 549422 226098 549604 226334
rect 549004 190654 549604 226098
rect 549004 190418 549186 190654
rect 549422 190418 549604 190654
rect 549004 190334 549604 190418
rect 549004 190098 549186 190334
rect 549422 190098 549604 190334
rect 549004 154654 549604 190098
rect 549004 154418 549186 154654
rect 549422 154418 549604 154654
rect 549004 154334 549604 154418
rect 549004 154098 549186 154334
rect 549422 154098 549604 154334
rect 549004 118654 549604 154098
rect 549004 118418 549186 118654
rect 549422 118418 549604 118654
rect 549004 118334 549604 118418
rect 549004 118098 549186 118334
rect 549422 118098 549604 118334
rect 549004 82654 549604 118098
rect 549004 82418 549186 82654
rect 549422 82418 549604 82654
rect 549004 82334 549604 82418
rect 549004 82098 549186 82334
rect 549422 82098 549604 82334
rect 549004 46654 549604 82098
rect 549004 46418 549186 46654
rect 549422 46418 549604 46654
rect 549004 46334 549604 46418
rect 549004 46098 549186 46334
rect 549422 46098 549604 46334
rect 549004 10654 549604 46098
rect 549004 10418 549186 10654
rect 549422 10418 549604 10654
rect 549004 10334 549604 10418
rect 549004 10098 549186 10334
rect 549422 10098 549604 10334
rect 549004 -4106 549604 10098
rect 549004 -4342 549186 -4106
rect 549422 -4342 549604 -4106
rect 549004 -4426 549604 -4342
rect 549004 -4662 549186 -4426
rect 549422 -4662 549604 -4426
rect 549004 -5624 549604 -4662
rect 552604 698254 553204 709922
rect 570604 711418 571204 711440
rect 570604 711182 570786 711418
rect 571022 711182 571204 711418
rect 570604 711098 571204 711182
rect 570604 710862 570786 711098
rect 571022 710862 571204 711098
rect 567004 709538 567604 709560
rect 567004 709302 567186 709538
rect 567422 709302 567604 709538
rect 567004 709218 567604 709302
rect 567004 708982 567186 709218
rect 567422 708982 567604 709218
rect 563404 707658 564004 707680
rect 563404 707422 563586 707658
rect 563822 707422 564004 707658
rect 563404 707338 564004 707422
rect 563404 707102 563586 707338
rect 563822 707102 564004 707338
rect 552604 698018 552786 698254
rect 553022 698018 553204 698254
rect 552604 697934 553204 698018
rect 552604 697698 552786 697934
rect 553022 697698 553204 697934
rect 552604 662254 553204 697698
rect 552604 662018 552786 662254
rect 553022 662018 553204 662254
rect 552604 661934 553204 662018
rect 552604 661698 552786 661934
rect 553022 661698 553204 661934
rect 552604 626254 553204 661698
rect 552604 626018 552786 626254
rect 553022 626018 553204 626254
rect 552604 625934 553204 626018
rect 552604 625698 552786 625934
rect 553022 625698 553204 625934
rect 552604 590254 553204 625698
rect 552604 590018 552786 590254
rect 553022 590018 553204 590254
rect 552604 589934 553204 590018
rect 552604 589698 552786 589934
rect 553022 589698 553204 589934
rect 552604 554254 553204 589698
rect 552604 554018 552786 554254
rect 553022 554018 553204 554254
rect 552604 553934 553204 554018
rect 552604 553698 552786 553934
rect 553022 553698 553204 553934
rect 552604 518254 553204 553698
rect 552604 518018 552786 518254
rect 553022 518018 553204 518254
rect 552604 517934 553204 518018
rect 552604 517698 552786 517934
rect 553022 517698 553204 517934
rect 552604 482254 553204 517698
rect 552604 482018 552786 482254
rect 553022 482018 553204 482254
rect 552604 481934 553204 482018
rect 552604 481698 552786 481934
rect 553022 481698 553204 481934
rect 552604 446254 553204 481698
rect 552604 446018 552786 446254
rect 553022 446018 553204 446254
rect 552604 445934 553204 446018
rect 552604 445698 552786 445934
rect 553022 445698 553204 445934
rect 552604 410254 553204 445698
rect 552604 410018 552786 410254
rect 553022 410018 553204 410254
rect 552604 409934 553204 410018
rect 552604 409698 552786 409934
rect 553022 409698 553204 409934
rect 552604 374254 553204 409698
rect 552604 374018 552786 374254
rect 553022 374018 553204 374254
rect 552604 373934 553204 374018
rect 552604 373698 552786 373934
rect 553022 373698 553204 373934
rect 552604 338254 553204 373698
rect 552604 338018 552786 338254
rect 553022 338018 553204 338254
rect 552604 337934 553204 338018
rect 552604 337698 552786 337934
rect 553022 337698 553204 337934
rect 552604 302254 553204 337698
rect 552604 302018 552786 302254
rect 553022 302018 553204 302254
rect 552604 301934 553204 302018
rect 552604 301698 552786 301934
rect 553022 301698 553204 301934
rect 552604 266254 553204 301698
rect 552604 266018 552786 266254
rect 553022 266018 553204 266254
rect 552604 265934 553204 266018
rect 552604 265698 552786 265934
rect 553022 265698 553204 265934
rect 552604 230254 553204 265698
rect 552604 230018 552786 230254
rect 553022 230018 553204 230254
rect 552604 229934 553204 230018
rect 552604 229698 552786 229934
rect 553022 229698 553204 229934
rect 552604 194254 553204 229698
rect 552604 194018 552786 194254
rect 553022 194018 553204 194254
rect 552604 193934 553204 194018
rect 552604 193698 552786 193934
rect 553022 193698 553204 193934
rect 552604 158254 553204 193698
rect 552604 158018 552786 158254
rect 553022 158018 553204 158254
rect 552604 157934 553204 158018
rect 552604 157698 552786 157934
rect 553022 157698 553204 157934
rect 552604 122254 553204 157698
rect 552604 122018 552786 122254
rect 553022 122018 553204 122254
rect 552604 121934 553204 122018
rect 552604 121698 552786 121934
rect 553022 121698 553204 121934
rect 552604 86254 553204 121698
rect 552604 86018 552786 86254
rect 553022 86018 553204 86254
rect 552604 85934 553204 86018
rect 552604 85698 552786 85934
rect 553022 85698 553204 85934
rect 552604 50254 553204 85698
rect 552604 50018 552786 50254
rect 553022 50018 553204 50254
rect 552604 49934 553204 50018
rect 552604 49698 552786 49934
rect 553022 49698 553204 49934
rect 552604 14254 553204 49698
rect 552604 14018 552786 14254
rect 553022 14018 553204 14254
rect 552604 13934 553204 14018
rect 552604 13698 552786 13934
rect 553022 13698 553204 13934
rect 534604 -7162 534786 -6926
rect 535022 -7162 535204 -6926
rect 534604 -7246 535204 -7162
rect 534604 -7482 534786 -7246
rect 535022 -7482 535204 -7246
rect 534604 -7504 535204 -7482
rect 552604 -5986 553204 13698
rect 559804 705778 560404 705800
rect 559804 705542 559986 705778
rect 560222 705542 560404 705778
rect 559804 705458 560404 705542
rect 559804 705222 559986 705458
rect 560222 705222 560404 705458
rect 559804 669454 560404 705222
rect 559804 669218 559986 669454
rect 560222 669218 560404 669454
rect 559804 669134 560404 669218
rect 559804 668898 559986 669134
rect 560222 668898 560404 669134
rect 559804 633454 560404 668898
rect 559804 633218 559986 633454
rect 560222 633218 560404 633454
rect 559804 633134 560404 633218
rect 559804 632898 559986 633134
rect 560222 632898 560404 633134
rect 559804 597454 560404 632898
rect 559804 597218 559986 597454
rect 560222 597218 560404 597454
rect 559804 597134 560404 597218
rect 559804 596898 559986 597134
rect 560222 596898 560404 597134
rect 559804 561454 560404 596898
rect 559804 561218 559986 561454
rect 560222 561218 560404 561454
rect 559804 561134 560404 561218
rect 559804 560898 559986 561134
rect 560222 560898 560404 561134
rect 559804 525454 560404 560898
rect 559804 525218 559986 525454
rect 560222 525218 560404 525454
rect 559804 525134 560404 525218
rect 559804 524898 559986 525134
rect 560222 524898 560404 525134
rect 559804 489454 560404 524898
rect 559804 489218 559986 489454
rect 560222 489218 560404 489454
rect 559804 489134 560404 489218
rect 559804 488898 559986 489134
rect 560222 488898 560404 489134
rect 559804 453454 560404 488898
rect 559804 453218 559986 453454
rect 560222 453218 560404 453454
rect 559804 453134 560404 453218
rect 559804 452898 559986 453134
rect 560222 452898 560404 453134
rect 559804 417454 560404 452898
rect 559804 417218 559986 417454
rect 560222 417218 560404 417454
rect 559804 417134 560404 417218
rect 559804 416898 559986 417134
rect 560222 416898 560404 417134
rect 559804 381454 560404 416898
rect 559804 381218 559986 381454
rect 560222 381218 560404 381454
rect 559804 381134 560404 381218
rect 559804 380898 559986 381134
rect 560222 380898 560404 381134
rect 559804 345454 560404 380898
rect 559804 345218 559986 345454
rect 560222 345218 560404 345454
rect 559804 345134 560404 345218
rect 559804 344898 559986 345134
rect 560222 344898 560404 345134
rect 559804 309454 560404 344898
rect 559804 309218 559986 309454
rect 560222 309218 560404 309454
rect 559804 309134 560404 309218
rect 559804 308898 559986 309134
rect 560222 308898 560404 309134
rect 559804 273454 560404 308898
rect 559804 273218 559986 273454
rect 560222 273218 560404 273454
rect 559804 273134 560404 273218
rect 559804 272898 559986 273134
rect 560222 272898 560404 273134
rect 559804 237454 560404 272898
rect 559804 237218 559986 237454
rect 560222 237218 560404 237454
rect 559804 237134 560404 237218
rect 559804 236898 559986 237134
rect 560222 236898 560404 237134
rect 559804 201454 560404 236898
rect 559804 201218 559986 201454
rect 560222 201218 560404 201454
rect 559804 201134 560404 201218
rect 559804 200898 559986 201134
rect 560222 200898 560404 201134
rect 559804 165454 560404 200898
rect 559804 165218 559986 165454
rect 560222 165218 560404 165454
rect 559804 165134 560404 165218
rect 559804 164898 559986 165134
rect 560222 164898 560404 165134
rect 559804 129454 560404 164898
rect 559804 129218 559986 129454
rect 560222 129218 560404 129454
rect 559804 129134 560404 129218
rect 559804 128898 559986 129134
rect 560222 128898 560404 129134
rect 559804 93454 560404 128898
rect 559804 93218 559986 93454
rect 560222 93218 560404 93454
rect 559804 93134 560404 93218
rect 559804 92898 559986 93134
rect 560222 92898 560404 93134
rect 559804 57454 560404 92898
rect 559804 57218 559986 57454
rect 560222 57218 560404 57454
rect 559804 57134 560404 57218
rect 559804 56898 559986 57134
rect 560222 56898 560404 57134
rect 559804 21454 560404 56898
rect 559804 21218 559986 21454
rect 560222 21218 560404 21454
rect 559804 21134 560404 21218
rect 559804 20898 559986 21134
rect 560222 20898 560404 21134
rect 559804 -1286 560404 20898
rect 559804 -1522 559986 -1286
rect 560222 -1522 560404 -1286
rect 559804 -1606 560404 -1522
rect 559804 -1842 559986 -1606
rect 560222 -1842 560404 -1606
rect 559804 -1864 560404 -1842
rect 563404 673054 564004 707102
rect 563404 672818 563586 673054
rect 563822 672818 564004 673054
rect 563404 672734 564004 672818
rect 563404 672498 563586 672734
rect 563822 672498 564004 672734
rect 563404 637054 564004 672498
rect 563404 636818 563586 637054
rect 563822 636818 564004 637054
rect 563404 636734 564004 636818
rect 563404 636498 563586 636734
rect 563822 636498 564004 636734
rect 563404 601054 564004 636498
rect 563404 600818 563586 601054
rect 563822 600818 564004 601054
rect 563404 600734 564004 600818
rect 563404 600498 563586 600734
rect 563822 600498 564004 600734
rect 563404 565054 564004 600498
rect 563404 564818 563586 565054
rect 563822 564818 564004 565054
rect 563404 564734 564004 564818
rect 563404 564498 563586 564734
rect 563822 564498 564004 564734
rect 563404 529054 564004 564498
rect 563404 528818 563586 529054
rect 563822 528818 564004 529054
rect 563404 528734 564004 528818
rect 563404 528498 563586 528734
rect 563822 528498 564004 528734
rect 563404 493054 564004 528498
rect 563404 492818 563586 493054
rect 563822 492818 564004 493054
rect 563404 492734 564004 492818
rect 563404 492498 563586 492734
rect 563822 492498 564004 492734
rect 563404 457054 564004 492498
rect 563404 456818 563586 457054
rect 563822 456818 564004 457054
rect 563404 456734 564004 456818
rect 563404 456498 563586 456734
rect 563822 456498 564004 456734
rect 563404 421054 564004 456498
rect 563404 420818 563586 421054
rect 563822 420818 564004 421054
rect 563404 420734 564004 420818
rect 563404 420498 563586 420734
rect 563822 420498 564004 420734
rect 563404 385054 564004 420498
rect 563404 384818 563586 385054
rect 563822 384818 564004 385054
rect 563404 384734 564004 384818
rect 563404 384498 563586 384734
rect 563822 384498 564004 384734
rect 563404 349054 564004 384498
rect 563404 348818 563586 349054
rect 563822 348818 564004 349054
rect 563404 348734 564004 348818
rect 563404 348498 563586 348734
rect 563822 348498 564004 348734
rect 563404 313054 564004 348498
rect 563404 312818 563586 313054
rect 563822 312818 564004 313054
rect 563404 312734 564004 312818
rect 563404 312498 563586 312734
rect 563822 312498 564004 312734
rect 563404 277054 564004 312498
rect 563404 276818 563586 277054
rect 563822 276818 564004 277054
rect 563404 276734 564004 276818
rect 563404 276498 563586 276734
rect 563822 276498 564004 276734
rect 563404 241054 564004 276498
rect 563404 240818 563586 241054
rect 563822 240818 564004 241054
rect 563404 240734 564004 240818
rect 563404 240498 563586 240734
rect 563822 240498 564004 240734
rect 563404 205054 564004 240498
rect 563404 204818 563586 205054
rect 563822 204818 564004 205054
rect 563404 204734 564004 204818
rect 563404 204498 563586 204734
rect 563822 204498 564004 204734
rect 563404 169054 564004 204498
rect 563404 168818 563586 169054
rect 563822 168818 564004 169054
rect 563404 168734 564004 168818
rect 563404 168498 563586 168734
rect 563822 168498 564004 168734
rect 563404 133054 564004 168498
rect 563404 132818 563586 133054
rect 563822 132818 564004 133054
rect 563404 132734 564004 132818
rect 563404 132498 563586 132734
rect 563822 132498 564004 132734
rect 563404 97054 564004 132498
rect 563404 96818 563586 97054
rect 563822 96818 564004 97054
rect 563404 96734 564004 96818
rect 563404 96498 563586 96734
rect 563822 96498 564004 96734
rect 563404 61054 564004 96498
rect 563404 60818 563586 61054
rect 563822 60818 564004 61054
rect 563404 60734 564004 60818
rect 563404 60498 563586 60734
rect 563822 60498 564004 60734
rect 563404 25054 564004 60498
rect 563404 24818 563586 25054
rect 563822 24818 564004 25054
rect 563404 24734 564004 24818
rect 563404 24498 563586 24734
rect 563822 24498 564004 24734
rect 563404 -3166 564004 24498
rect 563404 -3402 563586 -3166
rect 563822 -3402 564004 -3166
rect 563404 -3486 564004 -3402
rect 563404 -3722 563586 -3486
rect 563822 -3722 564004 -3486
rect 563404 -3744 564004 -3722
rect 567004 676654 567604 708982
rect 567004 676418 567186 676654
rect 567422 676418 567604 676654
rect 567004 676334 567604 676418
rect 567004 676098 567186 676334
rect 567422 676098 567604 676334
rect 567004 640654 567604 676098
rect 567004 640418 567186 640654
rect 567422 640418 567604 640654
rect 567004 640334 567604 640418
rect 567004 640098 567186 640334
rect 567422 640098 567604 640334
rect 567004 604654 567604 640098
rect 567004 604418 567186 604654
rect 567422 604418 567604 604654
rect 567004 604334 567604 604418
rect 567004 604098 567186 604334
rect 567422 604098 567604 604334
rect 567004 568654 567604 604098
rect 567004 568418 567186 568654
rect 567422 568418 567604 568654
rect 567004 568334 567604 568418
rect 567004 568098 567186 568334
rect 567422 568098 567604 568334
rect 567004 532654 567604 568098
rect 567004 532418 567186 532654
rect 567422 532418 567604 532654
rect 567004 532334 567604 532418
rect 567004 532098 567186 532334
rect 567422 532098 567604 532334
rect 567004 496654 567604 532098
rect 567004 496418 567186 496654
rect 567422 496418 567604 496654
rect 567004 496334 567604 496418
rect 567004 496098 567186 496334
rect 567422 496098 567604 496334
rect 567004 460654 567604 496098
rect 567004 460418 567186 460654
rect 567422 460418 567604 460654
rect 567004 460334 567604 460418
rect 567004 460098 567186 460334
rect 567422 460098 567604 460334
rect 567004 424654 567604 460098
rect 567004 424418 567186 424654
rect 567422 424418 567604 424654
rect 567004 424334 567604 424418
rect 567004 424098 567186 424334
rect 567422 424098 567604 424334
rect 567004 388654 567604 424098
rect 567004 388418 567186 388654
rect 567422 388418 567604 388654
rect 567004 388334 567604 388418
rect 567004 388098 567186 388334
rect 567422 388098 567604 388334
rect 567004 352654 567604 388098
rect 567004 352418 567186 352654
rect 567422 352418 567604 352654
rect 567004 352334 567604 352418
rect 567004 352098 567186 352334
rect 567422 352098 567604 352334
rect 567004 316654 567604 352098
rect 567004 316418 567186 316654
rect 567422 316418 567604 316654
rect 567004 316334 567604 316418
rect 567004 316098 567186 316334
rect 567422 316098 567604 316334
rect 567004 280654 567604 316098
rect 567004 280418 567186 280654
rect 567422 280418 567604 280654
rect 567004 280334 567604 280418
rect 567004 280098 567186 280334
rect 567422 280098 567604 280334
rect 567004 244654 567604 280098
rect 567004 244418 567186 244654
rect 567422 244418 567604 244654
rect 567004 244334 567604 244418
rect 567004 244098 567186 244334
rect 567422 244098 567604 244334
rect 567004 208654 567604 244098
rect 567004 208418 567186 208654
rect 567422 208418 567604 208654
rect 567004 208334 567604 208418
rect 567004 208098 567186 208334
rect 567422 208098 567604 208334
rect 567004 172654 567604 208098
rect 567004 172418 567186 172654
rect 567422 172418 567604 172654
rect 567004 172334 567604 172418
rect 567004 172098 567186 172334
rect 567422 172098 567604 172334
rect 567004 136654 567604 172098
rect 567004 136418 567186 136654
rect 567422 136418 567604 136654
rect 567004 136334 567604 136418
rect 567004 136098 567186 136334
rect 567422 136098 567604 136334
rect 567004 100654 567604 136098
rect 567004 100418 567186 100654
rect 567422 100418 567604 100654
rect 567004 100334 567604 100418
rect 567004 100098 567186 100334
rect 567422 100098 567604 100334
rect 567004 64654 567604 100098
rect 567004 64418 567186 64654
rect 567422 64418 567604 64654
rect 567004 64334 567604 64418
rect 567004 64098 567186 64334
rect 567422 64098 567604 64334
rect 567004 28654 567604 64098
rect 567004 28418 567186 28654
rect 567422 28418 567604 28654
rect 567004 28334 567604 28418
rect 567004 28098 567186 28334
rect 567422 28098 567604 28334
rect 567004 -5046 567604 28098
rect 567004 -5282 567186 -5046
rect 567422 -5282 567604 -5046
rect 567004 -5366 567604 -5282
rect 567004 -5602 567186 -5366
rect 567422 -5602 567604 -5366
rect 567004 -5624 567604 -5602
rect 570604 680254 571204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 581404 706718 582004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 581404 706482 581586 706718
rect 581822 706482 582004 706718
rect 581404 706398 582004 706482
rect 581404 706162 581586 706398
rect 581822 706162 582004 706398
rect 570604 680018 570786 680254
rect 571022 680018 571204 680254
rect 570604 679934 571204 680018
rect 570604 679698 570786 679934
rect 571022 679698 571204 679934
rect 570604 644254 571204 679698
rect 570604 644018 570786 644254
rect 571022 644018 571204 644254
rect 570604 643934 571204 644018
rect 570604 643698 570786 643934
rect 571022 643698 571204 643934
rect 570604 608254 571204 643698
rect 570604 608018 570786 608254
rect 571022 608018 571204 608254
rect 570604 607934 571204 608018
rect 570604 607698 570786 607934
rect 571022 607698 571204 607934
rect 570604 572254 571204 607698
rect 570604 572018 570786 572254
rect 571022 572018 571204 572254
rect 570604 571934 571204 572018
rect 570604 571698 570786 571934
rect 571022 571698 571204 571934
rect 570604 536254 571204 571698
rect 570604 536018 570786 536254
rect 571022 536018 571204 536254
rect 570604 535934 571204 536018
rect 570604 535698 570786 535934
rect 571022 535698 571204 535934
rect 570604 500254 571204 535698
rect 570604 500018 570786 500254
rect 571022 500018 571204 500254
rect 570604 499934 571204 500018
rect 570604 499698 570786 499934
rect 571022 499698 571204 499934
rect 570604 464254 571204 499698
rect 570604 464018 570786 464254
rect 571022 464018 571204 464254
rect 570604 463934 571204 464018
rect 570604 463698 570786 463934
rect 571022 463698 571204 463934
rect 570604 428254 571204 463698
rect 570604 428018 570786 428254
rect 571022 428018 571204 428254
rect 570604 427934 571204 428018
rect 570604 427698 570786 427934
rect 571022 427698 571204 427934
rect 570604 392254 571204 427698
rect 570604 392018 570786 392254
rect 571022 392018 571204 392254
rect 570604 391934 571204 392018
rect 570604 391698 570786 391934
rect 571022 391698 571204 391934
rect 570604 356254 571204 391698
rect 570604 356018 570786 356254
rect 571022 356018 571204 356254
rect 570604 355934 571204 356018
rect 570604 355698 570786 355934
rect 571022 355698 571204 355934
rect 570604 320254 571204 355698
rect 570604 320018 570786 320254
rect 571022 320018 571204 320254
rect 570604 319934 571204 320018
rect 570604 319698 570786 319934
rect 571022 319698 571204 319934
rect 570604 284254 571204 319698
rect 570604 284018 570786 284254
rect 571022 284018 571204 284254
rect 570604 283934 571204 284018
rect 570604 283698 570786 283934
rect 571022 283698 571204 283934
rect 570604 248254 571204 283698
rect 570604 248018 570786 248254
rect 571022 248018 571204 248254
rect 570604 247934 571204 248018
rect 570604 247698 570786 247934
rect 571022 247698 571204 247934
rect 570604 212254 571204 247698
rect 570604 212018 570786 212254
rect 571022 212018 571204 212254
rect 570604 211934 571204 212018
rect 570604 211698 570786 211934
rect 571022 211698 571204 211934
rect 570604 176254 571204 211698
rect 570604 176018 570786 176254
rect 571022 176018 571204 176254
rect 570604 175934 571204 176018
rect 570604 175698 570786 175934
rect 571022 175698 571204 175934
rect 570604 140254 571204 175698
rect 570604 140018 570786 140254
rect 571022 140018 571204 140254
rect 570604 139934 571204 140018
rect 570604 139698 570786 139934
rect 571022 139698 571204 139934
rect 570604 104254 571204 139698
rect 570604 104018 570786 104254
rect 571022 104018 571204 104254
rect 570604 103934 571204 104018
rect 570604 103698 570786 103934
rect 571022 103698 571204 103934
rect 570604 68254 571204 103698
rect 570604 68018 570786 68254
rect 571022 68018 571204 68254
rect 570604 67934 571204 68018
rect 570604 67698 570786 67934
rect 571022 67698 571204 67934
rect 570604 32254 571204 67698
rect 570604 32018 570786 32254
rect 571022 32018 571204 32254
rect 570604 31934 571204 32018
rect 570604 31698 570786 31934
rect 571022 31698 571204 31934
rect 552604 -6222 552786 -5986
rect 553022 -6222 553204 -5986
rect 552604 -6306 553204 -6222
rect 552604 -6542 552786 -6306
rect 553022 -6542 553204 -6306
rect 552604 -7504 553204 -6542
rect 570604 -6926 571204 31698
rect 577804 704838 578404 705800
rect 577804 704602 577986 704838
rect 578222 704602 578404 704838
rect 577804 704518 578404 704602
rect 577804 704282 577986 704518
rect 578222 704282 578404 704518
rect 577804 687454 578404 704282
rect 577804 687218 577986 687454
rect 578222 687218 578404 687454
rect 577804 687134 578404 687218
rect 577804 686898 577986 687134
rect 578222 686898 578404 687134
rect 577804 651454 578404 686898
rect 577804 651218 577986 651454
rect 578222 651218 578404 651454
rect 577804 651134 578404 651218
rect 577804 650898 577986 651134
rect 578222 650898 578404 651134
rect 577804 615454 578404 650898
rect 577804 615218 577986 615454
rect 578222 615218 578404 615454
rect 577804 615134 578404 615218
rect 577804 614898 577986 615134
rect 578222 614898 578404 615134
rect 577804 579454 578404 614898
rect 577804 579218 577986 579454
rect 578222 579218 578404 579454
rect 577804 579134 578404 579218
rect 577804 578898 577986 579134
rect 578222 578898 578404 579134
rect 577804 543454 578404 578898
rect 577804 543218 577986 543454
rect 578222 543218 578404 543454
rect 577804 543134 578404 543218
rect 577804 542898 577986 543134
rect 578222 542898 578404 543134
rect 577804 507454 578404 542898
rect 577804 507218 577986 507454
rect 578222 507218 578404 507454
rect 577804 507134 578404 507218
rect 577804 506898 577986 507134
rect 578222 506898 578404 507134
rect 577804 471454 578404 506898
rect 577804 471218 577986 471454
rect 578222 471218 578404 471454
rect 577804 471134 578404 471218
rect 577804 470898 577986 471134
rect 578222 470898 578404 471134
rect 577804 435454 578404 470898
rect 577804 435218 577986 435454
rect 578222 435218 578404 435454
rect 577804 435134 578404 435218
rect 577804 434898 577986 435134
rect 578222 434898 578404 435134
rect 577804 399454 578404 434898
rect 577804 399218 577986 399454
rect 578222 399218 578404 399454
rect 577804 399134 578404 399218
rect 577804 398898 577986 399134
rect 578222 398898 578404 399134
rect 577804 363454 578404 398898
rect 577804 363218 577986 363454
rect 578222 363218 578404 363454
rect 577804 363134 578404 363218
rect 577804 362898 577986 363134
rect 578222 362898 578404 363134
rect 577804 327454 578404 362898
rect 577804 327218 577986 327454
rect 578222 327218 578404 327454
rect 577804 327134 578404 327218
rect 577804 326898 577986 327134
rect 578222 326898 578404 327134
rect 577804 291454 578404 326898
rect 577804 291218 577986 291454
rect 578222 291218 578404 291454
rect 577804 291134 578404 291218
rect 577804 290898 577986 291134
rect 578222 290898 578404 291134
rect 577804 255454 578404 290898
rect 577804 255218 577986 255454
rect 578222 255218 578404 255454
rect 577804 255134 578404 255218
rect 577804 254898 577986 255134
rect 578222 254898 578404 255134
rect 577804 219454 578404 254898
rect 577804 219218 577986 219454
rect 578222 219218 578404 219454
rect 577804 219134 578404 219218
rect 577804 218898 577986 219134
rect 578222 218898 578404 219134
rect 577804 183454 578404 218898
rect 577804 183218 577986 183454
rect 578222 183218 578404 183454
rect 577804 183134 578404 183218
rect 577804 182898 577986 183134
rect 578222 182898 578404 183134
rect 577804 147454 578404 182898
rect 577804 147218 577986 147454
rect 578222 147218 578404 147454
rect 577804 147134 578404 147218
rect 577804 146898 577986 147134
rect 578222 146898 578404 147134
rect 577804 111454 578404 146898
rect 577804 111218 577986 111454
rect 578222 111218 578404 111454
rect 577804 111134 578404 111218
rect 577804 110898 577986 111134
rect 578222 110898 578404 111134
rect 577804 75454 578404 110898
rect 577804 75218 577986 75454
rect 578222 75218 578404 75454
rect 577804 75134 578404 75218
rect 577804 74898 577986 75134
rect 578222 74898 578404 75134
rect 577804 39454 578404 74898
rect 577804 39218 577986 39454
rect 578222 39218 578404 39454
rect 577804 39134 578404 39218
rect 577804 38898 577986 39134
rect 578222 38898 578404 39134
rect 577804 3454 578404 38898
rect 577804 3218 577986 3454
rect 578222 3218 578404 3454
rect 577804 3134 578404 3218
rect 577804 2898 577986 3134
rect 578222 2898 578404 3134
rect 577804 -346 578404 2898
rect 577804 -582 577986 -346
rect 578222 -582 578404 -346
rect 577804 -666 578404 -582
rect 577804 -902 577986 -666
rect 578222 -902 578404 -666
rect 577804 -1864 578404 -902
rect 581404 691054 582004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 581404 690818 581586 691054
rect 581822 690818 582004 691054
rect 581404 690734 582004 690818
rect 581404 690498 581586 690734
rect 581822 690498 582004 690734
rect 581404 655054 582004 690498
rect 581404 654818 581586 655054
rect 581822 654818 582004 655054
rect 581404 654734 582004 654818
rect 581404 654498 581586 654734
rect 581822 654498 582004 654734
rect 581404 619054 582004 654498
rect 581404 618818 581586 619054
rect 581822 618818 582004 619054
rect 581404 618734 582004 618818
rect 581404 618498 581586 618734
rect 581822 618498 582004 618734
rect 581404 583054 582004 618498
rect 581404 582818 581586 583054
rect 581822 582818 582004 583054
rect 581404 582734 582004 582818
rect 581404 582498 581586 582734
rect 581822 582498 582004 582734
rect 581404 547054 582004 582498
rect 581404 546818 581586 547054
rect 581822 546818 582004 547054
rect 581404 546734 582004 546818
rect 581404 546498 581586 546734
rect 581822 546498 582004 546734
rect 581404 511054 582004 546498
rect 581404 510818 581586 511054
rect 581822 510818 582004 511054
rect 581404 510734 582004 510818
rect 581404 510498 581586 510734
rect 581822 510498 582004 510734
rect 581404 475054 582004 510498
rect 581404 474818 581586 475054
rect 581822 474818 582004 475054
rect 581404 474734 582004 474818
rect 581404 474498 581586 474734
rect 581822 474498 582004 474734
rect 581404 439054 582004 474498
rect 581404 438818 581586 439054
rect 581822 438818 582004 439054
rect 581404 438734 582004 438818
rect 581404 438498 581586 438734
rect 581822 438498 582004 438734
rect 581404 403054 582004 438498
rect 581404 402818 581586 403054
rect 581822 402818 582004 403054
rect 581404 402734 582004 402818
rect 581404 402498 581586 402734
rect 581822 402498 582004 402734
rect 581404 367054 582004 402498
rect 581404 366818 581586 367054
rect 581822 366818 582004 367054
rect 581404 366734 582004 366818
rect 581404 366498 581586 366734
rect 581822 366498 582004 366734
rect 581404 331054 582004 366498
rect 581404 330818 581586 331054
rect 581822 330818 582004 331054
rect 581404 330734 582004 330818
rect 581404 330498 581586 330734
rect 581822 330498 582004 330734
rect 581404 295054 582004 330498
rect 581404 294818 581586 295054
rect 581822 294818 582004 295054
rect 581404 294734 582004 294818
rect 581404 294498 581586 294734
rect 581822 294498 582004 294734
rect 581404 259054 582004 294498
rect 581404 258818 581586 259054
rect 581822 258818 582004 259054
rect 581404 258734 582004 258818
rect 581404 258498 581586 258734
rect 581822 258498 582004 258734
rect 581404 223054 582004 258498
rect 581404 222818 581586 223054
rect 581822 222818 582004 223054
rect 581404 222734 582004 222818
rect 581404 222498 581586 222734
rect 581822 222498 582004 222734
rect 581404 187054 582004 222498
rect 581404 186818 581586 187054
rect 581822 186818 582004 187054
rect 581404 186734 582004 186818
rect 581404 186498 581586 186734
rect 581822 186498 582004 186734
rect 581404 151054 582004 186498
rect 581404 150818 581586 151054
rect 581822 150818 582004 151054
rect 581404 150734 582004 150818
rect 581404 150498 581586 150734
rect 581822 150498 582004 150734
rect 581404 115054 582004 150498
rect 581404 114818 581586 115054
rect 581822 114818 582004 115054
rect 581404 114734 582004 114818
rect 581404 114498 581586 114734
rect 581822 114498 582004 114734
rect 581404 79054 582004 114498
rect 581404 78818 581586 79054
rect 581822 78818 582004 79054
rect 581404 78734 582004 78818
rect 581404 78498 581586 78734
rect 581822 78498 582004 78734
rect 581404 43054 582004 78498
rect 581404 42818 581586 43054
rect 581822 42818 582004 43054
rect 581404 42734 582004 42818
rect 581404 42498 581586 42734
rect 581822 42498 582004 42734
rect 581404 7054 582004 42498
rect 581404 6818 581586 7054
rect 581822 6818 582004 7054
rect 581404 6734 582004 6818
rect 581404 6498 581586 6734
rect 581822 6498 582004 6734
rect 581404 -2226 582004 6498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 687454 585920 704282
rect 585320 687218 585502 687454
rect 585738 687218 585920 687454
rect 585320 687134 585920 687218
rect 585320 686898 585502 687134
rect 585738 686898 585920 687134
rect 585320 651454 585920 686898
rect 585320 651218 585502 651454
rect 585738 651218 585920 651454
rect 585320 651134 585920 651218
rect 585320 650898 585502 651134
rect 585738 650898 585920 651134
rect 585320 615454 585920 650898
rect 585320 615218 585502 615454
rect 585738 615218 585920 615454
rect 585320 615134 585920 615218
rect 585320 614898 585502 615134
rect 585738 614898 585920 615134
rect 585320 579454 585920 614898
rect 585320 579218 585502 579454
rect 585738 579218 585920 579454
rect 585320 579134 585920 579218
rect 585320 578898 585502 579134
rect 585738 578898 585920 579134
rect 585320 543454 585920 578898
rect 585320 543218 585502 543454
rect 585738 543218 585920 543454
rect 585320 543134 585920 543218
rect 585320 542898 585502 543134
rect 585738 542898 585920 543134
rect 585320 507454 585920 542898
rect 585320 507218 585502 507454
rect 585738 507218 585920 507454
rect 585320 507134 585920 507218
rect 585320 506898 585502 507134
rect 585738 506898 585920 507134
rect 585320 471454 585920 506898
rect 585320 471218 585502 471454
rect 585738 471218 585920 471454
rect 585320 471134 585920 471218
rect 585320 470898 585502 471134
rect 585738 470898 585920 471134
rect 585320 435454 585920 470898
rect 585320 435218 585502 435454
rect 585738 435218 585920 435454
rect 585320 435134 585920 435218
rect 585320 434898 585502 435134
rect 585738 434898 585920 435134
rect 585320 399454 585920 434898
rect 585320 399218 585502 399454
rect 585738 399218 585920 399454
rect 585320 399134 585920 399218
rect 585320 398898 585502 399134
rect 585738 398898 585920 399134
rect 585320 363454 585920 398898
rect 585320 363218 585502 363454
rect 585738 363218 585920 363454
rect 585320 363134 585920 363218
rect 585320 362898 585502 363134
rect 585738 362898 585920 363134
rect 585320 327454 585920 362898
rect 585320 327218 585502 327454
rect 585738 327218 585920 327454
rect 585320 327134 585920 327218
rect 585320 326898 585502 327134
rect 585738 326898 585920 327134
rect 585320 291454 585920 326898
rect 585320 291218 585502 291454
rect 585738 291218 585920 291454
rect 585320 291134 585920 291218
rect 585320 290898 585502 291134
rect 585738 290898 585920 291134
rect 585320 255454 585920 290898
rect 585320 255218 585502 255454
rect 585738 255218 585920 255454
rect 585320 255134 585920 255218
rect 585320 254898 585502 255134
rect 585738 254898 585920 255134
rect 585320 219454 585920 254898
rect 585320 219218 585502 219454
rect 585738 219218 585920 219454
rect 585320 219134 585920 219218
rect 585320 218898 585502 219134
rect 585738 218898 585920 219134
rect 585320 183454 585920 218898
rect 585320 183218 585502 183454
rect 585738 183218 585920 183454
rect 585320 183134 585920 183218
rect 585320 182898 585502 183134
rect 585738 182898 585920 183134
rect 585320 147454 585920 182898
rect 585320 147218 585502 147454
rect 585738 147218 585920 147454
rect 585320 147134 585920 147218
rect 585320 146898 585502 147134
rect 585738 146898 585920 147134
rect 585320 111454 585920 146898
rect 585320 111218 585502 111454
rect 585738 111218 585920 111454
rect 585320 111134 585920 111218
rect 585320 110898 585502 111134
rect 585738 110898 585920 111134
rect 585320 75454 585920 110898
rect 585320 75218 585502 75454
rect 585738 75218 585920 75454
rect 585320 75134 585920 75218
rect 585320 74898 585502 75134
rect 585738 74898 585920 75134
rect 585320 39454 585920 74898
rect 585320 39218 585502 39454
rect 585738 39218 585920 39454
rect 585320 39134 585920 39218
rect 585320 38898 585502 39134
rect 585738 38898 585920 39134
rect 585320 3454 585920 38898
rect 585320 3218 585502 3454
rect 585738 3218 585920 3454
rect 585320 3134 585920 3218
rect 585320 2898 585502 3134
rect 585738 2898 585920 3134
rect 585320 -346 585920 2898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 669454 586860 705222
rect 586260 669218 586442 669454
rect 586678 669218 586860 669454
rect 586260 669134 586860 669218
rect 586260 668898 586442 669134
rect 586678 668898 586860 669134
rect 586260 633454 586860 668898
rect 586260 633218 586442 633454
rect 586678 633218 586860 633454
rect 586260 633134 586860 633218
rect 586260 632898 586442 633134
rect 586678 632898 586860 633134
rect 586260 597454 586860 632898
rect 586260 597218 586442 597454
rect 586678 597218 586860 597454
rect 586260 597134 586860 597218
rect 586260 596898 586442 597134
rect 586678 596898 586860 597134
rect 586260 561454 586860 596898
rect 586260 561218 586442 561454
rect 586678 561218 586860 561454
rect 586260 561134 586860 561218
rect 586260 560898 586442 561134
rect 586678 560898 586860 561134
rect 586260 525454 586860 560898
rect 586260 525218 586442 525454
rect 586678 525218 586860 525454
rect 586260 525134 586860 525218
rect 586260 524898 586442 525134
rect 586678 524898 586860 525134
rect 586260 489454 586860 524898
rect 586260 489218 586442 489454
rect 586678 489218 586860 489454
rect 586260 489134 586860 489218
rect 586260 488898 586442 489134
rect 586678 488898 586860 489134
rect 586260 453454 586860 488898
rect 586260 453218 586442 453454
rect 586678 453218 586860 453454
rect 586260 453134 586860 453218
rect 586260 452898 586442 453134
rect 586678 452898 586860 453134
rect 586260 417454 586860 452898
rect 586260 417218 586442 417454
rect 586678 417218 586860 417454
rect 586260 417134 586860 417218
rect 586260 416898 586442 417134
rect 586678 416898 586860 417134
rect 586260 381454 586860 416898
rect 586260 381218 586442 381454
rect 586678 381218 586860 381454
rect 586260 381134 586860 381218
rect 586260 380898 586442 381134
rect 586678 380898 586860 381134
rect 586260 345454 586860 380898
rect 586260 345218 586442 345454
rect 586678 345218 586860 345454
rect 586260 345134 586860 345218
rect 586260 344898 586442 345134
rect 586678 344898 586860 345134
rect 586260 309454 586860 344898
rect 586260 309218 586442 309454
rect 586678 309218 586860 309454
rect 586260 309134 586860 309218
rect 586260 308898 586442 309134
rect 586678 308898 586860 309134
rect 586260 273454 586860 308898
rect 586260 273218 586442 273454
rect 586678 273218 586860 273454
rect 586260 273134 586860 273218
rect 586260 272898 586442 273134
rect 586678 272898 586860 273134
rect 586260 237454 586860 272898
rect 586260 237218 586442 237454
rect 586678 237218 586860 237454
rect 586260 237134 586860 237218
rect 586260 236898 586442 237134
rect 586678 236898 586860 237134
rect 586260 201454 586860 236898
rect 586260 201218 586442 201454
rect 586678 201218 586860 201454
rect 586260 201134 586860 201218
rect 586260 200898 586442 201134
rect 586678 200898 586860 201134
rect 586260 165454 586860 200898
rect 586260 165218 586442 165454
rect 586678 165218 586860 165454
rect 586260 165134 586860 165218
rect 586260 164898 586442 165134
rect 586678 164898 586860 165134
rect 586260 129454 586860 164898
rect 586260 129218 586442 129454
rect 586678 129218 586860 129454
rect 586260 129134 586860 129218
rect 586260 128898 586442 129134
rect 586678 128898 586860 129134
rect 586260 93454 586860 128898
rect 586260 93218 586442 93454
rect 586678 93218 586860 93454
rect 586260 93134 586860 93218
rect 586260 92898 586442 93134
rect 586678 92898 586860 93134
rect 586260 57454 586860 92898
rect 586260 57218 586442 57454
rect 586678 57218 586860 57454
rect 586260 57134 586860 57218
rect 586260 56898 586442 57134
rect 586678 56898 586860 57134
rect 586260 21454 586860 56898
rect 586260 21218 586442 21454
rect 586678 21218 586860 21454
rect 586260 21134 586860 21218
rect 586260 20898 586442 21134
rect 586678 20898 586860 21134
rect 586260 -1286 586860 20898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 691054 587800 706162
rect 587200 690818 587382 691054
rect 587618 690818 587800 691054
rect 587200 690734 587800 690818
rect 587200 690498 587382 690734
rect 587618 690498 587800 690734
rect 587200 655054 587800 690498
rect 587200 654818 587382 655054
rect 587618 654818 587800 655054
rect 587200 654734 587800 654818
rect 587200 654498 587382 654734
rect 587618 654498 587800 654734
rect 587200 619054 587800 654498
rect 587200 618818 587382 619054
rect 587618 618818 587800 619054
rect 587200 618734 587800 618818
rect 587200 618498 587382 618734
rect 587618 618498 587800 618734
rect 587200 583054 587800 618498
rect 587200 582818 587382 583054
rect 587618 582818 587800 583054
rect 587200 582734 587800 582818
rect 587200 582498 587382 582734
rect 587618 582498 587800 582734
rect 587200 547054 587800 582498
rect 587200 546818 587382 547054
rect 587618 546818 587800 547054
rect 587200 546734 587800 546818
rect 587200 546498 587382 546734
rect 587618 546498 587800 546734
rect 587200 511054 587800 546498
rect 587200 510818 587382 511054
rect 587618 510818 587800 511054
rect 587200 510734 587800 510818
rect 587200 510498 587382 510734
rect 587618 510498 587800 510734
rect 587200 475054 587800 510498
rect 587200 474818 587382 475054
rect 587618 474818 587800 475054
rect 587200 474734 587800 474818
rect 587200 474498 587382 474734
rect 587618 474498 587800 474734
rect 587200 439054 587800 474498
rect 587200 438818 587382 439054
rect 587618 438818 587800 439054
rect 587200 438734 587800 438818
rect 587200 438498 587382 438734
rect 587618 438498 587800 438734
rect 587200 403054 587800 438498
rect 587200 402818 587382 403054
rect 587618 402818 587800 403054
rect 587200 402734 587800 402818
rect 587200 402498 587382 402734
rect 587618 402498 587800 402734
rect 587200 367054 587800 402498
rect 587200 366818 587382 367054
rect 587618 366818 587800 367054
rect 587200 366734 587800 366818
rect 587200 366498 587382 366734
rect 587618 366498 587800 366734
rect 587200 331054 587800 366498
rect 587200 330818 587382 331054
rect 587618 330818 587800 331054
rect 587200 330734 587800 330818
rect 587200 330498 587382 330734
rect 587618 330498 587800 330734
rect 587200 295054 587800 330498
rect 587200 294818 587382 295054
rect 587618 294818 587800 295054
rect 587200 294734 587800 294818
rect 587200 294498 587382 294734
rect 587618 294498 587800 294734
rect 587200 259054 587800 294498
rect 587200 258818 587382 259054
rect 587618 258818 587800 259054
rect 587200 258734 587800 258818
rect 587200 258498 587382 258734
rect 587618 258498 587800 258734
rect 587200 223054 587800 258498
rect 587200 222818 587382 223054
rect 587618 222818 587800 223054
rect 587200 222734 587800 222818
rect 587200 222498 587382 222734
rect 587618 222498 587800 222734
rect 587200 187054 587800 222498
rect 587200 186818 587382 187054
rect 587618 186818 587800 187054
rect 587200 186734 587800 186818
rect 587200 186498 587382 186734
rect 587618 186498 587800 186734
rect 587200 151054 587800 186498
rect 587200 150818 587382 151054
rect 587618 150818 587800 151054
rect 587200 150734 587800 150818
rect 587200 150498 587382 150734
rect 587618 150498 587800 150734
rect 587200 115054 587800 150498
rect 587200 114818 587382 115054
rect 587618 114818 587800 115054
rect 587200 114734 587800 114818
rect 587200 114498 587382 114734
rect 587618 114498 587800 114734
rect 587200 79054 587800 114498
rect 587200 78818 587382 79054
rect 587618 78818 587800 79054
rect 587200 78734 587800 78818
rect 587200 78498 587382 78734
rect 587618 78498 587800 78734
rect 587200 43054 587800 78498
rect 587200 42818 587382 43054
rect 587618 42818 587800 43054
rect 587200 42734 587800 42818
rect 587200 42498 587382 42734
rect 587618 42498 587800 42734
rect 587200 7054 587800 42498
rect 587200 6818 587382 7054
rect 587618 6818 587800 7054
rect 587200 6734 587800 6818
rect 587200 6498 587382 6734
rect 587618 6498 587800 6734
rect 581404 -2462 581586 -2226
rect 581822 -2462 582004 -2226
rect 581404 -2546 582004 -2462
rect 581404 -2782 581586 -2546
rect 581822 -2782 582004 -2546
rect 581404 -3744 582004 -2782
rect 587200 -2226 587800 6498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 673054 588740 707102
rect 588140 672818 588322 673054
rect 588558 672818 588740 673054
rect 588140 672734 588740 672818
rect 588140 672498 588322 672734
rect 588558 672498 588740 672734
rect 588140 637054 588740 672498
rect 588140 636818 588322 637054
rect 588558 636818 588740 637054
rect 588140 636734 588740 636818
rect 588140 636498 588322 636734
rect 588558 636498 588740 636734
rect 588140 601054 588740 636498
rect 588140 600818 588322 601054
rect 588558 600818 588740 601054
rect 588140 600734 588740 600818
rect 588140 600498 588322 600734
rect 588558 600498 588740 600734
rect 588140 565054 588740 600498
rect 588140 564818 588322 565054
rect 588558 564818 588740 565054
rect 588140 564734 588740 564818
rect 588140 564498 588322 564734
rect 588558 564498 588740 564734
rect 588140 529054 588740 564498
rect 588140 528818 588322 529054
rect 588558 528818 588740 529054
rect 588140 528734 588740 528818
rect 588140 528498 588322 528734
rect 588558 528498 588740 528734
rect 588140 493054 588740 528498
rect 588140 492818 588322 493054
rect 588558 492818 588740 493054
rect 588140 492734 588740 492818
rect 588140 492498 588322 492734
rect 588558 492498 588740 492734
rect 588140 457054 588740 492498
rect 588140 456818 588322 457054
rect 588558 456818 588740 457054
rect 588140 456734 588740 456818
rect 588140 456498 588322 456734
rect 588558 456498 588740 456734
rect 588140 421054 588740 456498
rect 588140 420818 588322 421054
rect 588558 420818 588740 421054
rect 588140 420734 588740 420818
rect 588140 420498 588322 420734
rect 588558 420498 588740 420734
rect 588140 385054 588740 420498
rect 588140 384818 588322 385054
rect 588558 384818 588740 385054
rect 588140 384734 588740 384818
rect 588140 384498 588322 384734
rect 588558 384498 588740 384734
rect 588140 349054 588740 384498
rect 588140 348818 588322 349054
rect 588558 348818 588740 349054
rect 588140 348734 588740 348818
rect 588140 348498 588322 348734
rect 588558 348498 588740 348734
rect 588140 313054 588740 348498
rect 588140 312818 588322 313054
rect 588558 312818 588740 313054
rect 588140 312734 588740 312818
rect 588140 312498 588322 312734
rect 588558 312498 588740 312734
rect 588140 277054 588740 312498
rect 588140 276818 588322 277054
rect 588558 276818 588740 277054
rect 588140 276734 588740 276818
rect 588140 276498 588322 276734
rect 588558 276498 588740 276734
rect 588140 241054 588740 276498
rect 588140 240818 588322 241054
rect 588558 240818 588740 241054
rect 588140 240734 588740 240818
rect 588140 240498 588322 240734
rect 588558 240498 588740 240734
rect 588140 205054 588740 240498
rect 588140 204818 588322 205054
rect 588558 204818 588740 205054
rect 588140 204734 588740 204818
rect 588140 204498 588322 204734
rect 588558 204498 588740 204734
rect 588140 169054 588740 204498
rect 588140 168818 588322 169054
rect 588558 168818 588740 169054
rect 588140 168734 588740 168818
rect 588140 168498 588322 168734
rect 588558 168498 588740 168734
rect 588140 133054 588740 168498
rect 588140 132818 588322 133054
rect 588558 132818 588740 133054
rect 588140 132734 588740 132818
rect 588140 132498 588322 132734
rect 588558 132498 588740 132734
rect 588140 97054 588740 132498
rect 588140 96818 588322 97054
rect 588558 96818 588740 97054
rect 588140 96734 588740 96818
rect 588140 96498 588322 96734
rect 588558 96498 588740 96734
rect 588140 61054 588740 96498
rect 588140 60818 588322 61054
rect 588558 60818 588740 61054
rect 588140 60734 588740 60818
rect 588140 60498 588322 60734
rect 588558 60498 588740 60734
rect 588140 25054 588740 60498
rect 588140 24818 588322 25054
rect 588558 24818 588740 25054
rect 588140 24734 588740 24818
rect 588140 24498 588322 24734
rect 588558 24498 588740 24734
rect 588140 -3166 588740 24498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 694654 589680 708042
rect 589080 694418 589262 694654
rect 589498 694418 589680 694654
rect 589080 694334 589680 694418
rect 589080 694098 589262 694334
rect 589498 694098 589680 694334
rect 589080 658654 589680 694098
rect 589080 658418 589262 658654
rect 589498 658418 589680 658654
rect 589080 658334 589680 658418
rect 589080 658098 589262 658334
rect 589498 658098 589680 658334
rect 589080 622654 589680 658098
rect 589080 622418 589262 622654
rect 589498 622418 589680 622654
rect 589080 622334 589680 622418
rect 589080 622098 589262 622334
rect 589498 622098 589680 622334
rect 589080 586654 589680 622098
rect 589080 586418 589262 586654
rect 589498 586418 589680 586654
rect 589080 586334 589680 586418
rect 589080 586098 589262 586334
rect 589498 586098 589680 586334
rect 589080 550654 589680 586098
rect 589080 550418 589262 550654
rect 589498 550418 589680 550654
rect 589080 550334 589680 550418
rect 589080 550098 589262 550334
rect 589498 550098 589680 550334
rect 589080 514654 589680 550098
rect 589080 514418 589262 514654
rect 589498 514418 589680 514654
rect 589080 514334 589680 514418
rect 589080 514098 589262 514334
rect 589498 514098 589680 514334
rect 589080 478654 589680 514098
rect 589080 478418 589262 478654
rect 589498 478418 589680 478654
rect 589080 478334 589680 478418
rect 589080 478098 589262 478334
rect 589498 478098 589680 478334
rect 589080 442654 589680 478098
rect 589080 442418 589262 442654
rect 589498 442418 589680 442654
rect 589080 442334 589680 442418
rect 589080 442098 589262 442334
rect 589498 442098 589680 442334
rect 589080 406654 589680 442098
rect 589080 406418 589262 406654
rect 589498 406418 589680 406654
rect 589080 406334 589680 406418
rect 589080 406098 589262 406334
rect 589498 406098 589680 406334
rect 589080 370654 589680 406098
rect 589080 370418 589262 370654
rect 589498 370418 589680 370654
rect 589080 370334 589680 370418
rect 589080 370098 589262 370334
rect 589498 370098 589680 370334
rect 589080 334654 589680 370098
rect 589080 334418 589262 334654
rect 589498 334418 589680 334654
rect 589080 334334 589680 334418
rect 589080 334098 589262 334334
rect 589498 334098 589680 334334
rect 589080 298654 589680 334098
rect 589080 298418 589262 298654
rect 589498 298418 589680 298654
rect 589080 298334 589680 298418
rect 589080 298098 589262 298334
rect 589498 298098 589680 298334
rect 589080 262654 589680 298098
rect 589080 262418 589262 262654
rect 589498 262418 589680 262654
rect 589080 262334 589680 262418
rect 589080 262098 589262 262334
rect 589498 262098 589680 262334
rect 589080 226654 589680 262098
rect 589080 226418 589262 226654
rect 589498 226418 589680 226654
rect 589080 226334 589680 226418
rect 589080 226098 589262 226334
rect 589498 226098 589680 226334
rect 589080 190654 589680 226098
rect 589080 190418 589262 190654
rect 589498 190418 589680 190654
rect 589080 190334 589680 190418
rect 589080 190098 589262 190334
rect 589498 190098 589680 190334
rect 589080 154654 589680 190098
rect 589080 154418 589262 154654
rect 589498 154418 589680 154654
rect 589080 154334 589680 154418
rect 589080 154098 589262 154334
rect 589498 154098 589680 154334
rect 589080 118654 589680 154098
rect 589080 118418 589262 118654
rect 589498 118418 589680 118654
rect 589080 118334 589680 118418
rect 589080 118098 589262 118334
rect 589498 118098 589680 118334
rect 589080 82654 589680 118098
rect 589080 82418 589262 82654
rect 589498 82418 589680 82654
rect 589080 82334 589680 82418
rect 589080 82098 589262 82334
rect 589498 82098 589680 82334
rect 589080 46654 589680 82098
rect 589080 46418 589262 46654
rect 589498 46418 589680 46654
rect 589080 46334 589680 46418
rect 589080 46098 589262 46334
rect 589498 46098 589680 46334
rect 589080 10654 589680 46098
rect 589080 10418 589262 10654
rect 589498 10418 589680 10654
rect 589080 10334 589680 10418
rect 589080 10098 589262 10334
rect 589498 10098 589680 10334
rect 589080 -4106 589680 10098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 676654 590620 708982
rect 590020 676418 590202 676654
rect 590438 676418 590620 676654
rect 590020 676334 590620 676418
rect 590020 676098 590202 676334
rect 590438 676098 590620 676334
rect 590020 640654 590620 676098
rect 590020 640418 590202 640654
rect 590438 640418 590620 640654
rect 590020 640334 590620 640418
rect 590020 640098 590202 640334
rect 590438 640098 590620 640334
rect 590020 604654 590620 640098
rect 590020 604418 590202 604654
rect 590438 604418 590620 604654
rect 590020 604334 590620 604418
rect 590020 604098 590202 604334
rect 590438 604098 590620 604334
rect 590020 568654 590620 604098
rect 590020 568418 590202 568654
rect 590438 568418 590620 568654
rect 590020 568334 590620 568418
rect 590020 568098 590202 568334
rect 590438 568098 590620 568334
rect 590020 532654 590620 568098
rect 590020 532418 590202 532654
rect 590438 532418 590620 532654
rect 590020 532334 590620 532418
rect 590020 532098 590202 532334
rect 590438 532098 590620 532334
rect 590020 496654 590620 532098
rect 590020 496418 590202 496654
rect 590438 496418 590620 496654
rect 590020 496334 590620 496418
rect 590020 496098 590202 496334
rect 590438 496098 590620 496334
rect 590020 460654 590620 496098
rect 590020 460418 590202 460654
rect 590438 460418 590620 460654
rect 590020 460334 590620 460418
rect 590020 460098 590202 460334
rect 590438 460098 590620 460334
rect 590020 424654 590620 460098
rect 590020 424418 590202 424654
rect 590438 424418 590620 424654
rect 590020 424334 590620 424418
rect 590020 424098 590202 424334
rect 590438 424098 590620 424334
rect 590020 388654 590620 424098
rect 590020 388418 590202 388654
rect 590438 388418 590620 388654
rect 590020 388334 590620 388418
rect 590020 388098 590202 388334
rect 590438 388098 590620 388334
rect 590020 352654 590620 388098
rect 590020 352418 590202 352654
rect 590438 352418 590620 352654
rect 590020 352334 590620 352418
rect 590020 352098 590202 352334
rect 590438 352098 590620 352334
rect 590020 316654 590620 352098
rect 590020 316418 590202 316654
rect 590438 316418 590620 316654
rect 590020 316334 590620 316418
rect 590020 316098 590202 316334
rect 590438 316098 590620 316334
rect 590020 280654 590620 316098
rect 590020 280418 590202 280654
rect 590438 280418 590620 280654
rect 590020 280334 590620 280418
rect 590020 280098 590202 280334
rect 590438 280098 590620 280334
rect 590020 244654 590620 280098
rect 590020 244418 590202 244654
rect 590438 244418 590620 244654
rect 590020 244334 590620 244418
rect 590020 244098 590202 244334
rect 590438 244098 590620 244334
rect 590020 208654 590620 244098
rect 590020 208418 590202 208654
rect 590438 208418 590620 208654
rect 590020 208334 590620 208418
rect 590020 208098 590202 208334
rect 590438 208098 590620 208334
rect 590020 172654 590620 208098
rect 590020 172418 590202 172654
rect 590438 172418 590620 172654
rect 590020 172334 590620 172418
rect 590020 172098 590202 172334
rect 590438 172098 590620 172334
rect 590020 136654 590620 172098
rect 590020 136418 590202 136654
rect 590438 136418 590620 136654
rect 590020 136334 590620 136418
rect 590020 136098 590202 136334
rect 590438 136098 590620 136334
rect 590020 100654 590620 136098
rect 590020 100418 590202 100654
rect 590438 100418 590620 100654
rect 590020 100334 590620 100418
rect 590020 100098 590202 100334
rect 590438 100098 590620 100334
rect 590020 64654 590620 100098
rect 590020 64418 590202 64654
rect 590438 64418 590620 64654
rect 590020 64334 590620 64418
rect 590020 64098 590202 64334
rect 590438 64098 590620 64334
rect 590020 28654 590620 64098
rect 590020 28418 590202 28654
rect 590438 28418 590620 28654
rect 590020 28334 590620 28418
rect 590020 28098 590202 28334
rect 590438 28098 590620 28334
rect 590020 -5046 590620 28098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 698254 591560 709922
rect 590960 698018 591142 698254
rect 591378 698018 591560 698254
rect 590960 697934 591560 698018
rect 590960 697698 591142 697934
rect 591378 697698 591560 697934
rect 590960 662254 591560 697698
rect 590960 662018 591142 662254
rect 591378 662018 591560 662254
rect 590960 661934 591560 662018
rect 590960 661698 591142 661934
rect 591378 661698 591560 661934
rect 590960 626254 591560 661698
rect 590960 626018 591142 626254
rect 591378 626018 591560 626254
rect 590960 625934 591560 626018
rect 590960 625698 591142 625934
rect 591378 625698 591560 625934
rect 590960 590254 591560 625698
rect 590960 590018 591142 590254
rect 591378 590018 591560 590254
rect 590960 589934 591560 590018
rect 590960 589698 591142 589934
rect 591378 589698 591560 589934
rect 590960 554254 591560 589698
rect 590960 554018 591142 554254
rect 591378 554018 591560 554254
rect 590960 553934 591560 554018
rect 590960 553698 591142 553934
rect 591378 553698 591560 553934
rect 590960 518254 591560 553698
rect 590960 518018 591142 518254
rect 591378 518018 591560 518254
rect 590960 517934 591560 518018
rect 590960 517698 591142 517934
rect 591378 517698 591560 517934
rect 590960 482254 591560 517698
rect 590960 482018 591142 482254
rect 591378 482018 591560 482254
rect 590960 481934 591560 482018
rect 590960 481698 591142 481934
rect 591378 481698 591560 481934
rect 590960 446254 591560 481698
rect 590960 446018 591142 446254
rect 591378 446018 591560 446254
rect 590960 445934 591560 446018
rect 590960 445698 591142 445934
rect 591378 445698 591560 445934
rect 590960 410254 591560 445698
rect 590960 410018 591142 410254
rect 591378 410018 591560 410254
rect 590960 409934 591560 410018
rect 590960 409698 591142 409934
rect 591378 409698 591560 409934
rect 590960 374254 591560 409698
rect 590960 374018 591142 374254
rect 591378 374018 591560 374254
rect 590960 373934 591560 374018
rect 590960 373698 591142 373934
rect 591378 373698 591560 373934
rect 590960 338254 591560 373698
rect 590960 338018 591142 338254
rect 591378 338018 591560 338254
rect 590960 337934 591560 338018
rect 590960 337698 591142 337934
rect 591378 337698 591560 337934
rect 590960 302254 591560 337698
rect 590960 302018 591142 302254
rect 591378 302018 591560 302254
rect 590960 301934 591560 302018
rect 590960 301698 591142 301934
rect 591378 301698 591560 301934
rect 590960 266254 591560 301698
rect 590960 266018 591142 266254
rect 591378 266018 591560 266254
rect 590960 265934 591560 266018
rect 590960 265698 591142 265934
rect 591378 265698 591560 265934
rect 590960 230254 591560 265698
rect 590960 230018 591142 230254
rect 591378 230018 591560 230254
rect 590960 229934 591560 230018
rect 590960 229698 591142 229934
rect 591378 229698 591560 229934
rect 590960 194254 591560 229698
rect 590960 194018 591142 194254
rect 591378 194018 591560 194254
rect 590960 193934 591560 194018
rect 590960 193698 591142 193934
rect 591378 193698 591560 193934
rect 590960 158254 591560 193698
rect 590960 158018 591142 158254
rect 591378 158018 591560 158254
rect 590960 157934 591560 158018
rect 590960 157698 591142 157934
rect 591378 157698 591560 157934
rect 590960 122254 591560 157698
rect 590960 122018 591142 122254
rect 591378 122018 591560 122254
rect 590960 121934 591560 122018
rect 590960 121698 591142 121934
rect 591378 121698 591560 121934
rect 590960 86254 591560 121698
rect 590960 86018 591142 86254
rect 591378 86018 591560 86254
rect 590960 85934 591560 86018
rect 590960 85698 591142 85934
rect 591378 85698 591560 85934
rect 590960 50254 591560 85698
rect 590960 50018 591142 50254
rect 591378 50018 591560 50254
rect 590960 49934 591560 50018
rect 590960 49698 591142 49934
rect 591378 49698 591560 49934
rect 590960 14254 591560 49698
rect 590960 14018 591142 14254
rect 591378 14018 591560 14254
rect 590960 13934 591560 14018
rect 590960 13698 591142 13934
rect 591378 13698 591560 13934
rect 590960 -5986 591560 13698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 680254 592500 710862
rect 591900 680018 592082 680254
rect 592318 680018 592500 680254
rect 591900 679934 592500 680018
rect 591900 679698 592082 679934
rect 592318 679698 592500 679934
rect 591900 644254 592500 679698
rect 591900 644018 592082 644254
rect 592318 644018 592500 644254
rect 591900 643934 592500 644018
rect 591900 643698 592082 643934
rect 592318 643698 592500 643934
rect 591900 608254 592500 643698
rect 591900 608018 592082 608254
rect 592318 608018 592500 608254
rect 591900 607934 592500 608018
rect 591900 607698 592082 607934
rect 592318 607698 592500 607934
rect 591900 572254 592500 607698
rect 591900 572018 592082 572254
rect 592318 572018 592500 572254
rect 591900 571934 592500 572018
rect 591900 571698 592082 571934
rect 592318 571698 592500 571934
rect 591900 536254 592500 571698
rect 591900 536018 592082 536254
rect 592318 536018 592500 536254
rect 591900 535934 592500 536018
rect 591900 535698 592082 535934
rect 592318 535698 592500 535934
rect 591900 500254 592500 535698
rect 591900 500018 592082 500254
rect 592318 500018 592500 500254
rect 591900 499934 592500 500018
rect 591900 499698 592082 499934
rect 592318 499698 592500 499934
rect 591900 464254 592500 499698
rect 591900 464018 592082 464254
rect 592318 464018 592500 464254
rect 591900 463934 592500 464018
rect 591900 463698 592082 463934
rect 592318 463698 592500 463934
rect 591900 428254 592500 463698
rect 591900 428018 592082 428254
rect 592318 428018 592500 428254
rect 591900 427934 592500 428018
rect 591900 427698 592082 427934
rect 592318 427698 592500 427934
rect 591900 392254 592500 427698
rect 591900 392018 592082 392254
rect 592318 392018 592500 392254
rect 591900 391934 592500 392018
rect 591900 391698 592082 391934
rect 592318 391698 592500 391934
rect 591900 356254 592500 391698
rect 591900 356018 592082 356254
rect 592318 356018 592500 356254
rect 591900 355934 592500 356018
rect 591900 355698 592082 355934
rect 592318 355698 592500 355934
rect 591900 320254 592500 355698
rect 591900 320018 592082 320254
rect 592318 320018 592500 320254
rect 591900 319934 592500 320018
rect 591900 319698 592082 319934
rect 592318 319698 592500 319934
rect 591900 284254 592500 319698
rect 591900 284018 592082 284254
rect 592318 284018 592500 284254
rect 591900 283934 592500 284018
rect 591900 283698 592082 283934
rect 592318 283698 592500 283934
rect 591900 248254 592500 283698
rect 591900 248018 592082 248254
rect 592318 248018 592500 248254
rect 591900 247934 592500 248018
rect 591900 247698 592082 247934
rect 592318 247698 592500 247934
rect 591900 212254 592500 247698
rect 591900 212018 592082 212254
rect 592318 212018 592500 212254
rect 591900 211934 592500 212018
rect 591900 211698 592082 211934
rect 592318 211698 592500 211934
rect 591900 176254 592500 211698
rect 591900 176018 592082 176254
rect 592318 176018 592500 176254
rect 591900 175934 592500 176018
rect 591900 175698 592082 175934
rect 592318 175698 592500 175934
rect 591900 140254 592500 175698
rect 591900 140018 592082 140254
rect 592318 140018 592500 140254
rect 591900 139934 592500 140018
rect 591900 139698 592082 139934
rect 592318 139698 592500 139934
rect 591900 104254 592500 139698
rect 591900 104018 592082 104254
rect 592318 104018 592500 104254
rect 591900 103934 592500 104018
rect 591900 103698 592082 103934
rect 592318 103698 592500 103934
rect 591900 68254 592500 103698
rect 591900 68018 592082 68254
rect 592318 68018 592500 68254
rect 591900 67934 592500 68018
rect 591900 67698 592082 67934
rect 592318 67698 592500 67934
rect 591900 32254 592500 67698
rect 591900 32018 592082 32254
rect 592318 32018 592500 32254
rect 591900 31934 592500 32018
rect 591900 31698 592082 31934
rect 592318 31698 592500 31934
rect 570604 -7162 570786 -6926
rect 571022 -7162 571204 -6926
rect 570604 -7246 571204 -7162
rect 570604 -7482 570786 -7246
rect 571022 -7482 571204 -7246
rect 570604 -7504 571204 -7482
rect 591900 -6926 592500 31698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 680018 -8158 680254
rect -8394 679698 -8158 679934
rect -8394 644018 -8158 644254
rect -8394 643698 -8158 643934
rect -8394 608018 -8158 608254
rect -8394 607698 -8158 607934
rect -8394 572018 -8158 572254
rect -8394 571698 -8158 571934
rect -8394 536018 -8158 536254
rect -8394 535698 -8158 535934
rect -8394 500018 -8158 500254
rect -8394 499698 -8158 499934
rect -8394 464018 -8158 464254
rect -8394 463698 -8158 463934
rect -8394 428018 -8158 428254
rect -8394 427698 -8158 427934
rect -8394 392018 -8158 392254
rect -8394 391698 -8158 391934
rect -8394 356018 -8158 356254
rect -8394 355698 -8158 355934
rect -8394 320018 -8158 320254
rect -8394 319698 -8158 319934
rect -8394 284018 -8158 284254
rect -8394 283698 -8158 283934
rect -8394 248018 -8158 248254
rect -8394 247698 -8158 247934
rect -8394 212018 -8158 212254
rect -8394 211698 -8158 211934
rect -8394 176018 -8158 176254
rect -8394 175698 -8158 175934
rect -8394 140018 -8158 140254
rect -8394 139698 -8158 139934
rect -8394 104018 -8158 104254
rect -8394 103698 -8158 103934
rect -8394 68018 -8158 68254
rect -8394 67698 -8158 67934
rect -8394 32018 -8158 32254
rect -8394 31698 -8158 31934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 12786 710242 13022 710478
rect 12786 709922 13022 710158
rect -7454 698018 -7218 698254
rect -7454 697698 -7218 697934
rect -7454 662018 -7218 662254
rect -7454 661698 -7218 661934
rect -7454 626018 -7218 626254
rect -7454 625698 -7218 625934
rect -7454 590018 -7218 590254
rect -7454 589698 -7218 589934
rect -7454 554018 -7218 554254
rect -7454 553698 -7218 553934
rect -7454 518018 -7218 518254
rect -7454 517698 -7218 517934
rect -7454 482018 -7218 482254
rect -7454 481698 -7218 481934
rect -7454 446018 -7218 446254
rect -7454 445698 -7218 445934
rect -7454 410018 -7218 410254
rect -7454 409698 -7218 409934
rect -7454 374018 -7218 374254
rect -7454 373698 -7218 373934
rect -7454 338018 -7218 338254
rect -7454 337698 -7218 337934
rect -7454 302018 -7218 302254
rect -7454 301698 -7218 301934
rect -7454 266018 -7218 266254
rect -7454 265698 -7218 265934
rect -7454 230018 -7218 230254
rect -7454 229698 -7218 229934
rect -7454 194018 -7218 194254
rect -7454 193698 -7218 193934
rect -7454 158018 -7218 158254
rect -7454 157698 -7218 157934
rect -7454 122018 -7218 122254
rect -7454 121698 -7218 121934
rect -7454 86018 -7218 86254
rect -7454 85698 -7218 85934
rect -7454 50018 -7218 50254
rect -7454 49698 -7218 49934
rect -7454 14018 -7218 14254
rect -7454 13698 -7218 13934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 676418 -6278 676654
rect -6514 676098 -6278 676334
rect -6514 640418 -6278 640654
rect -6514 640098 -6278 640334
rect -6514 604418 -6278 604654
rect -6514 604098 -6278 604334
rect -6514 568418 -6278 568654
rect -6514 568098 -6278 568334
rect -6514 532418 -6278 532654
rect -6514 532098 -6278 532334
rect -6514 496418 -6278 496654
rect -6514 496098 -6278 496334
rect -6514 460418 -6278 460654
rect -6514 460098 -6278 460334
rect -6514 424418 -6278 424654
rect -6514 424098 -6278 424334
rect -6514 388418 -6278 388654
rect -6514 388098 -6278 388334
rect -6514 352418 -6278 352654
rect -6514 352098 -6278 352334
rect -6514 316418 -6278 316654
rect -6514 316098 -6278 316334
rect -6514 280418 -6278 280654
rect -6514 280098 -6278 280334
rect -6514 244418 -6278 244654
rect -6514 244098 -6278 244334
rect -6514 208418 -6278 208654
rect -6514 208098 -6278 208334
rect -6514 172418 -6278 172654
rect -6514 172098 -6278 172334
rect -6514 136418 -6278 136654
rect -6514 136098 -6278 136334
rect -6514 100418 -6278 100654
rect -6514 100098 -6278 100334
rect -6514 64418 -6278 64654
rect -6514 64098 -6278 64334
rect -6514 28418 -6278 28654
rect -6514 28098 -6278 28334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 9186 708362 9422 708598
rect 9186 708042 9422 708278
rect -5574 694418 -5338 694654
rect -5574 694098 -5338 694334
rect -5574 658418 -5338 658654
rect -5574 658098 -5338 658334
rect -5574 622418 -5338 622654
rect -5574 622098 -5338 622334
rect -5574 586418 -5338 586654
rect -5574 586098 -5338 586334
rect -5574 550418 -5338 550654
rect -5574 550098 -5338 550334
rect -5574 514418 -5338 514654
rect -5574 514098 -5338 514334
rect -5574 478418 -5338 478654
rect -5574 478098 -5338 478334
rect -5574 442418 -5338 442654
rect -5574 442098 -5338 442334
rect -5574 406418 -5338 406654
rect -5574 406098 -5338 406334
rect -5574 370418 -5338 370654
rect -5574 370098 -5338 370334
rect -5574 334418 -5338 334654
rect -5574 334098 -5338 334334
rect -5574 298418 -5338 298654
rect -5574 298098 -5338 298334
rect -5574 262418 -5338 262654
rect -5574 262098 -5338 262334
rect -5574 226418 -5338 226654
rect -5574 226098 -5338 226334
rect -5574 190418 -5338 190654
rect -5574 190098 -5338 190334
rect -5574 154418 -5338 154654
rect -5574 154098 -5338 154334
rect -5574 118418 -5338 118654
rect -5574 118098 -5338 118334
rect -5574 82418 -5338 82654
rect -5574 82098 -5338 82334
rect -5574 46418 -5338 46654
rect -5574 46098 -5338 46334
rect -5574 10418 -5338 10654
rect -5574 10098 -5338 10334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 672818 -4398 673054
rect -4634 672498 -4398 672734
rect -4634 636818 -4398 637054
rect -4634 636498 -4398 636734
rect -4634 600818 -4398 601054
rect -4634 600498 -4398 600734
rect -4634 564818 -4398 565054
rect -4634 564498 -4398 564734
rect -4634 528818 -4398 529054
rect -4634 528498 -4398 528734
rect -4634 492818 -4398 493054
rect -4634 492498 -4398 492734
rect -4634 456818 -4398 457054
rect -4634 456498 -4398 456734
rect -4634 420818 -4398 421054
rect -4634 420498 -4398 420734
rect -4634 384818 -4398 385054
rect -4634 384498 -4398 384734
rect -4634 348818 -4398 349054
rect -4634 348498 -4398 348734
rect -4634 312818 -4398 313054
rect -4634 312498 -4398 312734
rect -4634 276818 -4398 277054
rect -4634 276498 -4398 276734
rect -4634 240818 -4398 241054
rect -4634 240498 -4398 240734
rect -4634 204818 -4398 205054
rect -4634 204498 -4398 204734
rect -4634 168818 -4398 169054
rect -4634 168498 -4398 168734
rect -4634 132818 -4398 133054
rect -4634 132498 -4398 132734
rect -4634 96818 -4398 97054
rect -4634 96498 -4398 96734
rect -4634 60818 -4398 61054
rect -4634 60498 -4398 60734
rect -4634 24818 -4398 25054
rect -4634 24498 -4398 24734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 5586 706482 5822 706718
rect 5586 706162 5822 706398
rect -3694 690818 -3458 691054
rect -3694 690498 -3458 690734
rect -3694 654818 -3458 655054
rect -3694 654498 -3458 654734
rect -3694 618818 -3458 619054
rect -3694 618498 -3458 618734
rect -3694 582818 -3458 583054
rect -3694 582498 -3458 582734
rect -3694 546818 -3458 547054
rect -3694 546498 -3458 546734
rect -3694 510818 -3458 511054
rect -3694 510498 -3458 510734
rect -3694 474818 -3458 475054
rect -3694 474498 -3458 474734
rect -3694 438818 -3458 439054
rect -3694 438498 -3458 438734
rect -3694 402818 -3458 403054
rect -3694 402498 -3458 402734
rect -3694 366818 -3458 367054
rect -3694 366498 -3458 366734
rect -3694 330818 -3458 331054
rect -3694 330498 -3458 330734
rect -3694 294818 -3458 295054
rect -3694 294498 -3458 294734
rect -3694 258818 -3458 259054
rect -3694 258498 -3458 258734
rect -3694 222818 -3458 223054
rect -3694 222498 -3458 222734
rect -3694 186818 -3458 187054
rect -3694 186498 -3458 186734
rect -3694 150818 -3458 151054
rect -3694 150498 -3458 150734
rect -3694 114818 -3458 115054
rect -3694 114498 -3458 114734
rect -3694 78818 -3458 79054
rect -3694 78498 -3458 78734
rect -3694 42818 -3458 43054
rect -3694 42498 -3458 42734
rect -3694 6818 -3458 7054
rect -3694 6498 -3458 6734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 669218 -2518 669454
rect -2754 668898 -2518 669134
rect -2754 633218 -2518 633454
rect -2754 632898 -2518 633134
rect -2754 597218 -2518 597454
rect -2754 596898 -2518 597134
rect -2754 561218 -2518 561454
rect -2754 560898 -2518 561134
rect -2754 525218 -2518 525454
rect -2754 524898 -2518 525134
rect -2754 489218 -2518 489454
rect -2754 488898 -2518 489134
rect -2754 453218 -2518 453454
rect -2754 452898 -2518 453134
rect -2754 417218 -2518 417454
rect -2754 416898 -2518 417134
rect -2754 381218 -2518 381454
rect -2754 380898 -2518 381134
rect -2754 345218 -2518 345454
rect -2754 344898 -2518 345134
rect -2754 309218 -2518 309454
rect -2754 308898 -2518 309134
rect -2754 273218 -2518 273454
rect -2754 272898 -2518 273134
rect -2754 237218 -2518 237454
rect -2754 236898 -2518 237134
rect -2754 201218 -2518 201454
rect -2754 200898 -2518 201134
rect -2754 165218 -2518 165454
rect -2754 164898 -2518 165134
rect -2754 129218 -2518 129454
rect -2754 128898 -2518 129134
rect -2754 93218 -2518 93454
rect -2754 92898 -2518 93134
rect -2754 57218 -2518 57454
rect -2754 56898 -2518 57134
rect -2754 21218 -2518 21454
rect -2754 20898 -2518 21134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 687218 -1578 687454
rect -1814 686898 -1578 687134
rect -1814 651218 -1578 651454
rect -1814 650898 -1578 651134
rect -1814 615218 -1578 615454
rect -1814 614898 -1578 615134
rect -1814 579218 -1578 579454
rect -1814 578898 -1578 579134
rect -1814 543218 -1578 543454
rect -1814 542898 -1578 543134
rect -1814 507218 -1578 507454
rect -1814 506898 -1578 507134
rect -1814 471218 -1578 471454
rect -1814 470898 -1578 471134
rect -1814 435218 -1578 435454
rect -1814 434898 -1578 435134
rect -1814 399218 -1578 399454
rect -1814 398898 -1578 399134
rect -1814 363218 -1578 363454
rect -1814 362898 -1578 363134
rect -1814 327218 -1578 327454
rect -1814 326898 -1578 327134
rect -1814 291218 -1578 291454
rect -1814 290898 -1578 291134
rect -1814 255218 -1578 255454
rect -1814 254898 -1578 255134
rect -1814 219218 -1578 219454
rect -1814 218898 -1578 219134
rect -1814 183218 -1578 183454
rect -1814 182898 -1578 183134
rect -1814 147218 -1578 147454
rect -1814 146898 -1578 147134
rect -1814 111218 -1578 111454
rect -1814 110898 -1578 111134
rect -1814 75218 -1578 75454
rect -1814 74898 -1578 75134
rect -1814 39218 -1578 39454
rect -1814 38898 -1578 39134
rect -1814 3218 -1578 3454
rect -1814 2898 -1578 3134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 1986 704602 2222 704838
rect 1986 704282 2222 704518
rect 1986 687218 2222 687454
rect 1986 686898 2222 687134
rect 1986 651218 2222 651454
rect 1986 650898 2222 651134
rect 1986 615218 2222 615454
rect 1986 614898 2222 615134
rect 1986 579218 2222 579454
rect 1986 578898 2222 579134
rect 1986 543218 2222 543454
rect 1986 542898 2222 543134
rect 1986 507218 2222 507454
rect 1986 506898 2222 507134
rect 5586 690818 5822 691054
rect 5586 690498 5822 690734
rect 5586 654818 5822 655054
rect 5586 654498 5822 654734
rect 5586 618818 5822 619054
rect 5586 618498 5822 618734
rect 5586 582818 5822 583054
rect 5586 582498 5822 582734
rect 5586 546818 5822 547054
rect 5586 546498 5822 546734
rect 5586 510818 5822 511054
rect 5586 510498 5822 510734
rect 1986 471218 2222 471454
rect 1986 470898 2222 471134
rect 1986 435218 2222 435454
rect 1986 434898 2222 435134
rect 1986 399218 2222 399454
rect 1986 398898 2222 399134
rect 1986 363218 2222 363454
rect 1986 362898 2222 363134
rect 1986 327218 2222 327454
rect 1986 326898 2222 327134
rect 1986 291218 2222 291454
rect 1986 290898 2222 291134
rect 1986 255218 2222 255454
rect 1986 254898 2222 255134
rect 1986 219218 2222 219454
rect 1986 218898 2222 219134
rect 1986 183218 2222 183454
rect 1986 182898 2222 183134
rect 1986 147218 2222 147454
rect 1986 146898 2222 147134
rect 1986 111218 2222 111454
rect 1986 110898 2222 111134
rect 1986 75218 2222 75454
rect 1986 74898 2222 75134
rect 1986 39218 2222 39454
rect 1986 38898 2222 39134
rect 1986 3218 2222 3454
rect 1986 2898 2222 3134
rect 1986 -582 2222 -346
rect 1986 -902 2222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 5586 474818 5822 475054
rect 5586 474498 5822 474734
rect 5586 438818 5822 439054
rect 5586 438498 5822 438734
rect 5586 402818 5822 403054
rect 5586 402498 5822 402734
rect 5586 366818 5822 367054
rect 5586 366498 5822 366734
rect 5586 330818 5822 331054
rect 5586 330498 5822 330734
rect 5586 294818 5822 295054
rect 5586 294498 5822 294734
rect 5586 258818 5822 259054
rect 5586 258498 5822 258734
rect 5586 222818 5822 223054
rect 5586 222498 5822 222734
rect 5586 186818 5822 187054
rect 5586 186498 5822 186734
rect 5586 150818 5822 151054
rect 5586 150498 5822 150734
rect 5586 114818 5822 115054
rect 5586 114498 5822 114734
rect 5586 78818 5822 79054
rect 5586 78498 5822 78734
rect 5586 42818 5822 43054
rect 5586 42498 5822 42734
rect 5586 6818 5822 7054
rect 5586 6498 5822 6734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 5586 -2462 5822 -2226
rect 5586 -2782 5822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 9186 694418 9422 694654
rect 9186 694098 9422 694334
rect 9186 658418 9422 658654
rect 9186 658098 9422 658334
rect 9186 622418 9422 622654
rect 9186 622098 9422 622334
rect 9186 586418 9422 586654
rect 9186 586098 9422 586334
rect 9186 550418 9422 550654
rect 9186 550098 9422 550334
rect 9186 514418 9422 514654
rect 9186 514098 9422 514334
rect 9186 478418 9422 478654
rect 9186 478098 9422 478334
rect 9186 442418 9422 442654
rect 9186 442098 9422 442334
rect 9186 406418 9422 406654
rect 9186 406098 9422 406334
rect 9186 370418 9422 370654
rect 9186 370098 9422 370334
rect 9186 334418 9422 334654
rect 9186 334098 9422 334334
rect 9186 298418 9422 298654
rect 9186 298098 9422 298334
rect 9186 262418 9422 262654
rect 9186 262098 9422 262334
rect 9186 226418 9422 226654
rect 9186 226098 9422 226334
rect 9186 190418 9422 190654
rect 9186 190098 9422 190334
rect 9186 154418 9422 154654
rect 9186 154098 9422 154334
rect 9186 118418 9422 118654
rect 9186 118098 9422 118334
rect 9186 82418 9422 82654
rect 9186 82098 9422 82334
rect 9186 46418 9422 46654
rect 9186 46098 9422 46334
rect 9186 10418 9422 10654
rect 9186 10098 9422 10334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 9186 -4342 9422 -4106
rect 9186 -4662 9422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 30786 711182 31022 711418
rect 30786 710862 31022 711098
rect 27186 709302 27422 709538
rect 27186 708982 27422 709218
rect 23586 707422 23822 707658
rect 23586 707102 23822 707338
rect 12786 698018 13022 698254
rect 12786 697698 13022 697934
rect 12786 662018 13022 662254
rect 12786 661698 13022 661934
rect 12786 626018 13022 626254
rect 12786 625698 13022 625934
rect 12786 590018 13022 590254
rect 12786 589698 13022 589934
rect 12786 554018 13022 554254
rect 12786 553698 13022 553934
rect 12786 518018 13022 518254
rect 12786 517698 13022 517934
rect 12786 482018 13022 482254
rect 12786 481698 13022 481934
rect 12786 446018 13022 446254
rect 12786 445698 13022 445934
rect 12786 410018 13022 410254
rect 12786 409698 13022 409934
rect 12786 374018 13022 374254
rect 12786 373698 13022 373934
rect 12786 338018 13022 338254
rect 12786 337698 13022 337934
rect 12786 302018 13022 302254
rect 12786 301698 13022 301934
rect 12786 266018 13022 266254
rect 12786 265698 13022 265934
rect 12786 230018 13022 230254
rect 12786 229698 13022 229934
rect 12786 194018 13022 194254
rect 12786 193698 13022 193934
rect 12786 158018 13022 158254
rect 12786 157698 13022 157934
rect 12786 122018 13022 122254
rect 12786 121698 13022 121934
rect 12786 86018 13022 86254
rect 12786 85698 13022 85934
rect 12786 50018 13022 50254
rect 12786 49698 13022 49934
rect 12786 14018 13022 14254
rect 12786 13698 13022 13934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 19986 705542 20222 705778
rect 19986 705222 20222 705458
rect 19986 669218 20222 669454
rect 19986 668898 20222 669134
rect 19986 633218 20222 633454
rect 19986 632898 20222 633134
rect 19986 597218 20222 597454
rect 19986 596898 20222 597134
rect 19986 561218 20222 561454
rect 19986 560898 20222 561134
rect 19986 525218 20222 525454
rect 19986 524898 20222 525134
rect 19986 489218 20222 489454
rect 19986 488898 20222 489134
rect 19986 453218 20222 453454
rect 19986 452898 20222 453134
rect 19986 417218 20222 417454
rect 19986 416898 20222 417134
rect 19986 381218 20222 381454
rect 19986 380898 20222 381134
rect 19986 345218 20222 345454
rect 19986 344898 20222 345134
rect 19986 309218 20222 309454
rect 19986 308898 20222 309134
rect 19986 273218 20222 273454
rect 19986 272898 20222 273134
rect 19986 237218 20222 237454
rect 19986 236898 20222 237134
rect 19986 201218 20222 201454
rect 19986 200898 20222 201134
rect 19986 165218 20222 165454
rect 19986 164898 20222 165134
rect 19986 129218 20222 129454
rect 19986 128898 20222 129134
rect 19986 93218 20222 93454
rect 19986 92898 20222 93134
rect 19986 57218 20222 57454
rect 19986 56898 20222 57134
rect 19986 21218 20222 21454
rect 19986 20898 20222 21134
rect 19986 -1522 20222 -1286
rect 19986 -1842 20222 -1606
rect 23586 672818 23822 673054
rect 23586 672498 23822 672734
rect 23586 636818 23822 637054
rect 23586 636498 23822 636734
rect 23586 600818 23822 601054
rect 23586 600498 23822 600734
rect 23586 564818 23822 565054
rect 23586 564498 23822 564734
rect 23586 528818 23822 529054
rect 23586 528498 23822 528734
rect 23586 492818 23822 493054
rect 23586 492498 23822 492734
rect 23586 456818 23822 457054
rect 23586 456498 23822 456734
rect 23586 420818 23822 421054
rect 23586 420498 23822 420734
rect 23586 384818 23822 385054
rect 23586 384498 23822 384734
rect 23586 348818 23822 349054
rect 23586 348498 23822 348734
rect 23586 312818 23822 313054
rect 23586 312498 23822 312734
rect 23586 276818 23822 277054
rect 23586 276498 23822 276734
rect 23586 240818 23822 241054
rect 23586 240498 23822 240734
rect 23586 204818 23822 205054
rect 23586 204498 23822 204734
rect 23586 168818 23822 169054
rect 23586 168498 23822 168734
rect 23586 132818 23822 133054
rect 23586 132498 23822 132734
rect 23586 96818 23822 97054
rect 23586 96498 23822 96734
rect 23586 60818 23822 61054
rect 23586 60498 23822 60734
rect 23586 24818 23822 25054
rect 23586 24498 23822 24734
rect 23586 -3402 23822 -3166
rect 23586 -3722 23822 -3486
rect 27186 676418 27422 676654
rect 27186 676098 27422 676334
rect 27186 640418 27422 640654
rect 27186 640098 27422 640334
rect 27186 604418 27422 604654
rect 27186 604098 27422 604334
rect 27186 568418 27422 568654
rect 27186 568098 27422 568334
rect 27186 532418 27422 532654
rect 27186 532098 27422 532334
rect 27186 496418 27422 496654
rect 27186 496098 27422 496334
rect 27186 460418 27422 460654
rect 27186 460098 27422 460334
rect 27186 424418 27422 424654
rect 27186 424098 27422 424334
rect 27186 388418 27422 388654
rect 27186 388098 27422 388334
rect 27186 352418 27422 352654
rect 27186 352098 27422 352334
rect 27186 316418 27422 316654
rect 27186 316098 27422 316334
rect 27186 280418 27422 280654
rect 27186 280098 27422 280334
rect 27186 244418 27422 244654
rect 27186 244098 27422 244334
rect 27186 208418 27422 208654
rect 27186 208098 27422 208334
rect 27186 172418 27422 172654
rect 27186 172098 27422 172334
rect 27186 136418 27422 136654
rect 27186 136098 27422 136334
rect 27186 100418 27422 100654
rect 27186 100098 27422 100334
rect 27186 64418 27422 64654
rect 27186 64098 27422 64334
rect 27186 28418 27422 28654
rect 27186 28098 27422 28334
rect 27186 -5282 27422 -5046
rect 27186 -5602 27422 -5366
rect 48786 710242 49022 710478
rect 48786 709922 49022 710158
rect 45186 708362 45422 708598
rect 45186 708042 45422 708278
rect 41586 706482 41822 706718
rect 41586 706162 41822 706398
rect 30786 680018 31022 680254
rect 30786 679698 31022 679934
rect 30786 644018 31022 644254
rect 30786 643698 31022 643934
rect 30786 608018 31022 608254
rect 30786 607698 31022 607934
rect 30786 572018 31022 572254
rect 30786 571698 31022 571934
rect 30786 536018 31022 536254
rect 30786 535698 31022 535934
rect 30786 500018 31022 500254
rect 30786 499698 31022 499934
rect 30786 464018 31022 464254
rect 30786 463698 31022 463934
rect 30786 428018 31022 428254
rect 30786 427698 31022 427934
rect 30786 392018 31022 392254
rect 30786 391698 31022 391934
rect 30786 356018 31022 356254
rect 30786 355698 31022 355934
rect 30786 320018 31022 320254
rect 30786 319698 31022 319934
rect 30786 284018 31022 284254
rect 30786 283698 31022 283934
rect 30786 248018 31022 248254
rect 30786 247698 31022 247934
rect 30786 212018 31022 212254
rect 30786 211698 31022 211934
rect 30786 176018 31022 176254
rect 30786 175698 31022 175934
rect 30786 140018 31022 140254
rect 30786 139698 31022 139934
rect 30786 104018 31022 104254
rect 30786 103698 31022 103934
rect 30786 68018 31022 68254
rect 30786 67698 31022 67934
rect 30786 32018 31022 32254
rect 30786 31698 31022 31934
rect 12786 -6222 13022 -5986
rect 12786 -6542 13022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 37986 704602 38222 704838
rect 37986 704282 38222 704518
rect 37986 687218 38222 687454
rect 37986 686898 38222 687134
rect 37986 651218 38222 651454
rect 37986 650898 38222 651134
rect 37986 615218 38222 615454
rect 37986 614898 38222 615134
rect 37986 579218 38222 579454
rect 37986 578898 38222 579134
rect 37986 543218 38222 543454
rect 37986 542898 38222 543134
rect 37986 507218 38222 507454
rect 37986 506898 38222 507134
rect 37986 471218 38222 471454
rect 37986 470898 38222 471134
rect 37986 435218 38222 435454
rect 37986 434898 38222 435134
rect 37986 399218 38222 399454
rect 37986 398898 38222 399134
rect 37986 363218 38222 363454
rect 37986 362898 38222 363134
rect 37986 327218 38222 327454
rect 37986 326898 38222 327134
rect 37986 291218 38222 291454
rect 37986 290898 38222 291134
rect 37986 255218 38222 255454
rect 37986 254898 38222 255134
rect 37986 219218 38222 219454
rect 37986 218898 38222 219134
rect 37986 183218 38222 183454
rect 37986 182898 38222 183134
rect 37986 147218 38222 147454
rect 37986 146898 38222 147134
rect 37986 111218 38222 111454
rect 37986 110898 38222 111134
rect 37986 75218 38222 75454
rect 37986 74898 38222 75134
rect 37986 39218 38222 39454
rect 37986 38898 38222 39134
rect 37986 3218 38222 3454
rect 37986 2898 38222 3134
rect 37986 -582 38222 -346
rect 37986 -902 38222 -666
rect 41586 690818 41822 691054
rect 41586 690498 41822 690734
rect 41586 654818 41822 655054
rect 41586 654498 41822 654734
rect 41586 618818 41822 619054
rect 41586 618498 41822 618734
rect 41586 582818 41822 583054
rect 41586 582498 41822 582734
rect 41586 546818 41822 547054
rect 41586 546498 41822 546734
rect 41586 510818 41822 511054
rect 41586 510498 41822 510734
rect 41586 474818 41822 475054
rect 41586 474498 41822 474734
rect 41586 438818 41822 439054
rect 41586 438498 41822 438734
rect 41586 402818 41822 403054
rect 41586 402498 41822 402734
rect 41586 366818 41822 367054
rect 41586 366498 41822 366734
rect 41586 330818 41822 331054
rect 41586 330498 41822 330734
rect 41586 294818 41822 295054
rect 41586 294498 41822 294734
rect 41586 258818 41822 259054
rect 41586 258498 41822 258734
rect 41586 222818 41822 223054
rect 41586 222498 41822 222734
rect 41586 186818 41822 187054
rect 41586 186498 41822 186734
rect 41586 150818 41822 151054
rect 41586 150498 41822 150734
rect 41586 114818 41822 115054
rect 41586 114498 41822 114734
rect 41586 78818 41822 79054
rect 41586 78498 41822 78734
rect 41586 42818 41822 43054
rect 41586 42498 41822 42734
rect 41586 6818 41822 7054
rect 41586 6498 41822 6734
rect 41586 -2462 41822 -2226
rect 41586 -2782 41822 -2546
rect 45186 694418 45422 694654
rect 45186 694098 45422 694334
rect 45186 658418 45422 658654
rect 45186 658098 45422 658334
rect 45186 622418 45422 622654
rect 45186 622098 45422 622334
rect 45186 586418 45422 586654
rect 45186 586098 45422 586334
rect 45186 550418 45422 550654
rect 45186 550098 45422 550334
rect 45186 514418 45422 514654
rect 45186 514098 45422 514334
rect 45186 478418 45422 478654
rect 45186 478098 45422 478334
rect 45186 442418 45422 442654
rect 45186 442098 45422 442334
rect 45186 406418 45422 406654
rect 45186 406098 45422 406334
rect 45186 370418 45422 370654
rect 45186 370098 45422 370334
rect 45186 334418 45422 334654
rect 45186 334098 45422 334334
rect 45186 298418 45422 298654
rect 45186 298098 45422 298334
rect 45186 262418 45422 262654
rect 45186 262098 45422 262334
rect 45186 226418 45422 226654
rect 45186 226098 45422 226334
rect 45186 190418 45422 190654
rect 45186 190098 45422 190334
rect 45186 154418 45422 154654
rect 45186 154098 45422 154334
rect 45186 118418 45422 118654
rect 45186 118098 45422 118334
rect 45186 82418 45422 82654
rect 45186 82098 45422 82334
rect 45186 46418 45422 46654
rect 45186 46098 45422 46334
rect 45186 10418 45422 10654
rect 45186 10098 45422 10334
rect 45186 -4342 45422 -4106
rect 45186 -4662 45422 -4426
rect 66786 711182 67022 711418
rect 66786 710862 67022 711098
rect 63186 709302 63422 709538
rect 63186 708982 63422 709218
rect 59586 707422 59822 707658
rect 59586 707102 59822 707338
rect 48786 698018 49022 698254
rect 48786 697698 49022 697934
rect 48786 662018 49022 662254
rect 48786 661698 49022 661934
rect 48786 626018 49022 626254
rect 48786 625698 49022 625934
rect 48786 590018 49022 590254
rect 48786 589698 49022 589934
rect 48786 554018 49022 554254
rect 48786 553698 49022 553934
rect 48786 518018 49022 518254
rect 48786 517698 49022 517934
rect 48786 482018 49022 482254
rect 48786 481698 49022 481934
rect 48786 446018 49022 446254
rect 48786 445698 49022 445934
rect 48786 410018 49022 410254
rect 48786 409698 49022 409934
rect 48786 374018 49022 374254
rect 48786 373698 49022 373934
rect 48786 338018 49022 338254
rect 48786 337698 49022 337934
rect 48786 302018 49022 302254
rect 48786 301698 49022 301934
rect 48786 266018 49022 266254
rect 48786 265698 49022 265934
rect 48786 230018 49022 230254
rect 48786 229698 49022 229934
rect 48786 194018 49022 194254
rect 48786 193698 49022 193934
rect 48786 158018 49022 158254
rect 48786 157698 49022 157934
rect 48786 122018 49022 122254
rect 48786 121698 49022 121934
rect 48786 86018 49022 86254
rect 48786 85698 49022 85934
rect 48786 50018 49022 50254
rect 48786 49698 49022 49934
rect 48786 14018 49022 14254
rect 48786 13698 49022 13934
rect 30786 -7162 31022 -6926
rect 30786 -7482 31022 -7246
rect 55986 705542 56222 705778
rect 55986 705222 56222 705458
rect 55986 669218 56222 669454
rect 55986 668898 56222 669134
rect 55986 633218 56222 633454
rect 55986 632898 56222 633134
rect 55986 597218 56222 597454
rect 55986 596898 56222 597134
rect 55986 561218 56222 561454
rect 55986 560898 56222 561134
rect 55986 525218 56222 525454
rect 55986 524898 56222 525134
rect 55986 489218 56222 489454
rect 55986 488898 56222 489134
rect 55986 453218 56222 453454
rect 55986 452898 56222 453134
rect 55986 417218 56222 417454
rect 55986 416898 56222 417134
rect 55986 381218 56222 381454
rect 55986 380898 56222 381134
rect 55986 345218 56222 345454
rect 55986 344898 56222 345134
rect 55986 309218 56222 309454
rect 55986 308898 56222 309134
rect 55986 273218 56222 273454
rect 55986 272898 56222 273134
rect 55986 237218 56222 237454
rect 55986 236898 56222 237134
rect 55986 201218 56222 201454
rect 55986 200898 56222 201134
rect 55986 165218 56222 165454
rect 55986 164898 56222 165134
rect 55986 129218 56222 129454
rect 55986 128898 56222 129134
rect 55986 93218 56222 93454
rect 55986 92898 56222 93134
rect 55986 57218 56222 57454
rect 55986 56898 56222 57134
rect 55986 21218 56222 21454
rect 55986 20898 56222 21134
rect 55986 -1522 56222 -1286
rect 55986 -1842 56222 -1606
rect 59586 672818 59822 673054
rect 59586 672498 59822 672734
rect 59586 636818 59822 637054
rect 59586 636498 59822 636734
rect 59586 600818 59822 601054
rect 59586 600498 59822 600734
rect 59586 564818 59822 565054
rect 59586 564498 59822 564734
rect 59586 528818 59822 529054
rect 59586 528498 59822 528734
rect 59586 492818 59822 493054
rect 59586 492498 59822 492734
rect 59586 456818 59822 457054
rect 59586 456498 59822 456734
rect 59586 420818 59822 421054
rect 59586 420498 59822 420734
rect 59586 384818 59822 385054
rect 59586 384498 59822 384734
rect 59586 348818 59822 349054
rect 59586 348498 59822 348734
rect 59586 312818 59822 313054
rect 59586 312498 59822 312734
rect 59586 276818 59822 277054
rect 59586 276498 59822 276734
rect 59586 240818 59822 241054
rect 59586 240498 59822 240734
rect 59586 204818 59822 205054
rect 59586 204498 59822 204734
rect 59586 168818 59822 169054
rect 59586 168498 59822 168734
rect 59586 132818 59822 133054
rect 59586 132498 59822 132734
rect 59586 96818 59822 97054
rect 59586 96498 59822 96734
rect 59586 60818 59822 61054
rect 59586 60498 59822 60734
rect 59586 24818 59822 25054
rect 59586 24498 59822 24734
rect 59586 -3402 59822 -3166
rect 59586 -3722 59822 -3486
rect 63186 676418 63422 676654
rect 63186 676098 63422 676334
rect 63186 640418 63422 640654
rect 63186 640098 63422 640334
rect 63186 604418 63422 604654
rect 63186 604098 63422 604334
rect 63186 568418 63422 568654
rect 63186 568098 63422 568334
rect 63186 532418 63422 532654
rect 63186 532098 63422 532334
rect 63186 496418 63422 496654
rect 63186 496098 63422 496334
rect 63186 460418 63422 460654
rect 63186 460098 63422 460334
rect 63186 424418 63422 424654
rect 63186 424098 63422 424334
rect 63186 388418 63422 388654
rect 63186 388098 63422 388334
rect 63186 352418 63422 352654
rect 63186 352098 63422 352334
rect 63186 316418 63422 316654
rect 63186 316098 63422 316334
rect 63186 280418 63422 280654
rect 63186 280098 63422 280334
rect 63186 244418 63422 244654
rect 63186 244098 63422 244334
rect 63186 208418 63422 208654
rect 63186 208098 63422 208334
rect 63186 172418 63422 172654
rect 63186 172098 63422 172334
rect 63186 136418 63422 136654
rect 63186 136098 63422 136334
rect 63186 100418 63422 100654
rect 63186 100098 63422 100334
rect 63186 64418 63422 64654
rect 63186 64098 63422 64334
rect 63186 28418 63422 28654
rect 63186 28098 63422 28334
rect 63186 -5282 63422 -5046
rect 63186 -5602 63422 -5366
rect 84786 710242 85022 710478
rect 84786 709922 85022 710158
rect 81186 708362 81422 708598
rect 81186 708042 81422 708278
rect 77586 706482 77822 706718
rect 77586 706162 77822 706398
rect 66786 680018 67022 680254
rect 66786 679698 67022 679934
rect 66786 644018 67022 644254
rect 66786 643698 67022 643934
rect 66786 608018 67022 608254
rect 66786 607698 67022 607934
rect 66786 572018 67022 572254
rect 66786 571698 67022 571934
rect 66786 536018 67022 536254
rect 66786 535698 67022 535934
rect 66786 500018 67022 500254
rect 66786 499698 67022 499934
rect 66786 464018 67022 464254
rect 66786 463698 67022 463934
rect 66786 428018 67022 428254
rect 66786 427698 67022 427934
rect 66786 392018 67022 392254
rect 66786 391698 67022 391934
rect 66786 356018 67022 356254
rect 66786 355698 67022 355934
rect 66786 320018 67022 320254
rect 66786 319698 67022 319934
rect 66786 284018 67022 284254
rect 66786 283698 67022 283934
rect 66786 248018 67022 248254
rect 66786 247698 67022 247934
rect 66786 212018 67022 212254
rect 66786 211698 67022 211934
rect 66786 176018 67022 176254
rect 66786 175698 67022 175934
rect 66786 140018 67022 140254
rect 66786 139698 67022 139934
rect 66786 104018 67022 104254
rect 66786 103698 67022 103934
rect 66786 68018 67022 68254
rect 66786 67698 67022 67934
rect 66786 32018 67022 32254
rect 66786 31698 67022 31934
rect 48786 -6222 49022 -5986
rect 48786 -6542 49022 -6306
rect 73986 704602 74222 704838
rect 73986 704282 74222 704518
rect 73986 687218 74222 687454
rect 73986 686898 74222 687134
rect 73986 651218 74222 651454
rect 73986 650898 74222 651134
rect 73986 615218 74222 615454
rect 73986 614898 74222 615134
rect 73986 579218 74222 579454
rect 73986 578898 74222 579134
rect 73986 543218 74222 543454
rect 73986 542898 74222 543134
rect 73986 507218 74222 507454
rect 73986 506898 74222 507134
rect 73986 471218 74222 471454
rect 73986 470898 74222 471134
rect 73986 435218 74222 435454
rect 73986 434898 74222 435134
rect 73986 399218 74222 399454
rect 73986 398898 74222 399134
rect 73986 363218 74222 363454
rect 73986 362898 74222 363134
rect 73986 327218 74222 327454
rect 73986 326898 74222 327134
rect 73986 291218 74222 291454
rect 73986 290898 74222 291134
rect 73986 255218 74222 255454
rect 73986 254898 74222 255134
rect 73986 219218 74222 219454
rect 73986 218898 74222 219134
rect 73986 183218 74222 183454
rect 73986 182898 74222 183134
rect 73986 147218 74222 147454
rect 73986 146898 74222 147134
rect 73986 111218 74222 111454
rect 73986 110898 74222 111134
rect 73986 75218 74222 75454
rect 73986 74898 74222 75134
rect 73986 39218 74222 39454
rect 73986 38898 74222 39134
rect 73986 3218 74222 3454
rect 73986 2898 74222 3134
rect 73986 -582 74222 -346
rect 73986 -902 74222 -666
rect 77586 690818 77822 691054
rect 77586 690498 77822 690734
rect 77586 654818 77822 655054
rect 77586 654498 77822 654734
rect 77586 618818 77822 619054
rect 77586 618498 77822 618734
rect 77586 582818 77822 583054
rect 77586 582498 77822 582734
rect 77586 546818 77822 547054
rect 77586 546498 77822 546734
rect 77586 510818 77822 511054
rect 77586 510498 77822 510734
rect 77586 474818 77822 475054
rect 77586 474498 77822 474734
rect 77586 438818 77822 439054
rect 77586 438498 77822 438734
rect 77586 402818 77822 403054
rect 77586 402498 77822 402734
rect 77586 366818 77822 367054
rect 77586 366498 77822 366734
rect 77586 330818 77822 331054
rect 77586 330498 77822 330734
rect 77586 294818 77822 295054
rect 77586 294498 77822 294734
rect 77586 258818 77822 259054
rect 77586 258498 77822 258734
rect 77586 222818 77822 223054
rect 77586 222498 77822 222734
rect 77586 186818 77822 187054
rect 77586 186498 77822 186734
rect 77586 150818 77822 151054
rect 77586 150498 77822 150734
rect 77586 114818 77822 115054
rect 77586 114498 77822 114734
rect 77586 78818 77822 79054
rect 77586 78498 77822 78734
rect 77586 42818 77822 43054
rect 77586 42498 77822 42734
rect 77586 6818 77822 7054
rect 77586 6498 77822 6734
rect 77586 -2462 77822 -2226
rect 77586 -2782 77822 -2546
rect 81186 694418 81422 694654
rect 81186 694098 81422 694334
rect 81186 658418 81422 658654
rect 81186 658098 81422 658334
rect 81186 622418 81422 622654
rect 81186 622098 81422 622334
rect 81186 586418 81422 586654
rect 81186 586098 81422 586334
rect 81186 550418 81422 550654
rect 81186 550098 81422 550334
rect 81186 514418 81422 514654
rect 81186 514098 81422 514334
rect 81186 478418 81422 478654
rect 81186 478098 81422 478334
rect 81186 442418 81422 442654
rect 81186 442098 81422 442334
rect 81186 406418 81422 406654
rect 81186 406098 81422 406334
rect 81186 370418 81422 370654
rect 81186 370098 81422 370334
rect 81186 334418 81422 334654
rect 81186 334098 81422 334334
rect 81186 298418 81422 298654
rect 81186 298098 81422 298334
rect 81186 262418 81422 262654
rect 81186 262098 81422 262334
rect 81186 226418 81422 226654
rect 81186 226098 81422 226334
rect 81186 190418 81422 190654
rect 81186 190098 81422 190334
rect 81186 154418 81422 154654
rect 81186 154098 81422 154334
rect 81186 118418 81422 118654
rect 81186 118098 81422 118334
rect 81186 82418 81422 82654
rect 81186 82098 81422 82334
rect 81186 46418 81422 46654
rect 81186 46098 81422 46334
rect 81186 10418 81422 10654
rect 81186 10098 81422 10334
rect 81186 -4342 81422 -4106
rect 81186 -4662 81422 -4426
rect 102786 711182 103022 711418
rect 102786 710862 103022 711098
rect 99186 709302 99422 709538
rect 99186 708982 99422 709218
rect 95586 707422 95822 707658
rect 95586 707102 95822 707338
rect 84786 698018 85022 698254
rect 84786 697698 85022 697934
rect 84786 662018 85022 662254
rect 84786 661698 85022 661934
rect 84786 626018 85022 626254
rect 84786 625698 85022 625934
rect 84786 590018 85022 590254
rect 84786 589698 85022 589934
rect 84786 554018 85022 554254
rect 84786 553698 85022 553934
rect 84786 518018 85022 518254
rect 84786 517698 85022 517934
rect 84786 482018 85022 482254
rect 84786 481698 85022 481934
rect 84786 446018 85022 446254
rect 84786 445698 85022 445934
rect 84786 410018 85022 410254
rect 84786 409698 85022 409934
rect 84786 374018 85022 374254
rect 84786 373698 85022 373934
rect 84786 338018 85022 338254
rect 84786 337698 85022 337934
rect 84786 302018 85022 302254
rect 84786 301698 85022 301934
rect 84786 266018 85022 266254
rect 84786 265698 85022 265934
rect 84786 230018 85022 230254
rect 84786 229698 85022 229934
rect 84786 194018 85022 194254
rect 84786 193698 85022 193934
rect 84786 158018 85022 158254
rect 84786 157698 85022 157934
rect 84786 122018 85022 122254
rect 84786 121698 85022 121934
rect 84786 86018 85022 86254
rect 84786 85698 85022 85934
rect 84786 50018 85022 50254
rect 84786 49698 85022 49934
rect 84786 14018 85022 14254
rect 84786 13698 85022 13934
rect 66786 -7162 67022 -6926
rect 66786 -7482 67022 -7246
rect 91986 705542 92222 705778
rect 91986 705222 92222 705458
rect 91986 669218 92222 669454
rect 91986 668898 92222 669134
rect 91986 633218 92222 633454
rect 91986 632898 92222 633134
rect 91986 597218 92222 597454
rect 91986 596898 92222 597134
rect 91986 561218 92222 561454
rect 91986 560898 92222 561134
rect 91986 525218 92222 525454
rect 91986 524898 92222 525134
rect 91986 489218 92222 489454
rect 91986 488898 92222 489134
rect 91986 453218 92222 453454
rect 91986 452898 92222 453134
rect 91986 417218 92222 417454
rect 91986 416898 92222 417134
rect 91986 381218 92222 381454
rect 91986 380898 92222 381134
rect 91986 345218 92222 345454
rect 91986 344898 92222 345134
rect 91986 309218 92222 309454
rect 91986 308898 92222 309134
rect 91986 273218 92222 273454
rect 91986 272898 92222 273134
rect 91986 237218 92222 237454
rect 91986 236898 92222 237134
rect 91986 201218 92222 201454
rect 91986 200898 92222 201134
rect 91986 165218 92222 165454
rect 91986 164898 92222 165134
rect 91986 129218 92222 129454
rect 91986 128898 92222 129134
rect 91986 93218 92222 93454
rect 91986 92898 92222 93134
rect 91986 57218 92222 57454
rect 91986 56898 92222 57134
rect 91986 21218 92222 21454
rect 91986 20898 92222 21134
rect 91986 -1522 92222 -1286
rect 91986 -1842 92222 -1606
rect 95586 672818 95822 673054
rect 95586 672498 95822 672734
rect 95586 636818 95822 637054
rect 95586 636498 95822 636734
rect 95586 600818 95822 601054
rect 95586 600498 95822 600734
rect 95586 564818 95822 565054
rect 95586 564498 95822 564734
rect 95586 528818 95822 529054
rect 95586 528498 95822 528734
rect 95586 492818 95822 493054
rect 95586 492498 95822 492734
rect 95586 456818 95822 457054
rect 95586 456498 95822 456734
rect 95586 420818 95822 421054
rect 95586 420498 95822 420734
rect 95586 384818 95822 385054
rect 95586 384498 95822 384734
rect 95586 348818 95822 349054
rect 95586 348498 95822 348734
rect 95586 312818 95822 313054
rect 95586 312498 95822 312734
rect 95586 276818 95822 277054
rect 95586 276498 95822 276734
rect 95586 240818 95822 241054
rect 95586 240498 95822 240734
rect 95586 204818 95822 205054
rect 95586 204498 95822 204734
rect 95586 168818 95822 169054
rect 95586 168498 95822 168734
rect 95586 132818 95822 133054
rect 95586 132498 95822 132734
rect 95586 96818 95822 97054
rect 95586 96498 95822 96734
rect 95586 60818 95822 61054
rect 95586 60498 95822 60734
rect 95586 24818 95822 25054
rect 95586 24498 95822 24734
rect 95586 -3402 95822 -3166
rect 95586 -3722 95822 -3486
rect 99186 676418 99422 676654
rect 99186 676098 99422 676334
rect 99186 640418 99422 640654
rect 99186 640098 99422 640334
rect 99186 604418 99422 604654
rect 99186 604098 99422 604334
rect 99186 568418 99422 568654
rect 99186 568098 99422 568334
rect 99186 532418 99422 532654
rect 99186 532098 99422 532334
rect 99186 496418 99422 496654
rect 99186 496098 99422 496334
rect 99186 460418 99422 460654
rect 99186 460098 99422 460334
rect 99186 424418 99422 424654
rect 99186 424098 99422 424334
rect 99186 388418 99422 388654
rect 99186 388098 99422 388334
rect 99186 352418 99422 352654
rect 99186 352098 99422 352334
rect 99186 316418 99422 316654
rect 99186 316098 99422 316334
rect 99186 280418 99422 280654
rect 99186 280098 99422 280334
rect 99186 244418 99422 244654
rect 99186 244098 99422 244334
rect 99186 208418 99422 208654
rect 99186 208098 99422 208334
rect 99186 172418 99422 172654
rect 99186 172098 99422 172334
rect 99186 136418 99422 136654
rect 99186 136098 99422 136334
rect 99186 100418 99422 100654
rect 99186 100098 99422 100334
rect 99186 64418 99422 64654
rect 99186 64098 99422 64334
rect 99186 28418 99422 28654
rect 99186 28098 99422 28334
rect 99186 -5282 99422 -5046
rect 99186 -5602 99422 -5366
rect 120786 710242 121022 710478
rect 120786 709922 121022 710158
rect 117186 708362 117422 708598
rect 117186 708042 117422 708278
rect 113586 706482 113822 706718
rect 113586 706162 113822 706398
rect 102786 680018 103022 680254
rect 102786 679698 103022 679934
rect 102786 644018 103022 644254
rect 102786 643698 103022 643934
rect 102786 608018 103022 608254
rect 102786 607698 103022 607934
rect 102786 572018 103022 572254
rect 102786 571698 103022 571934
rect 102786 536018 103022 536254
rect 102786 535698 103022 535934
rect 102786 500018 103022 500254
rect 102786 499698 103022 499934
rect 102786 464018 103022 464254
rect 102786 463698 103022 463934
rect 102786 428018 103022 428254
rect 102786 427698 103022 427934
rect 102786 392018 103022 392254
rect 102786 391698 103022 391934
rect 102786 356018 103022 356254
rect 102786 355698 103022 355934
rect 102786 320018 103022 320254
rect 102786 319698 103022 319934
rect 102786 284018 103022 284254
rect 102786 283698 103022 283934
rect 102786 248018 103022 248254
rect 102786 247698 103022 247934
rect 102786 212018 103022 212254
rect 102786 211698 103022 211934
rect 102786 176018 103022 176254
rect 102786 175698 103022 175934
rect 102786 140018 103022 140254
rect 102786 139698 103022 139934
rect 102786 104018 103022 104254
rect 102786 103698 103022 103934
rect 102786 68018 103022 68254
rect 102786 67698 103022 67934
rect 102786 32018 103022 32254
rect 102786 31698 103022 31934
rect 84786 -6222 85022 -5986
rect 84786 -6542 85022 -6306
rect 109986 704602 110222 704838
rect 109986 704282 110222 704518
rect 109986 687218 110222 687454
rect 109986 686898 110222 687134
rect 109986 651218 110222 651454
rect 109986 650898 110222 651134
rect 109986 615218 110222 615454
rect 109986 614898 110222 615134
rect 109986 579218 110222 579454
rect 109986 578898 110222 579134
rect 109986 543218 110222 543454
rect 109986 542898 110222 543134
rect 109986 507218 110222 507454
rect 109986 506898 110222 507134
rect 109986 471218 110222 471454
rect 109986 470898 110222 471134
rect 109986 435218 110222 435454
rect 109986 434898 110222 435134
rect 109986 399218 110222 399454
rect 109986 398898 110222 399134
rect 109986 363218 110222 363454
rect 109986 362898 110222 363134
rect 109986 327218 110222 327454
rect 109986 326898 110222 327134
rect 109986 291218 110222 291454
rect 109986 290898 110222 291134
rect 109986 255218 110222 255454
rect 109986 254898 110222 255134
rect 109986 219218 110222 219454
rect 109986 218898 110222 219134
rect 109986 183218 110222 183454
rect 109986 182898 110222 183134
rect 109986 147218 110222 147454
rect 109986 146898 110222 147134
rect 109986 111218 110222 111454
rect 109986 110898 110222 111134
rect 109986 75218 110222 75454
rect 109986 74898 110222 75134
rect 109986 39218 110222 39454
rect 109986 38898 110222 39134
rect 109986 3218 110222 3454
rect 109986 2898 110222 3134
rect 109986 -582 110222 -346
rect 109986 -902 110222 -666
rect 113586 690818 113822 691054
rect 113586 690498 113822 690734
rect 113586 654818 113822 655054
rect 113586 654498 113822 654734
rect 113586 618818 113822 619054
rect 113586 618498 113822 618734
rect 113586 582818 113822 583054
rect 113586 582498 113822 582734
rect 113586 546818 113822 547054
rect 113586 546498 113822 546734
rect 113586 510818 113822 511054
rect 113586 510498 113822 510734
rect 113586 474818 113822 475054
rect 113586 474498 113822 474734
rect 113586 438818 113822 439054
rect 113586 438498 113822 438734
rect 113586 402818 113822 403054
rect 113586 402498 113822 402734
rect 113586 366818 113822 367054
rect 113586 366498 113822 366734
rect 113586 330818 113822 331054
rect 113586 330498 113822 330734
rect 113586 294818 113822 295054
rect 113586 294498 113822 294734
rect 113586 258818 113822 259054
rect 113586 258498 113822 258734
rect 113586 222818 113822 223054
rect 113586 222498 113822 222734
rect 113586 186818 113822 187054
rect 113586 186498 113822 186734
rect 113586 150818 113822 151054
rect 113586 150498 113822 150734
rect 113586 114818 113822 115054
rect 113586 114498 113822 114734
rect 113586 78818 113822 79054
rect 113586 78498 113822 78734
rect 113586 42818 113822 43054
rect 113586 42498 113822 42734
rect 113586 6818 113822 7054
rect 113586 6498 113822 6734
rect 113586 -2462 113822 -2226
rect 113586 -2782 113822 -2546
rect 117186 694418 117422 694654
rect 117186 694098 117422 694334
rect 117186 658418 117422 658654
rect 117186 658098 117422 658334
rect 117186 622418 117422 622654
rect 117186 622098 117422 622334
rect 117186 586418 117422 586654
rect 117186 586098 117422 586334
rect 117186 550418 117422 550654
rect 117186 550098 117422 550334
rect 117186 514418 117422 514654
rect 117186 514098 117422 514334
rect 117186 478418 117422 478654
rect 117186 478098 117422 478334
rect 117186 442418 117422 442654
rect 117186 442098 117422 442334
rect 117186 406418 117422 406654
rect 117186 406098 117422 406334
rect 117186 370418 117422 370654
rect 117186 370098 117422 370334
rect 117186 334418 117422 334654
rect 117186 334098 117422 334334
rect 117186 298418 117422 298654
rect 117186 298098 117422 298334
rect 117186 262418 117422 262654
rect 117186 262098 117422 262334
rect 117186 226418 117422 226654
rect 117186 226098 117422 226334
rect 117186 190418 117422 190654
rect 117186 190098 117422 190334
rect 117186 154418 117422 154654
rect 117186 154098 117422 154334
rect 117186 118418 117422 118654
rect 117186 118098 117422 118334
rect 117186 82418 117422 82654
rect 117186 82098 117422 82334
rect 117186 46418 117422 46654
rect 117186 46098 117422 46334
rect 117186 10418 117422 10654
rect 117186 10098 117422 10334
rect 117186 -4342 117422 -4106
rect 117186 -4662 117422 -4426
rect 138786 711182 139022 711418
rect 138786 710862 139022 711098
rect 135186 709302 135422 709538
rect 135186 708982 135422 709218
rect 131586 707422 131822 707658
rect 131586 707102 131822 707338
rect 120786 698018 121022 698254
rect 120786 697698 121022 697934
rect 120786 662018 121022 662254
rect 120786 661698 121022 661934
rect 120786 626018 121022 626254
rect 120786 625698 121022 625934
rect 120786 590018 121022 590254
rect 120786 589698 121022 589934
rect 120786 554018 121022 554254
rect 120786 553698 121022 553934
rect 120786 518018 121022 518254
rect 120786 517698 121022 517934
rect 120786 482018 121022 482254
rect 120786 481698 121022 481934
rect 120786 446018 121022 446254
rect 120786 445698 121022 445934
rect 120786 410018 121022 410254
rect 120786 409698 121022 409934
rect 120786 374018 121022 374254
rect 120786 373698 121022 373934
rect 120786 338018 121022 338254
rect 120786 337698 121022 337934
rect 120786 302018 121022 302254
rect 120786 301698 121022 301934
rect 120786 266018 121022 266254
rect 120786 265698 121022 265934
rect 120786 230018 121022 230254
rect 120786 229698 121022 229934
rect 120786 194018 121022 194254
rect 120786 193698 121022 193934
rect 120786 158018 121022 158254
rect 120786 157698 121022 157934
rect 120786 122018 121022 122254
rect 120786 121698 121022 121934
rect 120786 86018 121022 86254
rect 120786 85698 121022 85934
rect 120786 50018 121022 50254
rect 120786 49698 121022 49934
rect 120786 14018 121022 14254
rect 120786 13698 121022 13934
rect 102786 -7162 103022 -6926
rect 102786 -7482 103022 -7246
rect 127986 705542 128222 705778
rect 127986 705222 128222 705458
rect 127986 669218 128222 669454
rect 127986 668898 128222 669134
rect 127986 633218 128222 633454
rect 127986 632898 128222 633134
rect 127986 597218 128222 597454
rect 127986 596898 128222 597134
rect 127986 561218 128222 561454
rect 127986 560898 128222 561134
rect 127986 525218 128222 525454
rect 127986 524898 128222 525134
rect 127986 489218 128222 489454
rect 127986 488898 128222 489134
rect 127986 453218 128222 453454
rect 127986 452898 128222 453134
rect 127986 417218 128222 417454
rect 127986 416898 128222 417134
rect 127986 381218 128222 381454
rect 127986 380898 128222 381134
rect 127986 345218 128222 345454
rect 127986 344898 128222 345134
rect 127986 309218 128222 309454
rect 127986 308898 128222 309134
rect 127986 273218 128222 273454
rect 127986 272898 128222 273134
rect 127986 237218 128222 237454
rect 127986 236898 128222 237134
rect 127986 201218 128222 201454
rect 127986 200898 128222 201134
rect 127986 165218 128222 165454
rect 127986 164898 128222 165134
rect 127986 129218 128222 129454
rect 127986 128898 128222 129134
rect 127986 93218 128222 93454
rect 127986 92898 128222 93134
rect 127986 57218 128222 57454
rect 127986 56898 128222 57134
rect 127986 21218 128222 21454
rect 127986 20898 128222 21134
rect 127986 -1522 128222 -1286
rect 127986 -1842 128222 -1606
rect 131586 672818 131822 673054
rect 131586 672498 131822 672734
rect 131586 636818 131822 637054
rect 131586 636498 131822 636734
rect 131586 600818 131822 601054
rect 131586 600498 131822 600734
rect 131586 564818 131822 565054
rect 131586 564498 131822 564734
rect 131586 528818 131822 529054
rect 131586 528498 131822 528734
rect 131586 492818 131822 493054
rect 131586 492498 131822 492734
rect 131586 456818 131822 457054
rect 131586 456498 131822 456734
rect 131586 420818 131822 421054
rect 131586 420498 131822 420734
rect 131586 384818 131822 385054
rect 131586 384498 131822 384734
rect 131586 348818 131822 349054
rect 131586 348498 131822 348734
rect 131586 312818 131822 313054
rect 131586 312498 131822 312734
rect 131586 276818 131822 277054
rect 131586 276498 131822 276734
rect 131586 240818 131822 241054
rect 131586 240498 131822 240734
rect 131586 204818 131822 205054
rect 131586 204498 131822 204734
rect 131586 168818 131822 169054
rect 131586 168498 131822 168734
rect 131586 132818 131822 133054
rect 131586 132498 131822 132734
rect 131586 96818 131822 97054
rect 131586 96498 131822 96734
rect 131586 60818 131822 61054
rect 131586 60498 131822 60734
rect 131586 24818 131822 25054
rect 131586 24498 131822 24734
rect 131586 -3402 131822 -3166
rect 131586 -3722 131822 -3486
rect 135186 676418 135422 676654
rect 135186 676098 135422 676334
rect 135186 640418 135422 640654
rect 135186 640098 135422 640334
rect 135186 604418 135422 604654
rect 135186 604098 135422 604334
rect 135186 568418 135422 568654
rect 135186 568098 135422 568334
rect 135186 532418 135422 532654
rect 135186 532098 135422 532334
rect 135186 496418 135422 496654
rect 135186 496098 135422 496334
rect 135186 460418 135422 460654
rect 135186 460098 135422 460334
rect 135186 424418 135422 424654
rect 135186 424098 135422 424334
rect 135186 388418 135422 388654
rect 135186 388098 135422 388334
rect 135186 352418 135422 352654
rect 135186 352098 135422 352334
rect 135186 316418 135422 316654
rect 135186 316098 135422 316334
rect 135186 280418 135422 280654
rect 135186 280098 135422 280334
rect 135186 244418 135422 244654
rect 135186 244098 135422 244334
rect 135186 208418 135422 208654
rect 135186 208098 135422 208334
rect 135186 172418 135422 172654
rect 135186 172098 135422 172334
rect 135186 136418 135422 136654
rect 135186 136098 135422 136334
rect 135186 100418 135422 100654
rect 135186 100098 135422 100334
rect 135186 64418 135422 64654
rect 135186 64098 135422 64334
rect 135186 28418 135422 28654
rect 135186 28098 135422 28334
rect 135186 -5282 135422 -5046
rect 135186 -5602 135422 -5366
rect 156786 710242 157022 710478
rect 156786 709922 157022 710158
rect 153186 708362 153422 708598
rect 153186 708042 153422 708278
rect 149586 706482 149822 706718
rect 149586 706162 149822 706398
rect 138786 680018 139022 680254
rect 138786 679698 139022 679934
rect 138786 644018 139022 644254
rect 138786 643698 139022 643934
rect 138786 608018 139022 608254
rect 138786 607698 139022 607934
rect 138786 572018 139022 572254
rect 138786 571698 139022 571934
rect 138786 536018 139022 536254
rect 138786 535698 139022 535934
rect 138786 500018 139022 500254
rect 138786 499698 139022 499934
rect 138786 464018 139022 464254
rect 138786 463698 139022 463934
rect 138786 428018 139022 428254
rect 138786 427698 139022 427934
rect 138786 392018 139022 392254
rect 138786 391698 139022 391934
rect 138786 356018 139022 356254
rect 138786 355698 139022 355934
rect 138786 320018 139022 320254
rect 138786 319698 139022 319934
rect 138786 284018 139022 284254
rect 138786 283698 139022 283934
rect 138786 248018 139022 248254
rect 138786 247698 139022 247934
rect 138786 212018 139022 212254
rect 138786 211698 139022 211934
rect 138786 176018 139022 176254
rect 138786 175698 139022 175934
rect 138786 140018 139022 140254
rect 138786 139698 139022 139934
rect 138786 104018 139022 104254
rect 138786 103698 139022 103934
rect 138786 68018 139022 68254
rect 138786 67698 139022 67934
rect 138786 32018 139022 32254
rect 138786 31698 139022 31934
rect 120786 -6222 121022 -5986
rect 120786 -6542 121022 -6306
rect 145986 704602 146222 704838
rect 145986 704282 146222 704518
rect 145986 687218 146222 687454
rect 145986 686898 146222 687134
rect 145986 651218 146222 651454
rect 145986 650898 146222 651134
rect 145986 615218 146222 615454
rect 145986 614898 146222 615134
rect 145986 579218 146222 579454
rect 145986 578898 146222 579134
rect 145986 543218 146222 543454
rect 145986 542898 146222 543134
rect 145986 507218 146222 507454
rect 145986 506898 146222 507134
rect 145986 471218 146222 471454
rect 145986 470898 146222 471134
rect 145986 435218 146222 435454
rect 145986 434898 146222 435134
rect 145986 399218 146222 399454
rect 145986 398898 146222 399134
rect 145986 363218 146222 363454
rect 145986 362898 146222 363134
rect 145986 327218 146222 327454
rect 145986 326898 146222 327134
rect 145986 291218 146222 291454
rect 145986 290898 146222 291134
rect 145986 255218 146222 255454
rect 145986 254898 146222 255134
rect 145986 219218 146222 219454
rect 145986 218898 146222 219134
rect 145986 183218 146222 183454
rect 145986 182898 146222 183134
rect 145986 147218 146222 147454
rect 145986 146898 146222 147134
rect 145986 111218 146222 111454
rect 145986 110898 146222 111134
rect 145986 75218 146222 75454
rect 145986 74898 146222 75134
rect 145986 39218 146222 39454
rect 145986 38898 146222 39134
rect 145986 3218 146222 3454
rect 145986 2898 146222 3134
rect 145986 -582 146222 -346
rect 145986 -902 146222 -666
rect 149586 690818 149822 691054
rect 149586 690498 149822 690734
rect 149586 654818 149822 655054
rect 149586 654498 149822 654734
rect 149586 618818 149822 619054
rect 149586 618498 149822 618734
rect 149586 582818 149822 583054
rect 149586 582498 149822 582734
rect 149586 546818 149822 547054
rect 149586 546498 149822 546734
rect 149586 510818 149822 511054
rect 149586 510498 149822 510734
rect 149586 474818 149822 475054
rect 149586 474498 149822 474734
rect 149586 438818 149822 439054
rect 149586 438498 149822 438734
rect 149586 402818 149822 403054
rect 149586 402498 149822 402734
rect 149586 366818 149822 367054
rect 149586 366498 149822 366734
rect 149586 330818 149822 331054
rect 149586 330498 149822 330734
rect 149586 294818 149822 295054
rect 149586 294498 149822 294734
rect 149586 258818 149822 259054
rect 149586 258498 149822 258734
rect 149586 222818 149822 223054
rect 149586 222498 149822 222734
rect 149586 186818 149822 187054
rect 149586 186498 149822 186734
rect 149586 150818 149822 151054
rect 149586 150498 149822 150734
rect 149586 114818 149822 115054
rect 149586 114498 149822 114734
rect 149586 78818 149822 79054
rect 149586 78498 149822 78734
rect 149586 42818 149822 43054
rect 149586 42498 149822 42734
rect 149586 6818 149822 7054
rect 149586 6498 149822 6734
rect 149586 -2462 149822 -2226
rect 149586 -2782 149822 -2546
rect 153186 694418 153422 694654
rect 153186 694098 153422 694334
rect 153186 658418 153422 658654
rect 153186 658098 153422 658334
rect 153186 622418 153422 622654
rect 153186 622098 153422 622334
rect 153186 586418 153422 586654
rect 153186 586098 153422 586334
rect 153186 550418 153422 550654
rect 153186 550098 153422 550334
rect 153186 514418 153422 514654
rect 153186 514098 153422 514334
rect 174786 711182 175022 711418
rect 174786 710862 175022 711098
rect 171186 709302 171422 709538
rect 171186 708982 171422 709218
rect 167586 707422 167822 707658
rect 167586 707102 167822 707338
rect 156786 698018 157022 698254
rect 156786 697698 157022 697934
rect 156786 662018 157022 662254
rect 156786 661698 157022 661934
rect 156786 626018 157022 626254
rect 156786 625698 157022 625934
rect 156786 590018 157022 590254
rect 156786 589698 157022 589934
rect 156786 554018 157022 554254
rect 156786 553698 157022 553934
rect 156786 518018 157022 518254
rect 156786 517698 157022 517934
rect 163986 705542 164222 705778
rect 163986 705222 164222 705458
rect 163986 669218 164222 669454
rect 163986 668898 164222 669134
rect 163986 633218 164222 633454
rect 163986 632898 164222 633134
rect 163986 597218 164222 597454
rect 163986 596898 164222 597134
rect 163986 561218 164222 561454
rect 163986 560898 164222 561134
rect 163986 525218 164222 525454
rect 163986 524898 164222 525134
rect 167586 672818 167822 673054
rect 167586 672498 167822 672734
rect 167586 636818 167822 637054
rect 167586 636498 167822 636734
rect 167586 600818 167822 601054
rect 167586 600498 167822 600734
rect 167586 564818 167822 565054
rect 167586 564498 167822 564734
rect 167586 528818 167822 529054
rect 167586 528498 167822 528734
rect 171186 676418 171422 676654
rect 171186 676098 171422 676334
rect 171186 640418 171422 640654
rect 171186 640098 171422 640334
rect 171186 604418 171422 604654
rect 171186 604098 171422 604334
rect 171186 568418 171422 568654
rect 171186 568098 171422 568334
rect 171186 532418 171422 532654
rect 171186 532098 171422 532334
rect 192786 710242 193022 710478
rect 192786 709922 193022 710158
rect 189186 708362 189422 708598
rect 189186 708042 189422 708278
rect 185586 706482 185822 706718
rect 185586 706162 185822 706398
rect 174786 680018 175022 680254
rect 174786 679698 175022 679934
rect 174786 644018 175022 644254
rect 174786 643698 175022 643934
rect 174786 608018 175022 608254
rect 174786 607698 175022 607934
rect 174786 572018 175022 572254
rect 174786 571698 175022 571934
rect 174786 536018 175022 536254
rect 174786 535698 175022 535934
rect 181986 704602 182222 704838
rect 181986 704282 182222 704518
rect 181986 687218 182222 687454
rect 181986 686898 182222 687134
rect 181986 651218 182222 651454
rect 181986 650898 182222 651134
rect 181986 615218 182222 615454
rect 181986 614898 182222 615134
rect 181986 579218 182222 579454
rect 181986 578898 182222 579134
rect 181986 543218 182222 543454
rect 181986 542898 182222 543134
rect 185586 690818 185822 691054
rect 185586 690498 185822 690734
rect 185586 654818 185822 655054
rect 185586 654498 185822 654734
rect 185586 618818 185822 619054
rect 185586 618498 185822 618734
rect 185586 582818 185822 583054
rect 185586 582498 185822 582734
rect 185586 546818 185822 547054
rect 185586 546498 185822 546734
rect 185586 510818 185822 511054
rect 185586 510498 185822 510734
rect 189186 694418 189422 694654
rect 189186 694098 189422 694334
rect 189186 658418 189422 658654
rect 189186 658098 189422 658334
rect 189186 622418 189422 622654
rect 189186 622098 189422 622334
rect 189186 586418 189422 586654
rect 189186 586098 189422 586334
rect 189186 550418 189422 550654
rect 189186 550098 189422 550334
rect 189186 514418 189422 514654
rect 189186 514098 189422 514334
rect 210786 711182 211022 711418
rect 210786 710862 211022 711098
rect 207186 709302 207422 709538
rect 207186 708982 207422 709218
rect 203586 707422 203822 707658
rect 203586 707102 203822 707338
rect 192786 698018 193022 698254
rect 192786 697698 193022 697934
rect 192786 662018 193022 662254
rect 192786 661698 193022 661934
rect 192786 626018 193022 626254
rect 192786 625698 193022 625934
rect 192786 590018 193022 590254
rect 192786 589698 193022 589934
rect 192786 554018 193022 554254
rect 192786 553698 193022 553934
rect 192786 518018 193022 518254
rect 192786 517698 193022 517934
rect 199986 705542 200222 705778
rect 199986 705222 200222 705458
rect 199986 669218 200222 669454
rect 199986 668898 200222 669134
rect 199986 633218 200222 633454
rect 199986 632898 200222 633134
rect 199986 597218 200222 597454
rect 199986 596898 200222 597134
rect 199986 561218 200222 561454
rect 199986 560898 200222 561134
rect 199986 525218 200222 525454
rect 199986 524898 200222 525134
rect 203586 672818 203822 673054
rect 203586 672498 203822 672734
rect 203586 636818 203822 637054
rect 203586 636498 203822 636734
rect 203586 600818 203822 601054
rect 203586 600498 203822 600734
rect 203586 564818 203822 565054
rect 203586 564498 203822 564734
rect 203586 528818 203822 529054
rect 203586 528498 203822 528734
rect 207186 676418 207422 676654
rect 207186 676098 207422 676334
rect 207186 640418 207422 640654
rect 207186 640098 207422 640334
rect 207186 604418 207422 604654
rect 207186 604098 207422 604334
rect 207186 568418 207422 568654
rect 207186 568098 207422 568334
rect 207186 532418 207422 532654
rect 207186 532098 207422 532334
rect 228786 710242 229022 710478
rect 228786 709922 229022 710158
rect 225186 708362 225422 708598
rect 225186 708042 225422 708278
rect 221586 706482 221822 706718
rect 221586 706162 221822 706398
rect 210786 680018 211022 680254
rect 210786 679698 211022 679934
rect 210786 644018 211022 644254
rect 210786 643698 211022 643934
rect 210786 608018 211022 608254
rect 210786 607698 211022 607934
rect 210786 572018 211022 572254
rect 210786 571698 211022 571934
rect 210786 536018 211022 536254
rect 210786 535698 211022 535934
rect 217986 704602 218222 704838
rect 217986 704282 218222 704518
rect 217986 687218 218222 687454
rect 217986 686898 218222 687134
rect 217986 651218 218222 651454
rect 217986 650898 218222 651134
rect 217986 615218 218222 615454
rect 217986 614898 218222 615134
rect 217986 579218 218222 579454
rect 217986 578898 218222 579134
rect 217986 543218 218222 543454
rect 217986 542898 218222 543134
rect 221586 690818 221822 691054
rect 221586 690498 221822 690734
rect 221586 654818 221822 655054
rect 221586 654498 221822 654734
rect 221586 618818 221822 619054
rect 221586 618498 221822 618734
rect 221586 582818 221822 583054
rect 221586 582498 221822 582734
rect 221586 546818 221822 547054
rect 221586 546498 221822 546734
rect 221586 510818 221822 511054
rect 221586 510498 221822 510734
rect 225186 694418 225422 694654
rect 225186 694098 225422 694334
rect 225186 658418 225422 658654
rect 225186 658098 225422 658334
rect 225186 622418 225422 622654
rect 225186 622098 225422 622334
rect 225186 586418 225422 586654
rect 225186 586098 225422 586334
rect 225186 550418 225422 550654
rect 225186 550098 225422 550334
rect 225186 514418 225422 514654
rect 225186 514098 225422 514334
rect 246786 711182 247022 711418
rect 246786 710862 247022 711098
rect 243186 709302 243422 709538
rect 243186 708982 243422 709218
rect 239586 707422 239822 707658
rect 239586 707102 239822 707338
rect 228786 698018 229022 698254
rect 228786 697698 229022 697934
rect 228786 662018 229022 662254
rect 228786 661698 229022 661934
rect 228786 626018 229022 626254
rect 228786 625698 229022 625934
rect 228786 590018 229022 590254
rect 228786 589698 229022 589934
rect 228786 554018 229022 554254
rect 228786 553698 229022 553934
rect 228786 518018 229022 518254
rect 228786 517698 229022 517934
rect 235986 705542 236222 705778
rect 235986 705222 236222 705458
rect 235986 669218 236222 669454
rect 235986 668898 236222 669134
rect 235986 633218 236222 633454
rect 235986 632898 236222 633134
rect 235986 597218 236222 597454
rect 235986 596898 236222 597134
rect 235986 561218 236222 561454
rect 235986 560898 236222 561134
rect 235986 525218 236222 525454
rect 235986 524898 236222 525134
rect 239586 672818 239822 673054
rect 239586 672498 239822 672734
rect 239586 636818 239822 637054
rect 239586 636498 239822 636734
rect 239586 600818 239822 601054
rect 239586 600498 239822 600734
rect 239586 564818 239822 565054
rect 239586 564498 239822 564734
rect 239586 528818 239822 529054
rect 239586 528498 239822 528734
rect 243186 676418 243422 676654
rect 243186 676098 243422 676334
rect 243186 640418 243422 640654
rect 243186 640098 243422 640334
rect 243186 604418 243422 604654
rect 243186 604098 243422 604334
rect 243186 568418 243422 568654
rect 243186 568098 243422 568334
rect 243186 532418 243422 532654
rect 243186 532098 243422 532334
rect 264786 710242 265022 710478
rect 264786 709922 265022 710158
rect 261186 708362 261422 708598
rect 261186 708042 261422 708278
rect 257586 706482 257822 706718
rect 257586 706162 257822 706398
rect 246786 680018 247022 680254
rect 246786 679698 247022 679934
rect 246786 644018 247022 644254
rect 246786 643698 247022 643934
rect 246786 608018 247022 608254
rect 246786 607698 247022 607934
rect 246786 572018 247022 572254
rect 246786 571698 247022 571934
rect 246786 536018 247022 536254
rect 246786 535698 247022 535934
rect 253986 704602 254222 704838
rect 253986 704282 254222 704518
rect 253986 687218 254222 687454
rect 253986 686898 254222 687134
rect 253986 651218 254222 651454
rect 253986 650898 254222 651134
rect 253986 615218 254222 615454
rect 253986 614898 254222 615134
rect 253986 579218 254222 579454
rect 253986 578898 254222 579134
rect 253986 543218 254222 543454
rect 253986 542898 254222 543134
rect 257586 690818 257822 691054
rect 257586 690498 257822 690734
rect 257586 654818 257822 655054
rect 257586 654498 257822 654734
rect 257586 618818 257822 619054
rect 257586 618498 257822 618734
rect 257586 582818 257822 583054
rect 257586 582498 257822 582734
rect 257586 546818 257822 547054
rect 257586 546498 257822 546734
rect 257586 510818 257822 511054
rect 257586 510498 257822 510734
rect 261186 694418 261422 694654
rect 261186 694098 261422 694334
rect 261186 658418 261422 658654
rect 261186 658098 261422 658334
rect 261186 622418 261422 622654
rect 261186 622098 261422 622334
rect 261186 586418 261422 586654
rect 261186 586098 261422 586334
rect 261186 550418 261422 550654
rect 261186 550098 261422 550334
rect 261186 514418 261422 514654
rect 261186 514098 261422 514334
rect 282786 711182 283022 711418
rect 282786 710862 283022 711098
rect 279186 709302 279422 709538
rect 279186 708982 279422 709218
rect 275586 707422 275822 707658
rect 275586 707102 275822 707338
rect 264786 698018 265022 698254
rect 264786 697698 265022 697934
rect 264786 662018 265022 662254
rect 264786 661698 265022 661934
rect 264786 626018 265022 626254
rect 264786 625698 265022 625934
rect 264786 590018 265022 590254
rect 264786 589698 265022 589934
rect 264786 554018 265022 554254
rect 264786 553698 265022 553934
rect 264786 518018 265022 518254
rect 264786 517698 265022 517934
rect 271986 705542 272222 705778
rect 271986 705222 272222 705458
rect 271986 669218 272222 669454
rect 271986 668898 272222 669134
rect 271986 633218 272222 633454
rect 271986 632898 272222 633134
rect 271986 597218 272222 597454
rect 271986 596898 272222 597134
rect 271986 561218 272222 561454
rect 271986 560898 272222 561134
rect 271986 525218 272222 525454
rect 271986 524898 272222 525134
rect 275586 672818 275822 673054
rect 275586 672498 275822 672734
rect 275586 636818 275822 637054
rect 275586 636498 275822 636734
rect 275586 600818 275822 601054
rect 275586 600498 275822 600734
rect 275586 564818 275822 565054
rect 275586 564498 275822 564734
rect 275586 528818 275822 529054
rect 275586 528498 275822 528734
rect 279186 676418 279422 676654
rect 279186 676098 279422 676334
rect 279186 640418 279422 640654
rect 279186 640098 279422 640334
rect 279186 604418 279422 604654
rect 279186 604098 279422 604334
rect 279186 568418 279422 568654
rect 279186 568098 279422 568334
rect 279186 532418 279422 532654
rect 279186 532098 279422 532334
rect 300786 710242 301022 710478
rect 300786 709922 301022 710158
rect 297186 708362 297422 708598
rect 297186 708042 297422 708278
rect 293586 706482 293822 706718
rect 293586 706162 293822 706398
rect 282786 680018 283022 680254
rect 282786 679698 283022 679934
rect 282786 644018 283022 644254
rect 282786 643698 283022 643934
rect 282786 608018 283022 608254
rect 282786 607698 283022 607934
rect 282786 572018 283022 572254
rect 282786 571698 283022 571934
rect 282786 536018 283022 536254
rect 282786 535698 283022 535934
rect 289986 704602 290222 704838
rect 289986 704282 290222 704518
rect 289986 687218 290222 687454
rect 289986 686898 290222 687134
rect 289986 651218 290222 651454
rect 289986 650898 290222 651134
rect 289986 615218 290222 615454
rect 289986 614898 290222 615134
rect 289986 579218 290222 579454
rect 289986 578898 290222 579134
rect 289986 543218 290222 543454
rect 289986 542898 290222 543134
rect 293586 690818 293822 691054
rect 293586 690498 293822 690734
rect 293586 654818 293822 655054
rect 293586 654498 293822 654734
rect 293586 618818 293822 619054
rect 293586 618498 293822 618734
rect 293586 582818 293822 583054
rect 293586 582498 293822 582734
rect 293586 546818 293822 547054
rect 293586 546498 293822 546734
rect 293586 510818 293822 511054
rect 293586 510498 293822 510734
rect 297186 694418 297422 694654
rect 297186 694098 297422 694334
rect 297186 658418 297422 658654
rect 297186 658098 297422 658334
rect 297186 622418 297422 622654
rect 297186 622098 297422 622334
rect 297186 586418 297422 586654
rect 297186 586098 297422 586334
rect 297186 550418 297422 550654
rect 297186 550098 297422 550334
rect 297186 514418 297422 514654
rect 297186 514098 297422 514334
rect 318786 711182 319022 711418
rect 318786 710862 319022 711098
rect 315186 709302 315422 709538
rect 315186 708982 315422 709218
rect 311586 707422 311822 707658
rect 311586 707102 311822 707338
rect 300786 698018 301022 698254
rect 300786 697698 301022 697934
rect 300786 662018 301022 662254
rect 300786 661698 301022 661934
rect 300786 626018 301022 626254
rect 300786 625698 301022 625934
rect 300786 590018 301022 590254
rect 300786 589698 301022 589934
rect 300786 554018 301022 554254
rect 300786 553698 301022 553934
rect 300786 518018 301022 518254
rect 300786 517698 301022 517934
rect 307986 705542 308222 705778
rect 307986 705222 308222 705458
rect 307986 669218 308222 669454
rect 307986 668898 308222 669134
rect 307986 633218 308222 633454
rect 307986 632898 308222 633134
rect 307986 597218 308222 597454
rect 307986 596898 308222 597134
rect 307986 561218 308222 561454
rect 307986 560898 308222 561134
rect 307986 525218 308222 525454
rect 307986 524898 308222 525134
rect 311586 672818 311822 673054
rect 311586 672498 311822 672734
rect 311586 636818 311822 637054
rect 311586 636498 311822 636734
rect 311586 600818 311822 601054
rect 311586 600498 311822 600734
rect 311586 564818 311822 565054
rect 311586 564498 311822 564734
rect 311586 528818 311822 529054
rect 311586 528498 311822 528734
rect 315186 676418 315422 676654
rect 315186 676098 315422 676334
rect 315186 640418 315422 640654
rect 315186 640098 315422 640334
rect 315186 604418 315422 604654
rect 315186 604098 315422 604334
rect 315186 568418 315422 568654
rect 315186 568098 315422 568334
rect 315186 532418 315422 532654
rect 315186 532098 315422 532334
rect 336786 710242 337022 710478
rect 336786 709922 337022 710158
rect 333186 708362 333422 708598
rect 333186 708042 333422 708278
rect 329586 706482 329822 706718
rect 329586 706162 329822 706398
rect 318786 680018 319022 680254
rect 318786 679698 319022 679934
rect 318786 644018 319022 644254
rect 318786 643698 319022 643934
rect 318786 608018 319022 608254
rect 318786 607698 319022 607934
rect 318786 572018 319022 572254
rect 318786 571698 319022 571934
rect 318786 536018 319022 536254
rect 318786 535698 319022 535934
rect 325986 704602 326222 704838
rect 325986 704282 326222 704518
rect 325986 687218 326222 687454
rect 325986 686898 326222 687134
rect 325986 651218 326222 651454
rect 325986 650898 326222 651134
rect 325986 615218 326222 615454
rect 325986 614898 326222 615134
rect 325986 579218 326222 579454
rect 325986 578898 326222 579134
rect 325986 543218 326222 543454
rect 325986 542898 326222 543134
rect 329586 690818 329822 691054
rect 329586 690498 329822 690734
rect 329586 654818 329822 655054
rect 329586 654498 329822 654734
rect 329586 618818 329822 619054
rect 329586 618498 329822 618734
rect 329586 582818 329822 583054
rect 329586 582498 329822 582734
rect 329586 546818 329822 547054
rect 329586 546498 329822 546734
rect 329586 510818 329822 511054
rect 329586 510498 329822 510734
rect 333186 694418 333422 694654
rect 333186 694098 333422 694334
rect 333186 658418 333422 658654
rect 333186 658098 333422 658334
rect 333186 622418 333422 622654
rect 333186 622098 333422 622334
rect 333186 586418 333422 586654
rect 333186 586098 333422 586334
rect 333186 550418 333422 550654
rect 333186 550098 333422 550334
rect 333186 514418 333422 514654
rect 333186 514098 333422 514334
rect 354786 711182 355022 711418
rect 354786 710862 355022 711098
rect 351186 709302 351422 709538
rect 351186 708982 351422 709218
rect 347586 707422 347822 707658
rect 347586 707102 347822 707338
rect 336786 698018 337022 698254
rect 336786 697698 337022 697934
rect 336786 662018 337022 662254
rect 336786 661698 337022 661934
rect 336786 626018 337022 626254
rect 336786 625698 337022 625934
rect 336786 590018 337022 590254
rect 336786 589698 337022 589934
rect 336786 554018 337022 554254
rect 336786 553698 337022 553934
rect 336786 518018 337022 518254
rect 336786 517698 337022 517934
rect 343986 705542 344222 705778
rect 343986 705222 344222 705458
rect 343986 669218 344222 669454
rect 343986 668898 344222 669134
rect 343986 633218 344222 633454
rect 343986 632898 344222 633134
rect 343986 597218 344222 597454
rect 343986 596898 344222 597134
rect 343986 561218 344222 561454
rect 343986 560898 344222 561134
rect 343986 525218 344222 525454
rect 343986 524898 344222 525134
rect 347586 672818 347822 673054
rect 347586 672498 347822 672734
rect 347586 636818 347822 637054
rect 347586 636498 347822 636734
rect 347586 600818 347822 601054
rect 347586 600498 347822 600734
rect 347586 564818 347822 565054
rect 347586 564498 347822 564734
rect 347586 528818 347822 529054
rect 347586 528498 347822 528734
rect 351186 676418 351422 676654
rect 351186 676098 351422 676334
rect 351186 640418 351422 640654
rect 351186 640098 351422 640334
rect 351186 604418 351422 604654
rect 351186 604098 351422 604334
rect 351186 568418 351422 568654
rect 351186 568098 351422 568334
rect 351186 532418 351422 532654
rect 351186 532098 351422 532334
rect 372786 710242 373022 710478
rect 372786 709922 373022 710158
rect 369186 708362 369422 708598
rect 369186 708042 369422 708278
rect 365586 706482 365822 706718
rect 365586 706162 365822 706398
rect 354786 680018 355022 680254
rect 354786 679698 355022 679934
rect 354786 644018 355022 644254
rect 354786 643698 355022 643934
rect 354786 608018 355022 608254
rect 354786 607698 355022 607934
rect 354786 572018 355022 572254
rect 354786 571698 355022 571934
rect 354786 536018 355022 536254
rect 354786 535698 355022 535934
rect 361986 704602 362222 704838
rect 361986 704282 362222 704518
rect 361986 687218 362222 687454
rect 361986 686898 362222 687134
rect 361986 651218 362222 651454
rect 361986 650898 362222 651134
rect 361986 615218 362222 615454
rect 361986 614898 362222 615134
rect 361986 579218 362222 579454
rect 361986 578898 362222 579134
rect 361986 543218 362222 543454
rect 361986 542898 362222 543134
rect 365586 690818 365822 691054
rect 365586 690498 365822 690734
rect 365586 654818 365822 655054
rect 365586 654498 365822 654734
rect 365586 618818 365822 619054
rect 365586 618498 365822 618734
rect 365586 582818 365822 583054
rect 365586 582498 365822 582734
rect 365586 546818 365822 547054
rect 365586 546498 365822 546734
rect 365586 510818 365822 511054
rect 365586 510498 365822 510734
rect 369186 694418 369422 694654
rect 369186 694098 369422 694334
rect 369186 658418 369422 658654
rect 369186 658098 369422 658334
rect 369186 622418 369422 622654
rect 369186 622098 369422 622334
rect 369186 586418 369422 586654
rect 369186 586098 369422 586334
rect 369186 550418 369422 550654
rect 369186 550098 369422 550334
rect 369186 514418 369422 514654
rect 369186 514098 369422 514334
rect 390786 711182 391022 711418
rect 390786 710862 391022 711098
rect 387186 709302 387422 709538
rect 387186 708982 387422 709218
rect 383586 707422 383822 707658
rect 383586 707102 383822 707338
rect 372786 698018 373022 698254
rect 372786 697698 373022 697934
rect 372786 662018 373022 662254
rect 372786 661698 373022 661934
rect 372786 626018 373022 626254
rect 372786 625698 373022 625934
rect 372786 590018 373022 590254
rect 372786 589698 373022 589934
rect 372786 554018 373022 554254
rect 372786 553698 373022 553934
rect 372786 518018 373022 518254
rect 372786 517698 373022 517934
rect 379986 705542 380222 705778
rect 379986 705222 380222 705458
rect 379986 669218 380222 669454
rect 379986 668898 380222 669134
rect 379986 633218 380222 633454
rect 379986 632898 380222 633134
rect 379986 597218 380222 597454
rect 379986 596898 380222 597134
rect 379986 561218 380222 561454
rect 379986 560898 380222 561134
rect 379986 525218 380222 525454
rect 379986 524898 380222 525134
rect 383586 672818 383822 673054
rect 383586 672498 383822 672734
rect 383586 636818 383822 637054
rect 383586 636498 383822 636734
rect 383586 600818 383822 601054
rect 383586 600498 383822 600734
rect 383586 564818 383822 565054
rect 383586 564498 383822 564734
rect 383586 528818 383822 529054
rect 383586 528498 383822 528734
rect 387186 676418 387422 676654
rect 387186 676098 387422 676334
rect 387186 640418 387422 640654
rect 387186 640098 387422 640334
rect 387186 604418 387422 604654
rect 387186 604098 387422 604334
rect 387186 568418 387422 568654
rect 387186 568098 387422 568334
rect 387186 532418 387422 532654
rect 387186 532098 387422 532334
rect 408786 710242 409022 710478
rect 408786 709922 409022 710158
rect 405186 708362 405422 708598
rect 405186 708042 405422 708278
rect 401586 706482 401822 706718
rect 401586 706162 401822 706398
rect 390786 680018 391022 680254
rect 390786 679698 391022 679934
rect 390786 644018 391022 644254
rect 390786 643698 391022 643934
rect 390786 608018 391022 608254
rect 390786 607698 391022 607934
rect 390786 572018 391022 572254
rect 390786 571698 391022 571934
rect 390786 536018 391022 536254
rect 390786 535698 391022 535934
rect 397986 704602 398222 704838
rect 397986 704282 398222 704518
rect 397986 687218 398222 687454
rect 397986 686898 398222 687134
rect 397986 651218 398222 651454
rect 397986 650898 398222 651134
rect 397986 615218 398222 615454
rect 397986 614898 398222 615134
rect 397986 579218 398222 579454
rect 397986 578898 398222 579134
rect 397986 543218 398222 543454
rect 397986 542898 398222 543134
rect 401586 690818 401822 691054
rect 401586 690498 401822 690734
rect 401586 654818 401822 655054
rect 401586 654498 401822 654734
rect 401586 618818 401822 619054
rect 401586 618498 401822 618734
rect 401586 582818 401822 583054
rect 401586 582498 401822 582734
rect 401586 546818 401822 547054
rect 401586 546498 401822 546734
rect 401586 510818 401822 511054
rect 401586 510498 401822 510734
rect 405186 694418 405422 694654
rect 405186 694098 405422 694334
rect 405186 658418 405422 658654
rect 405186 658098 405422 658334
rect 405186 622418 405422 622654
rect 405186 622098 405422 622334
rect 405186 586418 405422 586654
rect 405186 586098 405422 586334
rect 405186 550418 405422 550654
rect 405186 550098 405422 550334
rect 405186 514418 405422 514654
rect 405186 514098 405422 514334
rect 426786 711182 427022 711418
rect 426786 710862 427022 711098
rect 423186 709302 423422 709538
rect 423186 708982 423422 709218
rect 419586 707422 419822 707658
rect 419586 707102 419822 707338
rect 408786 698018 409022 698254
rect 408786 697698 409022 697934
rect 408786 662018 409022 662254
rect 408786 661698 409022 661934
rect 408786 626018 409022 626254
rect 408786 625698 409022 625934
rect 408786 590018 409022 590254
rect 408786 589698 409022 589934
rect 408786 554018 409022 554254
rect 408786 553698 409022 553934
rect 408786 518018 409022 518254
rect 408786 517698 409022 517934
rect 415986 705542 416222 705778
rect 415986 705222 416222 705458
rect 415986 669218 416222 669454
rect 415986 668898 416222 669134
rect 415986 633218 416222 633454
rect 415986 632898 416222 633134
rect 415986 597218 416222 597454
rect 415986 596898 416222 597134
rect 415986 561218 416222 561454
rect 415986 560898 416222 561134
rect 415986 525218 416222 525454
rect 415986 524898 416222 525134
rect 419586 672818 419822 673054
rect 419586 672498 419822 672734
rect 419586 636818 419822 637054
rect 419586 636498 419822 636734
rect 419586 600818 419822 601054
rect 419586 600498 419822 600734
rect 419586 564818 419822 565054
rect 419586 564498 419822 564734
rect 419586 528818 419822 529054
rect 419586 528498 419822 528734
rect 423186 676418 423422 676654
rect 423186 676098 423422 676334
rect 423186 640418 423422 640654
rect 423186 640098 423422 640334
rect 423186 604418 423422 604654
rect 423186 604098 423422 604334
rect 423186 568418 423422 568654
rect 423186 568098 423422 568334
rect 423186 532418 423422 532654
rect 423186 532098 423422 532334
rect 444786 710242 445022 710478
rect 444786 709922 445022 710158
rect 441186 708362 441422 708598
rect 441186 708042 441422 708278
rect 437586 706482 437822 706718
rect 437586 706162 437822 706398
rect 426786 680018 427022 680254
rect 426786 679698 427022 679934
rect 426786 644018 427022 644254
rect 426786 643698 427022 643934
rect 426786 608018 427022 608254
rect 426786 607698 427022 607934
rect 426786 572018 427022 572254
rect 426786 571698 427022 571934
rect 426786 536018 427022 536254
rect 426786 535698 427022 535934
rect 433986 704602 434222 704838
rect 433986 704282 434222 704518
rect 433986 687218 434222 687454
rect 433986 686898 434222 687134
rect 433986 651218 434222 651454
rect 433986 650898 434222 651134
rect 433986 615218 434222 615454
rect 433986 614898 434222 615134
rect 433986 579218 434222 579454
rect 433986 578898 434222 579134
rect 433986 543218 434222 543454
rect 433986 542898 434222 543134
rect 437586 690818 437822 691054
rect 437586 690498 437822 690734
rect 437586 654818 437822 655054
rect 437586 654498 437822 654734
rect 437586 618818 437822 619054
rect 437586 618498 437822 618734
rect 437586 582818 437822 583054
rect 437586 582498 437822 582734
rect 437586 546818 437822 547054
rect 437586 546498 437822 546734
rect 437586 510818 437822 511054
rect 437586 510498 437822 510734
rect 441186 694418 441422 694654
rect 441186 694098 441422 694334
rect 441186 658418 441422 658654
rect 441186 658098 441422 658334
rect 441186 622418 441422 622654
rect 441186 622098 441422 622334
rect 441186 586418 441422 586654
rect 441186 586098 441422 586334
rect 441186 550418 441422 550654
rect 441186 550098 441422 550334
rect 441186 514418 441422 514654
rect 441186 514098 441422 514334
rect 153186 478418 153422 478654
rect 153186 478098 153422 478334
rect 153186 442418 153422 442654
rect 153186 442098 153422 442334
rect 153186 406418 153422 406654
rect 153186 406098 153422 406334
rect 153186 370418 153422 370654
rect 153186 370098 153422 370334
rect 441186 478418 441422 478654
rect 441186 478098 441422 478334
rect 441186 442418 441422 442654
rect 441186 442098 441422 442334
rect 441186 406418 441422 406654
rect 441186 406098 441422 406334
rect 441186 370418 441422 370654
rect 441186 370098 441422 370334
rect 153186 334418 153422 334654
rect 153186 334098 153422 334334
rect 153186 298418 153422 298654
rect 153186 298098 153422 298334
rect 153186 262418 153422 262654
rect 153186 262098 153422 262334
rect 153186 226418 153422 226654
rect 153186 226098 153422 226334
rect 153186 190418 153422 190654
rect 153186 190098 153422 190334
rect 153186 154418 153422 154654
rect 153186 154098 153422 154334
rect 153186 118418 153422 118654
rect 153186 118098 153422 118334
rect 153186 82418 153422 82654
rect 153186 82098 153422 82334
rect 153186 46418 153422 46654
rect 153186 46098 153422 46334
rect 153186 10418 153422 10654
rect 153186 10098 153422 10334
rect 153186 -4342 153422 -4106
rect 153186 -4662 153422 -4426
rect 156786 302018 157022 302254
rect 156786 301698 157022 301934
rect 156786 266018 157022 266254
rect 156786 265698 157022 265934
rect 156786 230018 157022 230254
rect 156786 229698 157022 229934
rect 156786 194018 157022 194254
rect 156786 193698 157022 193934
rect 156786 158018 157022 158254
rect 156786 157698 157022 157934
rect 156786 122018 157022 122254
rect 156786 121698 157022 121934
rect 156786 86018 157022 86254
rect 156786 85698 157022 85934
rect 156786 50018 157022 50254
rect 156786 49698 157022 49934
rect 156786 14018 157022 14254
rect 156786 13698 157022 13934
rect 138786 -7162 139022 -6926
rect 138786 -7482 139022 -7246
rect 163986 309218 164222 309454
rect 163986 308898 164222 309134
rect 163986 273218 164222 273454
rect 163986 272898 164222 273134
rect 163986 237218 164222 237454
rect 163986 236898 164222 237134
rect 163986 201218 164222 201454
rect 163986 200898 164222 201134
rect 163986 165218 164222 165454
rect 163986 164898 164222 165134
rect 163986 129218 164222 129454
rect 163986 128898 164222 129134
rect 163986 93218 164222 93454
rect 163986 92898 164222 93134
rect 163986 57218 164222 57454
rect 163986 56898 164222 57134
rect 163986 21218 164222 21454
rect 163986 20898 164222 21134
rect 163986 -1522 164222 -1286
rect 163986 -1842 164222 -1606
rect 167586 312818 167822 313054
rect 167586 312498 167822 312734
rect 167586 276818 167822 277054
rect 167586 276498 167822 276734
rect 167586 240818 167822 241054
rect 167586 240498 167822 240734
rect 167586 204818 167822 205054
rect 167586 204498 167822 204734
rect 167586 168818 167822 169054
rect 167586 168498 167822 168734
rect 167586 132818 167822 133054
rect 167586 132498 167822 132734
rect 167586 96818 167822 97054
rect 167586 96498 167822 96734
rect 167586 60818 167822 61054
rect 167586 60498 167822 60734
rect 167586 24818 167822 25054
rect 167586 24498 167822 24734
rect 167586 -3402 167822 -3166
rect 167586 -3722 167822 -3486
rect 171186 316418 171422 316654
rect 171186 316098 171422 316334
rect 171186 280418 171422 280654
rect 171186 280098 171422 280334
rect 171186 244418 171422 244654
rect 171186 244098 171422 244334
rect 171186 208418 171422 208654
rect 171186 208098 171422 208334
rect 171186 172418 171422 172654
rect 171186 172098 171422 172334
rect 171186 136418 171422 136654
rect 171186 136098 171422 136334
rect 171186 100418 171422 100654
rect 171186 100098 171422 100334
rect 171186 64418 171422 64654
rect 171186 64098 171422 64334
rect 171186 28418 171422 28654
rect 171186 28098 171422 28334
rect 171186 -5282 171422 -5046
rect 171186 -5602 171422 -5366
rect 174786 320018 175022 320254
rect 174786 319698 175022 319934
rect 174786 284018 175022 284254
rect 174786 283698 175022 283934
rect 174786 248018 175022 248254
rect 174786 247698 175022 247934
rect 174786 212018 175022 212254
rect 174786 211698 175022 211934
rect 174786 176018 175022 176254
rect 174786 175698 175022 175934
rect 174786 140018 175022 140254
rect 174786 139698 175022 139934
rect 174786 104018 175022 104254
rect 174786 103698 175022 103934
rect 174786 68018 175022 68254
rect 174786 67698 175022 67934
rect 174786 32018 175022 32254
rect 174786 31698 175022 31934
rect 156786 -6222 157022 -5986
rect 156786 -6542 157022 -6306
rect 181986 291218 182222 291454
rect 181986 290898 182222 291134
rect 181986 255218 182222 255454
rect 181986 254898 182222 255134
rect 181986 219218 182222 219454
rect 181986 218898 182222 219134
rect 181986 183218 182222 183454
rect 181986 182898 182222 183134
rect 181986 147218 182222 147454
rect 181986 146898 182222 147134
rect 181986 111218 182222 111454
rect 181986 110898 182222 111134
rect 181986 75218 182222 75454
rect 181986 74898 182222 75134
rect 181986 39218 182222 39454
rect 181986 38898 182222 39134
rect 181986 3218 182222 3454
rect 181986 2898 182222 3134
rect 181986 -582 182222 -346
rect 181986 -902 182222 -666
rect 185586 294818 185822 295054
rect 185586 294498 185822 294734
rect 185586 258818 185822 259054
rect 185586 258498 185822 258734
rect 185586 222818 185822 223054
rect 185586 222498 185822 222734
rect 185586 186818 185822 187054
rect 185586 186498 185822 186734
rect 185586 150818 185822 151054
rect 185586 150498 185822 150734
rect 185586 114818 185822 115054
rect 185586 114498 185822 114734
rect 185586 78818 185822 79054
rect 185586 78498 185822 78734
rect 185586 42818 185822 43054
rect 185586 42498 185822 42734
rect 185586 6818 185822 7054
rect 185586 6498 185822 6734
rect 185586 -2462 185822 -2226
rect 185586 -2782 185822 -2546
rect 189186 298418 189422 298654
rect 189186 298098 189422 298334
rect 189186 262418 189422 262654
rect 189186 262098 189422 262334
rect 189186 226418 189422 226654
rect 189186 226098 189422 226334
rect 189186 190418 189422 190654
rect 189186 190098 189422 190334
rect 189186 154418 189422 154654
rect 189186 154098 189422 154334
rect 189186 118418 189422 118654
rect 189186 118098 189422 118334
rect 189186 82418 189422 82654
rect 189186 82098 189422 82334
rect 189186 46418 189422 46654
rect 189186 46098 189422 46334
rect 189186 10418 189422 10654
rect 189186 10098 189422 10334
rect 189186 -4342 189422 -4106
rect 189186 -4662 189422 -4426
rect 192786 302018 193022 302254
rect 192786 301698 193022 301934
rect 192786 266018 193022 266254
rect 192786 265698 193022 265934
rect 192786 230018 193022 230254
rect 192786 229698 193022 229934
rect 192786 194018 193022 194254
rect 192786 193698 193022 193934
rect 192786 158018 193022 158254
rect 192786 157698 193022 157934
rect 192786 122018 193022 122254
rect 192786 121698 193022 121934
rect 192786 86018 193022 86254
rect 192786 85698 193022 85934
rect 192786 50018 193022 50254
rect 192786 49698 193022 49934
rect 192786 14018 193022 14254
rect 192786 13698 193022 13934
rect 174786 -7162 175022 -6926
rect 174786 -7482 175022 -7246
rect 199986 309218 200222 309454
rect 199986 308898 200222 309134
rect 199986 273218 200222 273454
rect 199986 272898 200222 273134
rect 199986 237218 200222 237454
rect 199986 236898 200222 237134
rect 199986 201218 200222 201454
rect 199986 200898 200222 201134
rect 199986 165218 200222 165454
rect 199986 164898 200222 165134
rect 199986 129218 200222 129454
rect 199986 128898 200222 129134
rect 199986 93218 200222 93454
rect 199986 92898 200222 93134
rect 199986 57218 200222 57454
rect 199986 56898 200222 57134
rect 199986 21218 200222 21454
rect 199986 20898 200222 21134
rect 199986 -1522 200222 -1286
rect 199986 -1842 200222 -1606
rect 203586 312818 203822 313054
rect 203586 312498 203822 312734
rect 203586 276818 203822 277054
rect 203586 276498 203822 276734
rect 203586 240818 203822 241054
rect 203586 240498 203822 240734
rect 203586 204818 203822 205054
rect 203586 204498 203822 204734
rect 203586 168818 203822 169054
rect 203586 168498 203822 168734
rect 203586 132818 203822 133054
rect 203586 132498 203822 132734
rect 203586 96818 203822 97054
rect 203586 96498 203822 96734
rect 203586 60818 203822 61054
rect 203586 60498 203822 60734
rect 203586 24818 203822 25054
rect 203586 24498 203822 24734
rect 203586 -3402 203822 -3166
rect 203586 -3722 203822 -3486
rect 207186 316418 207422 316654
rect 207186 316098 207422 316334
rect 207186 280418 207422 280654
rect 207186 280098 207422 280334
rect 207186 244418 207422 244654
rect 207186 244098 207422 244334
rect 207186 208418 207422 208654
rect 207186 208098 207422 208334
rect 207186 172418 207422 172654
rect 207186 172098 207422 172334
rect 207186 136418 207422 136654
rect 207186 136098 207422 136334
rect 207186 100418 207422 100654
rect 207186 100098 207422 100334
rect 207186 64418 207422 64654
rect 207186 64098 207422 64334
rect 207186 28418 207422 28654
rect 207186 28098 207422 28334
rect 207186 -5282 207422 -5046
rect 207186 -5602 207422 -5366
rect 210786 320018 211022 320254
rect 210786 319698 211022 319934
rect 210786 284018 211022 284254
rect 210786 283698 211022 283934
rect 210786 248018 211022 248254
rect 210786 247698 211022 247934
rect 210786 212018 211022 212254
rect 210786 211698 211022 211934
rect 210786 176018 211022 176254
rect 210786 175698 211022 175934
rect 210786 140018 211022 140254
rect 210786 139698 211022 139934
rect 210786 104018 211022 104254
rect 210786 103698 211022 103934
rect 210786 68018 211022 68254
rect 210786 67698 211022 67934
rect 210786 32018 211022 32254
rect 210786 31698 211022 31934
rect 192786 -6222 193022 -5986
rect 192786 -6542 193022 -6306
rect 217986 291218 218222 291454
rect 217986 290898 218222 291134
rect 217986 255218 218222 255454
rect 217986 254898 218222 255134
rect 217986 219218 218222 219454
rect 217986 218898 218222 219134
rect 217986 183218 218222 183454
rect 217986 182898 218222 183134
rect 217986 147218 218222 147454
rect 217986 146898 218222 147134
rect 217986 111218 218222 111454
rect 217986 110898 218222 111134
rect 217986 75218 218222 75454
rect 217986 74898 218222 75134
rect 217986 39218 218222 39454
rect 217986 38898 218222 39134
rect 217986 3218 218222 3454
rect 217986 2898 218222 3134
rect 217986 -582 218222 -346
rect 217986 -902 218222 -666
rect 221586 294818 221822 295054
rect 221586 294498 221822 294734
rect 221586 258818 221822 259054
rect 221586 258498 221822 258734
rect 221586 222818 221822 223054
rect 221586 222498 221822 222734
rect 221586 186818 221822 187054
rect 221586 186498 221822 186734
rect 221586 150818 221822 151054
rect 221586 150498 221822 150734
rect 221586 114818 221822 115054
rect 221586 114498 221822 114734
rect 221586 78818 221822 79054
rect 221586 78498 221822 78734
rect 221586 42818 221822 43054
rect 221586 42498 221822 42734
rect 221586 6818 221822 7054
rect 221586 6498 221822 6734
rect 221586 -2462 221822 -2226
rect 221586 -2782 221822 -2546
rect 225186 298418 225422 298654
rect 225186 298098 225422 298334
rect 225186 262418 225422 262654
rect 225186 262098 225422 262334
rect 225186 226418 225422 226654
rect 225186 226098 225422 226334
rect 225186 190418 225422 190654
rect 225186 190098 225422 190334
rect 225186 154418 225422 154654
rect 225186 154098 225422 154334
rect 225186 118418 225422 118654
rect 225186 118098 225422 118334
rect 225186 82418 225422 82654
rect 225186 82098 225422 82334
rect 225186 46418 225422 46654
rect 225186 46098 225422 46334
rect 225186 10418 225422 10654
rect 225186 10098 225422 10334
rect 225186 -4342 225422 -4106
rect 225186 -4662 225422 -4426
rect 228786 302018 229022 302254
rect 228786 301698 229022 301934
rect 228786 266018 229022 266254
rect 228786 265698 229022 265934
rect 228786 230018 229022 230254
rect 228786 229698 229022 229934
rect 228786 194018 229022 194254
rect 228786 193698 229022 193934
rect 228786 158018 229022 158254
rect 228786 157698 229022 157934
rect 228786 122018 229022 122254
rect 228786 121698 229022 121934
rect 228786 86018 229022 86254
rect 228786 85698 229022 85934
rect 228786 50018 229022 50254
rect 228786 49698 229022 49934
rect 228786 14018 229022 14254
rect 228786 13698 229022 13934
rect 210786 -7162 211022 -6926
rect 210786 -7482 211022 -7246
rect 235986 309218 236222 309454
rect 235986 308898 236222 309134
rect 235986 273218 236222 273454
rect 235986 272898 236222 273134
rect 235986 237218 236222 237454
rect 235986 236898 236222 237134
rect 235986 201218 236222 201454
rect 235986 200898 236222 201134
rect 235986 165218 236222 165454
rect 235986 164898 236222 165134
rect 235986 129218 236222 129454
rect 235986 128898 236222 129134
rect 235986 93218 236222 93454
rect 235986 92898 236222 93134
rect 235986 57218 236222 57454
rect 235986 56898 236222 57134
rect 235986 21218 236222 21454
rect 235986 20898 236222 21134
rect 235986 -1522 236222 -1286
rect 235986 -1842 236222 -1606
rect 239586 312818 239822 313054
rect 239586 312498 239822 312734
rect 239586 276818 239822 277054
rect 239586 276498 239822 276734
rect 239586 240818 239822 241054
rect 239586 240498 239822 240734
rect 239586 204818 239822 205054
rect 239586 204498 239822 204734
rect 239586 168818 239822 169054
rect 239586 168498 239822 168734
rect 239586 132818 239822 133054
rect 239586 132498 239822 132734
rect 239586 96818 239822 97054
rect 239586 96498 239822 96734
rect 239586 60818 239822 61054
rect 239586 60498 239822 60734
rect 239586 24818 239822 25054
rect 239586 24498 239822 24734
rect 239586 -3402 239822 -3166
rect 239586 -3722 239822 -3486
rect 243186 316418 243422 316654
rect 243186 316098 243422 316334
rect 243186 280418 243422 280654
rect 243186 280098 243422 280334
rect 243186 244418 243422 244654
rect 243186 244098 243422 244334
rect 243186 208418 243422 208654
rect 243186 208098 243422 208334
rect 243186 172418 243422 172654
rect 243186 172098 243422 172334
rect 243186 136418 243422 136654
rect 243186 136098 243422 136334
rect 243186 100418 243422 100654
rect 243186 100098 243422 100334
rect 243186 64418 243422 64654
rect 243186 64098 243422 64334
rect 243186 28418 243422 28654
rect 243186 28098 243422 28334
rect 243186 -5282 243422 -5046
rect 243186 -5602 243422 -5366
rect 246786 320018 247022 320254
rect 246786 319698 247022 319934
rect 246786 284018 247022 284254
rect 246786 283698 247022 283934
rect 246786 248018 247022 248254
rect 246786 247698 247022 247934
rect 246786 212018 247022 212254
rect 246786 211698 247022 211934
rect 246786 176018 247022 176254
rect 246786 175698 247022 175934
rect 246786 140018 247022 140254
rect 246786 139698 247022 139934
rect 246786 104018 247022 104254
rect 246786 103698 247022 103934
rect 246786 68018 247022 68254
rect 246786 67698 247022 67934
rect 246786 32018 247022 32254
rect 246786 31698 247022 31934
rect 228786 -6222 229022 -5986
rect 228786 -6542 229022 -6306
rect 253986 291218 254222 291454
rect 253986 290898 254222 291134
rect 253986 255218 254222 255454
rect 253986 254898 254222 255134
rect 253986 219218 254222 219454
rect 253986 218898 254222 219134
rect 253986 183218 254222 183454
rect 253986 182898 254222 183134
rect 253986 147218 254222 147454
rect 253986 146898 254222 147134
rect 253986 111218 254222 111454
rect 253986 110898 254222 111134
rect 253986 75218 254222 75454
rect 253986 74898 254222 75134
rect 253986 39218 254222 39454
rect 253986 38898 254222 39134
rect 253986 3218 254222 3454
rect 253986 2898 254222 3134
rect 253986 -582 254222 -346
rect 253986 -902 254222 -666
rect 257586 294818 257822 295054
rect 257586 294498 257822 294734
rect 257586 258818 257822 259054
rect 257586 258498 257822 258734
rect 257586 222818 257822 223054
rect 257586 222498 257822 222734
rect 257586 186818 257822 187054
rect 257586 186498 257822 186734
rect 257586 150818 257822 151054
rect 257586 150498 257822 150734
rect 257586 114818 257822 115054
rect 257586 114498 257822 114734
rect 257586 78818 257822 79054
rect 257586 78498 257822 78734
rect 257586 42818 257822 43054
rect 257586 42498 257822 42734
rect 257586 6818 257822 7054
rect 257586 6498 257822 6734
rect 257586 -2462 257822 -2226
rect 257586 -2782 257822 -2546
rect 261186 298418 261422 298654
rect 261186 298098 261422 298334
rect 261186 262418 261422 262654
rect 261186 262098 261422 262334
rect 261186 226418 261422 226654
rect 261186 226098 261422 226334
rect 261186 190418 261422 190654
rect 261186 190098 261422 190334
rect 261186 154418 261422 154654
rect 261186 154098 261422 154334
rect 261186 118418 261422 118654
rect 261186 118098 261422 118334
rect 261186 82418 261422 82654
rect 261186 82098 261422 82334
rect 261186 46418 261422 46654
rect 261186 46098 261422 46334
rect 261186 10418 261422 10654
rect 261186 10098 261422 10334
rect 261186 -4342 261422 -4106
rect 261186 -4662 261422 -4426
rect 264786 302018 265022 302254
rect 264786 301698 265022 301934
rect 264786 266018 265022 266254
rect 264786 265698 265022 265934
rect 264786 230018 265022 230254
rect 264786 229698 265022 229934
rect 264786 194018 265022 194254
rect 264786 193698 265022 193934
rect 264786 158018 265022 158254
rect 264786 157698 265022 157934
rect 264786 122018 265022 122254
rect 264786 121698 265022 121934
rect 264786 86018 265022 86254
rect 264786 85698 265022 85934
rect 264786 50018 265022 50254
rect 264786 49698 265022 49934
rect 264786 14018 265022 14254
rect 264786 13698 265022 13934
rect 246786 -7162 247022 -6926
rect 246786 -7482 247022 -7246
rect 271986 309218 272222 309454
rect 271986 308898 272222 309134
rect 271986 273218 272222 273454
rect 271986 272898 272222 273134
rect 271986 237218 272222 237454
rect 271986 236898 272222 237134
rect 271986 201218 272222 201454
rect 271986 200898 272222 201134
rect 271986 165218 272222 165454
rect 271986 164898 272222 165134
rect 271986 129218 272222 129454
rect 271986 128898 272222 129134
rect 271986 93218 272222 93454
rect 271986 92898 272222 93134
rect 271986 57218 272222 57454
rect 271986 56898 272222 57134
rect 271986 21218 272222 21454
rect 271986 20898 272222 21134
rect 271986 -1522 272222 -1286
rect 271986 -1842 272222 -1606
rect 275586 312818 275822 313054
rect 275586 312498 275822 312734
rect 275586 276818 275822 277054
rect 275586 276498 275822 276734
rect 275586 240818 275822 241054
rect 275586 240498 275822 240734
rect 275586 204818 275822 205054
rect 275586 204498 275822 204734
rect 275586 168818 275822 169054
rect 275586 168498 275822 168734
rect 275586 132818 275822 133054
rect 275586 132498 275822 132734
rect 275586 96818 275822 97054
rect 275586 96498 275822 96734
rect 275586 60818 275822 61054
rect 275586 60498 275822 60734
rect 275586 24818 275822 25054
rect 275586 24498 275822 24734
rect 275586 -3402 275822 -3166
rect 275586 -3722 275822 -3486
rect 279186 316418 279422 316654
rect 279186 316098 279422 316334
rect 279186 280418 279422 280654
rect 279186 280098 279422 280334
rect 279186 244418 279422 244654
rect 279186 244098 279422 244334
rect 279186 208418 279422 208654
rect 279186 208098 279422 208334
rect 279186 172418 279422 172654
rect 279186 172098 279422 172334
rect 279186 136418 279422 136654
rect 279186 136098 279422 136334
rect 279186 100418 279422 100654
rect 279186 100098 279422 100334
rect 279186 64418 279422 64654
rect 279186 64098 279422 64334
rect 279186 28418 279422 28654
rect 279186 28098 279422 28334
rect 279186 -5282 279422 -5046
rect 279186 -5602 279422 -5366
rect 282786 320018 283022 320254
rect 282786 319698 283022 319934
rect 282786 284018 283022 284254
rect 282786 283698 283022 283934
rect 282786 248018 283022 248254
rect 282786 247698 283022 247934
rect 282786 212018 283022 212254
rect 282786 211698 283022 211934
rect 282786 176018 283022 176254
rect 282786 175698 283022 175934
rect 282786 140018 283022 140254
rect 282786 139698 283022 139934
rect 282786 104018 283022 104254
rect 282786 103698 283022 103934
rect 282786 68018 283022 68254
rect 282786 67698 283022 67934
rect 282786 32018 283022 32254
rect 282786 31698 283022 31934
rect 264786 -6222 265022 -5986
rect 264786 -6542 265022 -6306
rect 289986 291218 290222 291454
rect 289986 290898 290222 291134
rect 289986 255218 290222 255454
rect 289986 254898 290222 255134
rect 289986 219218 290222 219454
rect 289986 218898 290222 219134
rect 289986 183218 290222 183454
rect 289986 182898 290222 183134
rect 289986 147218 290222 147454
rect 289986 146898 290222 147134
rect 289986 111218 290222 111454
rect 289986 110898 290222 111134
rect 289986 75218 290222 75454
rect 289986 74898 290222 75134
rect 289986 39218 290222 39454
rect 289986 38898 290222 39134
rect 289986 3218 290222 3454
rect 289986 2898 290222 3134
rect 289986 -582 290222 -346
rect 289986 -902 290222 -666
rect 293586 294818 293822 295054
rect 293586 294498 293822 294734
rect 293586 258818 293822 259054
rect 293586 258498 293822 258734
rect 293586 222818 293822 223054
rect 293586 222498 293822 222734
rect 293586 186818 293822 187054
rect 293586 186498 293822 186734
rect 293586 150818 293822 151054
rect 293586 150498 293822 150734
rect 293586 114818 293822 115054
rect 293586 114498 293822 114734
rect 293586 78818 293822 79054
rect 293586 78498 293822 78734
rect 293586 42818 293822 43054
rect 293586 42498 293822 42734
rect 293586 6818 293822 7054
rect 293586 6498 293822 6734
rect 293586 -2462 293822 -2226
rect 293586 -2782 293822 -2546
rect 297186 298418 297422 298654
rect 297186 298098 297422 298334
rect 297186 262418 297422 262654
rect 297186 262098 297422 262334
rect 297186 226418 297422 226654
rect 297186 226098 297422 226334
rect 297186 190418 297422 190654
rect 297186 190098 297422 190334
rect 297186 154418 297422 154654
rect 297186 154098 297422 154334
rect 297186 118418 297422 118654
rect 297186 118098 297422 118334
rect 297186 82418 297422 82654
rect 297186 82098 297422 82334
rect 297186 46418 297422 46654
rect 297186 46098 297422 46334
rect 297186 10418 297422 10654
rect 297186 10098 297422 10334
rect 297186 -4342 297422 -4106
rect 297186 -4662 297422 -4426
rect 300786 302018 301022 302254
rect 300786 301698 301022 301934
rect 300786 266018 301022 266254
rect 300786 265698 301022 265934
rect 300786 230018 301022 230254
rect 300786 229698 301022 229934
rect 300786 194018 301022 194254
rect 300786 193698 301022 193934
rect 300786 158018 301022 158254
rect 300786 157698 301022 157934
rect 300786 122018 301022 122254
rect 300786 121698 301022 121934
rect 300786 86018 301022 86254
rect 300786 85698 301022 85934
rect 300786 50018 301022 50254
rect 300786 49698 301022 49934
rect 300786 14018 301022 14254
rect 300786 13698 301022 13934
rect 282786 -7162 283022 -6926
rect 282786 -7482 283022 -7246
rect 307986 309218 308222 309454
rect 307986 308898 308222 309134
rect 307986 273218 308222 273454
rect 307986 272898 308222 273134
rect 307986 237218 308222 237454
rect 307986 236898 308222 237134
rect 307986 201218 308222 201454
rect 307986 200898 308222 201134
rect 307986 165218 308222 165454
rect 307986 164898 308222 165134
rect 307986 129218 308222 129454
rect 307986 128898 308222 129134
rect 307986 93218 308222 93454
rect 307986 92898 308222 93134
rect 307986 57218 308222 57454
rect 307986 56898 308222 57134
rect 307986 21218 308222 21454
rect 307986 20898 308222 21134
rect 307986 -1522 308222 -1286
rect 307986 -1842 308222 -1606
rect 311586 312818 311822 313054
rect 311586 312498 311822 312734
rect 311586 276818 311822 277054
rect 311586 276498 311822 276734
rect 311586 240818 311822 241054
rect 311586 240498 311822 240734
rect 311586 204818 311822 205054
rect 311586 204498 311822 204734
rect 311586 168818 311822 169054
rect 311586 168498 311822 168734
rect 311586 132818 311822 133054
rect 311586 132498 311822 132734
rect 311586 96818 311822 97054
rect 311586 96498 311822 96734
rect 311586 60818 311822 61054
rect 311586 60498 311822 60734
rect 311586 24818 311822 25054
rect 311586 24498 311822 24734
rect 311586 -3402 311822 -3166
rect 311586 -3722 311822 -3486
rect 315186 316418 315422 316654
rect 315186 316098 315422 316334
rect 315186 280418 315422 280654
rect 315186 280098 315422 280334
rect 315186 244418 315422 244654
rect 315186 244098 315422 244334
rect 315186 208418 315422 208654
rect 315186 208098 315422 208334
rect 315186 172418 315422 172654
rect 315186 172098 315422 172334
rect 315186 136418 315422 136654
rect 315186 136098 315422 136334
rect 315186 100418 315422 100654
rect 315186 100098 315422 100334
rect 315186 64418 315422 64654
rect 315186 64098 315422 64334
rect 315186 28418 315422 28654
rect 315186 28098 315422 28334
rect 315186 -5282 315422 -5046
rect 315186 -5602 315422 -5366
rect 318786 320018 319022 320254
rect 318786 319698 319022 319934
rect 318786 284018 319022 284254
rect 318786 283698 319022 283934
rect 318786 248018 319022 248254
rect 318786 247698 319022 247934
rect 318786 212018 319022 212254
rect 318786 211698 319022 211934
rect 318786 176018 319022 176254
rect 318786 175698 319022 175934
rect 318786 140018 319022 140254
rect 318786 139698 319022 139934
rect 318786 104018 319022 104254
rect 318786 103698 319022 103934
rect 318786 68018 319022 68254
rect 318786 67698 319022 67934
rect 318786 32018 319022 32254
rect 318786 31698 319022 31934
rect 300786 -6222 301022 -5986
rect 300786 -6542 301022 -6306
rect 325986 291218 326222 291454
rect 325986 290898 326222 291134
rect 325986 255218 326222 255454
rect 325986 254898 326222 255134
rect 325986 219218 326222 219454
rect 325986 218898 326222 219134
rect 325986 183218 326222 183454
rect 325986 182898 326222 183134
rect 325986 147218 326222 147454
rect 325986 146898 326222 147134
rect 325986 111218 326222 111454
rect 325986 110898 326222 111134
rect 325986 75218 326222 75454
rect 325986 74898 326222 75134
rect 325986 39218 326222 39454
rect 325986 38898 326222 39134
rect 325986 3218 326222 3454
rect 325986 2898 326222 3134
rect 325986 -582 326222 -346
rect 325986 -902 326222 -666
rect 329586 294818 329822 295054
rect 329586 294498 329822 294734
rect 329586 258818 329822 259054
rect 329586 258498 329822 258734
rect 329586 222818 329822 223054
rect 329586 222498 329822 222734
rect 329586 186818 329822 187054
rect 329586 186498 329822 186734
rect 329586 150818 329822 151054
rect 329586 150498 329822 150734
rect 329586 114818 329822 115054
rect 329586 114498 329822 114734
rect 329586 78818 329822 79054
rect 329586 78498 329822 78734
rect 329586 42818 329822 43054
rect 329586 42498 329822 42734
rect 329586 6818 329822 7054
rect 329586 6498 329822 6734
rect 329586 -2462 329822 -2226
rect 329586 -2782 329822 -2546
rect 333186 298418 333422 298654
rect 333186 298098 333422 298334
rect 333186 262418 333422 262654
rect 333186 262098 333422 262334
rect 333186 226418 333422 226654
rect 333186 226098 333422 226334
rect 333186 190418 333422 190654
rect 333186 190098 333422 190334
rect 333186 154418 333422 154654
rect 333186 154098 333422 154334
rect 333186 118418 333422 118654
rect 333186 118098 333422 118334
rect 333186 82418 333422 82654
rect 333186 82098 333422 82334
rect 333186 46418 333422 46654
rect 333186 46098 333422 46334
rect 333186 10418 333422 10654
rect 333186 10098 333422 10334
rect 333186 -4342 333422 -4106
rect 333186 -4662 333422 -4426
rect 336786 302018 337022 302254
rect 336786 301698 337022 301934
rect 336786 266018 337022 266254
rect 336786 265698 337022 265934
rect 336786 230018 337022 230254
rect 336786 229698 337022 229934
rect 336786 194018 337022 194254
rect 336786 193698 337022 193934
rect 336786 158018 337022 158254
rect 336786 157698 337022 157934
rect 336786 122018 337022 122254
rect 336786 121698 337022 121934
rect 336786 86018 337022 86254
rect 336786 85698 337022 85934
rect 336786 50018 337022 50254
rect 336786 49698 337022 49934
rect 336786 14018 337022 14254
rect 336786 13698 337022 13934
rect 318786 -7162 319022 -6926
rect 318786 -7482 319022 -7246
rect 343986 309218 344222 309454
rect 343986 308898 344222 309134
rect 343986 273218 344222 273454
rect 343986 272898 344222 273134
rect 343986 237218 344222 237454
rect 343986 236898 344222 237134
rect 343986 201218 344222 201454
rect 343986 200898 344222 201134
rect 343986 165218 344222 165454
rect 343986 164898 344222 165134
rect 343986 129218 344222 129454
rect 343986 128898 344222 129134
rect 343986 93218 344222 93454
rect 343986 92898 344222 93134
rect 343986 57218 344222 57454
rect 343986 56898 344222 57134
rect 343986 21218 344222 21454
rect 343986 20898 344222 21134
rect 343986 -1522 344222 -1286
rect 343986 -1842 344222 -1606
rect 347586 312818 347822 313054
rect 347586 312498 347822 312734
rect 347586 276818 347822 277054
rect 347586 276498 347822 276734
rect 347586 240818 347822 241054
rect 347586 240498 347822 240734
rect 347586 204818 347822 205054
rect 347586 204498 347822 204734
rect 347586 168818 347822 169054
rect 347586 168498 347822 168734
rect 347586 132818 347822 133054
rect 347586 132498 347822 132734
rect 347586 96818 347822 97054
rect 347586 96498 347822 96734
rect 347586 60818 347822 61054
rect 347586 60498 347822 60734
rect 347586 24818 347822 25054
rect 347586 24498 347822 24734
rect 347586 -3402 347822 -3166
rect 347586 -3722 347822 -3486
rect 351186 316418 351422 316654
rect 351186 316098 351422 316334
rect 351186 280418 351422 280654
rect 351186 280098 351422 280334
rect 351186 244418 351422 244654
rect 351186 244098 351422 244334
rect 351186 208418 351422 208654
rect 351186 208098 351422 208334
rect 351186 172418 351422 172654
rect 351186 172098 351422 172334
rect 351186 136418 351422 136654
rect 351186 136098 351422 136334
rect 351186 100418 351422 100654
rect 351186 100098 351422 100334
rect 351186 64418 351422 64654
rect 351186 64098 351422 64334
rect 351186 28418 351422 28654
rect 351186 28098 351422 28334
rect 351186 -5282 351422 -5046
rect 351186 -5602 351422 -5366
rect 354786 320018 355022 320254
rect 354786 319698 355022 319934
rect 354786 284018 355022 284254
rect 354786 283698 355022 283934
rect 354786 248018 355022 248254
rect 354786 247698 355022 247934
rect 354786 212018 355022 212254
rect 354786 211698 355022 211934
rect 354786 176018 355022 176254
rect 354786 175698 355022 175934
rect 354786 140018 355022 140254
rect 354786 139698 355022 139934
rect 354786 104018 355022 104254
rect 354786 103698 355022 103934
rect 354786 68018 355022 68254
rect 354786 67698 355022 67934
rect 354786 32018 355022 32254
rect 354786 31698 355022 31934
rect 336786 -6222 337022 -5986
rect 336786 -6542 337022 -6306
rect 361986 291218 362222 291454
rect 361986 290898 362222 291134
rect 361986 255218 362222 255454
rect 361986 254898 362222 255134
rect 361986 219218 362222 219454
rect 361986 218898 362222 219134
rect 361986 183218 362222 183454
rect 361986 182898 362222 183134
rect 361986 147218 362222 147454
rect 361986 146898 362222 147134
rect 361986 111218 362222 111454
rect 361986 110898 362222 111134
rect 361986 75218 362222 75454
rect 361986 74898 362222 75134
rect 361986 39218 362222 39454
rect 361986 38898 362222 39134
rect 361986 3218 362222 3454
rect 361986 2898 362222 3134
rect 361986 -582 362222 -346
rect 361986 -902 362222 -666
rect 365586 294818 365822 295054
rect 365586 294498 365822 294734
rect 365586 258818 365822 259054
rect 365586 258498 365822 258734
rect 365586 222818 365822 223054
rect 365586 222498 365822 222734
rect 365586 186818 365822 187054
rect 365586 186498 365822 186734
rect 365586 150818 365822 151054
rect 365586 150498 365822 150734
rect 365586 114818 365822 115054
rect 365586 114498 365822 114734
rect 365586 78818 365822 79054
rect 365586 78498 365822 78734
rect 365586 42818 365822 43054
rect 365586 42498 365822 42734
rect 365586 6818 365822 7054
rect 365586 6498 365822 6734
rect 365586 -2462 365822 -2226
rect 365586 -2782 365822 -2546
rect 369186 298418 369422 298654
rect 369186 298098 369422 298334
rect 369186 262418 369422 262654
rect 369186 262098 369422 262334
rect 369186 226418 369422 226654
rect 369186 226098 369422 226334
rect 369186 190418 369422 190654
rect 369186 190098 369422 190334
rect 369186 154418 369422 154654
rect 369186 154098 369422 154334
rect 369186 118418 369422 118654
rect 369186 118098 369422 118334
rect 369186 82418 369422 82654
rect 369186 82098 369422 82334
rect 369186 46418 369422 46654
rect 369186 46098 369422 46334
rect 369186 10418 369422 10654
rect 369186 10098 369422 10334
rect 369186 -4342 369422 -4106
rect 369186 -4662 369422 -4426
rect 372786 302018 373022 302254
rect 372786 301698 373022 301934
rect 372786 266018 373022 266254
rect 372786 265698 373022 265934
rect 372786 230018 373022 230254
rect 372786 229698 373022 229934
rect 372786 194018 373022 194254
rect 372786 193698 373022 193934
rect 372786 158018 373022 158254
rect 372786 157698 373022 157934
rect 372786 122018 373022 122254
rect 372786 121698 373022 121934
rect 372786 86018 373022 86254
rect 372786 85698 373022 85934
rect 372786 50018 373022 50254
rect 372786 49698 373022 49934
rect 372786 14018 373022 14254
rect 372786 13698 373022 13934
rect 354786 -7162 355022 -6926
rect 354786 -7482 355022 -7246
rect 379986 309218 380222 309454
rect 379986 308898 380222 309134
rect 379986 273218 380222 273454
rect 379986 272898 380222 273134
rect 379986 237218 380222 237454
rect 379986 236898 380222 237134
rect 379986 201218 380222 201454
rect 379986 200898 380222 201134
rect 379986 165218 380222 165454
rect 379986 164898 380222 165134
rect 379986 129218 380222 129454
rect 379986 128898 380222 129134
rect 379986 93218 380222 93454
rect 379986 92898 380222 93134
rect 379986 57218 380222 57454
rect 379986 56898 380222 57134
rect 379986 21218 380222 21454
rect 379986 20898 380222 21134
rect 379986 -1522 380222 -1286
rect 379986 -1842 380222 -1606
rect 383586 312818 383822 313054
rect 383586 312498 383822 312734
rect 383586 276818 383822 277054
rect 383586 276498 383822 276734
rect 383586 240818 383822 241054
rect 383586 240498 383822 240734
rect 383586 204818 383822 205054
rect 383586 204498 383822 204734
rect 383586 168818 383822 169054
rect 383586 168498 383822 168734
rect 383586 132818 383822 133054
rect 383586 132498 383822 132734
rect 383586 96818 383822 97054
rect 383586 96498 383822 96734
rect 383586 60818 383822 61054
rect 383586 60498 383822 60734
rect 383586 24818 383822 25054
rect 383586 24498 383822 24734
rect 383586 -3402 383822 -3166
rect 383586 -3722 383822 -3486
rect 387186 316418 387422 316654
rect 387186 316098 387422 316334
rect 387186 280418 387422 280654
rect 387186 280098 387422 280334
rect 387186 244418 387422 244654
rect 387186 244098 387422 244334
rect 387186 208418 387422 208654
rect 387186 208098 387422 208334
rect 387186 172418 387422 172654
rect 387186 172098 387422 172334
rect 387186 136418 387422 136654
rect 387186 136098 387422 136334
rect 387186 100418 387422 100654
rect 387186 100098 387422 100334
rect 387186 64418 387422 64654
rect 387186 64098 387422 64334
rect 387186 28418 387422 28654
rect 387186 28098 387422 28334
rect 387186 -5282 387422 -5046
rect 387186 -5602 387422 -5366
rect 390786 320018 391022 320254
rect 390786 319698 391022 319934
rect 390786 284018 391022 284254
rect 390786 283698 391022 283934
rect 390786 248018 391022 248254
rect 390786 247698 391022 247934
rect 390786 212018 391022 212254
rect 390786 211698 391022 211934
rect 390786 176018 391022 176254
rect 390786 175698 391022 175934
rect 390786 140018 391022 140254
rect 390786 139698 391022 139934
rect 390786 104018 391022 104254
rect 390786 103698 391022 103934
rect 390786 68018 391022 68254
rect 390786 67698 391022 67934
rect 390786 32018 391022 32254
rect 390786 31698 391022 31934
rect 372786 -6222 373022 -5986
rect 372786 -6542 373022 -6306
rect 397986 291218 398222 291454
rect 397986 290898 398222 291134
rect 397986 255218 398222 255454
rect 397986 254898 398222 255134
rect 397986 219218 398222 219454
rect 397986 218898 398222 219134
rect 397986 183218 398222 183454
rect 397986 182898 398222 183134
rect 397986 147218 398222 147454
rect 397986 146898 398222 147134
rect 397986 111218 398222 111454
rect 397986 110898 398222 111134
rect 397986 75218 398222 75454
rect 397986 74898 398222 75134
rect 397986 39218 398222 39454
rect 397986 38898 398222 39134
rect 397986 3218 398222 3454
rect 397986 2898 398222 3134
rect 397986 -582 398222 -346
rect 397986 -902 398222 -666
rect 401586 294818 401822 295054
rect 401586 294498 401822 294734
rect 401586 258818 401822 259054
rect 401586 258498 401822 258734
rect 401586 222818 401822 223054
rect 401586 222498 401822 222734
rect 401586 186818 401822 187054
rect 401586 186498 401822 186734
rect 401586 150818 401822 151054
rect 401586 150498 401822 150734
rect 401586 114818 401822 115054
rect 401586 114498 401822 114734
rect 401586 78818 401822 79054
rect 401586 78498 401822 78734
rect 401586 42818 401822 43054
rect 401586 42498 401822 42734
rect 401586 6818 401822 7054
rect 401586 6498 401822 6734
rect 401586 -2462 401822 -2226
rect 401586 -2782 401822 -2546
rect 405186 298418 405422 298654
rect 405186 298098 405422 298334
rect 405186 262418 405422 262654
rect 405186 262098 405422 262334
rect 405186 226418 405422 226654
rect 405186 226098 405422 226334
rect 405186 190418 405422 190654
rect 405186 190098 405422 190334
rect 405186 154418 405422 154654
rect 405186 154098 405422 154334
rect 405186 118418 405422 118654
rect 405186 118098 405422 118334
rect 405186 82418 405422 82654
rect 405186 82098 405422 82334
rect 405186 46418 405422 46654
rect 405186 46098 405422 46334
rect 405186 10418 405422 10654
rect 405186 10098 405422 10334
rect 405186 -4342 405422 -4106
rect 405186 -4662 405422 -4426
rect 408786 302018 409022 302254
rect 408786 301698 409022 301934
rect 408786 266018 409022 266254
rect 408786 265698 409022 265934
rect 408786 230018 409022 230254
rect 408786 229698 409022 229934
rect 408786 194018 409022 194254
rect 408786 193698 409022 193934
rect 408786 158018 409022 158254
rect 408786 157698 409022 157934
rect 408786 122018 409022 122254
rect 408786 121698 409022 121934
rect 408786 86018 409022 86254
rect 408786 85698 409022 85934
rect 408786 50018 409022 50254
rect 408786 49698 409022 49934
rect 408786 14018 409022 14254
rect 408786 13698 409022 13934
rect 390786 -7162 391022 -6926
rect 390786 -7482 391022 -7246
rect 415986 309218 416222 309454
rect 415986 308898 416222 309134
rect 415986 273218 416222 273454
rect 415986 272898 416222 273134
rect 415986 237218 416222 237454
rect 415986 236898 416222 237134
rect 415986 201218 416222 201454
rect 415986 200898 416222 201134
rect 415986 165218 416222 165454
rect 415986 164898 416222 165134
rect 415986 129218 416222 129454
rect 415986 128898 416222 129134
rect 415986 93218 416222 93454
rect 415986 92898 416222 93134
rect 415986 57218 416222 57454
rect 415986 56898 416222 57134
rect 415986 21218 416222 21454
rect 415986 20898 416222 21134
rect 415986 -1522 416222 -1286
rect 415986 -1842 416222 -1606
rect 419586 312818 419822 313054
rect 419586 312498 419822 312734
rect 419586 276818 419822 277054
rect 419586 276498 419822 276734
rect 419586 240818 419822 241054
rect 419586 240498 419822 240734
rect 419586 204818 419822 205054
rect 419586 204498 419822 204734
rect 419586 168818 419822 169054
rect 419586 168498 419822 168734
rect 419586 132818 419822 133054
rect 419586 132498 419822 132734
rect 419586 96818 419822 97054
rect 419586 96498 419822 96734
rect 419586 60818 419822 61054
rect 419586 60498 419822 60734
rect 419586 24818 419822 25054
rect 419586 24498 419822 24734
rect 419586 -3402 419822 -3166
rect 419586 -3722 419822 -3486
rect 423186 316418 423422 316654
rect 423186 316098 423422 316334
rect 423186 280418 423422 280654
rect 423186 280098 423422 280334
rect 423186 244418 423422 244654
rect 423186 244098 423422 244334
rect 423186 208418 423422 208654
rect 423186 208098 423422 208334
rect 423186 172418 423422 172654
rect 423186 172098 423422 172334
rect 423186 136418 423422 136654
rect 423186 136098 423422 136334
rect 423186 100418 423422 100654
rect 423186 100098 423422 100334
rect 423186 64418 423422 64654
rect 423186 64098 423422 64334
rect 423186 28418 423422 28654
rect 423186 28098 423422 28334
rect 423186 -5282 423422 -5046
rect 423186 -5602 423422 -5366
rect 426786 320018 427022 320254
rect 426786 319698 427022 319934
rect 426786 284018 427022 284254
rect 426786 283698 427022 283934
rect 426786 248018 427022 248254
rect 426786 247698 427022 247934
rect 426786 212018 427022 212254
rect 426786 211698 427022 211934
rect 426786 176018 427022 176254
rect 426786 175698 427022 175934
rect 426786 140018 427022 140254
rect 426786 139698 427022 139934
rect 426786 104018 427022 104254
rect 426786 103698 427022 103934
rect 426786 68018 427022 68254
rect 426786 67698 427022 67934
rect 426786 32018 427022 32254
rect 426786 31698 427022 31934
rect 408786 -6222 409022 -5986
rect 408786 -6542 409022 -6306
rect 441186 334418 441422 334654
rect 441186 334098 441422 334334
rect 433986 291218 434222 291454
rect 433986 290898 434222 291134
rect 433986 255218 434222 255454
rect 433986 254898 434222 255134
rect 433986 219218 434222 219454
rect 433986 218898 434222 219134
rect 433986 183218 434222 183454
rect 433986 182898 434222 183134
rect 433986 147218 434222 147454
rect 433986 146898 434222 147134
rect 433986 111218 434222 111454
rect 433986 110898 434222 111134
rect 433986 75218 434222 75454
rect 433986 74898 434222 75134
rect 433986 39218 434222 39454
rect 433986 38898 434222 39134
rect 433986 3218 434222 3454
rect 433986 2898 434222 3134
rect 433986 -582 434222 -346
rect 433986 -902 434222 -666
rect 437586 294818 437822 295054
rect 437586 294498 437822 294734
rect 437586 258818 437822 259054
rect 437586 258498 437822 258734
rect 437586 222818 437822 223054
rect 437586 222498 437822 222734
rect 437586 186818 437822 187054
rect 437586 186498 437822 186734
rect 437586 150818 437822 151054
rect 437586 150498 437822 150734
rect 437586 114818 437822 115054
rect 437586 114498 437822 114734
rect 437586 78818 437822 79054
rect 437586 78498 437822 78734
rect 437586 42818 437822 43054
rect 437586 42498 437822 42734
rect 437586 6818 437822 7054
rect 437586 6498 437822 6734
rect 437586 -2462 437822 -2226
rect 437586 -2782 437822 -2546
rect 441186 298418 441422 298654
rect 441186 298098 441422 298334
rect 441186 262418 441422 262654
rect 441186 262098 441422 262334
rect 441186 226418 441422 226654
rect 441186 226098 441422 226334
rect 441186 190418 441422 190654
rect 441186 190098 441422 190334
rect 441186 154418 441422 154654
rect 441186 154098 441422 154334
rect 441186 118418 441422 118654
rect 441186 118098 441422 118334
rect 441186 82418 441422 82654
rect 441186 82098 441422 82334
rect 441186 46418 441422 46654
rect 441186 46098 441422 46334
rect 441186 10418 441422 10654
rect 441186 10098 441422 10334
rect 441186 -4342 441422 -4106
rect 441186 -4662 441422 -4426
rect 462786 711182 463022 711418
rect 462786 710862 463022 711098
rect 459186 709302 459422 709538
rect 459186 708982 459422 709218
rect 455586 707422 455822 707658
rect 455586 707102 455822 707338
rect 444786 698018 445022 698254
rect 444786 697698 445022 697934
rect 444786 662018 445022 662254
rect 444786 661698 445022 661934
rect 444786 626018 445022 626254
rect 444786 625698 445022 625934
rect 444786 590018 445022 590254
rect 444786 589698 445022 589934
rect 444786 554018 445022 554254
rect 444786 553698 445022 553934
rect 444786 518018 445022 518254
rect 444786 517698 445022 517934
rect 444786 482018 445022 482254
rect 444786 481698 445022 481934
rect 444786 446018 445022 446254
rect 444786 445698 445022 445934
rect 444786 410018 445022 410254
rect 444786 409698 445022 409934
rect 444786 374018 445022 374254
rect 444786 373698 445022 373934
rect 444786 338018 445022 338254
rect 444786 337698 445022 337934
rect 444786 302018 445022 302254
rect 444786 301698 445022 301934
rect 444786 266018 445022 266254
rect 444786 265698 445022 265934
rect 444786 230018 445022 230254
rect 444786 229698 445022 229934
rect 444786 194018 445022 194254
rect 444786 193698 445022 193934
rect 444786 158018 445022 158254
rect 444786 157698 445022 157934
rect 444786 122018 445022 122254
rect 444786 121698 445022 121934
rect 444786 86018 445022 86254
rect 444786 85698 445022 85934
rect 444786 50018 445022 50254
rect 444786 49698 445022 49934
rect 444786 14018 445022 14254
rect 444786 13698 445022 13934
rect 426786 -7162 427022 -6926
rect 426786 -7482 427022 -7246
rect 451986 705542 452222 705778
rect 451986 705222 452222 705458
rect 451986 669218 452222 669454
rect 451986 668898 452222 669134
rect 451986 633218 452222 633454
rect 451986 632898 452222 633134
rect 451986 597218 452222 597454
rect 451986 596898 452222 597134
rect 451986 561218 452222 561454
rect 451986 560898 452222 561134
rect 451986 525218 452222 525454
rect 451986 524898 452222 525134
rect 451986 489218 452222 489454
rect 451986 488898 452222 489134
rect 451986 453218 452222 453454
rect 451986 452898 452222 453134
rect 451986 417218 452222 417454
rect 451986 416898 452222 417134
rect 451986 381218 452222 381454
rect 451986 380898 452222 381134
rect 451986 345218 452222 345454
rect 451986 344898 452222 345134
rect 451986 309218 452222 309454
rect 451986 308898 452222 309134
rect 451986 273218 452222 273454
rect 451986 272898 452222 273134
rect 451986 237218 452222 237454
rect 451986 236898 452222 237134
rect 451986 201218 452222 201454
rect 451986 200898 452222 201134
rect 451986 165218 452222 165454
rect 451986 164898 452222 165134
rect 451986 129218 452222 129454
rect 451986 128898 452222 129134
rect 451986 93218 452222 93454
rect 451986 92898 452222 93134
rect 451986 57218 452222 57454
rect 451986 56898 452222 57134
rect 451986 21218 452222 21454
rect 451986 20898 452222 21134
rect 451986 -1522 452222 -1286
rect 451986 -1842 452222 -1606
rect 455586 672818 455822 673054
rect 455586 672498 455822 672734
rect 455586 636818 455822 637054
rect 455586 636498 455822 636734
rect 455586 600818 455822 601054
rect 455586 600498 455822 600734
rect 455586 564818 455822 565054
rect 455586 564498 455822 564734
rect 455586 528818 455822 529054
rect 455586 528498 455822 528734
rect 455586 492818 455822 493054
rect 455586 492498 455822 492734
rect 455586 456818 455822 457054
rect 455586 456498 455822 456734
rect 455586 420818 455822 421054
rect 455586 420498 455822 420734
rect 455586 384818 455822 385054
rect 455586 384498 455822 384734
rect 455586 348818 455822 349054
rect 455586 348498 455822 348734
rect 455586 312818 455822 313054
rect 455586 312498 455822 312734
rect 455586 276818 455822 277054
rect 455586 276498 455822 276734
rect 455586 240818 455822 241054
rect 455586 240498 455822 240734
rect 455586 204818 455822 205054
rect 455586 204498 455822 204734
rect 455586 168818 455822 169054
rect 455586 168498 455822 168734
rect 455586 132818 455822 133054
rect 455586 132498 455822 132734
rect 455586 96818 455822 97054
rect 455586 96498 455822 96734
rect 455586 60818 455822 61054
rect 455586 60498 455822 60734
rect 455586 24818 455822 25054
rect 455586 24498 455822 24734
rect 455586 -3402 455822 -3166
rect 455586 -3722 455822 -3486
rect 459186 676418 459422 676654
rect 459186 676098 459422 676334
rect 459186 640418 459422 640654
rect 459186 640098 459422 640334
rect 459186 604418 459422 604654
rect 459186 604098 459422 604334
rect 459186 568418 459422 568654
rect 459186 568098 459422 568334
rect 459186 532418 459422 532654
rect 459186 532098 459422 532334
rect 459186 496418 459422 496654
rect 459186 496098 459422 496334
rect 459186 460418 459422 460654
rect 459186 460098 459422 460334
rect 459186 424418 459422 424654
rect 459186 424098 459422 424334
rect 459186 388418 459422 388654
rect 459186 388098 459422 388334
rect 459186 352418 459422 352654
rect 459186 352098 459422 352334
rect 459186 316418 459422 316654
rect 459186 316098 459422 316334
rect 459186 280418 459422 280654
rect 459186 280098 459422 280334
rect 459186 244418 459422 244654
rect 459186 244098 459422 244334
rect 459186 208418 459422 208654
rect 459186 208098 459422 208334
rect 459186 172418 459422 172654
rect 459186 172098 459422 172334
rect 459186 136418 459422 136654
rect 459186 136098 459422 136334
rect 459186 100418 459422 100654
rect 459186 100098 459422 100334
rect 459186 64418 459422 64654
rect 459186 64098 459422 64334
rect 459186 28418 459422 28654
rect 459186 28098 459422 28334
rect 459186 -5282 459422 -5046
rect 459186 -5602 459422 -5366
rect 480786 710242 481022 710478
rect 480786 709922 481022 710158
rect 477186 708362 477422 708598
rect 477186 708042 477422 708278
rect 473586 706482 473822 706718
rect 473586 706162 473822 706398
rect 462786 680018 463022 680254
rect 462786 679698 463022 679934
rect 462786 644018 463022 644254
rect 462786 643698 463022 643934
rect 462786 608018 463022 608254
rect 462786 607698 463022 607934
rect 462786 572018 463022 572254
rect 462786 571698 463022 571934
rect 462786 536018 463022 536254
rect 462786 535698 463022 535934
rect 462786 500018 463022 500254
rect 462786 499698 463022 499934
rect 462786 464018 463022 464254
rect 462786 463698 463022 463934
rect 462786 428018 463022 428254
rect 462786 427698 463022 427934
rect 462786 392018 463022 392254
rect 462786 391698 463022 391934
rect 462786 356018 463022 356254
rect 462786 355698 463022 355934
rect 462786 320018 463022 320254
rect 462786 319698 463022 319934
rect 462786 284018 463022 284254
rect 462786 283698 463022 283934
rect 462786 248018 463022 248254
rect 462786 247698 463022 247934
rect 462786 212018 463022 212254
rect 462786 211698 463022 211934
rect 462786 176018 463022 176254
rect 462786 175698 463022 175934
rect 462786 140018 463022 140254
rect 462786 139698 463022 139934
rect 462786 104018 463022 104254
rect 462786 103698 463022 103934
rect 462786 68018 463022 68254
rect 462786 67698 463022 67934
rect 462786 32018 463022 32254
rect 462786 31698 463022 31934
rect 444786 -6222 445022 -5986
rect 444786 -6542 445022 -6306
rect 469986 704602 470222 704838
rect 469986 704282 470222 704518
rect 469986 687218 470222 687454
rect 469986 686898 470222 687134
rect 469986 651218 470222 651454
rect 469986 650898 470222 651134
rect 469986 615218 470222 615454
rect 469986 614898 470222 615134
rect 469986 579218 470222 579454
rect 469986 578898 470222 579134
rect 469986 543218 470222 543454
rect 469986 542898 470222 543134
rect 469986 507218 470222 507454
rect 469986 506898 470222 507134
rect 469986 471218 470222 471454
rect 469986 470898 470222 471134
rect 469986 435218 470222 435454
rect 469986 434898 470222 435134
rect 469986 399218 470222 399454
rect 469986 398898 470222 399134
rect 469986 363218 470222 363454
rect 469986 362898 470222 363134
rect 469986 327218 470222 327454
rect 469986 326898 470222 327134
rect 469986 291218 470222 291454
rect 469986 290898 470222 291134
rect 469986 255218 470222 255454
rect 469986 254898 470222 255134
rect 469986 219218 470222 219454
rect 469986 218898 470222 219134
rect 469986 183218 470222 183454
rect 469986 182898 470222 183134
rect 469986 147218 470222 147454
rect 469986 146898 470222 147134
rect 469986 111218 470222 111454
rect 469986 110898 470222 111134
rect 469986 75218 470222 75454
rect 469986 74898 470222 75134
rect 469986 39218 470222 39454
rect 469986 38898 470222 39134
rect 469986 3218 470222 3454
rect 469986 2898 470222 3134
rect 469986 -582 470222 -346
rect 469986 -902 470222 -666
rect 473586 690818 473822 691054
rect 473586 690498 473822 690734
rect 473586 654818 473822 655054
rect 473586 654498 473822 654734
rect 473586 618818 473822 619054
rect 473586 618498 473822 618734
rect 473586 582818 473822 583054
rect 473586 582498 473822 582734
rect 473586 546818 473822 547054
rect 473586 546498 473822 546734
rect 473586 510818 473822 511054
rect 473586 510498 473822 510734
rect 473586 474818 473822 475054
rect 473586 474498 473822 474734
rect 473586 438818 473822 439054
rect 473586 438498 473822 438734
rect 473586 402818 473822 403054
rect 473586 402498 473822 402734
rect 473586 366818 473822 367054
rect 473586 366498 473822 366734
rect 473586 330818 473822 331054
rect 473586 330498 473822 330734
rect 473586 294818 473822 295054
rect 473586 294498 473822 294734
rect 473586 258818 473822 259054
rect 473586 258498 473822 258734
rect 473586 222818 473822 223054
rect 473586 222498 473822 222734
rect 473586 186818 473822 187054
rect 473586 186498 473822 186734
rect 473586 150818 473822 151054
rect 473586 150498 473822 150734
rect 473586 114818 473822 115054
rect 473586 114498 473822 114734
rect 473586 78818 473822 79054
rect 473586 78498 473822 78734
rect 473586 42818 473822 43054
rect 473586 42498 473822 42734
rect 473586 6818 473822 7054
rect 473586 6498 473822 6734
rect 473586 -2462 473822 -2226
rect 473586 -2782 473822 -2546
rect 477186 694418 477422 694654
rect 477186 694098 477422 694334
rect 477186 658418 477422 658654
rect 477186 658098 477422 658334
rect 477186 622418 477422 622654
rect 477186 622098 477422 622334
rect 477186 586418 477422 586654
rect 477186 586098 477422 586334
rect 477186 550418 477422 550654
rect 477186 550098 477422 550334
rect 477186 514418 477422 514654
rect 477186 514098 477422 514334
rect 477186 478418 477422 478654
rect 477186 478098 477422 478334
rect 477186 442418 477422 442654
rect 477186 442098 477422 442334
rect 477186 406418 477422 406654
rect 477186 406098 477422 406334
rect 477186 370418 477422 370654
rect 477186 370098 477422 370334
rect 477186 334418 477422 334654
rect 477186 334098 477422 334334
rect 477186 298418 477422 298654
rect 477186 298098 477422 298334
rect 477186 262418 477422 262654
rect 477186 262098 477422 262334
rect 477186 226418 477422 226654
rect 477186 226098 477422 226334
rect 477186 190418 477422 190654
rect 477186 190098 477422 190334
rect 477186 154418 477422 154654
rect 477186 154098 477422 154334
rect 477186 118418 477422 118654
rect 477186 118098 477422 118334
rect 477186 82418 477422 82654
rect 477186 82098 477422 82334
rect 477186 46418 477422 46654
rect 477186 46098 477422 46334
rect 477186 10418 477422 10654
rect 477186 10098 477422 10334
rect 477186 -4342 477422 -4106
rect 477186 -4662 477422 -4426
rect 498786 711182 499022 711418
rect 498786 710862 499022 711098
rect 495186 709302 495422 709538
rect 495186 708982 495422 709218
rect 491586 707422 491822 707658
rect 491586 707102 491822 707338
rect 480786 698018 481022 698254
rect 480786 697698 481022 697934
rect 480786 662018 481022 662254
rect 480786 661698 481022 661934
rect 480786 626018 481022 626254
rect 480786 625698 481022 625934
rect 480786 590018 481022 590254
rect 480786 589698 481022 589934
rect 480786 554018 481022 554254
rect 480786 553698 481022 553934
rect 480786 518018 481022 518254
rect 480786 517698 481022 517934
rect 480786 482018 481022 482254
rect 480786 481698 481022 481934
rect 480786 446018 481022 446254
rect 480786 445698 481022 445934
rect 480786 410018 481022 410254
rect 480786 409698 481022 409934
rect 480786 374018 481022 374254
rect 480786 373698 481022 373934
rect 480786 338018 481022 338254
rect 480786 337698 481022 337934
rect 480786 302018 481022 302254
rect 480786 301698 481022 301934
rect 480786 266018 481022 266254
rect 480786 265698 481022 265934
rect 480786 230018 481022 230254
rect 480786 229698 481022 229934
rect 480786 194018 481022 194254
rect 480786 193698 481022 193934
rect 480786 158018 481022 158254
rect 480786 157698 481022 157934
rect 480786 122018 481022 122254
rect 480786 121698 481022 121934
rect 480786 86018 481022 86254
rect 480786 85698 481022 85934
rect 480786 50018 481022 50254
rect 480786 49698 481022 49934
rect 480786 14018 481022 14254
rect 480786 13698 481022 13934
rect 462786 -7162 463022 -6926
rect 462786 -7482 463022 -7246
rect 487986 705542 488222 705778
rect 487986 705222 488222 705458
rect 487986 669218 488222 669454
rect 487986 668898 488222 669134
rect 487986 633218 488222 633454
rect 487986 632898 488222 633134
rect 487986 597218 488222 597454
rect 487986 596898 488222 597134
rect 487986 561218 488222 561454
rect 487986 560898 488222 561134
rect 487986 525218 488222 525454
rect 487986 524898 488222 525134
rect 487986 489218 488222 489454
rect 487986 488898 488222 489134
rect 487986 453218 488222 453454
rect 487986 452898 488222 453134
rect 487986 417218 488222 417454
rect 487986 416898 488222 417134
rect 487986 381218 488222 381454
rect 487986 380898 488222 381134
rect 487986 345218 488222 345454
rect 487986 344898 488222 345134
rect 487986 309218 488222 309454
rect 487986 308898 488222 309134
rect 487986 273218 488222 273454
rect 487986 272898 488222 273134
rect 487986 237218 488222 237454
rect 487986 236898 488222 237134
rect 487986 201218 488222 201454
rect 487986 200898 488222 201134
rect 487986 165218 488222 165454
rect 487986 164898 488222 165134
rect 487986 129218 488222 129454
rect 487986 128898 488222 129134
rect 487986 93218 488222 93454
rect 487986 92898 488222 93134
rect 487986 57218 488222 57454
rect 487986 56898 488222 57134
rect 487986 21218 488222 21454
rect 487986 20898 488222 21134
rect 487986 -1522 488222 -1286
rect 487986 -1842 488222 -1606
rect 491586 672818 491822 673054
rect 491586 672498 491822 672734
rect 491586 636818 491822 637054
rect 491586 636498 491822 636734
rect 491586 600818 491822 601054
rect 491586 600498 491822 600734
rect 491586 564818 491822 565054
rect 491586 564498 491822 564734
rect 491586 528818 491822 529054
rect 491586 528498 491822 528734
rect 491586 492818 491822 493054
rect 491586 492498 491822 492734
rect 491586 456818 491822 457054
rect 491586 456498 491822 456734
rect 491586 420818 491822 421054
rect 491586 420498 491822 420734
rect 491586 384818 491822 385054
rect 491586 384498 491822 384734
rect 491586 348818 491822 349054
rect 491586 348498 491822 348734
rect 491586 312818 491822 313054
rect 491586 312498 491822 312734
rect 491586 276818 491822 277054
rect 491586 276498 491822 276734
rect 491586 240818 491822 241054
rect 491586 240498 491822 240734
rect 491586 204818 491822 205054
rect 491586 204498 491822 204734
rect 491586 168818 491822 169054
rect 491586 168498 491822 168734
rect 491586 132818 491822 133054
rect 491586 132498 491822 132734
rect 491586 96818 491822 97054
rect 491586 96498 491822 96734
rect 491586 60818 491822 61054
rect 491586 60498 491822 60734
rect 491586 24818 491822 25054
rect 491586 24498 491822 24734
rect 491586 -3402 491822 -3166
rect 491586 -3722 491822 -3486
rect 495186 676418 495422 676654
rect 495186 676098 495422 676334
rect 495186 640418 495422 640654
rect 495186 640098 495422 640334
rect 495186 604418 495422 604654
rect 495186 604098 495422 604334
rect 495186 568418 495422 568654
rect 495186 568098 495422 568334
rect 495186 532418 495422 532654
rect 495186 532098 495422 532334
rect 495186 496418 495422 496654
rect 495186 496098 495422 496334
rect 495186 460418 495422 460654
rect 495186 460098 495422 460334
rect 495186 424418 495422 424654
rect 495186 424098 495422 424334
rect 495186 388418 495422 388654
rect 495186 388098 495422 388334
rect 495186 352418 495422 352654
rect 495186 352098 495422 352334
rect 495186 316418 495422 316654
rect 495186 316098 495422 316334
rect 495186 280418 495422 280654
rect 495186 280098 495422 280334
rect 495186 244418 495422 244654
rect 495186 244098 495422 244334
rect 495186 208418 495422 208654
rect 495186 208098 495422 208334
rect 495186 172418 495422 172654
rect 495186 172098 495422 172334
rect 495186 136418 495422 136654
rect 495186 136098 495422 136334
rect 495186 100418 495422 100654
rect 495186 100098 495422 100334
rect 495186 64418 495422 64654
rect 495186 64098 495422 64334
rect 495186 28418 495422 28654
rect 495186 28098 495422 28334
rect 495186 -5282 495422 -5046
rect 495186 -5602 495422 -5366
rect 516786 710242 517022 710478
rect 516786 709922 517022 710158
rect 513186 708362 513422 708598
rect 513186 708042 513422 708278
rect 509586 706482 509822 706718
rect 509586 706162 509822 706398
rect 498786 680018 499022 680254
rect 498786 679698 499022 679934
rect 498786 644018 499022 644254
rect 498786 643698 499022 643934
rect 498786 608018 499022 608254
rect 498786 607698 499022 607934
rect 498786 572018 499022 572254
rect 498786 571698 499022 571934
rect 498786 536018 499022 536254
rect 498786 535698 499022 535934
rect 498786 500018 499022 500254
rect 498786 499698 499022 499934
rect 498786 464018 499022 464254
rect 498786 463698 499022 463934
rect 498786 428018 499022 428254
rect 498786 427698 499022 427934
rect 498786 392018 499022 392254
rect 498786 391698 499022 391934
rect 498786 356018 499022 356254
rect 498786 355698 499022 355934
rect 498786 320018 499022 320254
rect 498786 319698 499022 319934
rect 498786 284018 499022 284254
rect 498786 283698 499022 283934
rect 498786 248018 499022 248254
rect 498786 247698 499022 247934
rect 498786 212018 499022 212254
rect 498786 211698 499022 211934
rect 498786 176018 499022 176254
rect 498786 175698 499022 175934
rect 498786 140018 499022 140254
rect 498786 139698 499022 139934
rect 498786 104018 499022 104254
rect 498786 103698 499022 103934
rect 498786 68018 499022 68254
rect 498786 67698 499022 67934
rect 498786 32018 499022 32254
rect 498786 31698 499022 31934
rect 480786 -6222 481022 -5986
rect 480786 -6542 481022 -6306
rect 505986 704602 506222 704838
rect 505986 704282 506222 704518
rect 505986 687218 506222 687454
rect 505986 686898 506222 687134
rect 505986 651218 506222 651454
rect 505986 650898 506222 651134
rect 505986 615218 506222 615454
rect 505986 614898 506222 615134
rect 505986 579218 506222 579454
rect 505986 578898 506222 579134
rect 505986 543218 506222 543454
rect 505986 542898 506222 543134
rect 505986 507218 506222 507454
rect 505986 506898 506222 507134
rect 505986 471218 506222 471454
rect 505986 470898 506222 471134
rect 505986 435218 506222 435454
rect 505986 434898 506222 435134
rect 505986 399218 506222 399454
rect 505986 398898 506222 399134
rect 505986 363218 506222 363454
rect 505986 362898 506222 363134
rect 505986 327218 506222 327454
rect 505986 326898 506222 327134
rect 505986 291218 506222 291454
rect 505986 290898 506222 291134
rect 505986 255218 506222 255454
rect 505986 254898 506222 255134
rect 505986 219218 506222 219454
rect 505986 218898 506222 219134
rect 505986 183218 506222 183454
rect 505986 182898 506222 183134
rect 505986 147218 506222 147454
rect 505986 146898 506222 147134
rect 505986 111218 506222 111454
rect 505986 110898 506222 111134
rect 505986 75218 506222 75454
rect 505986 74898 506222 75134
rect 505986 39218 506222 39454
rect 505986 38898 506222 39134
rect 505986 3218 506222 3454
rect 505986 2898 506222 3134
rect 505986 -582 506222 -346
rect 505986 -902 506222 -666
rect 509586 690818 509822 691054
rect 509586 690498 509822 690734
rect 509586 654818 509822 655054
rect 509586 654498 509822 654734
rect 509586 618818 509822 619054
rect 509586 618498 509822 618734
rect 509586 582818 509822 583054
rect 509586 582498 509822 582734
rect 509586 546818 509822 547054
rect 509586 546498 509822 546734
rect 509586 510818 509822 511054
rect 509586 510498 509822 510734
rect 509586 474818 509822 475054
rect 509586 474498 509822 474734
rect 509586 438818 509822 439054
rect 509586 438498 509822 438734
rect 509586 402818 509822 403054
rect 509586 402498 509822 402734
rect 509586 366818 509822 367054
rect 509586 366498 509822 366734
rect 509586 330818 509822 331054
rect 509586 330498 509822 330734
rect 509586 294818 509822 295054
rect 509586 294498 509822 294734
rect 509586 258818 509822 259054
rect 509586 258498 509822 258734
rect 509586 222818 509822 223054
rect 509586 222498 509822 222734
rect 509586 186818 509822 187054
rect 509586 186498 509822 186734
rect 509586 150818 509822 151054
rect 509586 150498 509822 150734
rect 509586 114818 509822 115054
rect 509586 114498 509822 114734
rect 509586 78818 509822 79054
rect 509586 78498 509822 78734
rect 509586 42818 509822 43054
rect 509586 42498 509822 42734
rect 509586 6818 509822 7054
rect 509586 6498 509822 6734
rect 509586 -2462 509822 -2226
rect 509586 -2782 509822 -2546
rect 513186 694418 513422 694654
rect 513186 694098 513422 694334
rect 513186 658418 513422 658654
rect 513186 658098 513422 658334
rect 513186 622418 513422 622654
rect 513186 622098 513422 622334
rect 513186 586418 513422 586654
rect 513186 586098 513422 586334
rect 513186 550418 513422 550654
rect 513186 550098 513422 550334
rect 513186 514418 513422 514654
rect 513186 514098 513422 514334
rect 513186 478418 513422 478654
rect 513186 478098 513422 478334
rect 513186 442418 513422 442654
rect 513186 442098 513422 442334
rect 513186 406418 513422 406654
rect 513186 406098 513422 406334
rect 513186 370418 513422 370654
rect 513186 370098 513422 370334
rect 513186 334418 513422 334654
rect 513186 334098 513422 334334
rect 513186 298418 513422 298654
rect 513186 298098 513422 298334
rect 513186 262418 513422 262654
rect 513186 262098 513422 262334
rect 513186 226418 513422 226654
rect 513186 226098 513422 226334
rect 513186 190418 513422 190654
rect 513186 190098 513422 190334
rect 513186 154418 513422 154654
rect 513186 154098 513422 154334
rect 513186 118418 513422 118654
rect 513186 118098 513422 118334
rect 513186 82418 513422 82654
rect 513186 82098 513422 82334
rect 513186 46418 513422 46654
rect 513186 46098 513422 46334
rect 513186 10418 513422 10654
rect 513186 10098 513422 10334
rect 513186 -4342 513422 -4106
rect 513186 -4662 513422 -4426
rect 534786 711182 535022 711418
rect 534786 710862 535022 711098
rect 531186 709302 531422 709538
rect 531186 708982 531422 709218
rect 527586 707422 527822 707658
rect 527586 707102 527822 707338
rect 516786 698018 517022 698254
rect 516786 697698 517022 697934
rect 516786 662018 517022 662254
rect 516786 661698 517022 661934
rect 516786 626018 517022 626254
rect 516786 625698 517022 625934
rect 516786 590018 517022 590254
rect 516786 589698 517022 589934
rect 516786 554018 517022 554254
rect 516786 553698 517022 553934
rect 516786 518018 517022 518254
rect 516786 517698 517022 517934
rect 516786 482018 517022 482254
rect 516786 481698 517022 481934
rect 516786 446018 517022 446254
rect 516786 445698 517022 445934
rect 516786 410018 517022 410254
rect 516786 409698 517022 409934
rect 516786 374018 517022 374254
rect 516786 373698 517022 373934
rect 516786 338018 517022 338254
rect 516786 337698 517022 337934
rect 516786 302018 517022 302254
rect 516786 301698 517022 301934
rect 516786 266018 517022 266254
rect 516786 265698 517022 265934
rect 516786 230018 517022 230254
rect 516786 229698 517022 229934
rect 516786 194018 517022 194254
rect 516786 193698 517022 193934
rect 516786 158018 517022 158254
rect 516786 157698 517022 157934
rect 516786 122018 517022 122254
rect 516786 121698 517022 121934
rect 516786 86018 517022 86254
rect 516786 85698 517022 85934
rect 516786 50018 517022 50254
rect 516786 49698 517022 49934
rect 516786 14018 517022 14254
rect 516786 13698 517022 13934
rect 498786 -7162 499022 -6926
rect 498786 -7482 499022 -7246
rect 523986 705542 524222 705778
rect 523986 705222 524222 705458
rect 523986 669218 524222 669454
rect 523986 668898 524222 669134
rect 523986 633218 524222 633454
rect 523986 632898 524222 633134
rect 523986 597218 524222 597454
rect 523986 596898 524222 597134
rect 523986 561218 524222 561454
rect 523986 560898 524222 561134
rect 523986 525218 524222 525454
rect 523986 524898 524222 525134
rect 523986 489218 524222 489454
rect 523986 488898 524222 489134
rect 523986 453218 524222 453454
rect 523986 452898 524222 453134
rect 523986 417218 524222 417454
rect 523986 416898 524222 417134
rect 523986 381218 524222 381454
rect 523986 380898 524222 381134
rect 523986 345218 524222 345454
rect 523986 344898 524222 345134
rect 523986 309218 524222 309454
rect 523986 308898 524222 309134
rect 523986 273218 524222 273454
rect 523986 272898 524222 273134
rect 523986 237218 524222 237454
rect 523986 236898 524222 237134
rect 523986 201218 524222 201454
rect 523986 200898 524222 201134
rect 523986 165218 524222 165454
rect 523986 164898 524222 165134
rect 523986 129218 524222 129454
rect 523986 128898 524222 129134
rect 523986 93218 524222 93454
rect 523986 92898 524222 93134
rect 523986 57218 524222 57454
rect 523986 56898 524222 57134
rect 523986 21218 524222 21454
rect 523986 20898 524222 21134
rect 523986 -1522 524222 -1286
rect 523986 -1842 524222 -1606
rect 527586 672818 527822 673054
rect 527586 672498 527822 672734
rect 527586 636818 527822 637054
rect 527586 636498 527822 636734
rect 527586 600818 527822 601054
rect 527586 600498 527822 600734
rect 527586 564818 527822 565054
rect 527586 564498 527822 564734
rect 527586 528818 527822 529054
rect 527586 528498 527822 528734
rect 527586 492818 527822 493054
rect 527586 492498 527822 492734
rect 527586 456818 527822 457054
rect 527586 456498 527822 456734
rect 527586 420818 527822 421054
rect 527586 420498 527822 420734
rect 527586 384818 527822 385054
rect 527586 384498 527822 384734
rect 527586 348818 527822 349054
rect 527586 348498 527822 348734
rect 527586 312818 527822 313054
rect 527586 312498 527822 312734
rect 527586 276818 527822 277054
rect 527586 276498 527822 276734
rect 527586 240818 527822 241054
rect 527586 240498 527822 240734
rect 527586 204818 527822 205054
rect 527586 204498 527822 204734
rect 527586 168818 527822 169054
rect 527586 168498 527822 168734
rect 527586 132818 527822 133054
rect 527586 132498 527822 132734
rect 527586 96818 527822 97054
rect 527586 96498 527822 96734
rect 527586 60818 527822 61054
rect 527586 60498 527822 60734
rect 527586 24818 527822 25054
rect 527586 24498 527822 24734
rect 527586 -3402 527822 -3166
rect 527586 -3722 527822 -3486
rect 531186 676418 531422 676654
rect 531186 676098 531422 676334
rect 531186 640418 531422 640654
rect 531186 640098 531422 640334
rect 531186 604418 531422 604654
rect 531186 604098 531422 604334
rect 531186 568418 531422 568654
rect 531186 568098 531422 568334
rect 531186 532418 531422 532654
rect 531186 532098 531422 532334
rect 531186 496418 531422 496654
rect 531186 496098 531422 496334
rect 531186 460418 531422 460654
rect 531186 460098 531422 460334
rect 531186 424418 531422 424654
rect 531186 424098 531422 424334
rect 531186 388418 531422 388654
rect 531186 388098 531422 388334
rect 531186 352418 531422 352654
rect 531186 352098 531422 352334
rect 531186 316418 531422 316654
rect 531186 316098 531422 316334
rect 531186 280418 531422 280654
rect 531186 280098 531422 280334
rect 531186 244418 531422 244654
rect 531186 244098 531422 244334
rect 531186 208418 531422 208654
rect 531186 208098 531422 208334
rect 531186 172418 531422 172654
rect 531186 172098 531422 172334
rect 531186 136418 531422 136654
rect 531186 136098 531422 136334
rect 531186 100418 531422 100654
rect 531186 100098 531422 100334
rect 531186 64418 531422 64654
rect 531186 64098 531422 64334
rect 531186 28418 531422 28654
rect 531186 28098 531422 28334
rect 531186 -5282 531422 -5046
rect 531186 -5602 531422 -5366
rect 552786 710242 553022 710478
rect 552786 709922 553022 710158
rect 549186 708362 549422 708598
rect 549186 708042 549422 708278
rect 545586 706482 545822 706718
rect 545586 706162 545822 706398
rect 534786 680018 535022 680254
rect 534786 679698 535022 679934
rect 534786 644018 535022 644254
rect 534786 643698 535022 643934
rect 534786 608018 535022 608254
rect 534786 607698 535022 607934
rect 534786 572018 535022 572254
rect 534786 571698 535022 571934
rect 534786 536018 535022 536254
rect 534786 535698 535022 535934
rect 534786 500018 535022 500254
rect 534786 499698 535022 499934
rect 534786 464018 535022 464254
rect 534786 463698 535022 463934
rect 534786 428018 535022 428254
rect 534786 427698 535022 427934
rect 534786 392018 535022 392254
rect 534786 391698 535022 391934
rect 534786 356018 535022 356254
rect 534786 355698 535022 355934
rect 534786 320018 535022 320254
rect 534786 319698 535022 319934
rect 534786 284018 535022 284254
rect 534786 283698 535022 283934
rect 534786 248018 535022 248254
rect 534786 247698 535022 247934
rect 534786 212018 535022 212254
rect 534786 211698 535022 211934
rect 534786 176018 535022 176254
rect 534786 175698 535022 175934
rect 534786 140018 535022 140254
rect 534786 139698 535022 139934
rect 534786 104018 535022 104254
rect 534786 103698 535022 103934
rect 534786 68018 535022 68254
rect 534786 67698 535022 67934
rect 534786 32018 535022 32254
rect 534786 31698 535022 31934
rect 516786 -6222 517022 -5986
rect 516786 -6542 517022 -6306
rect 541986 704602 542222 704838
rect 541986 704282 542222 704518
rect 541986 687218 542222 687454
rect 541986 686898 542222 687134
rect 541986 651218 542222 651454
rect 541986 650898 542222 651134
rect 541986 615218 542222 615454
rect 541986 614898 542222 615134
rect 541986 579218 542222 579454
rect 541986 578898 542222 579134
rect 541986 543218 542222 543454
rect 541986 542898 542222 543134
rect 541986 507218 542222 507454
rect 541986 506898 542222 507134
rect 541986 471218 542222 471454
rect 541986 470898 542222 471134
rect 541986 435218 542222 435454
rect 541986 434898 542222 435134
rect 541986 399218 542222 399454
rect 541986 398898 542222 399134
rect 541986 363218 542222 363454
rect 541986 362898 542222 363134
rect 541986 327218 542222 327454
rect 541986 326898 542222 327134
rect 541986 291218 542222 291454
rect 541986 290898 542222 291134
rect 541986 255218 542222 255454
rect 541986 254898 542222 255134
rect 541986 219218 542222 219454
rect 541986 218898 542222 219134
rect 541986 183218 542222 183454
rect 541986 182898 542222 183134
rect 541986 147218 542222 147454
rect 541986 146898 542222 147134
rect 541986 111218 542222 111454
rect 541986 110898 542222 111134
rect 541986 75218 542222 75454
rect 541986 74898 542222 75134
rect 541986 39218 542222 39454
rect 541986 38898 542222 39134
rect 541986 3218 542222 3454
rect 541986 2898 542222 3134
rect 541986 -582 542222 -346
rect 541986 -902 542222 -666
rect 545586 690818 545822 691054
rect 545586 690498 545822 690734
rect 545586 654818 545822 655054
rect 545586 654498 545822 654734
rect 545586 618818 545822 619054
rect 545586 618498 545822 618734
rect 545586 582818 545822 583054
rect 545586 582498 545822 582734
rect 545586 546818 545822 547054
rect 545586 546498 545822 546734
rect 545586 510818 545822 511054
rect 545586 510498 545822 510734
rect 545586 474818 545822 475054
rect 545586 474498 545822 474734
rect 545586 438818 545822 439054
rect 545586 438498 545822 438734
rect 545586 402818 545822 403054
rect 545586 402498 545822 402734
rect 545586 366818 545822 367054
rect 545586 366498 545822 366734
rect 545586 330818 545822 331054
rect 545586 330498 545822 330734
rect 545586 294818 545822 295054
rect 545586 294498 545822 294734
rect 545586 258818 545822 259054
rect 545586 258498 545822 258734
rect 545586 222818 545822 223054
rect 545586 222498 545822 222734
rect 545586 186818 545822 187054
rect 545586 186498 545822 186734
rect 545586 150818 545822 151054
rect 545586 150498 545822 150734
rect 545586 114818 545822 115054
rect 545586 114498 545822 114734
rect 545586 78818 545822 79054
rect 545586 78498 545822 78734
rect 545586 42818 545822 43054
rect 545586 42498 545822 42734
rect 545586 6818 545822 7054
rect 545586 6498 545822 6734
rect 545586 -2462 545822 -2226
rect 545586 -2782 545822 -2546
rect 549186 694418 549422 694654
rect 549186 694098 549422 694334
rect 549186 658418 549422 658654
rect 549186 658098 549422 658334
rect 549186 622418 549422 622654
rect 549186 622098 549422 622334
rect 549186 586418 549422 586654
rect 549186 586098 549422 586334
rect 549186 550418 549422 550654
rect 549186 550098 549422 550334
rect 549186 514418 549422 514654
rect 549186 514098 549422 514334
rect 549186 478418 549422 478654
rect 549186 478098 549422 478334
rect 549186 442418 549422 442654
rect 549186 442098 549422 442334
rect 549186 406418 549422 406654
rect 549186 406098 549422 406334
rect 549186 370418 549422 370654
rect 549186 370098 549422 370334
rect 549186 334418 549422 334654
rect 549186 334098 549422 334334
rect 549186 298418 549422 298654
rect 549186 298098 549422 298334
rect 549186 262418 549422 262654
rect 549186 262098 549422 262334
rect 549186 226418 549422 226654
rect 549186 226098 549422 226334
rect 549186 190418 549422 190654
rect 549186 190098 549422 190334
rect 549186 154418 549422 154654
rect 549186 154098 549422 154334
rect 549186 118418 549422 118654
rect 549186 118098 549422 118334
rect 549186 82418 549422 82654
rect 549186 82098 549422 82334
rect 549186 46418 549422 46654
rect 549186 46098 549422 46334
rect 549186 10418 549422 10654
rect 549186 10098 549422 10334
rect 549186 -4342 549422 -4106
rect 549186 -4662 549422 -4426
rect 570786 711182 571022 711418
rect 570786 710862 571022 711098
rect 567186 709302 567422 709538
rect 567186 708982 567422 709218
rect 563586 707422 563822 707658
rect 563586 707102 563822 707338
rect 552786 698018 553022 698254
rect 552786 697698 553022 697934
rect 552786 662018 553022 662254
rect 552786 661698 553022 661934
rect 552786 626018 553022 626254
rect 552786 625698 553022 625934
rect 552786 590018 553022 590254
rect 552786 589698 553022 589934
rect 552786 554018 553022 554254
rect 552786 553698 553022 553934
rect 552786 518018 553022 518254
rect 552786 517698 553022 517934
rect 552786 482018 553022 482254
rect 552786 481698 553022 481934
rect 552786 446018 553022 446254
rect 552786 445698 553022 445934
rect 552786 410018 553022 410254
rect 552786 409698 553022 409934
rect 552786 374018 553022 374254
rect 552786 373698 553022 373934
rect 552786 338018 553022 338254
rect 552786 337698 553022 337934
rect 552786 302018 553022 302254
rect 552786 301698 553022 301934
rect 552786 266018 553022 266254
rect 552786 265698 553022 265934
rect 552786 230018 553022 230254
rect 552786 229698 553022 229934
rect 552786 194018 553022 194254
rect 552786 193698 553022 193934
rect 552786 158018 553022 158254
rect 552786 157698 553022 157934
rect 552786 122018 553022 122254
rect 552786 121698 553022 121934
rect 552786 86018 553022 86254
rect 552786 85698 553022 85934
rect 552786 50018 553022 50254
rect 552786 49698 553022 49934
rect 552786 14018 553022 14254
rect 552786 13698 553022 13934
rect 534786 -7162 535022 -6926
rect 534786 -7482 535022 -7246
rect 559986 705542 560222 705778
rect 559986 705222 560222 705458
rect 559986 669218 560222 669454
rect 559986 668898 560222 669134
rect 559986 633218 560222 633454
rect 559986 632898 560222 633134
rect 559986 597218 560222 597454
rect 559986 596898 560222 597134
rect 559986 561218 560222 561454
rect 559986 560898 560222 561134
rect 559986 525218 560222 525454
rect 559986 524898 560222 525134
rect 559986 489218 560222 489454
rect 559986 488898 560222 489134
rect 559986 453218 560222 453454
rect 559986 452898 560222 453134
rect 559986 417218 560222 417454
rect 559986 416898 560222 417134
rect 559986 381218 560222 381454
rect 559986 380898 560222 381134
rect 559986 345218 560222 345454
rect 559986 344898 560222 345134
rect 559986 309218 560222 309454
rect 559986 308898 560222 309134
rect 559986 273218 560222 273454
rect 559986 272898 560222 273134
rect 559986 237218 560222 237454
rect 559986 236898 560222 237134
rect 559986 201218 560222 201454
rect 559986 200898 560222 201134
rect 559986 165218 560222 165454
rect 559986 164898 560222 165134
rect 559986 129218 560222 129454
rect 559986 128898 560222 129134
rect 559986 93218 560222 93454
rect 559986 92898 560222 93134
rect 559986 57218 560222 57454
rect 559986 56898 560222 57134
rect 559986 21218 560222 21454
rect 559986 20898 560222 21134
rect 559986 -1522 560222 -1286
rect 559986 -1842 560222 -1606
rect 563586 672818 563822 673054
rect 563586 672498 563822 672734
rect 563586 636818 563822 637054
rect 563586 636498 563822 636734
rect 563586 600818 563822 601054
rect 563586 600498 563822 600734
rect 563586 564818 563822 565054
rect 563586 564498 563822 564734
rect 563586 528818 563822 529054
rect 563586 528498 563822 528734
rect 563586 492818 563822 493054
rect 563586 492498 563822 492734
rect 563586 456818 563822 457054
rect 563586 456498 563822 456734
rect 563586 420818 563822 421054
rect 563586 420498 563822 420734
rect 563586 384818 563822 385054
rect 563586 384498 563822 384734
rect 563586 348818 563822 349054
rect 563586 348498 563822 348734
rect 563586 312818 563822 313054
rect 563586 312498 563822 312734
rect 563586 276818 563822 277054
rect 563586 276498 563822 276734
rect 563586 240818 563822 241054
rect 563586 240498 563822 240734
rect 563586 204818 563822 205054
rect 563586 204498 563822 204734
rect 563586 168818 563822 169054
rect 563586 168498 563822 168734
rect 563586 132818 563822 133054
rect 563586 132498 563822 132734
rect 563586 96818 563822 97054
rect 563586 96498 563822 96734
rect 563586 60818 563822 61054
rect 563586 60498 563822 60734
rect 563586 24818 563822 25054
rect 563586 24498 563822 24734
rect 563586 -3402 563822 -3166
rect 563586 -3722 563822 -3486
rect 567186 676418 567422 676654
rect 567186 676098 567422 676334
rect 567186 640418 567422 640654
rect 567186 640098 567422 640334
rect 567186 604418 567422 604654
rect 567186 604098 567422 604334
rect 567186 568418 567422 568654
rect 567186 568098 567422 568334
rect 567186 532418 567422 532654
rect 567186 532098 567422 532334
rect 567186 496418 567422 496654
rect 567186 496098 567422 496334
rect 567186 460418 567422 460654
rect 567186 460098 567422 460334
rect 567186 424418 567422 424654
rect 567186 424098 567422 424334
rect 567186 388418 567422 388654
rect 567186 388098 567422 388334
rect 567186 352418 567422 352654
rect 567186 352098 567422 352334
rect 567186 316418 567422 316654
rect 567186 316098 567422 316334
rect 567186 280418 567422 280654
rect 567186 280098 567422 280334
rect 567186 244418 567422 244654
rect 567186 244098 567422 244334
rect 567186 208418 567422 208654
rect 567186 208098 567422 208334
rect 567186 172418 567422 172654
rect 567186 172098 567422 172334
rect 567186 136418 567422 136654
rect 567186 136098 567422 136334
rect 567186 100418 567422 100654
rect 567186 100098 567422 100334
rect 567186 64418 567422 64654
rect 567186 64098 567422 64334
rect 567186 28418 567422 28654
rect 567186 28098 567422 28334
rect 567186 -5282 567422 -5046
rect 567186 -5602 567422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 581586 706482 581822 706718
rect 581586 706162 581822 706398
rect 570786 680018 571022 680254
rect 570786 679698 571022 679934
rect 570786 644018 571022 644254
rect 570786 643698 571022 643934
rect 570786 608018 571022 608254
rect 570786 607698 571022 607934
rect 570786 572018 571022 572254
rect 570786 571698 571022 571934
rect 570786 536018 571022 536254
rect 570786 535698 571022 535934
rect 570786 500018 571022 500254
rect 570786 499698 571022 499934
rect 570786 464018 571022 464254
rect 570786 463698 571022 463934
rect 570786 428018 571022 428254
rect 570786 427698 571022 427934
rect 570786 392018 571022 392254
rect 570786 391698 571022 391934
rect 570786 356018 571022 356254
rect 570786 355698 571022 355934
rect 570786 320018 571022 320254
rect 570786 319698 571022 319934
rect 570786 284018 571022 284254
rect 570786 283698 571022 283934
rect 570786 248018 571022 248254
rect 570786 247698 571022 247934
rect 570786 212018 571022 212254
rect 570786 211698 571022 211934
rect 570786 176018 571022 176254
rect 570786 175698 571022 175934
rect 570786 140018 571022 140254
rect 570786 139698 571022 139934
rect 570786 104018 571022 104254
rect 570786 103698 571022 103934
rect 570786 68018 571022 68254
rect 570786 67698 571022 67934
rect 570786 32018 571022 32254
rect 570786 31698 571022 31934
rect 552786 -6222 553022 -5986
rect 552786 -6542 553022 -6306
rect 577986 704602 578222 704838
rect 577986 704282 578222 704518
rect 577986 687218 578222 687454
rect 577986 686898 578222 687134
rect 577986 651218 578222 651454
rect 577986 650898 578222 651134
rect 577986 615218 578222 615454
rect 577986 614898 578222 615134
rect 577986 579218 578222 579454
rect 577986 578898 578222 579134
rect 577986 543218 578222 543454
rect 577986 542898 578222 543134
rect 577986 507218 578222 507454
rect 577986 506898 578222 507134
rect 577986 471218 578222 471454
rect 577986 470898 578222 471134
rect 577986 435218 578222 435454
rect 577986 434898 578222 435134
rect 577986 399218 578222 399454
rect 577986 398898 578222 399134
rect 577986 363218 578222 363454
rect 577986 362898 578222 363134
rect 577986 327218 578222 327454
rect 577986 326898 578222 327134
rect 577986 291218 578222 291454
rect 577986 290898 578222 291134
rect 577986 255218 578222 255454
rect 577986 254898 578222 255134
rect 577986 219218 578222 219454
rect 577986 218898 578222 219134
rect 577986 183218 578222 183454
rect 577986 182898 578222 183134
rect 577986 147218 578222 147454
rect 577986 146898 578222 147134
rect 577986 111218 578222 111454
rect 577986 110898 578222 111134
rect 577986 75218 578222 75454
rect 577986 74898 578222 75134
rect 577986 39218 578222 39454
rect 577986 38898 578222 39134
rect 577986 3218 578222 3454
rect 577986 2898 578222 3134
rect 577986 -582 578222 -346
rect 577986 -902 578222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 581586 690818 581822 691054
rect 581586 690498 581822 690734
rect 581586 654818 581822 655054
rect 581586 654498 581822 654734
rect 581586 618818 581822 619054
rect 581586 618498 581822 618734
rect 581586 582818 581822 583054
rect 581586 582498 581822 582734
rect 581586 546818 581822 547054
rect 581586 546498 581822 546734
rect 581586 510818 581822 511054
rect 581586 510498 581822 510734
rect 581586 474818 581822 475054
rect 581586 474498 581822 474734
rect 581586 438818 581822 439054
rect 581586 438498 581822 438734
rect 581586 402818 581822 403054
rect 581586 402498 581822 402734
rect 581586 366818 581822 367054
rect 581586 366498 581822 366734
rect 581586 330818 581822 331054
rect 581586 330498 581822 330734
rect 581586 294818 581822 295054
rect 581586 294498 581822 294734
rect 581586 258818 581822 259054
rect 581586 258498 581822 258734
rect 581586 222818 581822 223054
rect 581586 222498 581822 222734
rect 581586 186818 581822 187054
rect 581586 186498 581822 186734
rect 581586 150818 581822 151054
rect 581586 150498 581822 150734
rect 581586 114818 581822 115054
rect 581586 114498 581822 114734
rect 581586 78818 581822 79054
rect 581586 78498 581822 78734
rect 581586 42818 581822 43054
rect 581586 42498 581822 42734
rect 581586 6818 581822 7054
rect 581586 6498 581822 6734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 687218 585738 687454
rect 585502 686898 585738 687134
rect 585502 651218 585738 651454
rect 585502 650898 585738 651134
rect 585502 615218 585738 615454
rect 585502 614898 585738 615134
rect 585502 579218 585738 579454
rect 585502 578898 585738 579134
rect 585502 543218 585738 543454
rect 585502 542898 585738 543134
rect 585502 507218 585738 507454
rect 585502 506898 585738 507134
rect 585502 471218 585738 471454
rect 585502 470898 585738 471134
rect 585502 435218 585738 435454
rect 585502 434898 585738 435134
rect 585502 399218 585738 399454
rect 585502 398898 585738 399134
rect 585502 363218 585738 363454
rect 585502 362898 585738 363134
rect 585502 327218 585738 327454
rect 585502 326898 585738 327134
rect 585502 291218 585738 291454
rect 585502 290898 585738 291134
rect 585502 255218 585738 255454
rect 585502 254898 585738 255134
rect 585502 219218 585738 219454
rect 585502 218898 585738 219134
rect 585502 183218 585738 183454
rect 585502 182898 585738 183134
rect 585502 147218 585738 147454
rect 585502 146898 585738 147134
rect 585502 111218 585738 111454
rect 585502 110898 585738 111134
rect 585502 75218 585738 75454
rect 585502 74898 585738 75134
rect 585502 39218 585738 39454
rect 585502 38898 585738 39134
rect 585502 3218 585738 3454
rect 585502 2898 585738 3134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 669218 586678 669454
rect 586442 668898 586678 669134
rect 586442 633218 586678 633454
rect 586442 632898 586678 633134
rect 586442 597218 586678 597454
rect 586442 596898 586678 597134
rect 586442 561218 586678 561454
rect 586442 560898 586678 561134
rect 586442 525218 586678 525454
rect 586442 524898 586678 525134
rect 586442 489218 586678 489454
rect 586442 488898 586678 489134
rect 586442 453218 586678 453454
rect 586442 452898 586678 453134
rect 586442 417218 586678 417454
rect 586442 416898 586678 417134
rect 586442 381218 586678 381454
rect 586442 380898 586678 381134
rect 586442 345218 586678 345454
rect 586442 344898 586678 345134
rect 586442 309218 586678 309454
rect 586442 308898 586678 309134
rect 586442 273218 586678 273454
rect 586442 272898 586678 273134
rect 586442 237218 586678 237454
rect 586442 236898 586678 237134
rect 586442 201218 586678 201454
rect 586442 200898 586678 201134
rect 586442 165218 586678 165454
rect 586442 164898 586678 165134
rect 586442 129218 586678 129454
rect 586442 128898 586678 129134
rect 586442 93218 586678 93454
rect 586442 92898 586678 93134
rect 586442 57218 586678 57454
rect 586442 56898 586678 57134
rect 586442 21218 586678 21454
rect 586442 20898 586678 21134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 690818 587618 691054
rect 587382 690498 587618 690734
rect 587382 654818 587618 655054
rect 587382 654498 587618 654734
rect 587382 618818 587618 619054
rect 587382 618498 587618 618734
rect 587382 582818 587618 583054
rect 587382 582498 587618 582734
rect 587382 546818 587618 547054
rect 587382 546498 587618 546734
rect 587382 510818 587618 511054
rect 587382 510498 587618 510734
rect 587382 474818 587618 475054
rect 587382 474498 587618 474734
rect 587382 438818 587618 439054
rect 587382 438498 587618 438734
rect 587382 402818 587618 403054
rect 587382 402498 587618 402734
rect 587382 366818 587618 367054
rect 587382 366498 587618 366734
rect 587382 330818 587618 331054
rect 587382 330498 587618 330734
rect 587382 294818 587618 295054
rect 587382 294498 587618 294734
rect 587382 258818 587618 259054
rect 587382 258498 587618 258734
rect 587382 222818 587618 223054
rect 587382 222498 587618 222734
rect 587382 186818 587618 187054
rect 587382 186498 587618 186734
rect 587382 150818 587618 151054
rect 587382 150498 587618 150734
rect 587382 114818 587618 115054
rect 587382 114498 587618 114734
rect 587382 78818 587618 79054
rect 587382 78498 587618 78734
rect 587382 42818 587618 43054
rect 587382 42498 587618 42734
rect 587382 6818 587618 7054
rect 587382 6498 587618 6734
rect 581586 -2462 581822 -2226
rect 581586 -2782 581822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 672818 588558 673054
rect 588322 672498 588558 672734
rect 588322 636818 588558 637054
rect 588322 636498 588558 636734
rect 588322 600818 588558 601054
rect 588322 600498 588558 600734
rect 588322 564818 588558 565054
rect 588322 564498 588558 564734
rect 588322 528818 588558 529054
rect 588322 528498 588558 528734
rect 588322 492818 588558 493054
rect 588322 492498 588558 492734
rect 588322 456818 588558 457054
rect 588322 456498 588558 456734
rect 588322 420818 588558 421054
rect 588322 420498 588558 420734
rect 588322 384818 588558 385054
rect 588322 384498 588558 384734
rect 588322 348818 588558 349054
rect 588322 348498 588558 348734
rect 588322 312818 588558 313054
rect 588322 312498 588558 312734
rect 588322 276818 588558 277054
rect 588322 276498 588558 276734
rect 588322 240818 588558 241054
rect 588322 240498 588558 240734
rect 588322 204818 588558 205054
rect 588322 204498 588558 204734
rect 588322 168818 588558 169054
rect 588322 168498 588558 168734
rect 588322 132818 588558 133054
rect 588322 132498 588558 132734
rect 588322 96818 588558 97054
rect 588322 96498 588558 96734
rect 588322 60818 588558 61054
rect 588322 60498 588558 60734
rect 588322 24818 588558 25054
rect 588322 24498 588558 24734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 694418 589498 694654
rect 589262 694098 589498 694334
rect 589262 658418 589498 658654
rect 589262 658098 589498 658334
rect 589262 622418 589498 622654
rect 589262 622098 589498 622334
rect 589262 586418 589498 586654
rect 589262 586098 589498 586334
rect 589262 550418 589498 550654
rect 589262 550098 589498 550334
rect 589262 514418 589498 514654
rect 589262 514098 589498 514334
rect 589262 478418 589498 478654
rect 589262 478098 589498 478334
rect 589262 442418 589498 442654
rect 589262 442098 589498 442334
rect 589262 406418 589498 406654
rect 589262 406098 589498 406334
rect 589262 370418 589498 370654
rect 589262 370098 589498 370334
rect 589262 334418 589498 334654
rect 589262 334098 589498 334334
rect 589262 298418 589498 298654
rect 589262 298098 589498 298334
rect 589262 262418 589498 262654
rect 589262 262098 589498 262334
rect 589262 226418 589498 226654
rect 589262 226098 589498 226334
rect 589262 190418 589498 190654
rect 589262 190098 589498 190334
rect 589262 154418 589498 154654
rect 589262 154098 589498 154334
rect 589262 118418 589498 118654
rect 589262 118098 589498 118334
rect 589262 82418 589498 82654
rect 589262 82098 589498 82334
rect 589262 46418 589498 46654
rect 589262 46098 589498 46334
rect 589262 10418 589498 10654
rect 589262 10098 589498 10334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 676418 590438 676654
rect 590202 676098 590438 676334
rect 590202 640418 590438 640654
rect 590202 640098 590438 640334
rect 590202 604418 590438 604654
rect 590202 604098 590438 604334
rect 590202 568418 590438 568654
rect 590202 568098 590438 568334
rect 590202 532418 590438 532654
rect 590202 532098 590438 532334
rect 590202 496418 590438 496654
rect 590202 496098 590438 496334
rect 590202 460418 590438 460654
rect 590202 460098 590438 460334
rect 590202 424418 590438 424654
rect 590202 424098 590438 424334
rect 590202 388418 590438 388654
rect 590202 388098 590438 388334
rect 590202 352418 590438 352654
rect 590202 352098 590438 352334
rect 590202 316418 590438 316654
rect 590202 316098 590438 316334
rect 590202 280418 590438 280654
rect 590202 280098 590438 280334
rect 590202 244418 590438 244654
rect 590202 244098 590438 244334
rect 590202 208418 590438 208654
rect 590202 208098 590438 208334
rect 590202 172418 590438 172654
rect 590202 172098 590438 172334
rect 590202 136418 590438 136654
rect 590202 136098 590438 136334
rect 590202 100418 590438 100654
rect 590202 100098 590438 100334
rect 590202 64418 590438 64654
rect 590202 64098 590438 64334
rect 590202 28418 590438 28654
rect 590202 28098 590438 28334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 698018 591378 698254
rect 591142 697698 591378 697934
rect 591142 662018 591378 662254
rect 591142 661698 591378 661934
rect 591142 626018 591378 626254
rect 591142 625698 591378 625934
rect 591142 590018 591378 590254
rect 591142 589698 591378 589934
rect 591142 554018 591378 554254
rect 591142 553698 591378 553934
rect 591142 518018 591378 518254
rect 591142 517698 591378 517934
rect 591142 482018 591378 482254
rect 591142 481698 591378 481934
rect 591142 446018 591378 446254
rect 591142 445698 591378 445934
rect 591142 410018 591378 410254
rect 591142 409698 591378 409934
rect 591142 374018 591378 374254
rect 591142 373698 591378 373934
rect 591142 338018 591378 338254
rect 591142 337698 591378 337934
rect 591142 302018 591378 302254
rect 591142 301698 591378 301934
rect 591142 266018 591378 266254
rect 591142 265698 591378 265934
rect 591142 230018 591378 230254
rect 591142 229698 591378 229934
rect 591142 194018 591378 194254
rect 591142 193698 591378 193934
rect 591142 158018 591378 158254
rect 591142 157698 591378 157934
rect 591142 122018 591378 122254
rect 591142 121698 591378 121934
rect 591142 86018 591378 86254
rect 591142 85698 591378 85934
rect 591142 50018 591378 50254
rect 591142 49698 591378 49934
rect 591142 14018 591378 14254
rect 591142 13698 591378 13934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 680018 592318 680254
rect 592082 679698 592318 679934
rect 592082 644018 592318 644254
rect 592082 643698 592318 643934
rect 592082 608018 592318 608254
rect 592082 607698 592318 607934
rect 592082 572018 592318 572254
rect 592082 571698 592318 571934
rect 592082 536018 592318 536254
rect 592082 535698 592318 535934
rect 592082 500018 592318 500254
rect 592082 499698 592318 499934
rect 592082 464018 592318 464254
rect 592082 463698 592318 463934
rect 592082 428018 592318 428254
rect 592082 427698 592318 427934
rect 592082 392018 592318 392254
rect 592082 391698 592318 391934
rect 592082 356018 592318 356254
rect 592082 355698 592318 355934
rect 592082 320018 592318 320254
rect 592082 319698 592318 319934
rect 592082 284018 592318 284254
rect 592082 283698 592318 283934
rect 592082 248018 592318 248254
rect 592082 247698 592318 247934
rect 592082 212018 592318 212254
rect 592082 211698 592318 211934
rect 592082 176018 592318 176254
rect 592082 175698 592318 175934
rect 592082 140018 592318 140254
rect 592082 139698 592318 139934
rect 592082 104018 592318 104254
rect 592082 103698 592318 103934
rect 592082 68018 592318 68254
rect 592082 67698 592318 67934
rect 592082 32018 592318 32254
rect 592082 31698 592318 31934
rect 570786 -7162 571022 -6926
rect 570786 -7482 571022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 30786 711418
rect 31022 711182 66786 711418
rect 67022 711182 102786 711418
rect 103022 711182 138786 711418
rect 139022 711182 174786 711418
rect 175022 711182 210786 711418
rect 211022 711182 246786 711418
rect 247022 711182 282786 711418
rect 283022 711182 318786 711418
rect 319022 711182 354786 711418
rect 355022 711182 390786 711418
rect 391022 711182 426786 711418
rect 427022 711182 462786 711418
rect 463022 711182 498786 711418
rect 499022 711182 534786 711418
rect 535022 711182 570786 711418
rect 571022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 30786 711098
rect 31022 710862 66786 711098
rect 67022 710862 102786 711098
rect 103022 710862 138786 711098
rect 139022 710862 174786 711098
rect 175022 710862 210786 711098
rect 211022 710862 246786 711098
rect 247022 710862 282786 711098
rect 283022 710862 318786 711098
rect 319022 710862 354786 711098
rect 355022 710862 390786 711098
rect 391022 710862 426786 711098
rect 427022 710862 462786 711098
rect 463022 710862 498786 711098
rect 499022 710862 534786 711098
rect 535022 710862 570786 711098
rect 571022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 12786 710478
rect 13022 710242 48786 710478
rect 49022 710242 84786 710478
rect 85022 710242 120786 710478
rect 121022 710242 156786 710478
rect 157022 710242 192786 710478
rect 193022 710242 228786 710478
rect 229022 710242 264786 710478
rect 265022 710242 300786 710478
rect 301022 710242 336786 710478
rect 337022 710242 372786 710478
rect 373022 710242 408786 710478
rect 409022 710242 444786 710478
rect 445022 710242 480786 710478
rect 481022 710242 516786 710478
rect 517022 710242 552786 710478
rect 553022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 12786 710158
rect 13022 709922 48786 710158
rect 49022 709922 84786 710158
rect 85022 709922 120786 710158
rect 121022 709922 156786 710158
rect 157022 709922 192786 710158
rect 193022 709922 228786 710158
rect 229022 709922 264786 710158
rect 265022 709922 300786 710158
rect 301022 709922 336786 710158
rect 337022 709922 372786 710158
rect 373022 709922 408786 710158
rect 409022 709922 444786 710158
rect 445022 709922 480786 710158
rect 481022 709922 516786 710158
rect 517022 709922 552786 710158
rect 553022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 27186 709538
rect 27422 709302 63186 709538
rect 63422 709302 99186 709538
rect 99422 709302 135186 709538
rect 135422 709302 171186 709538
rect 171422 709302 207186 709538
rect 207422 709302 243186 709538
rect 243422 709302 279186 709538
rect 279422 709302 315186 709538
rect 315422 709302 351186 709538
rect 351422 709302 387186 709538
rect 387422 709302 423186 709538
rect 423422 709302 459186 709538
rect 459422 709302 495186 709538
rect 495422 709302 531186 709538
rect 531422 709302 567186 709538
rect 567422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 27186 709218
rect 27422 708982 63186 709218
rect 63422 708982 99186 709218
rect 99422 708982 135186 709218
rect 135422 708982 171186 709218
rect 171422 708982 207186 709218
rect 207422 708982 243186 709218
rect 243422 708982 279186 709218
rect 279422 708982 315186 709218
rect 315422 708982 351186 709218
rect 351422 708982 387186 709218
rect 387422 708982 423186 709218
rect 423422 708982 459186 709218
rect 459422 708982 495186 709218
rect 495422 708982 531186 709218
rect 531422 708982 567186 709218
rect 567422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 9186 708598
rect 9422 708362 45186 708598
rect 45422 708362 81186 708598
rect 81422 708362 117186 708598
rect 117422 708362 153186 708598
rect 153422 708362 189186 708598
rect 189422 708362 225186 708598
rect 225422 708362 261186 708598
rect 261422 708362 297186 708598
rect 297422 708362 333186 708598
rect 333422 708362 369186 708598
rect 369422 708362 405186 708598
rect 405422 708362 441186 708598
rect 441422 708362 477186 708598
rect 477422 708362 513186 708598
rect 513422 708362 549186 708598
rect 549422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 9186 708278
rect 9422 708042 45186 708278
rect 45422 708042 81186 708278
rect 81422 708042 117186 708278
rect 117422 708042 153186 708278
rect 153422 708042 189186 708278
rect 189422 708042 225186 708278
rect 225422 708042 261186 708278
rect 261422 708042 297186 708278
rect 297422 708042 333186 708278
rect 333422 708042 369186 708278
rect 369422 708042 405186 708278
rect 405422 708042 441186 708278
rect 441422 708042 477186 708278
rect 477422 708042 513186 708278
rect 513422 708042 549186 708278
rect 549422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 23586 707658
rect 23822 707422 59586 707658
rect 59822 707422 95586 707658
rect 95822 707422 131586 707658
rect 131822 707422 167586 707658
rect 167822 707422 203586 707658
rect 203822 707422 239586 707658
rect 239822 707422 275586 707658
rect 275822 707422 311586 707658
rect 311822 707422 347586 707658
rect 347822 707422 383586 707658
rect 383822 707422 419586 707658
rect 419822 707422 455586 707658
rect 455822 707422 491586 707658
rect 491822 707422 527586 707658
rect 527822 707422 563586 707658
rect 563822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 23586 707338
rect 23822 707102 59586 707338
rect 59822 707102 95586 707338
rect 95822 707102 131586 707338
rect 131822 707102 167586 707338
rect 167822 707102 203586 707338
rect 203822 707102 239586 707338
rect 239822 707102 275586 707338
rect 275822 707102 311586 707338
rect 311822 707102 347586 707338
rect 347822 707102 383586 707338
rect 383822 707102 419586 707338
rect 419822 707102 455586 707338
rect 455822 707102 491586 707338
rect 491822 707102 527586 707338
rect 527822 707102 563586 707338
rect 563822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 5586 706718
rect 5822 706482 41586 706718
rect 41822 706482 77586 706718
rect 77822 706482 113586 706718
rect 113822 706482 149586 706718
rect 149822 706482 185586 706718
rect 185822 706482 221586 706718
rect 221822 706482 257586 706718
rect 257822 706482 293586 706718
rect 293822 706482 329586 706718
rect 329822 706482 365586 706718
rect 365822 706482 401586 706718
rect 401822 706482 437586 706718
rect 437822 706482 473586 706718
rect 473822 706482 509586 706718
rect 509822 706482 545586 706718
rect 545822 706482 581586 706718
rect 581822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 5586 706398
rect 5822 706162 41586 706398
rect 41822 706162 77586 706398
rect 77822 706162 113586 706398
rect 113822 706162 149586 706398
rect 149822 706162 185586 706398
rect 185822 706162 221586 706398
rect 221822 706162 257586 706398
rect 257822 706162 293586 706398
rect 293822 706162 329586 706398
rect 329822 706162 365586 706398
rect 365822 706162 401586 706398
rect 401822 706162 437586 706398
rect 437822 706162 473586 706398
rect 473822 706162 509586 706398
rect 509822 706162 545586 706398
rect 545822 706162 581586 706398
rect 581822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 19986 705778
rect 20222 705542 55986 705778
rect 56222 705542 91986 705778
rect 92222 705542 127986 705778
rect 128222 705542 163986 705778
rect 164222 705542 199986 705778
rect 200222 705542 235986 705778
rect 236222 705542 271986 705778
rect 272222 705542 307986 705778
rect 308222 705542 343986 705778
rect 344222 705542 379986 705778
rect 380222 705542 415986 705778
rect 416222 705542 451986 705778
rect 452222 705542 487986 705778
rect 488222 705542 523986 705778
rect 524222 705542 559986 705778
rect 560222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 19986 705458
rect 20222 705222 55986 705458
rect 56222 705222 91986 705458
rect 92222 705222 127986 705458
rect 128222 705222 163986 705458
rect 164222 705222 199986 705458
rect 200222 705222 235986 705458
rect 236222 705222 271986 705458
rect 272222 705222 307986 705458
rect 308222 705222 343986 705458
rect 344222 705222 379986 705458
rect 380222 705222 415986 705458
rect 416222 705222 451986 705458
rect 452222 705222 487986 705458
rect 488222 705222 523986 705458
rect 524222 705222 559986 705458
rect 560222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 1986 704838
rect 2222 704602 37986 704838
rect 38222 704602 73986 704838
rect 74222 704602 109986 704838
rect 110222 704602 145986 704838
rect 146222 704602 181986 704838
rect 182222 704602 217986 704838
rect 218222 704602 253986 704838
rect 254222 704602 289986 704838
rect 290222 704602 325986 704838
rect 326222 704602 361986 704838
rect 362222 704602 397986 704838
rect 398222 704602 433986 704838
rect 434222 704602 469986 704838
rect 470222 704602 505986 704838
rect 506222 704602 541986 704838
rect 542222 704602 577986 704838
rect 578222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 1986 704518
rect 2222 704282 37986 704518
rect 38222 704282 73986 704518
rect 74222 704282 109986 704518
rect 110222 704282 145986 704518
rect 146222 704282 181986 704518
rect 182222 704282 217986 704518
rect 218222 704282 253986 704518
rect 254222 704282 289986 704518
rect 290222 704282 325986 704518
rect 326222 704282 361986 704518
rect 362222 704282 397986 704518
rect 398222 704282 433986 704518
rect 434222 704282 469986 704518
rect 470222 704282 505986 704518
rect 506222 704282 541986 704518
rect 542222 704282 577986 704518
rect 578222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect -7636 698276 -7036 698278
rect 12604 698276 13204 698278
rect 48604 698276 49204 698278
rect 84604 698276 85204 698278
rect 120604 698276 121204 698278
rect 156604 698276 157204 698278
rect 192604 698276 193204 698278
rect 228604 698276 229204 698278
rect 264604 698276 265204 698278
rect 300604 698276 301204 698278
rect 336604 698276 337204 698278
rect 372604 698276 373204 698278
rect 408604 698276 409204 698278
rect 444604 698276 445204 698278
rect 480604 698276 481204 698278
rect 516604 698276 517204 698278
rect 552604 698276 553204 698278
rect 590960 698276 591560 698278
rect -8576 698254 592500 698276
rect -8576 698018 -7454 698254
rect -7218 698018 12786 698254
rect 13022 698018 48786 698254
rect 49022 698018 84786 698254
rect 85022 698018 120786 698254
rect 121022 698018 156786 698254
rect 157022 698018 192786 698254
rect 193022 698018 228786 698254
rect 229022 698018 264786 698254
rect 265022 698018 300786 698254
rect 301022 698018 336786 698254
rect 337022 698018 372786 698254
rect 373022 698018 408786 698254
rect 409022 698018 444786 698254
rect 445022 698018 480786 698254
rect 481022 698018 516786 698254
rect 517022 698018 552786 698254
rect 553022 698018 591142 698254
rect 591378 698018 592500 698254
rect -8576 697934 592500 698018
rect -8576 697698 -7454 697934
rect -7218 697698 12786 697934
rect 13022 697698 48786 697934
rect 49022 697698 84786 697934
rect 85022 697698 120786 697934
rect 121022 697698 156786 697934
rect 157022 697698 192786 697934
rect 193022 697698 228786 697934
rect 229022 697698 264786 697934
rect 265022 697698 300786 697934
rect 301022 697698 336786 697934
rect 337022 697698 372786 697934
rect 373022 697698 408786 697934
rect 409022 697698 444786 697934
rect 445022 697698 480786 697934
rect 481022 697698 516786 697934
rect 517022 697698 552786 697934
rect 553022 697698 591142 697934
rect 591378 697698 592500 697934
rect -8576 697676 592500 697698
rect -7636 697674 -7036 697676
rect 12604 697674 13204 697676
rect 48604 697674 49204 697676
rect 84604 697674 85204 697676
rect 120604 697674 121204 697676
rect 156604 697674 157204 697676
rect 192604 697674 193204 697676
rect 228604 697674 229204 697676
rect 264604 697674 265204 697676
rect 300604 697674 301204 697676
rect 336604 697674 337204 697676
rect 372604 697674 373204 697676
rect 408604 697674 409204 697676
rect 444604 697674 445204 697676
rect 480604 697674 481204 697676
rect 516604 697674 517204 697676
rect 552604 697674 553204 697676
rect 590960 697674 591560 697676
rect -5756 694676 -5156 694678
rect 9004 694676 9604 694678
rect 45004 694676 45604 694678
rect 81004 694676 81604 694678
rect 117004 694676 117604 694678
rect 153004 694676 153604 694678
rect 189004 694676 189604 694678
rect 225004 694676 225604 694678
rect 261004 694676 261604 694678
rect 297004 694676 297604 694678
rect 333004 694676 333604 694678
rect 369004 694676 369604 694678
rect 405004 694676 405604 694678
rect 441004 694676 441604 694678
rect 477004 694676 477604 694678
rect 513004 694676 513604 694678
rect 549004 694676 549604 694678
rect 589080 694676 589680 694678
rect -6696 694654 590620 694676
rect -6696 694418 -5574 694654
rect -5338 694418 9186 694654
rect 9422 694418 45186 694654
rect 45422 694418 81186 694654
rect 81422 694418 117186 694654
rect 117422 694418 153186 694654
rect 153422 694418 189186 694654
rect 189422 694418 225186 694654
rect 225422 694418 261186 694654
rect 261422 694418 297186 694654
rect 297422 694418 333186 694654
rect 333422 694418 369186 694654
rect 369422 694418 405186 694654
rect 405422 694418 441186 694654
rect 441422 694418 477186 694654
rect 477422 694418 513186 694654
rect 513422 694418 549186 694654
rect 549422 694418 589262 694654
rect 589498 694418 590620 694654
rect -6696 694334 590620 694418
rect -6696 694098 -5574 694334
rect -5338 694098 9186 694334
rect 9422 694098 45186 694334
rect 45422 694098 81186 694334
rect 81422 694098 117186 694334
rect 117422 694098 153186 694334
rect 153422 694098 189186 694334
rect 189422 694098 225186 694334
rect 225422 694098 261186 694334
rect 261422 694098 297186 694334
rect 297422 694098 333186 694334
rect 333422 694098 369186 694334
rect 369422 694098 405186 694334
rect 405422 694098 441186 694334
rect 441422 694098 477186 694334
rect 477422 694098 513186 694334
rect 513422 694098 549186 694334
rect 549422 694098 589262 694334
rect 589498 694098 590620 694334
rect -6696 694076 590620 694098
rect -5756 694074 -5156 694076
rect 9004 694074 9604 694076
rect 45004 694074 45604 694076
rect 81004 694074 81604 694076
rect 117004 694074 117604 694076
rect 153004 694074 153604 694076
rect 189004 694074 189604 694076
rect 225004 694074 225604 694076
rect 261004 694074 261604 694076
rect 297004 694074 297604 694076
rect 333004 694074 333604 694076
rect 369004 694074 369604 694076
rect 405004 694074 405604 694076
rect 441004 694074 441604 694076
rect 477004 694074 477604 694076
rect 513004 694074 513604 694076
rect 549004 694074 549604 694076
rect 589080 694074 589680 694076
rect -3876 691076 -3276 691078
rect 5404 691076 6004 691078
rect 41404 691076 42004 691078
rect 77404 691076 78004 691078
rect 113404 691076 114004 691078
rect 149404 691076 150004 691078
rect 185404 691076 186004 691078
rect 221404 691076 222004 691078
rect 257404 691076 258004 691078
rect 293404 691076 294004 691078
rect 329404 691076 330004 691078
rect 365404 691076 366004 691078
rect 401404 691076 402004 691078
rect 437404 691076 438004 691078
rect 473404 691076 474004 691078
rect 509404 691076 510004 691078
rect 545404 691076 546004 691078
rect 581404 691076 582004 691078
rect 587200 691076 587800 691078
rect -4816 691054 588740 691076
rect -4816 690818 -3694 691054
rect -3458 690818 5586 691054
rect 5822 690818 41586 691054
rect 41822 690818 77586 691054
rect 77822 690818 113586 691054
rect 113822 690818 149586 691054
rect 149822 690818 185586 691054
rect 185822 690818 221586 691054
rect 221822 690818 257586 691054
rect 257822 690818 293586 691054
rect 293822 690818 329586 691054
rect 329822 690818 365586 691054
rect 365822 690818 401586 691054
rect 401822 690818 437586 691054
rect 437822 690818 473586 691054
rect 473822 690818 509586 691054
rect 509822 690818 545586 691054
rect 545822 690818 581586 691054
rect 581822 690818 587382 691054
rect 587618 690818 588740 691054
rect -4816 690734 588740 690818
rect -4816 690498 -3694 690734
rect -3458 690498 5586 690734
rect 5822 690498 41586 690734
rect 41822 690498 77586 690734
rect 77822 690498 113586 690734
rect 113822 690498 149586 690734
rect 149822 690498 185586 690734
rect 185822 690498 221586 690734
rect 221822 690498 257586 690734
rect 257822 690498 293586 690734
rect 293822 690498 329586 690734
rect 329822 690498 365586 690734
rect 365822 690498 401586 690734
rect 401822 690498 437586 690734
rect 437822 690498 473586 690734
rect 473822 690498 509586 690734
rect 509822 690498 545586 690734
rect 545822 690498 581586 690734
rect 581822 690498 587382 690734
rect 587618 690498 588740 690734
rect -4816 690476 588740 690498
rect -3876 690474 -3276 690476
rect 5404 690474 6004 690476
rect 41404 690474 42004 690476
rect 77404 690474 78004 690476
rect 113404 690474 114004 690476
rect 149404 690474 150004 690476
rect 185404 690474 186004 690476
rect 221404 690474 222004 690476
rect 257404 690474 258004 690476
rect 293404 690474 294004 690476
rect 329404 690474 330004 690476
rect 365404 690474 366004 690476
rect 401404 690474 402004 690476
rect 437404 690474 438004 690476
rect 473404 690474 474004 690476
rect 509404 690474 510004 690476
rect 545404 690474 546004 690476
rect 581404 690474 582004 690476
rect 587200 690474 587800 690476
rect -1996 687476 -1396 687478
rect 1804 687476 2404 687478
rect 37804 687476 38404 687478
rect 73804 687476 74404 687478
rect 109804 687476 110404 687478
rect 145804 687476 146404 687478
rect 181804 687476 182404 687478
rect 217804 687476 218404 687478
rect 253804 687476 254404 687478
rect 289804 687476 290404 687478
rect 325804 687476 326404 687478
rect 361804 687476 362404 687478
rect 397804 687476 398404 687478
rect 433804 687476 434404 687478
rect 469804 687476 470404 687478
rect 505804 687476 506404 687478
rect 541804 687476 542404 687478
rect 577804 687476 578404 687478
rect 585320 687476 585920 687478
rect -2936 687454 586860 687476
rect -2936 687218 -1814 687454
rect -1578 687218 1986 687454
rect 2222 687218 37986 687454
rect 38222 687218 73986 687454
rect 74222 687218 109986 687454
rect 110222 687218 145986 687454
rect 146222 687218 181986 687454
rect 182222 687218 217986 687454
rect 218222 687218 253986 687454
rect 254222 687218 289986 687454
rect 290222 687218 325986 687454
rect 326222 687218 361986 687454
rect 362222 687218 397986 687454
rect 398222 687218 433986 687454
rect 434222 687218 469986 687454
rect 470222 687218 505986 687454
rect 506222 687218 541986 687454
rect 542222 687218 577986 687454
rect 578222 687218 585502 687454
rect 585738 687218 586860 687454
rect -2936 687134 586860 687218
rect -2936 686898 -1814 687134
rect -1578 686898 1986 687134
rect 2222 686898 37986 687134
rect 38222 686898 73986 687134
rect 74222 686898 109986 687134
rect 110222 686898 145986 687134
rect 146222 686898 181986 687134
rect 182222 686898 217986 687134
rect 218222 686898 253986 687134
rect 254222 686898 289986 687134
rect 290222 686898 325986 687134
rect 326222 686898 361986 687134
rect 362222 686898 397986 687134
rect 398222 686898 433986 687134
rect 434222 686898 469986 687134
rect 470222 686898 505986 687134
rect 506222 686898 541986 687134
rect 542222 686898 577986 687134
rect 578222 686898 585502 687134
rect 585738 686898 586860 687134
rect -2936 686876 586860 686898
rect -1996 686874 -1396 686876
rect 1804 686874 2404 686876
rect 37804 686874 38404 686876
rect 73804 686874 74404 686876
rect 109804 686874 110404 686876
rect 145804 686874 146404 686876
rect 181804 686874 182404 686876
rect 217804 686874 218404 686876
rect 253804 686874 254404 686876
rect 289804 686874 290404 686876
rect 325804 686874 326404 686876
rect 361804 686874 362404 686876
rect 397804 686874 398404 686876
rect 433804 686874 434404 686876
rect 469804 686874 470404 686876
rect 505804 686874 506404 686876
rect 541804 686874 542404 686876
rect 577804 686874 578404 686876
rect 585320 686874 585920 686876
rect -8576 680276 -7976 680278
rect 30604 680276 31204 680278
rect 66604 680276 67204 680278
rect 102604 680276 103204 680278
rect 138604 680276 139204 680278
rect 174604 680276 175204 680278
rect 210604 680276 211204 680278
rect 246604 680276 247204 680278
rect 282604 680276 283204 680278
rect 318604 680276 319204 680278
rect 354604 680276 355204 680278
rect 390604 680276 391204 680278
rect 426604 680276 427204 680278
rect 462604 680276 463204 680278
rect 498604 680276 499204 680278
rect 534604 680276 535204 680278
rect 570604 680276 571204 680278
rect 591900 680276 592500 680278
rect -8576 680254 592500 680276
rect -8576 680018 -8394 680254
rect -8158 680018 30786 680254
rect 31022 680018 66786 680254
rect 67022 680018 102786 680254
rect 103022 680018 138786 680254
rect 139022 680018 174786 680254
rect 175022 680018 210786 680254
rect 211022 680018 246786 680254
rect 247022 680018 282786 680254
rect 283022 680018 318786 680254
rect 319022 680018 354786 680254
rect 355022 680018 390786 680254
rect 391022 680018 426786 680254
rect 427022 680018 462786 680254
rect 463022 680018 498786 680254
rect 499022 680018 534786 680254
rect 535022 680018 570786 680254
rect 571022 680018 592082 680254
rect 592318 680018 592500 680254
rect -8576 679934 592500 680018
rect -8576 679698 -8394 679934
rect -8158 679698 30786 679934
rect 31022 679698 66786 679934
rect 67022 679698 102786 679934
rect 103022 679698 138786 679934
rect 139022 679698 174786 679934
rect 175022 679698 210786 679934
rect 211022 679698 246786 679934
rect 247022 679698 282786 679934
rect 283022 679698 318786 679934
rect 319022 679698 354786 679934
rect 355022 679698 390786 679934
rect 391022 679698 426786 679934
rect 427022 679698 462786 679934
rect 463022 679698 498786 679934
rect 499022 679698 534786 679934
rect 535022 679698 570786 679934
rect 571022 679698 592082 679934
rect 592318 679698 592500 679934
rect -8576 679676 592500 679698
rect -8576 679674 -7976 679676
rect 30604 679674 31204 679676
rect 66604 679674 67204 679676
rect 102604 679674 103204 679676
rect 138604 679674 139204 679676
rect 174604 679674 175204 679676
rect 210604 679674 211204 679676
rect 246604 679674 247204 679676
rect 282604 679674 283204 679676
rect 318604 679674 319204 679676
rect 354604 679674 355204 679676
rect 390604 679674 391204 679676
rect 426604 679674 427204 679676
rect 462604 679674 463204 679676
rect 498604 679674 499204 679676
rect 534604 679674 535204 679676
rect 570604 679674 571204 679676
rect 591900 679674 592500 679676
rect -6696 676676 -6096 676678
rect 27004 676676 27604 676678
rect 63004 676676 63604 676678
rect 99004 676676 99604 676678
rect 135004 676676 135604 676678
rect 171004 676676 171604 676678
rect 207004 676676 207604 676678
rect 243004 676676 243604 676678
rect 279004 676676 279604 676678
rect 315004 676676 315604 676678
rect 351004 676676 351604 676678
rect 387004 676676 387604 676678
rect 423004 676676 423604 676678
rect 459004 676676 459604 676678
rect 495004 676676 495604 676678
rect 531004 676676 531604 676678
rect 567004 676676 567604 676678
rect 590020 676676 590620 676678
rect -6696 676654 590620 676676
rect -6696 676418 -6514 676654
rect -6278 676418 27186 676654
rect 27422 676418 63186 676654
rect 63422 676418 99186 676654
rect 99422 676418 135186 676654
rect 135422 676418 171186 676654
rect 171422 676418 207186 676654
rect 207422 676418 243186 676654
rect 243422 676418 279186 676654
rect 279422 676418 315186 676654
rect 315422 676418 351186 676654
rect 351422 676418 387186 676654
rect 387422 676418 423186 676654
rect 423422 676418 459186 676654
rect 459422 676418 495186 676654
rect 495422 676418 531186 676654
rect 531422 676418 567186 676654
rect 567422 676418 590202 676654
rect 590438 676418 590620 676654
rect -6696 676334 590620 676418
rect -6696 676098 -6514 676334
rect -6278 676098 27186 676334
rect 27422 676098 63186 676334
rect 63422 676098 99186 676334
rect 99422 676098 135186 676334
rect 135422 676098 171186 676334
rect 171422 676098 207186 676334
rect 207422 676098 243186 676334
rect 243422 676098 279186 676334
rect 279422 676098 315186 676334
rect 315422 676098 351186 676334
rect 351422 676098 387186 676334
rect 387422 676098 423186 676334
rect 423422 676098 459186 676334
rect 459422 676098 495186 676334
rect 495422 676098 531186 676334
rect 531422 676098 567186 676334
rect 567422 676098 590202 676334
rect 590438 676098 590620 676334
rect -6696 676076 590620 676098
rect -6696 676074 -6096 676076
rect 27004 676074 27604 676076
rect 63004 676074 63604 676076
rect 99004 676074 99604 676076
rect 135004 676074 135604 676076
rect 171004 676074 171604 676076
rect 207004 676074 207604 676076
rect 243004 676074 243604 676076
rect 279004 676074 279604 676076
rect 315004 676074 315604 676076
rect 351004 676074 351604 676076
rect 387004 676074 387604 676076
rect 423004 676074 423604 676076
rect 459004 676074 459604 676076
rect 495004 676074 495604 676076
rect 531004 676074 531604 676076
rect 567004 676074 567604 676076
rect 590020 676074 590620 676076
rect -4816 673076 -4216 673078
rect 23404 673076 24004 673078
rect 59404 673076 60004 673078
rect 95404 673076 96004 673078
rect 131404 673076 132004 673078
rect 167404 673076 168004 673078
rect 203404 673076 204004 673078
rect 239404 673076 240004 673078
rect 275404 673076 276004 673078
rect 311404 673076 312004 673078
rect 347404 673076 348004 673078
rect 383404 673076 384004 673078
rect 419404 673076 420004 673078
rect 455404 673076 456004 673078
rect 491404 673076 492004 673078
rect 527404 673076 528004 673078
rect 563404 673076 564004 673078
rect 588140 673076 588740 673078
rect -4816 673054 588740 673076
rect -4816 672818 -4634 673054
rect -4398 672818 23586 673054
rect 23822 672818 59586 673054
rect 59822 672818 95586 673054
rect 95822 672818 131586 673054
rect 131822 672818 167586 673054
rect 167822 672818 203586 673054
rect 203822 672818 239586 673054
rect 239822 672818 275586 673054
rect 275822 672818 311586 673054
rect 311822 672818 347586 673054
rect 347822 672818 383586 673054
rect 383822 672818 419586 673054
rect 419822 672818 455586 673054
rect 455822 672818 491586 673054
rect 491822 672818 527586 673054
rect 527822 672818 563586 673054
rect 563822 672818 588322 673054
rect 588558 672818 588740 673054
rect -4816 672734 588740 672818
rect -4816 672498 -4634 672734
rect -4398 672498 23586 672734
rect 23822 672498 59586 672734
rect 59822 672498 95586 672734
rect 95822 672498 131586 672734
rect 131822 672498 167586 672734
rect 167822 672498 203586 672734
rect 203822 672498 239586 672734
rect 239822 672498 275586 672734
rect 275822 672498 311586 672734
rect 311822 672498 347586 672734
rect 347822 672498 383586 672734
rect 383822 672498 419586 672734
rect 419822 672498 455586 672734
rect 455822 672498 491586 672734
rect 491822 672498 527586 672734
rect 527822 672498 563586 672734
rect 563822 672498 588322 672734
rect 588558 672498 588740 672734
rect -4816 672476 588740 672498
rect -4816 672474 -4216 672476
rect 23404 672474 24004 672476
rect 59404 672474 60004 672476
rect 95404 672474 96004 672476
rect 131404 672474 132004 672476
rect 167404 672474 168004 672476
rect 203404 672474 204004 672476
rect 239404 672474 240004 672476
rect 275404 672474 276004 672476
rect 311404 672474 312004 672476
rect 347404 672474 348004 672476
rect 383404 672474 384004 672476
rect 419404 672474 420004 672476
rect 455404 672474 456004 672476
rect 491404 672474 492004 672476
rect 527404 672474 528004 672476
rect 563404 672474 564004 672476
rect 588140 672474 588740 672476
rect -2936 669476 -2336 669478
rect 19804 669476 20404 669478
rect 55804 669476 56404 669478
rect 91804 669476 92404 669478
rect 127804 669476 128404 669478
rect 163804 669476 164404 669478
rect 199804 669476 200404 669478
rect 235804 669476 236404 669478
rect 271804 669476 272404 669478
rect 307804 669476 308404 669478
rect 343804 669476 344404 669478
rect 379804 669476 380404 669478
rect 415804 669476 416404 669478
rect 451804 669476 452404 669478
rect 487804 669476 488404 669478
rect 523804 669476 524404 669478
rect 559804 669476 560404 669478
rect 586260 669476 586860 669478
rect -2936 669454 586860 669476
rect -2936 669218 -2754 669454
rect -2518 669218 19986 669454
rect 20222 669218 55986 669454
rect 56222 669218 91986 669454
rect 92222 669218 127986 669454
rect 128222 669218 163986 669454
rect 164222 669218 199986 669454
rect 200222 669218 235986 669454
rect 236222 669218 271986 669454
rect 272222 669218 307986 669454
rect 308222 669218 343986 669454
rect 344222 669218 379986 669454
rect 380222 669218 415986 669454
rect 416222 669218 451986 669454
rect 452222 669218 487986 669454
rect 488222 669218 523986 669454
rect 524222 669218 559986 669454
rect 560222 669218 586442 669454
rect 586678 669218 586860 669454
rect -2936 669134 586860 669218
rect -2936 668898 -2754 669134
rect -2518 668898 19986 669134
rect 20222 668898 55986 669134
rect 56222 668898 91986 669134
rect 92222 668898 127986 669134
rect 128222 668898 163986 669134
rect 164222 668898 199986 669134
rect 200222 668898 235986 669134
rect 236222 668898 271986 669134
rect 272222 668898 307986 669134
rect 308222 668898 343986 669134
rect 344222 668898 379986 669134
rect 380222 668898 415986 669134
rect 416222 668898 451986 669134
rect 452222 668898 487986 669134
rect 488222 668898 523986 669134
rect 524222 668898 559986 669134
rect 560222 668898 586442 669134
rect 586678 668898 586860 669134
rect -2936 668876 586860 668898
rect -2936 668874 -2336 668876
rect 19804 668874 20404 668876
rect 55804 668874 56404 668876
rect 91804 668874 92404 668876
rect 127804 668874 128404 668876
rect 163804 668874 164404 668876
rect 199804 668874 200404 668876
rect 235804 668874 236404 668876
rect 271804 668874 272404 668876
rect 307804 668874 308404 668876
rect 343804 668874 344404 668876
rect 379804 668874 380404 668876
rect 415804 668874 416404 668876
rect 451804 668874 452404 668876
rect 487804 668874 488404 668876
rect 523804 668874 524404 668876
rect 559804 668874 560404 668876
rect 586260 668874 586860 668876
rect -7636 662276 -7036 662278
rect 12604 662276 13204 662278
rect 48604 662276 49204 662278
rect 84604 662276 85204 662278
rect 120604 662276 121204 662278
rect 156604 662276 157204 662278
rect 192604 662276 193204 662278
rect 228604 662276 229204 662278
rect 264604 662276 265204 662278
rect 300604 662276 301204 662278
rect 336604 662276 337204 662278
rect 372604 662276 373204 662278
rect 408604 662276 409204 662278
rect 444604 662276 445204 662278
rect 480604 662276 481204 662278
rect 516604 662276 517204 662278
rect 552604 662276 553204 662278
rect 590960 662276 591560 662278
rect -8576 662254 592500 662276
rect -8576 662018 -7454 662254
rect -7218 662018 12786 662254
rect 13022 662018 48786 662254
rect 49022 662018 84786 662254
rect 85022 662018 120786 662254
rect 121022 662018 156786 662254
rect 157022 662018 192786 662254
rect 193022 662018 228786 662254
rect 229022 662018 264786 662254
rect 265022 662018 300786 662254
rect 301022 662018 336786 662254
rect 337022 662018 372786 662254
rect 373022 662018 408786 662254
rect 409022 662018 444786 662254
rect 445022 662018 480786 662254
rect 481022 662018 516786 662254
rect 517022 662018 552786 662254
rect 553022 662018 591142 662254
rect 591378 662018 592500 662254
rect -8576 661934 592500 662018
rect -8576 661698 -7454 661934
rect -7218 661698 12786 661934
rect 13022 661698 48786 661934
rect 49022 661698 84786 661934
rect 85022 661698 120786 661934
rect 121022 661698 156786 661934
rect 157022 661698 192786 661934
rect 193022 661698 228786 661934
rect 229022 661698 264786 661934
rect 265022 661698 300786 661934
rect 301022 661698 336786 661934
rect 337022 661698 372786 661934
rect 373022 661698 408786 661934
rect 409022 661698 444786 661934
rect 445022 661698 480786 661934
rect 481022 661698 516786 661934
rect 517022 661698 552786 661934
rect 553022 661698 591142 661934
rect 591378 661698 592500 661934
rect -8576 661676 592500 661698
rect -7636 661674 -7036 661676
rect 12604 661674 13204 661676
rect 48604 661674 49204 661676
rect 84604 661674 85204 661676
rect 120604 661674 121204 661676
rect 156604 661674 157204 661676
rect 192604 661674 193204 661676
rect 228604 661674 229204 661676
rect 264604 661674 265204 661676
rect 300604 661674 301204 661676
rect 336604 661674 337204 661676
rect 372604 661674 373204 661676
rect 408604 661674 409204 661676
rect 444604 661674 445204 661676
rect 480604 661674 481204 661676
rect 516604 661674 517204 661676
rect 552604 661674 553204 661676
rect 590960 661674 591560 661676
rect -5756 658676 -5156 658678
rect 9004 658676 9604 658678
rect 45004 658676 45604 658678
rect 81004 658676 81604 658678
rect 117004 658676 117604 658678
rect 153004 658676 153604 658678
rect 189004 658676 189604 658678
rect 225004 658676 225604 658678
rect 261004 658676 261604 658678
rect 297004 658676 297604 658678
rect 333004 658676 333604 658678
rect 369004 658676 369604 658678
rect 405004 658676 405604 658678
rect 441004 658676 441604 658678
rect 477004 658676 477604 658678
rect 513004 658676 513604 658678
rect 549004 658676 549604 658678
rect 589080 658676 589680 658678
rect -6696 658654 590620 658676
rect -6696 658418 -5574 658654
rect -5338 658418 9186 658654
rect 9422 658418 45186 658654
rect 45422 658418 81186 658654
rect 81422 658418 117186 658654
rect 117422 658418 153186 658654
rect 153422 658418 189186 658654
rect 189422 658418 225186 658654
rect 225422 658418 261186 658654
rect 261422 658418 297186 658654
rect 297422 658418 333186 658654
rect 333422 658418 369186 658654
rect 369422 658418 405186 658654
rect 405422 658418 441186 658654
rect 441422 658418 477186 658654
rect 477422 658418 513186 658654
rect 513422 658418 549186 658654
rect 549422 658418 589262 658654
rect 589498 658418 590620 658654
rect -6696 658334 590620 658418
rect -6696 658098 -5574 658334
rect -5338 658098 9186 658334
rect 9422 658098 45186 658334
rect 45422 658098 81186 658334
rect 81422 658098 117186 658334
rect 117422 658098 153186 658334
rect 153422 658098 189186 658334
rect 189422 658098 225186 658334
rect 225422 658098 261186 658334
rect 261422 658098 297186 658334
rect 297422 658098 333186 658334
rect 333422 658098 369186 658334
rect 369422 658098 405186 658334
rect 405422 658098 441186 658334
rect 441422 658098 477186 658334
rect 477422 658098 513186 658334
rect 513422 658098 549186 658334
rect 549422 658098 589262 658334
rect 589498 658098 590620 658334
rect -6696 658076 590620 658098
rect -5756 658074 -5156 658076
rect 9004 658074 9604 658076
rect 45004 658074 45604 658076
rect 81004 658074 81604 658076
rect 117004 658074 117604 658076
rect 153004 658074 153604 658076
rect 189004 658074 189604 658076
rect 225004 658074 225604 658076
rect 261004 658074 261604 658076
rect 297004 658074 297604 658076
rect 333004 658074 333604 658076
rect 369004 658074 369604 658076
rect 405004 658074 405604 658076
rect 441004 658074 441604 658076
rect 477004 658074 477604 658076
rect 513004 658074 513604 658076
rect 549004 658074 549604 658076
rect 589080 658074 589680 658076
rect -3876 655076 -3276 655078
rect 5404 655076 6004 655078
rect 41404 655076 42004 655078
rect 77404 655076 78004 655078
rect 113404 655076 114004 655078
rect 149404 655076 150004 655078
rect 185404 655076 186004 655078
rect 221404 655076 222004 655078
rect 257404 655076 258004 655078
rect 293404 655076 294004 655078
rect 329404 655076 330004 655078
rect 365404 655076 366004 655078
rect 401404 655076 402004 655078
rect 437404 655076 438004 655078
rect 473404 655076 474004 655078
rect 509404 655076 510004 655078
rect 545404 655076 546004 655078
rect 581404 655076 582004 655078
rect 587200 655076 587800 655078
rect -4816 655054 588740 655076
rect -4816 654818 -3694 655054
rect -3458 654818 5586 655054
rect 5822 654818 41586 655054
rect 41822 654818 77586 655054
rect 77822 654818 113586 655054
rect 113822 654818 149586 655054
rect 149822 654818 185586 655054
rect 185822 654818 221586 655054
rect 221822 654818 257586 655054
rect 257822 654818 293586 655054
rect 293822 654818 329586 655054
rect 329822 654818 365586 655054
rect 365822 654818 401586 655054
rect 401822 654818 437586 655054
rect 437822 654818 473586 655054
rect 473822 654818 509586 655054
rect 509822 654818 545586 655054
rect 545822 654818 581586 655054
rect 581822 654818 587382 655054
rect 587618 654818 588740 655054
rect -4816 654734 588740 654818
rect -4816 654498 -3694 654734
rect -3458 654498 5586 654734
rect 5822 654498 41586 654734
rect 41822 654498 77586 654734
rect 77822 654498 113586 654734
rect 113822 654498 149586 654734
rect 149822 654498 185586 654734
rect 185822 654498 221586 654734
rect 221822 654498 257586 654734
rect 257822 654498 293586 654734
rect 293822 654498 329586 654734
rect 329822 654498 365586 654734
rect 365822 654498 401586 654734
rect 401822 654498 437586 654734
rect 437822 654498 473586 654734
rect 473822 654498 509586 654734
rect 509822 654498 545586 654734
rect 545822 654498 581586 654734
rect 581822 654498 587382 654734
rect 587618 654498 588740 654734
rect -4816 654476 588740 654498
rect -3876 654474 -3276 654476
rect 5404 654474 6004 654476
rect 41404 654474 42004 654476
rect 77404 654474 78004 654476
rect 113404 654474 114004 654476
rect 149404 654474 150004 654476
rect 185404 654474 186004 654476
rect 221404 654474 222004 654476
rect 257404 654474 258004 654476
rect 293404 654474 294004 654476
rect 329404 654474 330004 654476
rect 365404 654474 366004 654476
rect 401404 654474 402004 654476
rect 437404 654474 438004 654476
rect 473404 654474 474004 654476
rect 509404 654474 510004 654476
rect 545404 654474 546004 654476
rect 581404 654474 582004 654476
rect 587200 654474 587800 654476
rect -1996 651476 -1396 651478
rect 1804 651476 2404 651478
rect 37804 651476 38404 651478
rect 73804 651476 74404 651478
rect 109804 651476 110404 651478
rect 145804 651476 146404 651478
rect 181804 651476 182404 651478
rect 217804 651476 218404 651478
rect 253804 651476 254404 651478
rect 289804 651476 290404 651478
rect 325804 651476 326404 651478
rect 361804 651476 362404 651478
rect 397804 651476 398404 651478
rect 433804 651476 434404 651478
rect 469804 651476 470404 651478
rect 505804 651476 506404 651478
rect 541804 651476 542404 651478
rect 577804 651476 578404 651478
rect 585320 651476 585920 651478
rect -2936 651454 586860 651476
rect -2936 651218 -1814 651454
rect -1578 651218 1986 651454
rect 2222 651218 37986 651454
rect 38222 651218 73986 651454
rect 74222 651218 109986 651454
rect 110222 651218 145986 651454
rect 146222 651218 181986 651454
rect 182222 651218 217986 651454
rect 218222 651218 253986 651454
rect 254222 651218 289986 651454
rect 290222 651218 325986 651454
rect 326222 651218 361986 651454
rect 362222 651218 397986 651454
rect 398222 651218 433986 651454
rect 434222 651218 469986 651454
rect 470222 651218 505986 651454
rect 506222 651218 541986 651454
rect 542222 651218 577986 651454
rect 578222 651218 585502 651454
rect 585738 651218 586860 651454
rect -2936 651134 586860 651218
rect -2936 650898 -1814 651134
rect -1578 650898 1986 651134
rect 2222 650898 37986 651134
rect 38222 650898 73986 651134
rect 74222 650898 109986 651134
rect 110222 650898 145986 651134
rect 146222 650898 181986 651134
rect 182222 650898 217986 651134
rect 218222 650898 253986 651134
rect 254222 650898 289986 651134
rect 290222 650898 325986 651134
rect 326222 650898 361986 651134
rect 362222 650898 397986 651134
rect 398222 650898 433986 651134
rect 434222 650898 469986 651134
rect 470222 650898 505986 651134
rect 506222 650898 541986 651134
rect 542222 650898 577986 651134
rect 578222 650898 585502 651134
rect 585738 650898 586860 651134
rect -2936 650876 586860 650898
rect -1996 650874 -1396 650876
rect 1804 650874 2404 650876
rect 37804 650874 38404 650876
rect 73804 650874 74404 650876
rect 109804 650874 110404 650876
rect 145804 650874 146404 650876
rect 181804 650874 182404 650876
rect 217804 650874 218404 650876
rect 253804 650874 254404 650876
rect 289804 650874 290404 650876
rect 325804 650874 326404 650876
rect 361804 650874 362404 650876
rect 397804 650874 398404 650876
rect 433804 650874 434404 650876
rect 469804 650874 470404 650876
rect 505804 650874 506404 650876
rect 541804 650874 542404 650876
rect 577804 650874 578404 650876
rect 585320 650874 585920 650876
rect -8576 644276 -7976 644278
rect 30604 644276 31204 644278
rect 66604 644276 67204 644278
rect 102604 644276 103204 644278
rect 138604 644276 139204 644278
rect 174604 644276 175204 644278
rect 210604 644276 211204 644278
rect 246604 644276 247204 644278
rect 282604 644276 283204 644278
rect 318604 644276 319204 644278
rect 354604 644276 355204 644278
rect 390604 644276 391204 644278
rect 426604 644276 427204 644278
rect 462604 644276 463204 644278
rect 498604 644276 499204 644278
rect 534604 644276 535204 644278
rect 570604 644276 571204 644278
rect 591900 644276 592500 644278
rect -8576 644254 592500 644276
rect -8576 644018 -8394 644254
rect -8158 644018 30786 644254
rect 31022 644018 66786 644254
rect 67022 644018 102786 644254
rect 103022 644018 138786 644254
rect 139022 644018 174786 644254
rect 175022 644018 210786 644254
rect 211022 644018 246786 644254
rect 247022 644018 282786 644254
rect 283022 644018 318786 644254
rect 319022 644018 354786 644254
rect 355022 644018 390786 644254
rect 391022 644018 426786 644254
rect 427022 644018 462786 644254
rect 463022 644018 498786 644254
rect 499022 644018 534786 644254
rect 535022 644018 570786 644254
rect 571022 644018 592082 644254
rect 592318 644018 592500 644254
rect -8576 643934 592500 644018
rect -8576 643698 -8394 643934
rect -8158 643698 30786 643934
rect 31022 643698 66786 643934
rect 67022 643698 102786 643934
rect 103022 643698 138786 643934
rect 139022 643698 174786 643934
rect 175022 643698 210786 643934
rect 211022 643698 246786 643934
rect 247022 643698 282786 643934
rect 283022 643698 318786 643934
rect 319022 643698 354786 643934
rect 355022 643698 390786 643934
rect 391022 643698 426786 643934
rect 427022 643698 462786 643934
rect 463022 643698 498786 643934
rect 499022 643698 534786 643934
rect 535022 643698 570786 643934
rect 571022 643698 592082 643934
rect 592318 643698 592500 643934
rect -8576 643676 592500 643698
rect -8576 643674 -7976 643676
rect 30604 643674 31204 643676
rect 66604 643674 67204 643676
rect 102604 643674 103204 643676
rect 138604 643674 139204 643676
rect 174604 643674 175204 643676
rect 210604 643674 211204 643676
rect 246604 643674 247204 643676
rect 282604 643674 283204 643676
rect 318604 643674 319204 643676
rect 354604 643674 355204 643676
rect 390604 643674 391204 643676
rect 426604 643674 427204 643676
rect 462604 643674 463204 643676
rect 498604 643674 499204 643676
rect 534604 643674 535204 643676
rect 570604 643674 571204 643676
rect 591900 643674 592500 643676
rect -6696 640676 -6096 640678
rect 27004 640676 27604 640678
rect 63004 640676 63604 640678
rect 99004 640676 99604 640678
rect 135004 640676 135604 640678
rect 171004 640676 171604 640678
rect 207004 640676 207604 640678
rect 243004 640676 243604 640678
rect 279004 640676 279604 640678
rect 315004 640676 315604 640678
rect 351004 640676 351604 640678
rect 387004 640676 387604 640678
rect 423004 640676 423604 640678
rect 459004 640676 459604 640678
rect 495004 640676 495604 640678
rect 531004 640676 531604 640678
rect 567004 640676 567604 640678
rect 590020 640676 590620 640678
rect -6696 640654 590620 640676
rect -6696 640418 -6514 640654
rect -6278 640418 27186 640654
rect 27422 640418 63186 640654
rect 63422 640418 99186 640654
rect 99422 640418 135186 640654
rect 135422 640418 171186 640654
rect 171422 640418 207186 640654
rect 207422 640418 243186 640654
rect 243422 640418 279186 640654
rect 279422 640418 315186 640654
rect 315422 640418 351186 640654
rect 351422 640418 387186 640654
rect 387422 640418 423186 640654
rect 423422 640418 459186 640654
rect 459422 640418 495186 640654
rect 495422 640418 531186 640654
rect 531422 640418 567186 640654
rect 567422 640418 590202 640654
rect 590438 640418 590620 640654
rect -6696 640334 590620 640418
rect -6696 640098 -6514 640334
rect -6278 640098 27186 640334
rect 27422 640098 63186 640334
rect 63422 640098 99186 640334
rect 99422 640098 135186 640334
rect 135422 640098 171186 640334
rect 171422 640098 207186 640334
rect 207422 640098 243186 640334
rect 243422 640098 279186 640334
rect 279422 640098 315186 640334
rect 315422 640098 351186 640334
rect 351422 640098 387186 640334
rect 387422 640098 423186 640334
rect 423422 640098 459186 640334
rect 459422 640098 495186 640334
rect 495422 640098 531186 640334
rect 531422 640098 567186 640334
rect 567422 640098 590202 640334
rect 590438 640098 590620 640334
rect -6696 640076 590620 640098
rect -6696 640074 -6096 640076
rect 27004 640074 27604 640076
rect 63004 640074 63604 640076
rect 99004 640074 99604 640076
rect 135004 640074 135604 640076
rect 171004 640074 171604 640076
rect 207004 640074 207604 640076
rect 243004 640074 243604 640076
rect 279004 640074 279604 640076
rect 315004 640074 315604 640076
rect 351004 640074 351604 640076
rect 387004 640074 387604 640076
rect 423004 640074 423604 640076
rect 459004 640074 459604 640076
rect 495004 640074 495604 640076
rect 531004 640074 531604 640076
rect 567004 640074 567604 640076
rect 590020 640074 590620 640076
rect -4816 637076 -4216 637078
rect 23404 637076 24004 637078
rect 59404 637076 60004 637078
rect 95404 637076 96004 637078
rect 131404 637076 132004 637078
rect 167404 637076 168004 637078
rect 203404 637076 204004 637078
rect 239404 637076 240004 637078
rect 275404 637076 276004 637078
rect 311404 637076 312004 637078
rect 347404 637076 348004 637078
rect 383404 637076 384004 637078
rect 419404 637076 420004 637078
rect 455404 637076 456004 637078
rect 491404 637076 492004 637078
rect 527404 637076 528004 637078
rect 563404 637076 564004 637078
rect 588140 637076 588740 637078
rect -4816 637054 588740 637076
rect -4816 636818 -4634 637054
rect -4398 636818 23586 637054
rect 23822 636818 59586 637054
rect 59822 636818 95586 637054
rect 95822 636818 131586 637054
rect 131822 636818 167586 637054
rect 167822 636818 203586 637054
rect 203822 636818 239586 637054
rect 239822 636818 275586 637054
rect 275822 636818 311586 637054
rect 311822 636818 347586 637054
rect 347822 636818 383586 637054
rect 383822 636818 419586 637054
rect 419822 636818 455586 637054
rect 455822 636818 491586 637054
rect 491822 636818 527586 637054
rect 527822 636818 563586 637054
rect 563822 636818 588322 637054
rect 588558 636818 588740 637054
rect -4816 636734 588740 636818
rect -4816 636498 -4634 636734
rect -4398 636498 23586 636734
rect 23822 636498 59586 636734
rect 59822 636498 95586 636734
rect 95822 636498 131586 636734
rect 131822 636498 167586 636734
rect 167822 636498 203586 636734
rect 203822 636498 239586 636734
rect 239822 636498 275586 636734
rect 275822 636498 311586 636734
rect 311822 636498 347586 636734
rect 347822 636498 383586 636734
rect 383822 636498 419586 636734
rect 419822 636498 455586 636734
rect 455822 636498 491586 636734
rect 491822 636498 527586 636734
rect 527822 636498 563586 636734
rect 563822 636498 588322 636734
rect 588558 636498 588740 636734
rect -4816 636476 588740 636498
rect -4816 636474 -4216 636476
rect 23404 636474 24004 636476
rect 59404 636474 60004 636476
rect 95404 636474 96004 636476
rect 131404 636474 132004 636476
rect 167404 636474 168004 636476
rect 203404 636474 204004 636476
rect 239404 636474 240004 636476
rect 275404 636474 276004 636476
rect 311404 636474 312004 636476
rect 347404 636474 348004 636476
rect 383404 636474 384004 636476
rect 419404 636474 420004 636476
rect 455404 636474 456004 636476
rect 491404 636474 492004 636476
rect 527404 636474 528004 636476
rect 563404 636474 564004 636476
rect 588140 636474 588740 636476
rect -2936 633476 -2336 633478
rect 19804 633476 20404 633478
rect 55804 633476 56404 633478
rect 91804 633476 92404 633478
rect 127804 633476 128404 633478
rect 163804 633476 164404 633478
rect 199804 633476 200404 633478
rect 235804 633476 236404 633478
rect 271804 633476 272404 633478
rect 307804 633476 308404 633478
rect 343804 633476 344404 633478
rect 379804 633476 380404 633478
rect 415804 633476 416404 633478
rect 451804 633476 452404 633478
rect 487804 633476 488404 633478
rect 523804 633476 524404 633478
rect 559804 633476 560404 633478
rect 586260 633476 586860 633478
rect -2936 633454 586860 633476
rect -2936 633218 -2754 633454
rect -2518 633218 19986 633454
rect 20222 633218 55986 633454
rect 56222 633218 91986 633454
rect 92222 633218 127986 633454
rect 128222 633218 163986 633454
rect 164222 633218 199986 633454
rect 200222 633218 235986 633454
rect 236222 633218 271986 633454
rect 272222 633218 307986 633454
rect 308222 633218 343986 633454
rect 344222 633218 379986 633454
rect 380222 633218 415986 633454
rect 416222 633218 451986 633454
rect 452222 633218 487986 633454
rect 488222 633218 523986 633454
rect 524222 633218 559986 633454
rect 560222 633218 586442 633454
rect 586678 633218 586860 633454
rect -2936 633134 586860 633218
rect -2936 632898 -2754 633134
rect -2518 632898 19986 633134
rect 20222 632898 55986 633134
rect 56222 632898 91986 633134
rect 92222 632898 127986 633134
rect 128222 632898 163986 633134
rect 164222 632898 199986 633134
rect 200222 632898 235986 633134
rect 236222 632898 271986 633134
rect 272222 632898 307986 633134
rect 308222 632898 343986 633134
rect 344222 632898 379986 633134
rect 380222 632898 415986 633134
rect 416222 632898 451986 633134
rect 452222 632898 487986 633134
rect 488222 632898 523986 633134
rect 524222 632898 559986 633134
rect 560222 632898 586442 633134
rect 586678 632898 586860 633134
rect -2936 632876 586860 632898
rect -2936 632874 -2336 632876
rect 19804 632874 20404 632876
rect 55804 632874 56404 632876
rect 91804 632874 92404 632876
rect 127804 632874 128404 632876
rect 163804 632874 164404 632876
rect 199804 632874 200404 632876
rect 235804 632874 236404 632876
rect 271804 632874 272404 632876
rect 307804 632874 308404 632876
rect 343804 632874 344404 632876
rect 379804 632874 380404 632876
rect 415804 632874 416404 632876
rect 451804 632874 452404 632876
rect 487804 632874 488404 632876
rect 523804 632874 524404 632876
rect 559804 632874 560404 632876
rect 586260 632874 586860 632876
rect -7636 626276 -7036 626278
rect 12604 626276 13204 626278
rect 48604 626276 49204 626278
rect 84604 626276 85204 626278
rect 120604 626276 121204 626278
rect 156604 626276 157204 626278
rect 192604 626276 193204 626278
rect 228604 626276 229204 626278
rect 264604 626276 265204 626278
rect 300604 626276 301204 626278
rect 336604 626276 337204 626278
rect 372604 626276 373204 626278
rect 408604 626276 409204 626278
rect 444604 626276 445204 626278
rect 480604 626276 481204 626278
rect 516604 626276 517204 626278
rect 552604 626276 553204 626278
rect 590960 626276 591560 626278
rect -8576 626254 592500 626276
rect -8576 626018 -7454 626254
rect -7218 626018 12786 626254
rect 13022 626018 48786 626254
rect 49022 626018 84786 626254
rect 85022 626018 120786 626254
rect 121022 626018 156786 626254
rect 157022 626018 192786 626254
rect 193022 626018 228786 626254
rect 229022 626018 264786 626254
rect 265022 626018 300786 626254
rect 301022 626018 336786 626254
rect 337022 626018 372786 626254
rect 373022 626018 408786 626254
rect 409022 626018 444786 626254
rect 445022 626018 480786 626254
rect 481022 626018 516786 626254
rect 517022 626018 552786 626254
rect 553022 626018 591142 626254
rect 591378 626018 592500 626254
rect -8576 625934 592500 626018
rect -8576 625698 -7454 625934
rect -7218 625698 12786 625934
rect 13022 625698 48786 625934
rect 49022 625698 84786 625934
rect 85022 625698 120786 625934
rect 121022 625698 156786 625934
rect 157022 625698 192786 625934
rect 193022 625698 228786 625934
rect 229022 625698 264786 625934
rect 265022 625698 300786 625934
rect 301022 625698 336786 625934
rect 337022 625698 372786 625934
rect 373022 625698 408786 625934
rect 409022 625698 444786 625934
rect 445022 625698 480786 625934
rect 481022 625698 516786 625934
rect 517022 625698 552786 625934
rect 553022 625698 591142 625934
rect 591378 625698 592500 625934
rect -8576 625676 592500 625698
rect -7636 625674 -7036 625676
rect 12604 625674 13204 625676
rect 48604 625674 49204 625676
rect 84604 625674 85204 625676
rect 120604 625674 121204 625676
rect 156604 625674 157204 625676
rect 192604 625674 193204 625676
rect 228604 625674 229204 625676
rect 264604 625674 265204 625676
rect 300604 625674 301204 625676
rect 336604 625674 337204 625676
rect 372604 625674 373204 625676
rect 408604 625674 409204 625676
rect 444604 625674 445204 625676
rect 480604 625674 481204 625676
rect 516604 625674 517204 625676
rect 552604 625674 553204 625676
rect 590960 625674 591560 625676
rect -5756 622676 -5156 622678
rect 9004 622676 9604 622678
rect 45004 622676 45604 622678
rect 81004 622676 81604 622678
rect 117004 622676 117604 622678
rect 153004 622676 153604 622678
rect 189004 622676 189604 622678
rect 225004 622676 225604 622678
rect 261004 622676 261604 622678
rect 297004 622676 297604 622678
rect 333004 622676 333604 622678
rect 369004 622676 369604 622678
rect 405004 622676 405604 622678
rect 441004 622676 441604 622678
rect 477004 622676 477604 622678
rect 513004 622676 513604 622678
rect 549004 622676 549604 622678
rect 589080 622676 589680 622678
rect -6696 622654 590620 622676
rect -6696 622418 -5574 622654
rect -5338 622418 9186 622654
rect 9422 622418 45186 622654
rect 45422 622418 81186 622654
rect 81422 622418 117186 622654
rect 117422 622418 153186 622654
rect 153422 622418 189186 622654
rect 189422 622418 225186 622654
rect 225422 622418 261186 622654
rect 261422 622418 297186 622654
rect 297422 622418 333186 622654
rect 333422 622418 369186 622654
rect 369422 622418 405186 622654
rect 405422 622418 441186 622654
rect 441422 622418 477186 622654
rect 477422 622418 513186 622654
rect 513422 622418 549186 622654
rect 549422 622418 589262 622654
rect 589498 622418 590620 622654
rect -6696 622334 590620 622418
rect -6696 622098 -5574 622334
rect -5338 622098 9186 622334
rect 9422 622098 45186 622334
rect 45422 622098 81186 622334
rect 81422 622098 117186 622334
rect 117422 622098 153186 622334
rect 153422 622098 189186 622334
rect 189422 622098 225186 622334
rect 225422 622098 261186 622334
rect 261422 622098 297186 622334
rect 297422 622098 333186 622334
rect 333422 622098 369186 622334
rect 369422 622098 405186 622334
rect 405422 622098 441186 622334
rect 441422 622098 477186 622334
rect 477422 622098 513186 622334
rect 513422 622098 549186 622334
rect 549422 622098 589262 622334
rect 589498 622098 590620 622334
rect -6696 622076 590620 622098
rect -5756 622074 -5156 622076
rect 9004 622074 9604 622076
rect 45004 622074 45604 622076
rect 81004 622074 81604 622076
rect 117004 622074 117604 622076
rect 153004 622074 153604 622076
rect 189004 622074 189604 622076
rect 225004 622074 225604 622076
rect 261004 622074 261604 622076
rect 297004 622074 297604 622076
rect 333004 622074 333604 622076
rect 369004 622074 369604 622076
rect 405004 622074 405604 622076
rect 441004 622074 441604 622076
rect 477004 622074 477604 622076
rect 513004 622074 513604 622076
rect 549004 622074 549604 622076
rect 589080 622074 589680 622076
rect -3876 619076 -3276 619078
rect 5404 619076 6004 619078
rect 41404 619076 42004 619078
rect 77404 619076 78004 619078
rect 113404 619076 114004 619078
rect 149404 619076 150004 619078
rect 185404 619076 186004 619078
rect 221404 619076 222004 619078
rect 257404 619076 258004 619078
rect 293404 619076 294004 619078
rect 329404 619076 330004 619078
rect 365404 619076 366004 619078
rect 401404 619076 402004 619078
rect 437404 619076 438004 619078
rect 473404 619076 474004 619078
rect 509404 619076 510004 619078
rect 545404 619076 546004 619078
rect 581404 619076 582004 619078
rect 587200 619076 587800 619078
rect -4816 619054 588740 619076
rect -4816 618818 -3694 619054
rect -3458 618818 5586 619054
rect 5822 618818 41586 619054
rect 41822 618818 77586 619054
rect 77822 618818 113586 619054
rect 113822 618818 149586 619054
rect 149822 618818 185586 619054
rect 185822 618818 221586 619054
rect 221822 618818 257586 619054
rect 257822 618818 293586 619054
rect 293822 618818 329586 619054
rect 329822 618818 365586 619054
rect 365822 618818 401586 619054
rect 401822 618818 437586 619054
rect 437822 618818 473586 619054
rect 473822 618818 509586 619054
rect 509822 618818 545586 619054
rect 545822 618818 581586 619054
rect 581822 618818 587382 619054
rect 587618 618818 588740 619054
rect -4816 618734 588740 618818
rect -4816 618498 -3694 618734
rect -3458 618498 5586 618734
rect 5822 618498 41586 618734
rect 41822 618498 77586 618734
rect 77822 618498 113586 618734
rect 113822 618498 149586 618734
rect 149822 618498 185586 618734
rect 185822 618498 221586 618734
rect 221822 618498 257586 618734
rect 257822 618498 293586 618734
rect 293822 618498 329586 618734
rect 329822 618498 365586 618734
rect 365822 618498 401586 618734
rect 401822 618498 437586 618734
rect 437822 618498 473586 618734
rect 473822 618498 509586 618734
rect 509822 618498 545586 618734
rect 545822 618498 581586 618734
rect 581822 618498 587382 618734
rect 587618 618498 588740 618734
rect -4816 618476 588740 618498
rect -3876 618474 -3276 618476
rect 5404 618474 6004 618476
rect 41404 618474 42004 618476
rect 77404 618474 78004 618476
rect 113404 618474 114004 618476
rect 149404 618474 150004 618476
rect 185404 618474 186004 618476
rect 221404 618474 222004 618476
rect 257404 618474 258004 618476
rect 293404 618474 294004 618476
rect 329404 618474 330004 618476
rect 365404 618474 366004 618476
rect 401404 618474 402004 618476
rect 437404 618474 438004 618476
rect 473404 618474 474004 618476
rect 509404 618474 510004 618476
rect 545404 618474 546004 618476
rect 581404 618474 582004 618476
rect 587200 618474 587800 618476
rect -1996 615476 -1396 615478
rect 1804 615476 2404 615478
rect 37804 615476 38404 615478
rect 73804 615476 74404 615478
rect 109804 615476 110404 615478
rect 145804 615476 146404 615478
rect 181804 615476 182404 615478
rect 217804 615476 218404 615478
rect 253804 615476 254404 615478
rect 289804 615476 290404 615478
rect 325804 615476 326404 615478
rect 361804 615476 362404 615478
rect 397804 615476 398404 615478
rect 433804 615476 434404 615478
rect 469804 615476 470404 615478
rect 505804 615476 506404 615478
rect 541804 615476 542404 615478
rect 577804 615476 578404 615478
rect 585320 615476 585920 615478
rect -2936 615454 586860 615476
rect -2936 615218 -1814 615454
rect -1578 615218 1986 615454
rect 2222 615218 37986 615454
rect 38222 615218 73986 615454
rect 74222 615218 109986 615454
rect 110222 615218 145986 615454
rect 146222 615218 181986 615454
rect 182222 615218 217986 615454
rect 218222 615218 253986 615454
rect 254222 615218 289986 615454
rect 290222 615218 325986 615454
rect 326222 615218 361986 615454
rect 362222 615218 397986 615454
rect 398222 615218 433986 615454
rect 434222 615218 469986 615454
rect 470222 615218 505986 615454
rect 506222 615218 541986 615454
rect 542222 615218 577986 615454
rect 578222 615218 585502 615454
rect 585738 615218 586860 615454
rect -2936 615134 586860 615218
rect -2936 614898 -1814 615134
rect -1578 614898 1986 615134
rect 2222 614898 37986 615134
rect 38222 614898 73986 615134
rect 74222 614898 109986 615134
rect 110222 614898 145986 615134
rect 146222 614898 181986 615134
rect 182222 614898 217986 615134
rect 218222 614898 253986 615134
rect 254222 614898 289986 615134
rect 290222 614898 325986 615134
rect 326222 614898 361986 615134
rect 362222 614898 397986 615134
rect 398222 614898 433986 615134
rect 434222 614898 469986 615134
rect 470222 614898 505986 615134
rect 506222 614898 541986 615134
rect 542222 614898 577986 615134
rect 578222 614898 585502 615134
rect 585738 614898 586860 615134
rect -2936 614876 586860 614898
rect -1996 614874 -1396 614876
rect 1804 614874 2404 614876
rect 37804 614874 38404 614876
rect 73804 614874 74404 614876
rect 109804 614874 110404 614876
rect 145804 614874 146404 614876
rect 181804 614874 182404 614876
rect 217804 614874 218404 614876
rect 253804 614874 254404 614876
rect 289804 614874 290404 614876
rect 325804 614874 326404 614876
rect 361804 614874 362404 614876
rect 397804 614874 398404 614876
rect 433804 614874 434404 614876
rect 469804 614874 470404 614876
rect 505804 614874 506404 614876
rect 541804 614874 542404 614876
rect 577804 614874 578404 614876
rect 585320 614874 585920 614876
rect -8576 608276 -7976 608278
rect 30604 608276 31204 608278
rect 66604 608276 67204 608278
rect 102604 608276 103204 608278
rect 138604 608276 139204 608278
rect 174604 608276 175204 608278
rect 210604 608276 211204 608278
rect 246604 608276 247204 608278
rect 282604 608276 283204 608278
rect 318604 608276 319204 608278
rect 354604 608276 355204 608278
rect 390604 608276 391204 608278
rect 426604 608276 427204 608278
rect 462604 608276 463204 608278
rect 498604 608276 499204 608278
rect 534604 608276 535204 608278
rect 570604 608276 571204 608278
rect 591900 608276 592500 608278
rect -8576 608254 592500 608276
rect -8576 608018 -8394 608254
rect -8158 608018 30786 608254
rect 31022 608018 66786 608254
rect 67022 608018 102786 608254
rect 103022 608018 138786 608254
rect 139022 608018 174786 608254
rect 175022 608018 210786 608254
rect 211022 608018 246786 608254
rect 247022 608018 282786 608254
rect 283022 608018 318786 608254
rect 319022 608018 354786 608254
rect 355022 608018 390786 608254
rect 391022 608018 426786 608254
rect 427022 608018 462786 608254
rect 463022 608018 498786 608254
rect 499022 608018 534786 608254
rect 535022 608018 570786 608254
rect 571022 608018 592082 608254
rect 592318 608018 592500 608254
rect -8576 607934 592500 608018
rect -8576 607698 -8394 607934
rect -8158 607698 30786 607934
rect 31022 607698 66786 607934
rect 67022 607698 102786 607934
rect 103022 607698 138786 607934
rect 139022 607698 174786 607934
rect 175022 607698 210786 607934
rect 211022 607698 246786 607934
rect 247022 607698 282786 607934
rect 283022 607698 318786 607934
rect 319022 607698 354786 607934
rect 355022 607698 390786 607934
rect 391022 607698 426786 607934
rect 427022 607698 462786 607934
rect 463022 607698 498786 607934
rect 499022 607698 534786 607934
rect 535022 607698 570786 607934
rect 571022 607698 592082 607934
rect 592318 607698 592500 607934
rect -8576 607676 592500 607698
rect -8576 607674 -7976 607676
rect 30604 607674 31204 607676
rect 66604 607674 67204 607676
rect 102604 607674 103204 607676
rect 138604 607674 139204 607676
rect 174604 607674 175204 607676
rect 210604 607674 211204 607676
rect 246604 607674 247204 607676
rect 282604 607674 283204 607676
rect 318604 607674 319204 607676
rect 354604 607674 355204 607676
rect 390604 607674 391204 607676
rect 426604 607674 427204 607676
rect 462604 607674 463204 607676
rect 498604 607674 499204 607676
rect 534604 607674 535204 607676
rect 570604 607674 571204 607676
rect 591900 607674 592500 607676
rect -6696 604676 -6096 604678
rect 27004 604676 27604 604678
rect 63004 604676 63604 604678
rect 99004 604676 99604 604678
rect 135004 604676 135604 604678
rect 171004 604676 171604 604678
rect 207004 604676 207604 604678
rect 243004 604676 243604 604678
rect 279004 604676 279604 604678
rect 315004 604676 315604 604678
rect 351004 604676 351604 604678
rect 387004 604676 387604 604678
rect 423004 604676 423604 604678
rect 459004 604676 459604 604678
rect 495004 604676 495604 604678
rect 531004 604676 531604 604678
rect 567004 604676 567604 604678
rect 590020 604676 590620 604678
rect -6696 604654 590620 604676
rect -6696 604418 -6514 604654
rect -6278 604418 27186 604654
rect 27422 604418 63186 604654
rect 63422 604418 99186 604654
rect 99422 604418 135186 604654
rect 135422 604418 171186 604654
rect 171422 604418 207186 604654
rect 207422 604418 243186 604654
rect 243422 604418 279186 604654
rect 279422 604418 315186 604654
rect 315422 604418 351186 604654
rect 351422 604418 387186 604654
rect 387422 604418 423186 604654
rect 423422 604418 459186 604654
rect 459422 604418 495186 604654
rect 495422 604418 531186 604654
rect 531422 604418 567186 604654
rect 567422 604418 590202 604654
rect 590438 604418 590620 604654
rect -6696 604334 590620 604418
rect -6696 604098 -6514 604334
rect -6278 604098 27186 604334
rect 27422 604098 63186 604334
rect 63422 604098 99186 604334
rect 99422 604098 135186 604334
rect 135422 604098 171186 604334
rect 171422 604098 207186 604334
rect 207422 604098 243186 604334
rect 243422 604098 279186 604334
rect 279422 604098 315186 604334
rect 315422 604098 351186 604334
rect 351422 604098 387186 604334
rect 387422 604098 423186 604334
rect 423422 604098 459186 604334
rect 459422 604098 495186 604334
rect 495422 604098 531186 604334
rect 531422 604098 567186 604334
rect 567422 604098 590202 604334
rect 590438 604098 590620 604334
rect -6696 604076 590620 604098
rect -6696 604074 -6096 604076
rect 27004 604074 27604 604076
rect 63004 604074 63604 604076
rect 99004 604074 99604 604076
rect 135004 604074 135604 604076
rect 171004 604074 171604 604076
rect 207004 604074 207604 604076
rect 243004 604074 243604 604076
rect 279004 604074 279604 604076
rect 315004 604074 315604 604076
rect 351004 604074 351604 604076
rect 387004 604074 387604 604076
rect 423004 604074 423604 604076
rect 459004 604074 459604 604076
rect 495004 604074 495604 604076
rect 531004 604074 531604 604076
rect 567004 604074 567604 604076
rect 590020 604074 590620 604076
rect -4816 601076 -4216 601078
rect 23404 601076 24004 601078
rect 59404 601076 60004 601078
rect 95404 601076 96004 601078
rect 131404 601076 132004 601078
rect 167404 601076 168004 601078
rect 203404 601076 204004 601078
rect 239404 601076 240004 601078
rect 275404 601076 276004 601078
rect 311404 601076 312004 601078
rect 347404 601076 348004 601078
rect 383404 601076 384004 601078
rect 419404 601076 420004 601078
rect 455404 601076 456004 601078
rect 491404 601076 492004 601078
rect 527404 601076 528004 601078
rect 563404 601076 564004 601078
rect 588140 601076 588740 601078
rect -4816 601054 588740 601076
rect -4816 600818 -4634 601054
rect -4398 600818 23586 601054
rect 23822 600818 59586 601054
rect 59822 600818 95586 601054
rect 95822 600818 131586 601054
rect 131822 600818 167586 601054
rect 167822 600818 203586 601054
rect 203822 600818 239586 601054
rect 239822 600818 275586 601054
rect 275822 600818 311586 601054
rect 311822 600818 347586 601054
rect 347822 600818 383586 601054
rect 383822 600818 419586 601054
rect 419822 600818 455586 601054
rect 455822 600818 491586 601054
rect 491822 600818 527586 601054
rect 527822 600818 563586 601054
rect 563822 600818 588322 601054
rect 588558 600818 588740 601054
rect -4816 600734 588740 600818
rect -4816 600498 -4634 600734
rect -4398 600498 23586 600734
rect 23822 600498 59586 600734
rect 59822 600498 95586 600734
rect 95822 600498 131586 600734
rect 131822 600498 167586 600734
rect 167822 600498 203586 600734
rect 203822 600498 239586 600734
rect 239822 600498 275586 600734
rect 275822 600498 311586 600734
rect 311822 600498 347586 600734
rect 347822 600498 383586 600734
rect 383822 600498 419586 600734
rect 419822 600498 455586 600734
rect 455822 600498 491586 600734
rect 491822 600498 527586 600734
rect 527822 600498 563586 600734
rect 563822 600498 588322 600734
rect 588558 600498 588740 600734
rect -4816 600476 588740 600498
rect -4816 600474 -4216 600476
rect 23404 600474 24004 600476
rect 59404 600474 60004 600476
rect 95404 600474 96004 600476
rect 131404 600474 132004 600476
rect 167404 600474 168004 600476
rect 203404 600474 204004 600476
rect 239404 600474 240004 600476
rect 275404 600474 276004 600476
rect 311404 600474 312004 600476
rect 347404 600474 348004 600476
rect 383404 600474 384004 600476
rect 419404 600474 420004 600476
rect 455404 600474 456004 600476
rect 491404 600474 492004 600476
rect 527404 600474 528004 600476
rect 563404 600474 564004 600476
rect 588140 600474 588740 600476
rect -2936 597476 -2336 597478
rect 19804 597476 20404 597478
rect 55804 597476 56404 597478
rect 91804 597476 92404 597478
rect 127804 597476 128404 597478
rect 163804 597476 164404 597478
rect 199804 597476 200404 597478
rect 235804 597476 236404 597478
rect 271804 597476 272404 597478
rect 307804 597476 308404 597478
rect 343804 597476 344404 597478
rect 379804 597476 380404 597478
rect 415804 597476 416404 597478
rect 451804 597476 452404 597478
rect 487804 597476 488404 597478
rect 523804 597476 524404 597478
rect 559804 597476 560404 597478
rect 586260 597476 586860 597478
rect -2936 597454 586860 597476
rect -2936 597218 -2754 597454
rect -2518 597218 19986 597454
rect 20222 597218 55986 597454
rect 56222 597218 91986 597454
rect 92222 597218 127986 597454
rect 128222 597218 163986 597454
rect 164222 597218 199986 597454
rect 200222 597218 235986 597454
rect 236222 597218 271986 597454
rect 272222 597218 307986 597454
rect 308222 597218 343986 597454
rect 344222 597218 379986 597454
rect 380222 597218 415986 597454
rect 416222 597218 451986 597454
rect 452222 597218 487986 597454
rect 488222 597218 523986 597454
rect 524222 597218 559986 597454
rect 560222 597218 586442 597454
rect 586678 597218 586860 597454
rect -2936 597134 586860 597218
rect -2936 596898 -2754 597134
rect -2518 596898 19986 597134
rect 20222 596898 55986 597134
rect 56222 596898 91986 597134
rect 92222 596898 127986 597134
rect 128222 596898 163986 597134
rect 164222 596898 199986 597134
rect 200222 596898 235986 597134
rect 236222 596898 271986 597134
rect 272222 596898 307986 597134
rect 308222 596898 343986 597134
rect 344222 596898 379986 597134
rect 380222 596898 415986 597134
rect 416222 596898 451986 597134
rect 452222 596898 487986 597134
rect 488222 596898 523986 597134
rect 524222 596898 559986 597134
rect 560222 596898 586442 597134
rect 586678 596898 586860 597134
rect -2936 596876 586860 596898
rect -2936 596874 -2336 596876
rect 19804 596874 20404 596876
rect 55804 596874 56404 596876
rect 91804 596874 92404 596876
rect 127804 596874 128404 596876
rect 163804 596874 164404 596876
rect 199804 596874 200404 596876
rect 235804 596874 236404 596876
rect 271804 596874 272404 596876
rect 307804 596874 308404 596876
rect 343804 596874 344404 596876
rect 379804 596874 380404 596876
rect 415804 596874 416404 596876
rect 451804 596874 452404 596876
rect 487804 596874 488404 596876
rect 523804 596874 524404 596876
rect 559804 596874 560404 596876
rect 586260 596874 586860 596876
rect -7636 590276 -7036 590278
rect 12604 590276 13204 590278
rect 48604 590276 49204 590278
rect 84604 590276 85204 590278
rect 120604 590276 121204 590278
rect 156604 590276 157204 590278
rect 192604 590276 193204 590278
rect 228604 590276 229204 590278
rect 264604 590276 265204 590278
rect 300604 590276 301204 590278
rect 336604 590276 337204 590278
rect 372604 590276 373204 590278
rect 408604 590276 409204 590278
rect 444604 590276 445204 590278
rect 480604 590276 481204 590278
rect 516604 590276 517204 590278
rect 552604 590276 553204 590278
rect 590960 590276 591560 590278
rect -8576 590254 592500 590276
rect -8576 590018 -7454 590254
rect -7218 590018 12786 590254
rect 13022 590018 48786 590254
rect 49022 590018 84786 590254
rect 85022 590018 120786 590254
rect 121022 590018 156786 590254
rect 157022 590018 192786 590254
rect 193022 590018 228786 590254
rect 229022 590018 264786 590254
rect 265022 590018 300786 590254
rect 301022 590018 336786 590254
rect 337022 590018 372786 590254
rect 373022 590018 408786 590254
rect 409022 590018 444786 590254
rect 445022 590018 480786 590254
rect 481022 590018 516786 590254
rect 517022 590018 552786 590254
rect 553022 590018 591142 590254
rect 591378 590018 592500 590254
rect -8576 589934 592500 590018
rect -8576 589698 -7454 589934
rect -7218 589698 12786 589934
rect 13022 589698 48786 589934
rect 49022 589698 84786 589934
rect 85022 589698 120786 589934
rect 121022 589698 156786 589934
rect 157022 589698 192786 589934
rect 193022 589698 228786 589934
rect 229022 589698 264786 589934
rect 265022 589698 300786 589934
rect 301022 589698 336786 589934
rect 337022 589698 372786 589934
rect 373022 589698 408786 589934
rect 409022 589698 444786 589934
rect 445022 589698 480786 589934
rect 481022 589698 516786 589934
rect 517022 589698 552786 589934
rect 553022 589698 591142 589934
rect 591378 589698 592500 589934
rect -8576 589676 592500 589698
rect -7636 589674 -7036 589676
rect 12604 589674 13204 589676
rect 48604 589674 49204 589676
rect 84604 589674 85204 589676
rect 120604 589674 121204 589676
rect 156604 589674 157204 589676
rect 192604 589674 193204 589676
rect 228604 589674 229204 589676
rect 264604 589674 265204 589676
rect 300604 589674 301204 589676
rect 336604 589674 337204 589676
rect 372604 589674 373204 589676
rect 408604 589674 409204 589676
rect 444604 589674 445204 589676
rect 480604 589674 481204 589676
rect 516604 589674 517204 589676
rect 552604 589674 553204 589676
rect 590960 589674 591560 589676
rect -5756 586676 -5156 586678
rect 9004 586676 9604 586678
rect 45004 586676 45604 586678
rect 81004 586676 81604 586678
rect 117004 586676 117604 586678
rect 153004 586676 153604 586678
rect 189004 586676 189604 586678
rect 225004 586676 225604 586678
rect 261004 586676 261604 586678
rect 297004 586676 297604 586678
rect 333004 586676 333604 586678
rect 369004 586676 369604 586678
rect 405004 586676 405604 586678
rect 441004 586676 441604 586678
rect 477004 586676 477604 586678
rect 513004 586676 513604 586678
rect 549004 586676 549604 586678
rect 589080 586676 589680 586678
rect -6696 586654 590620 586676
rect -6696 586418 -5574 586654
rect -5338 586418 9186 586654
rect 9422 586418 45186 586654
rect 45422 586418 81186 586654
rect 81422 586418 117186 586654
rect 117422 586418 153186 586654
rect 153422 586418 189186 586654
rect 189422 586418 225186 586654
rect 225422 586418 261186 586654
rect 261422 586418 297186 586654
rect 297422 586418 333186 586654
rect 333422 586418 369186 586654
rect 369422 586418 405186 586654
rect 405422 586418 441186 586654
rect 441422 586418 477186 586654
rect 477422 586418 513186 586654
rect 513422 586418 549186 586654
rect 549422 586418 589262 586654
rect 589498 586418 590620 586654
rect -6696 586334 590620 586418
rect -6696 586098 -5574 586334
rect -5338 586098 9186 586334
rect 9422 586098 45186 586334
rect 45422 586098 81186 586334
rect 81422 586098 117186 586334
rect 117422 586098 153186 586334
rect 153422 586098 189186 586334
rect 189422 586098 225186 586334
rect 225422 586098 261186 586334
rect 261422 586098 297186 586334
rect 297422 586098 333186 586334
rect 333422 586098 369186 586334
rect 369422 586098 405186 586334
rect 405422 586098 441186 586334
rect 441422 586098 477186 586334
rect 477422 586098 513186 586334
rect 513422 586098 549186 586334
rect 549422 586098 589262 586334
rect 589498 586098 590620 586334
rect -6696 586076 590620 586098
rect -5756 586074 -5156 586076
rect 9004 586074 9604 586076
rect 45004 586074 45604 586076
rect 81004 586074 81604 586076
rect 117004 586074 117604 586076
rect 153004 586074 153604 586076
rect 189004 586074 189604 586076
rect 225004 586074 225604 586076
rect 261004 586074 261604 586076
rect 297004 586074 297604 586076
rect 333004 586074 333604 586076
rect 369004 586074 369604 586076
rect 405004 586074 405604 586076
rect 441004 586074 441604 586076
rect 477004 586074 477604 586076
rect 513004 586074 513604 586076
rect 549004 586074 549604 586076
rect 589080 586074 589680 586076
rect -3876 583076 -3276 583078
rect 5404 583076 6004 583078
rect 41404 583076 42004 583078
rect 77404 583076 78004 583078
rect 113404 583076 114004 583078
rect 149404 583076 150004 583078
rect 185404 583076 186004 583078
rect 221404 583076 222004 583078
rect 257404 583076 258004 583078
rect 293404 583076 294004 583078
rect 329404 583076 330004 583078
rect 365404 583076 366004 583078
rect 401404 583076 402004 583078
rect 437404 583076 438004 583078
rect 473404 583076 474004 583078
rect 509404 583076 510004 583078
rect 545404 583076 546004 583078
rect 581404 583076 582004 583078
rect 587200 583076 587800 583078
rect -4816 583054 588740 583076
rect -4816 582818 -3694 583054
rect -3458 582818 5586 583054
rect 5822 582818 41586 583054
rect 41822 582818 77586 583054
rect 77822 582818 113586 583054
rect 113822 582818 149586 583054
rect 149822 582818 185586 583054
rect 185822 582818 221586 583054
rect 221822 582818 257586 583054
rect 257822 582818 293586 583054
rect 293822 582818 329586 583054
rect 329822 582818 365586 583054
rect 365822 582818 401586 583054
rect 401822 582818 437586 583054
rect 437822 582818 473586 583054
rect 473822 582818 509586 583054
rect 509822 582818 545586 583054
rect 545822 582818 581586 583054
rect 581822 582818 587382 583054
rect 587618 582818 588740 583054
rect -4816 582734 588740 582818
rect -4816 582498 -3694 582734
rect -3458 582498 5586 582734
rect 5822 582498 41586 582734
rect 41822 582498 77586 582734
rect 77822 582498 113586 582734
rect 113822 582498 149586 582734
rect 149822 582498 185586 582734
rect 185822 582498 221586 582734
rect 221822 582498 257586 582734
rect 257822 582498 293586 582734
rect 293822 582498 329586 582734
rect 329822 582498 365586 582734
rect 365822 582498 401586 582734
rect 401822 582498 437586 582734
rect 437822 582498 473586 582734
rect 473822 582498 509586 582734
rect 509822 582498 545586 582734
rect 545822 582498 581586 582734
rect 581822 582498 587382 582734
rect 587618 582498 588740 582734
rect -4816 582476 588740 582498
rect -3876 582474 -3276 582476
rect 5404 582474 6004 582476
rect 41404 582474 42004 582476
rect 77404 582474 78004 582476
rect 113404 582474 114004 582476
rect 149404 582474 150004 582476
rect 185404 582474 186004 582476
rect 221404 582474 222004 582476
rect 257404 582474 258004 582476
rect 293404 582474 294004 582476
rect 329404 582474 330004 582476
rect 365404 582474 366004 582476
rect 401404 582474 402004 582476
rect 437404 582474 438004 582476
rect 473404 582474 474004 582476
rect 509404 582474 510004 582476
rect 545404 582474 546004 582476
rect 581404 582474 582004 582476
rect 587200 582474 587800 582476
rect -1996 579476 -1396 579478
rect 1804 579476 2404 579478
rect 37804 579476 38404 579478
rect 73804 579476 74404 579478
rect 109804 579476 110404 579478
rect 145804 579476 146404 579478
rect 181804 579476 182404 579478
rect 217804 579476 218404 579478
rect 253804 579476 254404 579478
rect 289804 579476 290404 579478
rect 325804 579476 326404 579478
rect 361804 579476 362404 579478
rect 397804 579476 398404 579478
rect 433804 579476 434404 579478
rect 469804 579476 470404 579478
rect 505804 579476 506404 579478
rect 541804 579476 542404 579478
rect 577804 579476 578404 579478
rect 585320 579476 585920 579478
rect -2936 579454 586860 579476
rect -2936 579218 -1814 579454
rect -1578 579218 1986 579454
rect 2222 579218 37986 579454
rect 38222 579218 73986 579454
rect 74222 579218 109986 579454
rect 110222 579218 145986 579454
rect 146222 579218 181986 579454
rect 182222 579218 217986 579454
rect 218222 579218 253986 579454
rect 254222 579218 289986 579454
rect 290222 579218 325986 579454
rect 326222 579218 361986 579454
rect 362222 579218 397986 579454
rect 398222 579218 433986 579454
rect 434222 579218 469986 579454
rect 470222 579218 505986 579454
rect 506222 579218 541986 579454
rect 542222 579218 577986 579454
rect 578222 579218 585502 579454
rect 585738 579218 586860 579454
rect -2936 579134 586860 579218
rect -2936 578898 -1814 579134
rect -1578 578898 1986 579134
rect 2222 578898 37986 579134
rect 38222 578898 73986 579134
rect 74222 578898 109986 579134
rect 110222 578898 145986 579134
rect 146222 578898 181986 579134
rect 182222 578898 217986 579134
rect 218222 578898 253986 579134
rect 254222 578898 289986 579134
rect 290222 578898 325986 579134
rect 326222 578898 361986 579134
rect 362222 578898 397986 579134
rect 398222 578898 433986 579134
rect 434222 578898 469986 579134
rect 470222 578898 505986 579134
rect 506222 578898 541986 579134
rect 542222 578898 577986 579134
rect 578222 578898 585502 579134
rect 585738 578898 586860 579134
rect -2936 578876 586860 578898
rect -1996 578874 -1396 578876
rect 1804 578874 2404 578876
rect 37804 578874 38404 578876
rect 73804 578874 74404 578876
rect 109804 578874 110404 578876
rect 145804 578874 146404 578876
rect 181804 578874 182404 578876
rect 217804 578874 218404 578876
rect 253804 578874 254404 578876
rect 289804 578874 290404 578876
rect 325804 578874 326404 578876
rect 361804 578874 362404 578876
rect 397804 578874 398404 578876
rect 433804 578874 434404 578876
rect 469804 578874 470404 578876
rect 505804 578874 506404 578876
rect 541804 578874 542404 578876
rect 577804 578874 578404 578876
rect 585320 578874 585920 578876
rect -8576 572276 -7976 572278
rect 30604 572276 31204 572278
rect 66604 572276 67204 572278
rect 102604 572276 103204 572278
rect 138604 572276 139204 572278
rect 174604 572276 175204 572278
rect 210604 572276 211204 572278
rect 246604 572276 247204 572278
rect 282604 572276 283204 572278
rect 318604 572276 319204 572278
rect 354604 572276 355204 572278
rect 390604 572276 391204 572278
rect 426604 572276 427204 572278
rect 462604 572276 463204 572278
rect 498604 572276 499204 572278
rect 534604 572276 535204 572278
rect 570604 572276 571204 572278
rect 591900 572276 592500 572278
rect -8576 572254 592500 572276
rect -8576 572018 -8394 572254
rect -8158 572018 30786 572254
rect 31022 572018 66786 572254
rect 67022 572018 102786 572254
rect 103022 572018 138786 572254
rect 139022 572018 174786 572254
rect 175022 572018 210786 572254
rect 211022 572018 246786 572254
rect 247022 572018 282786 572254
rect 283022 572018 318786 572254
rect 319022 572018 354786 572254
rect 355022 572018 390786 572254
rect 391022 572018 426786 572254
rect 427022 572018 462786 572254
rect 463022 572018 498786 572254
rect 499022 572018 534786 572254
rect 535022 572018 570786 572254
rect 571022 572018 592082 572254
rect 592318 572018 592500 572254
rect -8576 571934 592500 572018
rect -8576 571698 -8394 571934
rect -8158 571698 30786 571934
rect 31022 571698 66786 571934
rect 67022 571698 102786 571934
rect 103022 571698 138786 571934
rect 139022 571698 174786 571934
rect 175022 571698 210786 571934
rect 211022 571698 246786 571934
rect 247022 571698 282786 571934
rect 283022 571698 318786 571934
rect 319022 571698 354786 571934
rect 355022 571698 390786 571934
rect 391022 571698 426786 571934
rect 427022 571698 462786 571934
rect 463022 571698 498786 571934
rect 499022 571698 534786 571934
rect 535022 571698 570786 571934
rect 571022 571698 592082 571934
rect 592318 571698 592500 571934
rect -8576 571676 592500 571698
rect -8576 571674 -7976 571676
rect 30604 571674 31204 571676
rect 66604 571674 67204 571676
rect 102604 571674 103204 571676
rect 138604 571674 139204 571676
rect 174604 571674 175204 571676
rect 210604 571674 211204 571676
rect 246604 571674 247204 571676
rect 282604 571674 283204 571676
rect 318604 571674 319204 571676
rect 354604 571674 355204 571676
rect 390604 571674 391204 571676
rect 426604 571674 427204 571676
rect 462604 571674 463204 571676
rect 498604 571674 499204 571676
rect 534604 571674 535204 571676
rect 570604 571674 571204 571676
rect 591900 571674 592500 571676
rect -6696 568676 -6096 568678
rect 27004 568676 27604 568678
rect 63004 568676 63604 568678
rect 99004 568676 99604 568678
rect 135004 568676 135604 568678
rect 171004 568676 171604 568678
rect 207004 568676 207604 568678
rect 243004 568676 243604 568678
rect 279004 568676 279604 568678
rect 315004 568676 315604 568678
rect 351004 568676 351604 568678
rect 387004 568676 387604 568678
rect 423004 568676 423604 568678
rect 459004 568676 459604 568678
rect 495004 568676 495604 568678
rect 531004 568676 531604 568678
rect 567004 568676 567604 568678
rect 590020 568676 590620 568678
rect -6696 568654 590620 568676
rect -6696 568418 -6514 568654
rect -6278 568418 27186 568654
rect 27422 568418 63186 568654
rect 63422 568418 99186 568654
rect 99422 568418 135186 568654
rect 135422 568418 171186 568654
rect 171422 568418 207186 568654
rect 207422 568418 243186 568654
rect 243422 568418 279186 568654
rect 279422 568418 315186 568654
rect 315422 568418 351186 568654
rect 351422 568418 387186 568654
rect 387422 568418 423186 568654
rect 423422 568418 459186 568654
rect 459422 568418 495186 568654
rect 495422 568418 531186 568654
rect 531422 568418 567186 568654
rect 567422 568418 590202 568654
rect 590438 568418 590620 568654
rect -6696 568334 590620 568418
rect -6696 568098 -6514 568334
rect -6278 568098 27186 568334
rect 27422 568098 63186 568334
rect 63422 568098 99186 568334
rect 99422 568098 135186 568334
rect 135422 568098 171186 568334
rect 171422 568098 207186 568334
rect 207422 568098 243186 568334
rect 243422 568098 279186 568334
rect 279422 568098 315186 568334
rect 315422 568098 351186 568334
rect 351422 568098 387186 568334
rect 387422 568098 423186 568334
rect 423422 568098 459186 568334
rect 459422 568098 495186 568334
rect 495422 568098 531186 568334
rect 531422 568098 567186 568334
rect 567422 568098 590202 568334
rect 590438 568098 590620 568334
rect -6696 568076 590620 568098
rect -6696 568074 -6096 568076
rect 27004 568074 27604 568076
rect 63004 568074 63604 568076
rect 99004 568074 99604 568076
rect 135004 568074 135604 568076
rect 171004 568074 171604 568076
rect 207004 568074 207604 568076
rect 243004 568074 243604 568076
rect 279004 568074 279604 568076
rect 315004 568074 315604 568076
rect 351004 568074 351604 568076
rect 387004 568074 387604 568076
rect 423004 568074 423604 568076
rect 459004 568074 459604 568076
rect 495004 568074 495604 568076
rect 531004 568074 531604 568076
rect 567004 568074 567604 568076
rect 590020 568074 590620 568076
rect -4816 565076 -4216 565078
rect 23404 565076 24004 565078
rect 59404 565076 60004 565078
rect 95404 565076 96004 565078
rect 131404 565076 132004 565078
rect 167404 565076 168004 565078
rect 203404 565076 204004 565078
rect 239404 565076 240004 565078
rect 275404 565076 276004 565078
rect 311404 565076 312004 565078
rect 347404 565076 348004 565078
rect 383404 565076 384004 565078
rect 419404 565076 420004 565078
rect 455404 565076 456004 565078
rect 491404 565076 492004 565078
rect 527404 565076 528004 565078
rect 563404 565076 564004 565078
rect 588140 565076 588740 565078
rect -4816 565054 588740 565076
rect -4816 564818 -4634 565054
rect -4398 564818 23586 565054
rect 23822 564818 59586 565054
rect 59822 564818 95586 565054
rect 95822 564818 131586 565054
rect 131822 564818 167586 565054
rect 167822 564818 203586 565054
rect 203822 564818 239586 565054
rect 239822 564818 275586 565054
rect 275822 564818 311586 565054
rect 311822 564818 347586 565054
rect 347822 564818 383586 565054
rect 383822 564818 419586 565054
rect 419822 564818 455586 565054
rect 455822 564818 491586 565054
rect 491822 564818 527586 565054
rect 527822 564818 563586 565054
rect 563822 564818 588322 565054
rect 588558 564818 588740 565054
rect -4816 564734 588740 564818
rect -4816 564498 -4634 564734
rect -4398 564498 23586 564734
rect 23822 564498 59586 564734
rect 59822 564498 95586 564734
rect 95822 564498 131586 564734
rect 131822 564498 167586 564734
rect 167822 564498 203586 564734
rect 203822 564498 239586 564734
rect 239822 564498 275586 564734
rect 275822 564498 311586 564734
rect 311822 564498 347586 564734
rect 347822 564498 383586 564734
rect 383822 564498 419586 564734
rect 419822 564498 455586 564734
rect 455822 564498 491586 564734
rect 491822 564498 527586 564734
rect 527822 564498 563586 564734
rect 563822 564498 588322 564734
rect 588558 564498 588740 564734
rect -4816 564476 588740 564498
rect -4816 564474 -4216 564476
rect 23404 564474 24004 564476
rect 59404 564474 60004 564476
rect 95404 564474 96004 564476
rect 131404 564474 132004 564476
rect 167404 564474 168004 564476
rect 203404 564474 204004 564476
rect 239404 564474 240004 564476
rect 275404 564474 276004 564476
rect 311404 564474 312004 564476
rect 347404 564474 348004 564476
rect 383404 564474 384004 564476
rect 419404 564474 420004 564476
rect 455404 564474 456004 564476
rect 491404 564474 492004 564476
rect 527404 564474 528004 564476
rect 563404 564474 564004 564476
rect 588140 564474 588740 564476
rect -2936 561476 -2336 561478
rect 19804 561476 20404 561478
rect 55804 561476 56404 561478
rect 91804 561476 92404 561478
rect 127804 561476 128404 561478
rect 163804 561476 164404 561478
rect 199804 561476 200404 561478
rect 235804 561476 236404 561478
rect 271804 561476 272404 561478
rect 307804 561476 308404 561478
rect 343804 561476 344404 561478
rect 379804 561476 380404 561478
rect 415804 561476 416404 561478
rect 451804 561476 452404 561478
rect 487804 561476 488404 561478
rect 523804 561476 524404 561478
rect 559804 561476 560404 561478
rect 586260 561476 586860 561478
rect -2936 561454 586860 561476
rect -2936 561218 -2754 561454
rect -2518 561218 19986 561454
rect 20222 561218 55986 561454
rect 56222 561218 91986 561454
rect 92222 561218 127986 561454
rect 128222 561218 163986 561454
rect 164222 561218 199986 561454
rect 200222 561218 235986 561454
rect 236222 561218 271986 561454
rect 272222 561218 307986 561454
rect 308222 561218 343986 561454
rect 344222 561218 379986 561454
rect 380222 561218 415986 561454
rect 416222 561218 451986 561454
rect 452222 561218 487986 561454
rect 488222 561218 523986 561454
rect 524222 561218 559986 561454
rect 560222 561218 586442 561454
rect 586678 561218 586860 561454
rect -2936 561134 586860 561218
rect -2936 560898 -2754 561134
rect -2518 560898 19986 561134
rect 20222 560898 55986 561134
rect 56222 560898 91986 561134
rect 92222 560898 127986 561134
rect 128222 560898 163986 561134
rect 164222 560898 199986 561134
rect 200222 560898 235986 561134
rect 236222 560898 271986 561134
rect 272222 560898 307986 561134
rect 308222 560898 343986 561134
rect 344222 560898 379986 561134
rect 380222 560898 415986 561134
rect 416222 560898 451986 561134
rect 452222 560898 487986 561134
rect 488222 560898 523986 561134
rect 524222 560898 559986 561134
rect 560222 560898 586442 561134
rect 586678 560898 586860 561134
rect -2936 560876 586860 560898
rect -2936 560874 -2336 560876
rect 19804 560874 20404 560876
rect 55804 560874 56404 560876
rect 91804 560874 92404 560876
rect 127804 560874 128404 560876
rect 163804 560874 164404 560876
rect 199804 560874 200404 560876
rect 235804 560874 236404 560876
rect 271804 560874 272404 560876
rect 307804 560874 308404 560876
rect 343804 560874 344404 560876
rect 379804 560874 380404 560876
rect 415804 560874 416404 560876
rect 451804 560874 452404 560876
rect 487804 560874 488404 560876
rect 523804 560874 524404 560876
rect 559804 560874 560404 560876
rect 586260 560874 586860 560876
rect -7636 554276 -7036 554278
rect 12604 554276 13204 554278
rect 48604 554276 49204 554278
rect 84604 554276 85204 554278
rect 120604 554276 121204 554278
rect 156604 554276 157204 554278
rect 192604 554276 193204 554278
rect 228604 554276 229204 554278
rect 264604 554276 265204 554278
rect 300604 554276 301204 554278
rect 336604 554276 337204 554278
rect 372604 554276 373204 554278
rect 408604 554276 409204 554278
rect 444604 554276 445204 554278
rect 480604 554276 481204 554278
rect 516604 554276 517204 554278
rect 552604 554276 553204 554278
rect 590960 554276 591560 554278
rect -8576 554254 592500 554276
rect -8576 554018 -7454 554254
rect -7218 554018 12786 554254
rect 13022 554018 48786 554254
rect 49022 554018 84786 554254
rect 85022 554018 120786 554254
rect 121022 554018 156786 554254
rect 157022 554018 192786 554254
rect 193022 554018 228786 554254
rect 229022 554018 264786 554254
rect 265022 554018 300786 554254
rect 301022 554018 336786 554254
rect 337022 554018 372786 554254
rect 373022 554018 408786 554254
rect 409022 554018 444786 554254
rect 445022 554018 480786 554254
rect 481022 554018 516786 554254
rect 517022 554018 552786 554254
rect 553022 554018 591142 554254
rect 591378 554018 592500 554254
rect -8576 553934 592500 554018
rect -8576 553698 -7454 553934
rect -7218 553698 12786 553934
rect 13022 553698 48786 553934
rect 49022 553698 84786 553934
rect 85022 553698 120786 553934
rect 121022 553698 156786 553934
rect 157022 553698 192786 553934
rect 193022 553698 228786 553934
rect 229022 553698 264786 553934
rect 265022 553698 300786 553934
rect 301022 553698 336786 553934
rect 337022 553698 372786 553934
rect 373022 553698 408786 553934
rect 409022 553698 444786 553934
rect 445022 553698 480786 553934
rect 481022 553698 516786 553934
rect 517022 553698 552786 553934
rect 553022 553698 591142 553934
rect 591378 553698 592500 553934
rect -8576 553676 592500 553698
rect -7636 553674 -7036 553676
rect 12604 553674 13204 553676
rect 48604 553674 49204 553676
rect 84604 553674 85204 553676
rect 120604 553674 121204 553676
rect 156604 553674 157204 553676
rect 192604 553674 193204 553676
rect 228604 553674 229204 553676
rect 264604 553674 265204 553676
rect 300604 553674 301204 553676
rect 336604 553674 337204 553676
rect 372604 553674 373204 553676
rect 408604 553674 409204 553676
rect 444604 553674 445204 553676
rect 480604 553674 481204 553676
rect 516604 553674 517204 553676
rect 552604 553674 553204 553676
rect 590960 553674 591560 553676
rect -5756 550676 -5156 550678
rect 9004 550676 9604 550678
rect 45004 550676 45604 550678
rect 81004 550676 81604 550678
rect 117004 550676 117604 550678
rect 153004 550676 153604 550678
rect 189004 550676 189604 550678
rect 225004 550676 225604 550678
rect 261004 550676 261604 550678
rect 297004 550676 297604 550678
rect 333004 550676 333604 550678
rect 369004 550676 369604 550678
rect 405004 550676 405604 550678
rect 441004 550676 441604 550678
rect 477004 550676 477604 550678
rect 513004 550676 513604 550678
rect 549004 550676 549604 550678
rect 589080 550676 589680 550678
rect -6696 550654 590620 550676
rect -6696 550418 -5574 550654
rect -5338 550418 9186 550654
rect 9422 550418 45186 550654
rect 45422 550418 81186 550654
rect 81422 550418 117186 550654
rect 117422 550418 153186 550654
rect 153422 550418 189186 550654
rect 189422 550418 225186 550654
rect 225422 550418 261186 550654
rect 261422 550418 297186 550654
rect 297422 550418 333186 550654
rect 333422 550418 369186 550654
rect 369422 550418 405186 550654
rect 405422 550418 441186 550654
rect 441422 550418 477186 550654
rect 477422 550418 513186 550654
rect 513422 550418 549186 550654
rect 549422 550418 589262 550654
rect 589498 550418 590620 550654
rect -6696 550334 590620 550418
rect -6696 550098 -5574 550334
rect -5338 550098 9186 550334
rect 9422 550098 45186 550334
rect 45422 550098 81186 550334
rect 81422 550098 117186 550334
rect 117422 550098 153186 550334
rect 153422 550098 189186 550334
rect 189422 550098 225186 550334
rect 225422 550098 261186 550334
rect 261422 550098 297186 550334
rect 297422 550098 333186 550334
rect 333422 550098 369186 550334
rect 369422 550098 405186 550334
rect 405422 550098 441186 550334
rect 441422 550098 477186 550334
rect 477422 550098 513186 550334
rect 513422 550098 549186 550334
rect 549422 550098 589262 550334
rect 589498 550098 590620 550334
rect -6696 550076 590620 550098
rect -5756 550074 -5156 550076
rect 9004 550074 9604 550076
rect 45004 550074 45604 550076
rect 81004 550074 81604 550076
rect 117004 550074 117604 550076
rect 153004 550074 153604 550076
rect 189004 550074 189604 550076
rect 225004 550074 225604 550076
rect 261004 550074 261604 550076
rect 297004 550074 297604 550076
rect 333004 550074 333604 550076
rect 369004 550074 369604 550076
rect 405004 550074 405604 550076
rect 441004 550074 441604 550076
rect 477004 550074 477604 550076
rect 513004 550074 513604 550076
rect 549004 550074 549604 550076
rect 589080 550074 589680 550076
rect -3876 547076 -3276 547078
rect 5404 547076 6004 547078
rect 41404 547076 42004 547078
rect 77404 547076 78004 547078
rect 113404 547076 114004 547078
rect 149404 547076 150004 547078
rect 185404 547076 186004 547078
rect 221404 547076 222004 547078
rect 257404 547076 258004 547078
rect 293404 547076 294004 547078
rect 329404 547076 330004 547078
rect 365404 547076 366004 547078
rect 401404 547076 402004 547078
rect 437404 547076 438004 547078
rect 473404 547076 474004 547078
rect 509404 547076 510004 547078
rect 545404 547076 546004 547078
rect 581404 547076 582004 547078
rect 587200 547076 587800 547078
rect -4816 547054 588740 547076
rect -4816 546818 -3694 547054
rect -3458 546818 5586 547054
rect 5822 546818 41586 547054
rect 41822 546818 77586 547054
rect 77822 546818 113586 547054
rect 113822 546818 149586 547054
rect 149822 546818 185586 547054
rect 185822 546818 221586 547054
rect 221822 546818 257586 547054
rect 257822 546818 293586 547054
rect 293822 546818 329586 547054
rect 329822 546818 365586 547054
rect 365822 546818 401586 547054
rect 401822 546818 437586 547054
rect 437822 546818 473586 547054
rect 473822 546818 509586 547054
rect 509822 546818 545586 547054
rect 545822 546818 581586 547054
rect 581822 546818 587382 547054
rect 587618 546818 588740 547054
rect -4816 546734 588740 546818
rect -4816 546498 -3694 546734
rect -3458 546498 5586 546734
rect 5822 546498 41586 546734
rect 41822 546498 77586 546734
rect 77822 546498 113586 546734
rect 113822 546498 149586 546734
rect 149822 546498 185586 546734
rect 185822 546498 221586 546734
rect 221822 546498 257586 546734
rect 257822 546498 293586 546734
rect 293822 546498 329586 546734
rect 329822 546498 365586 546734
rect 365822 546498 401586 546734
rect 401822 546498 437586 546734
rect 437822 546498 473586 546734
rect 473822 546498 509586 546734
rect 509822 546498 545586 546734
rect 545822 546498 581586 546734
rect 581822 546498 587382 546734
rect 587618 546498 588740 546734
rect -4816 546476 588740 546498
rect -3876 546474 -3276 546476
rect 5404 546474 6004 546476
rect 41404 546474 42004 546476
rect 77404 546474 78004 546476
rect 113404 546474 114004 546476
rect 149404 546474 150004 546476
rect 185404 546474 186004 546476
rect 221404 546474 222004 546476
rect 257404 546474 258004 546476
rect 293404 546474 294004 546476
rect 329404 546474 330004 546476
rect 365404 546474 366004 546476
rect 401404 546474 402004 546476
rect 437404 546474 438004 546476
rect 473404 546474 474004 546476
rect 509404 546474 510004 546476
rect 545404 546474 546004 546476
rect 581404 546474 582004 546476
rect 587200 546474 587800 546476
rect -1996 543476 -1396 543478
rect 1804 543476 2404 543478
rect 37804 543476 38404 543478
rect 73804 543476 74404 543478
rect 109804 543476 110404 543478
rect 145804 543476 146404 543478
rect 181804 543476 182404 543478
rect 217804 543476 218404 543478
rect 253804 543476 254404 543478
rect 289804 543476 290404 543478
rect 325804 543476 326404 543478
rect 361804 543476 362404 543478
rect 397804 543476 398404 543478
rect 433804 543476 434404 543478
rect 469804 543476 470404 543478
rect 505804 543476 506404 543478
rect 541804 543476 542404 543478
rect 577804 543476 578404 543478
rect 585320 543476 585920 543478
rect -2936 543454 586860 543476
rect -2936 543218 -1814 543454
rect -1578 543218 1986 543454
rect 2222 543218 37986 543454
rect 38222 543218 73986 543454
rect 74222 543218 109986 543454
rect 110222 543218 145986 543454
rect 146222 543218 181986 543454
rect 182222 543218 217986 543454
rect 218222 543218 253986 543454
rect 254222 543218 289986 543454
rect 290222 543218 325986 543454
rect 326222 543218 361986 543454
rect 362222 543218 397986 543454
rect 398222 543218 433986 543454
rect 434222 543218 469986 543454
rect 470222 543218 505986 543454
rect 506222 543218 541986 543454
rect 542222 543218 577986 543454
rect 578222 543218 585502 543454
rect 585738 543218 586860 543454
rect -2936 543134 586860 543218
rect -2936 542898 -1814 543134
rect -1578 542898 1986 543134
rect 2222 542898 37986 543134
rect 38222 542898 73986 543134
rect 74222 542898 109986 543134
rect 110222 542898 145986 543134
rect 146222 542898 181986 543134
rect 182222 542898 217986 543134
rect 218222 542898 253986 543134
rect 254222 542898 289986 543134
rect 290222 542898 325986 543134
rect 326222 542898 361986 543134
rect 362222 542898 397986 543134
rect 398222 542898 433986 543134
rect 434222 542898 469986 543134
rect 470222 542898 505986 543134
rect 506222 542898 541986 543134
rect 542222 542898 577986 543134
rect 578222 542898 585502 543134
rect 585738 542898 586860 543134
rect -2936 542876 586860 542898
rect -1996 542874 -1396 542876
rect 1804 542874 2404 542876
rect 37804 542874 38404 542876
rect 73804 542874 74404 542876
rect 109804 542874 110404 542876
rect 145804 542874 146404 542876
rect 181804 542874 182404 542876
rect 217804 542874 218404 542876
rect 253804 542874 254404 542876
rect 289804 542874 290404 542876
rect 325804 542874 326404 542876
rect 361804 542874 362404 542876
rect 397804 542874 398404 542876
rect 433804 542874 434404 542876
rect 469804 542874 470404 542876
rect 505804 542874 506404 542876
rect 541804 542874 542404 542876
rect 577804 542874 578404 542876
rect 585320 542874 585920 542876
rect -8576 536276 -7976 536278
rect 30604 536276 31204 536278
rect 66604 536276 67204 536278
rect 102604 536276 103204 536278
rect 138604 536276 139204 536278
rect 174604 536276 175204 536278
rect 210604 536276 211204 536278
rect 246604 536276 247204 536278
rect 282604 536276 283204 536278
rect 318604 536276 319204 536278
rect 354604 536276 355204 536278
rect 390604 536276 391204 536278
rect 426604 536276 427204 536278
rect 462604 536276 463204 536278
rect 498604 536276 499204 536278
rect 534604 536276 535204 536278
rect 570604 536276 571204 536278
rect 591900 536276 592500 536278
rect -8576 536254 592500 536276
rect -8576 536018 -8394 536254
rect -8158 536018 30786 536254
rect 31022 536018 66786 536254
rect 67022 536018 102786 536254
rect 103022 536018 138786 536254
rect 139022 536018 174786 536254
rect 175022 536018 210786 536254
rect 211022 536018 246786 536254
rect 247022 536018 282786 536254
rect 283022 536018 318786 536254
rect 319022 536018 354786 536254
rect 355022 536018 390786 536254
rect 391022 536018 426786 536254
rect 427022 536018 462786 536254
rect 463022 536018 498786 536254
rect 499022 536018 534786 536254
rect 535022 536018 570786 536254
rect 571022 536018 592082 536254
rect 592318 536018 592500 536254
rect -8576 535934 592500 536018
rect -8576 535698 -8394 535934
rect -8158 535698 30786 535934
rect 31022 535698 66786 535934
rect 67022 535698 102786 535934
rect 103022 535698 138786 535934
rect 139022 535698 174786 535934
rect 175022 535698 210786 535934
rect 211022 535698 246786 535934
rect 247022 535698 282786 535934
rect 283022 535698 318786 535934
rect 319022 535698 354786 535934
rect 355022 535698 390786 535934
rect 391022 535698 426786 535934
rect 427022 535698 462786 535934
rect 463022 535698 498786 535934
rect 499022 535698 534786 535934
rect 535022 535698 570786 535934
rect 571022 535698 592082 535934
rect 592318 535698 592500 535934
rect -8576 535676 592500 535698
rect -8576 535674 -7976 535676
rect 30604 535674 31204 535676
rect 66604 535674 67204 535676
rect 102604 535674 103204 535676
rect 138604 535674 139204 535676
rect 174604 535674 175204 535676
rect 210604 535674 211204 535676
rect 246604 535674 247204 535676
rect 282604 535674 283204 535676
rect 318604 535674 319204 535676
rect 354604 535674 355204 535676
rect 390604 535674 391204 535676
rect 426604 535674 427204 535676
rect 462604 535674 463204 535676
rect 498604 535674 499204 535676
rect 534604 535674 535204 535676
rect 570604 535674 571204 535676
rect 591900 535674 592500 535676
rect -6696 532676 -6096 532678
rect 27004 532676 27604 532678
rect 63004 532676 63604 532678
rect 99004 532676 99604 532678
rect 135004 532676 135604 532678
rect 171004 532676 171604 532678
rect 207004 532676 207604 532678
rect 243004 532676 243604 532678
rect 279004 532676 279604 532678
rect 315004 532676 315604 532678
rect 351004 532676 351604 532678
rect 387004 532676 387604 532678
rect 423004 532676 423604 532678
rect 459004 532676 459604 532678
rect 495004 532676 495604 532678
rect 531004 532676 531604 532678
rect 567004 532676 567604 532678
rect 590020 532676 590620 532678
rect -6696 532654 590620 532676
rect -6696 532418 -6514 532654
rect -6278 532418 27186 532654
rect 27422 532418 63186 532654
rect 63422 532418 99186 532654
rect 99422 532418 135186 532654
rect 135422 532418 171186 532654
rect 171422 532418 207186 532654
rect 207422 532418 243186 532654
rect 243422 532418 279186 532654
rect 279422 532418 315186 532654
rect 315422 532418 351186 532654
rect 351422 532418 387186 532654
rect 387422 532418 423186 532654
rect 423422 532418 459186 532654
rect 459422 532418 495186 532654
rect 495422 532418 531186 532654
rect 531422 532418 567186 532654
rect 567422 532418 590202 532654
rect 590438 532418 590620 532654
rect -6696 532334 590620 532418
rect -6696 532098 -6514 532334
rect -6278 532098 27186 532334
rect 27422 532098 63186 532334
rect 63422 532098 99186 532334
rect 99422 532098 135186 532334
rect 135422 532098 171186 532334
rect 171422 532098 207186 532334
rect 207422 532098 243186 532334
rect 243422 532098 279186 532334
rect 279422 532098 315186 532334
rect 315422 532098 351186 532334
rect 351422 532098 387186 532334
rect 387422 532098 423186 532334
rect 423422 532098 459186 532334
rect 459422 532098 495186 532334
rect 495422 532098 531186 532334
rect 531422 532098 567186 532334
rect 567422 532098 590202 532334
rect 590438 532098 590620 532334
rect -6696 532076 590620 532098
rect -6696 532074 -6096 532076
rect 27004 532074 27604 532076
rect 63004 532074 63604 532076
rect 99004 532074 99604 532076
rect 135004 532074 135604 532076
rect 171004 532074 171604 532076
rect 207004 532074 207604 532076
rect 243004 532074 243604 532076
rect 279004 532074 279604 532076
rect 315004 532074 315604 532076
rect 351004 532074 351604 532076
rect 387004 532074 387604 532076
rect 423004 532074 423604 532076
rect 459004 532074 459604 532076
rect 495004 532074 495604 532076
rect 531004 532074 531604 532076
rect 567004 532074 567604 532076
rect 590020 532074 590620 532076
rect -4816 529076 -4216 529078
rect 23404 529076 24004 529078
rect 59404 529076 60004 529078
rect 95404 529076 96004 529078
rect 131404 529076 132004 529078
rect 167404 529076 168004 529078
rect 203404 529076 204004 529078
rect 239404 529076 240004 529078
rect 275404 529076 276004 529078
rect 311404 529076 312004 529078
rect 347404 529076 348004 529078
rect 383404 529076 384004 529078
rect 419404 529076 420004 529078
rect 455404 529076 456004 529078
rect 491404 529076 492004 529078
rect 527404 529076 528004 529078
rect 563404 529076 564004 529078
rect 588140 529076 588740 529078
rect -4816 529054 588740 529076
rect -4816 528818 -4634 529054
rect -4398 528818 23586 529054
rect 23822 528818 59586 529054
rect 59822 528818 95586 529054
rect 95822 528818 131586 529054
rect 131822 528818 167586 529054
rect 167822 528818 203586 529054
rect 203822 528818 239586 529054
rect 239822 528818 275586 529054
rect 275822 528818 311586 529054
rect 311822 528818 347586 529054
rect 347822 528818 383586 529054
rect 383822 528818 419586 529054
rect 419822 528818 455586 529054
rect 455822 528818 491586 529054
rect 491822 528818 527586 529054
rect 527822 528818 563586 529054
rect 563822 528818 588322 529054
rect 588558 528818 588740 529054
rect -4816 528734 588740 528818
rect -4816 528498 -4634 528734
rect -4398 528498 23586 528734
rect 23822 528498 59586 528734
rect 59822 528498 95586 528734
rect 95822 528498 131586 528734
rect 131822 528498 167586 528734
rect 167822 528498 203586 528734
rect 203822 528498 239586 528734
rect 239822 528498 275586 528734
rect 275822 528498 311586 528734
rect 311822 528498 347586 528734
rect 347822 528498 383586 528734
rect 383822 528498 419586 528734
rect 419822 528498 455586 528734
rect 455822 528498 491586 528734
rect 491822 528498 527586 528734
rect 527822 528498 563586 528734
rect 563822 528498 588322 528734
rect 588558 528498 588740 528734
rect -4816 528476 588740 528498
rect -4816 528474 -4216 528476
rect 23404 528474 24004 528476
rect 59404 528474 60004 528476
rect 95404 528474 96004 528476
rect 131404 528474 132004 528476
rect 167404 528474 168004 528476
rect 203404 528474 204004 528476
rect 239404 528474 240004 528476
rect 275404 528474 276004 528476
rect 311404 528474 312004 528476
rect 347404 528474 348004 528476
rect 383404 528474 384004 528476
rect 419404 528474 420004 528476
rect 455404 528474 456004 528476
rect 491404 528474 492004 528476
rect 527404 528474 528004 528476
rect 563404 528474 564004 528476
rect 588140 528474 588740 528476
rect -2936 525476 -2336 525478
rect 19804 525476 20404 525478
rect 55804 525476 56404 525478
rect 91804 525476 92404 525478
rect 127804 525476 128404 525478
rect 163804 525476 164404 525478
rect 199804 525476 200404 525478
rect 235804 525476 236404 525478
rect 271804 525476 272404 525478
rect 307804 525476 308404 525478
rect 343804 525476 344404 525478
rect 379804 525476 380404 525478
rect 415804 525476 416404 525478
rect 451804 525476 452404 525478
rect 487804 525476 488404 525478
rect 523804 525476 524404 525478
rect 559804 525476 560404 525478
rect 586260 525476 586860 525478
rect -2936 525454 586860 525476
rect -2936 525218 -2754 525454
rect -2518 525218 19986 525454
rect 20222 525218 55986 525454
rect 56222 525218 91986 525454
rect 92222 525218 127986 525454
rect 128222 525218 163986 525454
rect 164222 525218 199986 525454
rect 200222 525218 235986 525454
rect 236222 525218 271986 525454
rect 272222 525218 307986 525454
rect 308222 525218 343986 525454
rect 344222 525218 379986 525454
rect 380222 525218 415986 525454
rect 416222 525218 451986 525454
rect 452222 525218 487986 525454
rect 488222 525218 523986 525454
rect 524222 525218 559986 525454
rect 560222 525218 586442 525454
rect 586678 525218 586860 525454
rect -2936 525134 586860 525218
rect -2936 524898 -2754 525134
rect -2518 524898 19986 525134
rect 20222 524898 55986 525134
rect 56222 524898 91986 525134
rect 92222 524898 127986 525134
rect 128222 524898 163986 525134
rect 164222 524898 199986 525134
rect 200222 524898 235986 525134
rect 236222 524898 271986 525134
rect 272222 524898 307986 525134
rect 308222 524898 343986 525134
rect 344222 524898 379986 525134
rect 380222 524898 415986 525134
rect 416222 524898 451986 525134
rect 452222 524898 487986 525134
rect 488222 524898 523986 525134
rect 524222 524898 559986 525134
rect 560222 524898 586442 525134
rect 586678 524898 586860 525134
rect -2936 524876 586860 524898
rect -2936 524874 -2336 524876
rect 19804 524874 20404 524876
rect 55804 524874 56404 524876
rect 91804 524874 92404 524876
rect 127804 524874 128404 524876
rect 163804 524874 164404 524876
rect 199804 524874 200404 524876
rect 235804 524874 236404 524876
rect 271804 524874 272404 524876
rect 307804 524874 308404 524876
rect 343804 524874 344404 524876
rect 379804 524874 380404 524876
rect 415804 524874 416404 524876
rect 451804 524874 452404 524876
rect 487804 524874 488404 524876
rect 523804 524874 524404 524876
rect 559804 524874 560404 524876
rect 586260 524874 586860 524876
rect -7636 518276 -7036 518278
rect 12604 518276 13204 518278
rect 48604 518276 49204 518278
rect 84604 518276 85204 518278
rect 120604 518276 121204 518278
rect 156604 518276 157204 518278
rect 192604 518276 193204 518278
rect 228604 518276 229204 518278
rect 264604 518276 265204 518278
rect 300604 518276 301204 518278
rect 336604 518276 337204 518278
rect 372604 518276 373204 518278
rect 408604 518276 409204 518278
rect 444604 518276 445204 518278
rect 480604 518276 481204 518278
rect 516604 518276 517204 518278
rect 552604 518276 553204 518278
rect 590960 518276 591560 518278
rect -8576 518254 592500 518276
rect -8576 518018 -7454 518254
rect -7218 518018 12786 518254
rect 13022 518018 48786 518254
rect 49022 518018 84786 518254
rect 85022 518018 120786 518254
rect 121022 518018 156786 518254
rect 157022 518018 192786 518254
rect 193022 518018 228786 518254
rect 229022 518018 264786 518254
rect 265022 518018 300786 518254
rect 301022 518018 336786 518254
rect 337022 518018 372786 518254
rect 373022 518018 408786 518254
rect 409022 518018 444786 518254
rect 445022 518018 480786 518254
rect 481022 518018 516786 518254
rect 517022 518018 552786 518254
rect 553022 518018 591142 518254
rect 591378 518018 592500 518254
rect -8576 517934 592500 518018
rect -8576 517698 -7454 517934
rect -7218 517698 12786 517934
rect 13022 517698 48786 517934
rect 49022 517698 84786 517934
rect 85022 517698 120786 517934
rect 121022 517698 156786 517934
rect 157022 517698 192786 517934
rect 193022 517698 228786 517934
rect 229022 517698 264786 517934
rect 265022 517698 300786 517934
rect 301022 517698 336786 517934
rect 337022 517698 372786 517934
rect 373022 517698 408786 517934
rect 409022 517698 444786 517934
rect 445022 517698 480786 517934
rect 481022 517698 516786 517934
rect 517022 517698 552786 517934
rect 553022 517698 591142 517934
rect 591378 517698 592500 517934
rect -8576 517676 592500 517698
rect -7636 517674 -7036 517676
rect 12604 517674 13204 517676
rect 48604 517674 49204 517676
rect 84604 517674 85204 517676
rect 120604 517674 121204 517676
rect 156604 517674 157204 517676
rect 192604 517674 193204 517676
rect 228604 517674 229204 517676
rect 264604 517674 265204 517676
rect 300604 517674 301204 517676
rect 336604 517674 337204 517676
rect 372604 517674 373204 517676
rect 408604 517674 409204 517676
rect 444604 517674 445204 517676
rect 480604 517674 481204 517676
rect 516604 517674 517204 517676
rect 552604 517674 553204 517676
rect 590960 517674 591560 517676
rect -5756 514676 -5156 514678
rect 9004 514676 9604 514678
rect 45004 514676 45604 514678
rect 81004 514676 81604 514678
rect 117004 514676 117604 514678
rect 153004 514676 153604 514678
rect 189004 514676 189604 514678
rect 225004 514676 225604 514678
rect 261004 514676 261604 514678
rect 297004 514676 297604 514678
rect 333004 514676 333604 514678
rect 369004 514676 369604 514678
rect 405004 514676 405604 514678
rect 441004 514676 441604 514678
rect 477004 514676 477604 514678
rect 513004 514676 513604 514678
rect 549004 514676 549604 514678
rect 589080 514676 589680 514678
rect -6696 514654 590620 514676
rect -6696 514418 -5574 514654
rect -5338 514418 9186 514654
rect 9422 514418 45186 514654
rect 45422 514418 81186 514654
rect 81422 514418 117186 514654
rect 117422 514418 153186 514654
rect 153422 514418 189186 514654
rect 189422 514418 225186 514654
rect 225422 514418 261186 514654
rect 261422 514418 297186 514654
rect 297422 514418 333186 514654
rect 333422 514418 369186 514654
rect 369422 514418 405186 514654
rect 405422 514418 441186 514654
rect 441422 514418 477186 514654
rect 477422 514418 513186 514654
rect 513422 514418 549186 514654
rect 549422 514418 589262 514654
rect 589498 514418 590620 514654
rect -6696 514334 590620 514418
rect -6696 514098 -5574 514334
rect -5338 514098 9186 514334
rect 9422 514098 45186 514334
rect 45422 514098 81186 514334
rect 81422 514098 117186 514334
rect 117422 514098 153186 514334
rect 153422 514098 189186 514334
rect 189422 514098 225186 514334
rect 225422 514098 261186 514334
rect 261422 514098 297186 514334
rect 297422 514098 333186 514334
rect 333422 514098 369186 514334
rect 369422 514098 405186 514334
rect 405422 514098 441186 514334
rect 441422 514098 477186 514334
rect 477422 514098 513186 514334
rect 513422 514098 549186 514334
rect 549422 514098 589262 514334
rect 589498 514098 590620 514334
rect -6696 514076 590620 514098
rect -5756 514074 -5156 514076
rect 9004 514074 9604 514076
rect 45004 514074 45604 514076
rect 81004 514074 81604 514076
rect 117004 514074 117604 514076
rect 153004 514074 153604 514076
rect 189004 514074 189604 514076
rect 225004 514074 225604 514076
rect 261004 514074 261604 514076
rect 297004 514074 297604 514076
rect 333004 514074 333604 514076
rect 369004 514074 369604 514076
rect 405004 514074 405604 514076
rect 441004 514074 441604 514076
rect 477004 514074 477604 514076
rect 513004 514074 513604 514076
rect 549004 514074 549604 514076
rect 589080 514074 589680 514076
rect -3876 511076 -3276 511078
rect 5404 511076 6004 511078
rect 41404 511076 42004 511078
rect 77404 511076 78004 511078
rect 113404 511076 114004 511078
rect 149404 511076 150004 511078
rect 185404 511076 186004 511078
rect 221404 511076 222004 511078
rect 257404 511076 258004 511078
rect 293404 511076 294004 511078
rect 329404 511076 330004 511078
rect 365404 511076 366004 511078
rect 401404 511076 402004 511078
rect 437404 511076 438004 511078
rect 473404 511076 474004 511078
rect 509404 511076 510004 511078
rect 545404 511076 546004 511078
rect 581404 511076 582004 511078
rect 587200 511076 587800 511078
rect -4816 511054 588740 511076
rect -4816 510818 -3694 511054
rect -3458 510818 5586 511054
rect 5822 510818 41586 511054
rect 41822 510818 77586 511054
rect 77822 510818 113586 511054
rect 113822 510818 149586 511054
rect 149822 510818 185586 511054
rect 185822 510818 221586 511054
rect 221822 510818 257586 511054
rect 257822 510818 293586 511054
rect 293822 510818 329586 511054
rect 329822 510818 365586 511054
rect 365822 510818 401586 511054
rect 401822 510818 437586 511054
rect 437822 510818 473586 511054
rect 473822 510818 509586 511054
rect 509822 510818 545586 511054
rect 545822 510818 581586 511054
rect 581822 510818 587382 511054
rect 587618 510818 588740 511054
rect -4816 510734 588740 510818
rect -4816 510498 -3694 510734
rect -3458 510498 5586 510734
rect 5822 510498 41586 510734
rect 41822 510498 77586 510734
rect 77822 510498 113586 510734
rect 113822 510498 149586 510734
rect 149822 510498 185586 510734
rect 185822 510498 221586 510734
rect 221822 510498 257586 510734
rect 257822 510498 293586 510734
rect 293822 510498 329586 510734
rect 329822 510498 365586 510734
rect 365822 510498 401586 510734
rect 401822 510498 437586 510734
rect 437822 510498 473586 510734
rect 473822 510498 509586 510734
rect 509822 510498 545586 510734
rect 545822 510498 581586 510734
rect 581822 510498 587382 510734
rect 587618 510498 588740 510734
rect -4816 510476 588740 510498
rect -3876 510474 -3276 510476
rect 5404 510474 6004 510476
rect 41404 510474 42004 510476
rect 77404 510474 78004 510476
rect 113404 510474 114004 510476
rect 149404 510474 150004 510476
rect 185404 510474 186004 510476
rect 221404 510474 222004 510476
rect 257404 510474 258004 510476
rect 293404 510474 294004 510476
rect 329404 510474 330004 510476
rect 365404 510474 366004 510476
rect 401404 510474 402004 510476
rect 437404 510474 438004 510476
rect 473404 510474 474004 510476
rect 509404 510474 510004 510476
rect 545404 510474 546004 510476
rect 581404 510474 582004 510476
rect 587200 510474 587800 510476
rect -1996 507476 -1396 507478
rect 1804 507476 2404 507478
rect 37804 507476 38404 507478
rect 73804 507476 74404 507478
rect 109804 507476 110404 507478
rect 145804 507476 146404 507478
rect 469804 507476 470404 507478
rect 505804 507476 506404 507478
rect 541804 507476 542404 507478
rect 577804 507476 578404 507478
rect 585320 507476 585920 507478
rect -2936 507454 156000 507476
rect -2936 507218 -1814 507454
rect -1578 507218 1986 507454
rect 2222 507218 37986 507454
rect 38222 507218 73986 507454
rect 74222 507218 109986 507454
rect 110222 507218 145986 507454
rect 146222 507218 156000 507454
rect -2936 507134 156000 507218
rect -2936 506898 -1814 507134
rect -1578 506898 1986 507134
rect 2222 506898 37986 507134
rect 38222 506898 73986 507134
rect 74222 506898 109986 507134
rect 110222 506898 145986 507134
rect 146222 506898 156000 507134
rect -2936 506876 156000 506898
rect 440000 507454 586860 507476
rect 440000 507218 469986 507454
rect 470222 507218 505986 507454
rect 506222 507218 541986 507454
rect 542222 507218 577986 507454
rect 578222 507218 585502 507454
rect 585738 507218 586860 507454
rect 440000 507134 586860 507218
rect 440000 506898 469986 507134
rect 470222 506898 505986 507134
rect 506222 506898 541986 507134
rect 542222 506898 577986 507134
rect 578222 506898 585502 507134
rect 585738 506898 586860 507134
rect 440000 506876 586860 506898
rect -1996 506874 -1396 506876
rect 1804 506874 2404 506876
rect 37804 506874 38404 506876
rect 73804 506874 74404 506876
rect 109804 506874 110404 506876
rect 145804 506874 146404 506876
rect 469804 506874 470404 506876
rect 505804 506874 506404 506876
rect 541804 506874 542404 506876
rect 577804 506874 578404 506876
rect 585320 506874 585920 506876
rect -8576 500276 -7976 500278
rect 30604 500276 31204 500278
rect 66604 500276 67204 500278
rect 102604 500276 103204 500278
rect 138604 500276 139204 500278
rect 462604 500276 463204 500278
rect 498604 500276 499204 500278
rect 534604 500276 535204 500278
rect 570604 500276 571204 500278
rect 591900 500276 592500 500278
rect -8576 500254 156000 500276
rect -8576 500018 -8394 500254
rect -8158 500018 30786 500254
rect 31022 500018 66786 500254
rect 67022 500018 102786 500254
rect 103022 500018 138786 500254
rect 139022 500018 156000 500254
rect -8576 499934 156000 500018
rect -8576 499698 -8394 499934
rect -8158 499698 30786 499934
rect 31022 499698 66786 499934
rect 67022 499698 102786 499934
rect 103022 499698 138786 499934
rect 139022 499698 156000 499934
rect -8576 499676 156000 499698
rect 440000 500254 592500 500276
rect 440000 500018 462786 500254
rect 463022 500018 498786 500254
rect 499022 500018 534786 500254
rect 535022 500018 570786 500254
rect 571022 500018 592082 500254
rect 592318 500018 592500 500254
rect 440000 499934 592500 500018
rect 440000 499698 462786 499934
rect 463022 499698 498786 499934
rect 499022 499698 534786 499934
rect 535022 499698 570786 499934
rect 571022 499698 592082 499934
rect 592318 499698 592500 499934
rect 440000 499676 592500 499698
rect -8576 499674 -7976 499676
rect 30604 499674 31204 499676
rect 66604 499674 67204 499676
rect 102604 499674 103204 499676
rect 138604 499674 139204 499676
rect 462604 499674 463204 499676
rect 498604 499674 499204 499676
rect 534604 499674 535204 499676
rect 570604 499674 571204 499676
rect 591900 499674 592500 499676
rect -6696 496676 -6096 496678
rect 27004 496676 27604 496678
rect 63004 496676 63604 496678
rect 99004 496676 99604 496678
rect 135004 496676 135604 496678
rect 459004 496676 459604 496678
rect 495004 496676 495604 496678
rect 531004 496676 531604 496678
rect 567004 496676 567604 496678
rect 590020 496676 590620 496678
rect -6696 496654 156000 496676
rect -6696 496418 -6514 496654
rect -6278 496418 27186 496654
rect 27422 496418 63186 496654
rect 63422 496418 99186 496654
rect 99422 496418 135186 496654
rect 135422 496418 156000 496654
rect -6696 496334 156000 496418
rect -6696 496098 -6514 496334
rect -6278 496098 27186 496334
rect 27422 496098 63186 496334
rect 63422 496098 99186 496334
rect 99422 496098 135186 496334
rect 135422 496098 156000 496334
rect -6696 496076 156000 496098
rect 440000 496654 590620 496676
rect 440000 496418 459186 496654
rect 459422 496418 495186 496654
rect 495422 496418 531186 496654
rect 531422 496418 567186 496654
rect 567422 496418 590202 496654
rect 590438 496418 590620 496654
rect 440000 496334 590620 496418
rect 440000 496098 459186 496334
rect 459422 496098 495186 496334
rect 495422 496098 531186 496334
rect 531422 496098 567186 496334
rect 567422 496098 590202 496334
rect 590438 496098 590620 496334
rect 440000 496076 590620 496098
rect -6696 496074 -6096 496076
rect 27004 496074 27604 496076
rect 63004 496074 63604 496076
rect 99004 496074 99604 496076
rect 135004 496074 135604 496076
rect 459004 496074 459604 496076
rect 495004 496074 495604 496076
rect 531004 496074 531604 496076
rect 567004 496074 567604 496076
rect 590020 496074 590620 496076
rect -4816 493076 -4216 493078
rect 23404 493076 24004 493078
rect 59404 493076 60004 493078
rect 95404 493076 96004 493078
rect 131404 493076 132004 493078
rect 455404 493076 456004 493078
rect 491404 493076 492004 493078
rect 527404 493076 528004 493078
rect 563404 493076 564004 493078
rect 588140 493076 588740 493078
rect -4816 493054 156000 493076
rect -4816 492818 -4634 493054
rect -4398 492818 23586 493054
rect 23822 492818 59586 493054
rect 59822 492818 95586 493054
rect 95822 492818 131586 493054
rect 131822 492818 156000 493054
rect -4816 492734 156000 492818
rect -4816 492498 -4634 492734
rect -4398 492498 23586 492734
rect 23822 492498 59586 492734
rect 59822 492498 95586 492734
rect 95822 492498 131586 492734
rect 131822 492498 156000 492734
rect -4816 492476 156000 492498
rect 440000 493054 588740 493076
rect 440000 492818 455586 493054
rect 455822 492818 491586 493054
rect 491822 492818 527586 493054
rect 527822 492818 563586 493054
rect 563822 492818 588322 493054
rect 588558 492818 588740 493054
rect 440000 492734 588740 492818
rect 440000 492498 455586 492734
rect 455822 492498 491586 492734
rect 491822 492498 527586 492734
rect 527822 492498 563586 492734
rect 563822 492498 588322 492734
rect 588558 492498 588740 492734
rect 440000 492476 588740 492498
rect -4816 492474 -4216 492476
rect 23404 492474 24004 492476
rect 59404 492474 60004 492476
rect 95404 492474 96004 492476
rect 131404 492474 132004 492476
rect 455404 492474 456004 492476
rect 491404 492474 492004 492476
rect 527404 492474 528004 492476
rect 563404 492474 564004 492476
rect 588140 492474 588740 492476
rect -2936 489476 -2336 489478
rect 19804 489476 20404 489478
rect 55804 489476 56404 489478
rect 91804 489476 92404 489478
rect 127804 489476 128404 489478
rect 451804 489476 452404 489478
rect 487804 489476 488404 489478
rect 523804 489476 524404 489478
rect 559804 489476 560404 489478
rect 586260 489476 586860 489478
rect -2936 489454 156000 489476
rect -2936 489218 -2754 489454
rect -2518 489218 19986 489454
rect 20222 489218 55986 489454
rect 56222 489218 91986 489454
rect 92222 489218 127986 489454
rect 128222 489218 156000 489454
rect -2936 489134 156000 489218
rect -2936 488898 -2754 489134
rect -2518 488898 19986 489134
rect 20222 488898 55986 489134
rect 56222 488898 91986 489134
rect 92222 488898 127986 489134
rect 128222 488898 156000 489134
rect -2936 488876 156000 488898
rect 440000 489454 586860 489476
rect 440000 489218 451986 489454
rect 452222 489218 487986 489454
rect 488222 489218 523986 489454
rect 524222 489218 559986 489454
rect 560222 489218 586442 489454
rect 586678 489218 586860 489454
rect 440000 489134 586860 489218
rect 440000 488898 451986 489134
rect 452222 488898 487986 489134
rect 488222 488898 523986 489134
rect 524222 488898 559986 489134
rect 560222 488898 586442 489134
rect 586678 488898 586860 489134
rect 440000 488876 586860 488898
rect -2936 488874 -2336 488876
rect 19804 488874 20404 488876
rect 55804 488874 56404 488876
rect 91804 488874 92404 488876
rect 127804 488874 128404 488876
rect 451804 488874 452404 488876
rect 487804 488874 488404 488876
rect 523804 488874 524404 488876
rect 559804 488874 560404 488876
rect 586260 488874 586860 488876
rect -7636 482276 -7036 482278
rect 12604 482276 13204 482278
rect 48604 482276 49204 482278
rect 84604 482276 85204 482278
rect 120604 482276 121204 482278
rect 444604 482276 445204 482278
rect 480604 482276 481204 482278
rect 516604 482276 517204 482278
rect 552604 482276 553204 482278
rect 590960 482276 591560 482278
rect -8576 482254 156000 482276
rect -8576 482018 -7454 482254
rect -7218 482018 12786 482254
rect 13022 482018 48786 482254
rect 49022 482018 84786 482254
rect 85022 482018 120786 482254
rect 121022 482018 156000 482254
rect -8576 481934 156000 482018
rect -8576 481698 -7454 481934
rect -7218 481698 12786 481934
rect 13022 481698 48786 481934
rect 49022 481698 84786 481934
rect 85022 481698 120786 481934
rect 121022 481698 156000 481934
rect -8576 481676 156000 481698
rect 440000 482254 592500 482276
rect 440000 482018 444786 482254
rect 445022 482018 480786 482254
rect 481022 482018 516786 482254
rect 517022 482018 552786 482254
rect 553022 482018 591142 482254
rect 591378 482018 592500 482254
rect 440000 481934 592500 482018
rect 440000 481698 444786 481934
rect 445022 481698 480786 481934
rect 481022 481698 516786 481934
rect 517022 481698 552786 481934
rect 553022 481698 591142 481934
rect 591378 481698 592500 481934
rect 440000 481676 592500 481698
rect -7636 481674 -7036 481676
rect 12604 481674 13204 481676
rect 48604 481674 49204 481676
rect 84604 481674 85204 481676
rect 120604 481674 121204 481676
rect 444604 481674 445204 481676
rect 480604 481674 481204 481676
rect 516604 481674 517204 481676
rect 552604 481674 553204 481676
rect 590960 481674 591560 481676
rect -5756 478676 -5156 478678
rect 9004 478676 9604 478678
rect 45004 478676 45604 478678
rect 81004 478676 81604 478678
rect 117004 478676 117604 478678
rect 153004 478676 153604 478678
rect 441004 478676 441604 478678
rect 477004 478676 477604 478678
rect 513004 478676 513604 478678
rect 549004 478676 549604 478678
rect 589080 478676 589680 478678
rect -6696 478654 156000 478676
rect -6696 478418 -5574 478654
rect -5338 478418 9186 478654
rect 9422 478418 45186 478654
rect 45422 478418 81186 478654
rect 81422 478418 117186 478654
rect 117422 478418 153186 478654
rect 153422 478418 156000 478654
rect -6696 478334 156000 478418
rect -6696 478098 -5574 478334
rect -5338 478098 9186 478334
rect 9422 478098 45186 478334
rect 45422 478098 81186 478334
rect 81422 478098 117186 478334
rect 117422 478098 153186 478334
rect 153422 478098 156000 478334
rect -6696 478076 156000 478098
rect 440000 478654 590620 478676
rect 440000 478418 441186 478654
rect 441422 478418 477186 478654
rect 477422 478418 513186 478654
rect 513422 478418 549186 478654
rect 549422 478418 589262 478654
rect 589498 478418 590620 478654
rect 440000 478334 590620 478418
rect 440000 478098 441186 478334
rect 441422 478098 477186 478334
rect 477422 478098 513186 478334
rect 513422 478098 549186 478334
rect 549422 478098 589262 478334
rect 589498 478098 590620 478334
rect 440000 478076 590620 478098
rect -5756 478074 -5156 478076
rect 9004 478074 9604 478076
rect 45004 478074 45604 478076
rect 81004 478074 81604 478076
rect 117004 478074 117604 478076
rect 153004 478074 153604 478076
rect 441004 478074 441604 478076
rect 477004 478074 477604 478076
rect 513004 478074 513604 478076
rect 549004 478074 549604 478076
rect 589080 478074 589680 478076
rect -3876 475076 -3276 475078
rect 5404 475076 6004 475078
rect 41404 475076 42004 475078
rect 77404 475076 78004 475078
rect 113404 475076 114004 475078
rect 149404 475076 150004 475078
rect 473404 475076 474004 475078
rect 509404 475076 510004 475078
rect 545404 475076 546004 475078
rect 581404 475076 582004 475078
rect 587200 475076 587800 475078
rect -4816 475054 156000 475076
rect -4816 474818 -3694 475054
rect -3458 474818 5586 475054
rect 5822 474818 41586 475054
rect 41822 474818 77586 475054
rect 77822 474818 113586 475054
rect 113822 474818 149586 475054
rect 149822 474818 156000 475054
rect -4816 474734 156000 474818
rect -4816 474498 -3694 474734
rect -3458 474498 5586 474734
rect 5822 474498 41586 474734
rect 41822 474498 77586 474734
rect 77822 474498 113586 474734
rect 113822 474498 149586 474734
rect 149822 474498 156000 474734
rect -4816 474476 156000 474498
rect 440000 475054 588740 475076
rect 440000 474818 473586 475054
rect 473822 474818 509586 475054
rect 509822 474818 545586 475054
rect 545822 474818 581586 475054
rect 581822 474818 587382 475054
rect 587618 474818 588740 475054
rect 440000 474734 588740 474818
rect 440000 474498 473586 474734
rect 473822 474498 509586 474734
rect 509822 474498 545586 474734
rect 545822 474498 581586 474734
rect 581822 474498 587382 474734
rect 587618 474498 588740 474734
rect 440000 474476 588740 474498
rect -3876 474474 -3276 474476
rect 5404 474474 6004 474476
rect 41404 474474 42004 474476
rect 77404 474474 78004 474476
rect 113404 474474 114004 474476
rect 149404 474474 150004 474476
rect 473404 474474 474004 474476
rect 509404 474474 510004 474476
rect 545404 474474 546004 474476
rect 581404 474474 582004 474476
rect 587200 474474 587800 474476
rect -1996 471476 -1396 471478
rect 1804 471476 2404 471478
rect 37804 471476 38404 471478
rect 73804 471476 74404 471478
rect 109804 471476 110404 471478
rect 145804 471476 146404 471478
rect 469804 471476 470404 471478
rect 505804 471476 506404 471478
rect 541804 471476 542404 471478
rect 577804 471476 578404 471478
rect 585320 471476 585920 471478
rect -2936 471454 156000 471476
rect -2936 471218 -1814 471454
rect -1578 471218 1986 471454
rect 2222 471218 37986 471454
rect 38222 471218 73986 471454
rect 74222 471218 109986 471454
rect 110222 471218 145986 471454
rect 146222 471218 156000 471454
rect -2936 471134 156000 471218
rect -2936 470898 -1814 471134
rect -1578 470898 1986 471134
rect 2222 470898 37986 471134
rect 38222 470898 73986 471134
rect 74222 470898 109986 471134
rect 110222 470898 145986 471134
rect 146222 470898 156000 471134
rect -2936 470876 156000 470898
rect 440000 471454 586860 471476
rect 440000 471218 469986 471454
rect 470222 471218 505986 471454
rect 506222 471218 541986 471454
rect 542222 471218 577986 471454
rect 578222 471218 585502 471454
rect 585738 471218 586860 471454
rect 440000 471134 586860 471218
rect 440000 470898 469986 471134
rect 470222 470898 505986 471134
rect 506222 470898 541986 471134
rect 542222 470898 577986 471134
rect 578222 470898 585502 471134
rect 585738 470898 586860 471134
rect 440000 470876 586860 470898
rect -1996 470874 -1396 470876
rect 1804 470874 2404 470876
rect 37804 470874 38404 470876
rect 73804 470874 74404 470876
rect 109804 470874 110404 470876
rect 145804 470874 146404 470876
rect 469804 470874 470404 470876
rect 505804 470874 506404 470876
rect 541804 470874 542404 470876
rect 577804 470874 578404 470876
rect 585320 470874 585920 470876
rect -8576 464276 -7976 464278
rect 30604 464276 31204 464278
rect 66604 464276 67204 464278
rect 102604 464276 103204 464278
rect 138604 464276 139204 464278
rect 462604 464276 463204 464278
rect 498604 464276 499204 464278
rect 534604 464276 535204 464278
rect 570604 464276 571204 464278
rect 591900 464276 592500 464278
rect -8576 464254 156000 464276
rect -8576 464018 -8394 464254
rect -8158 464018 30786 464254
rect 31022 464018 66786 464254
rect 67022 464018 102786 464254
rect 103022 464018 138786 464254
rect 139022 464018 156000 464254
rect -8576 463934 156000 464018
rect -8576 463698 -8394 463934
rect -8158 463698 30786 463934
rect 31022 463698 66786 463934
rect 67022 463698 102786 463934
rect 103022 463698 138786 463934
rect 139022 463698 156000 463934
rect -8576 463676 156000 463698
rect 440000 464254 592500 464276
rect 440000 464018 462786 464254
rect 463022 464018 498786 464254
rect 499022 464018 534786 464254
rect 535022 464018 570786 464254
rect 571022 464018 592082 464254
rect 592318 464018 592500 464254
rect 440000 463934 592500 464018
rect 440000 463698 462786 463934
rect 463022 463698 498786 463934
rect 499022 463698 534786 463934
rect 535022 463698 570786 463934
rect 571022 463698 592082 463934
rect 592318 463698 592500 463934
rect 440000 463676 592500 463698
rect -8576 463674 -7976 463676
rect 30604 463674 31204 463676
rect 66604 463674 67204 463676
rect 102604 463674 103204 463676
rect 138604 463674 139204 463676
rect 462604 463674 463204 463676
rect 498604 463674 499204 463676
rect 534604 463674 535204 463676
rect 570604 463674 571204 463676
rect 591900 463674 592500 463676
rect -6696 460676 -6096 460678
rect 27004 460676 27604 460678
rect 63004 460676 63604 460678
rect 99004 460676 99604 460678
rect 135004 460676 135604 460678
rect 459004 460676 459604 460678
rect 495004 460676 495604 460678
rect 531004 460676 531604 460678
rect 567004 460676 567604 460678
rect 590020 460676 590620 460678
rect -6696 460654 156000 460676
rect -6696 460418 -6514 460654
rect -6278 460418 27186 460654
rect 27422 460418 63186 460654
rect 63422 460418 99186 460654
rect 99422 460418 135186 460654
rect 135422 460418 156000 460654
rect -6696 460334 156000 460418
rect -6696 460098 -6514 460334
rect -6278 460098 27186 460334
rect 27422 460098 63186 460334
rect 63422 460098 99186 460334
rect 99422 460098 135186 460334
rect 135422 460098 156000 460334
rect -6696 460076 156000 460098
rect 440000 460654 590620 460676
rect 440000 460418 459186 460654
rect 459422 460418 495186 460654
rect 495422 460418 531186 460654
rect 531422 460418 567186 460654
rect 567422 460418 590202 460654
rect 590438 460418 590620 460654
rect 440000 460334 590620 460418
rect 440000 460098 459186 460334
rect 459422 460098 495186 460334
rect 495422 460098 531186 460334
rect 531422 460098 567186 460334
rect 567422 460098 590202 460334
rect 590438 460098 590620 460334
rect 440000 460076 590620 460098
rect -6696 460074 -6096 460076
rect 27004 460074 27604 460076
rect 63004 460074 63604 460076
rect 99004 460074 99604 460076
rect 135004 460074 135604 460076
rect 459004 460074 459604 460076
rect 495004 460074 495604 460076
rect 531004 460074 531604 460076
rect 567004 460074 567604 460076
rect 590020 460074 590620 460076
rect -4816 457076 -4216 457078
rect 23404 457076 24004 457078
rect 59404 457076 60004 457078
rect 95404 457076 96004 457078
rect 131404 457076 132004 457078
rect 455404 457076 456004 457078
rect 491404 457076 492004 457078
rect 527404 457076 528004 457078
rect 563404 457076 564004 457078
rect 588140 457076 588740 457078
rect -4816 457054 156000 457076
rect -4816 456818 -4634 457054
rect -4398 456818 23586 457054
rect 23822 456818 59586 457054
rect 59822 456818 95586 457054
rect 95822 456818 131586 457054
rect 131822 456818 156000 457054
rect -4816 456734 156000 456818
rect -4816 456498 -4634 456734
rect -4398 456498 23586 456734
rect 23822 456498 59586 456734
rect 59822 456498 95586 456734
rect 95822 456498 131586 456734
rect 131822 456498 156000 456734
rect -4816 456476 156000 456498
rect 440000 457054 588740 457076
rect 440000 456818 455586 457054
rect 455822 456818 491586 457054
rect 491822 456818 527586 457054
rect 527822 456818 563586 457054
rect 563822 456818 588322 457054
rect 588558 456818 588740 457054
rect 440000 456734 588740 456818
rect 440000 456498 455586 456734
rect 455822 456498 491586 456734
rect 491822 456498 527586 456734
rect 527822 456498 563586 456734
rect 563822 456498 588322 456734
rect 588558 456498 588740 456734
rect 440000 456476 588740 456498
rect -4816 456474 -4216 456476
rect 23404 456474 24004 456476
rect 59404 456474 60004 456476
rect 95404 456474 96004 456476
rect 131404 456474 132004 456476
rect 455404 456474 456004 456476
rect 491404 456474 492004 456476
rect 527404 456474 528004 456476
rect 563404 456474 564004 456476
rect 588140 456474 588740 456476
rect -2936 453476 -2336 453478
rect 19804 453476 20404 453478
rect 55804 453476 56404 453478
rect 91804 453476 92404 453478
rect 127804 453476 128404 453478
rect 451804 453476 452404 453478
rect 487804 453476 488404 453478
rect 523804 453476 524404 453478
rect 559804 453476 560404 453478
rect 586260 453476 586860 453478
rect -2936 453454 156000 453476
rect -2936 453218 -2754 453454
rect -2518 453218 19986 453454
rect 20222 453218 55986 453454
rect 56222 453218 91986 453454
rect 92222 453218 127986 453454
rect 128222 453218 156000 453454
rect -2936 453134 156000 453218
rect -2936 452898 -2754 453134
rect -2518 452898 19986 453134
rect 20222 452898 55986 453134
rect 56222 452898 91986 453134
rect 92222 452898 127986 453134
rect 128222 452898 156000 453134
rect -2936 452876 156000 452898
rect 440000 453454 586860 453476
rect 440000 453218 451986 453454
rect 452222 453218 487986 453454
rect 488222 453218 523986 453454
rect 524222 453218 559986 453454
rect 560222 453218 586442 453454
rect 586678 453218 586860 453454
rect 440000 453134 586860 453218
rect 440000 452898 451986 453134
rect 452222 452898 487986 453134
rect 488222 452898 523986 453134
rect 524222 452898 559986 453134
rect 560222 452898 586442 453134
rect 586678 452898 586860 453134
rect 440000 452876 586860 452898
rect -2936 452874 -2336 452876
rect 19804 452874 20404 452876
rect 55804 452874 56404 452876
rect 91804 452874 92404 452876
rect 127804 452874 128404 452876
rect 451804 452874 452404 452876
rect 487804 452874 488404 452876
rect 523804 452874 524404 452876
rect 559804 452874 560404 452876
rect 586260 452874 586860 452876
rect -7636 446276 -7036 446278
rect 12604 446276 13204 446278
rect 48604 446276 49204 446278
rect 84604 446276 85204 446278
rect 120604 446276 121204 446278
rect 444604 446276 445204 446278
rect 480604 446276 481204 446278
rect 516604 446276 517204 446278
rect 552604 446276 553204 446278
rect 590960 446276 591560 446278
rect -8576 446254 156000 446276
rect -8576 446018 -7454 446254
rect -7218 446018 12786 446254
rect 13022 446018 48786 446254
rect 49022 446018 84786 446254
rect 85022 446018 120786 446254
rect 121022 446018 156000 446254
rect -8576 445934 156000 446018
rect -8576 445698 -7454 445934
rect -7218 445698 12786 445934
rect 13022 445698 48786 445934
rect 49022 445698 84786 445934
rect 85022 445698 120786 445934
rect 121022 445698 156000 445934
rect -8576 445676 156000 445698
rect 440000 446254 592500 446276
rect 440000 446018 444786 446254
rect 445022 446018 480786 446254
rect 481022 446018 516786 446254
rect 517022 446018 552786 446254
rect 553022 446018 591142 446254
rect 591378 446018 592500 446254
rect 440000 445934 592500 446018
rect 440000 445698 444786 445934
rect 445022 445698 480786 445934
rect 481022 445698 516786 445934
rect 517022 445698 552786 445934
rect 553022 445698 591142 445934
rect 591378 445698 592500 445934
rect 440000 445676 592500 445698
rect -7636 445674 -7036 445676
rect 12604 445674 13204 445676
rect 48604 445674 49204 445676
rect 84604 445674 85204 445676
rect 120604 445674 121204 445676
rect 444604 445674 445204 445676
rect 480604 445674 481204 445676
rect 516604 445674 517204 445676
rect 552604 445674 553204 445676
rect 590960 445674 591560 445676
rect -5756 442676 -5156 442678
rect 9004 442676 9604 442678
rect 45004 442676 45604 442678
rect 81004 442676 81604 442678
rect 117004 442676 117604 442678
rect 153004 442676 153604 442678
rect 441004 442676 441604 442678
rect 477004 442676 477604 442678
rect 513004 442676 513604 442678
rect 549004 442676 549604 442678
rect 589080 442676 589680 442678
rect -6696 442654 156000 442676
rect -6696 442418 -5574 442654
rect -5338 442418 9186 442654
rect 9422 442418 45186 442654
rect 45422 442418 81186 442654
rect 81422 442418 117186 442654
rect 117422 442418 153186 442654
rect 153422 442418 156000 442654
rect -6696 442334 156000 442418
rect -6696 442098 -5574 442334
rect -5338 442098 9186 442334
rect 9422 442098 45186 442334
rect 45422 442098 81186 442334
rect 81422 442098 117186 442334
rect 117422 442098 153186 442334
rect 153422 442098 156000 442334
rect -6696 442076 156000 442098
rect 440000 442654 590620 442676
rect 440000 442418 441186 442654
rect 441422 442418 477186 442654
rect 477422 442418 513186 442654
rect 513422 442418 549186 442654
rect 549422 442418 589262 442654
rect 589498 442418 590620 442654
rect 440000 442334 590620 442418
rect 440000 442098 441186 442334
rect 441422 442098 477186 442334
rect 477422 442098 513186 442334
rect 513422 442098 549186 442334
rect 549422 442098 589262 442334
rect 589498 442098 590620 442334
rect 440000 442076 590620 442098
rect -5756 442074 -5156 442076
rect 9004 442074 9604 442076
rect 45004 442074 45604 442076
rect 81004 442074 81604 442076
rect 117004 442074 117604 442076
rect 153004 442074 153604 442076
rect 441004 442074 441604 442076
rect 477004 442074 477604 442076
rect 513004 442074 513604 442076
rect 549004 442074 549604 442076
rect 589080 442074 589680 442076
rect -3876 439076 -3276 439078
rect 5404 439076 6004 439078
rect 41404 439076 42004 439078
rect 77404 439076 78004 439078
rect 113404 439076 114004 439078
rect 149404 439076 150004 439078
rect 473404 439076 474004 439078
rect 509404 439076 510004 439078
rect 545404 439076 546004 439078
rect 581404 439076 582004 439078
rect 587200 439076 587800 439078
rect -4816 439054 156000 439076
rect -4816 438818 -3694 439054
rect -3458 438818 5586 439054
rect 5822 438818 41586 439054
rect 41822 438818 77586 439054
rect 77822 438818 113586 439054
rect 113822 438818 149586 439054
rect 149822 438818 156000 439054
rect -4816 438734 156000 438818
rect -4816 438498 -3694 438734
rect -3458 438498 5586 438734
rect 5822 438498 41586 438734
rect 41822 438498 77586 438734
rect 77822 438498 113586 438734
rect 113822 438498 149586 438734
rect 149822 438498 156000 438734
rect -4816 438476 156000 438498
rect 440000 439054 588740 439076
rect 440000 438818 473586 439054
rect 473822 438818 509586 439054
rect 509822 438818 545586 439054
rect 545822 438818 581586 439054
rect 581822 438818 587382 439054
rect 587618 438818 588740 439054
rect 440000 438734 588740 438818
rect 440000 438498 473586 438734
rect 473822 438498 509586 438734
rect 509822 438498 545586 438734
rect 545822 438498 581586 438734
rect 581822 438498 587382 438734
rect 587618 438498 588740 438734
rect 440000 438476 588740 438498
rect -3876 438474 -3276 438476
rect 5404 438474 6004 438476
rect 41404 438474 42004 438476
rect 77404 438474 78004 438476
rect 113404 438474 114004 438476
rect 149404 438474 150004 438476
rect 473404 438474 474004 438476
rect 509404 438474 510004 438476
rect 545404 438474 546004 438476
rect 581404 438474 582004 438476
rect 587200 438474 587800 438476
rect -1996 435476 -1396 435478
rect 1804 435476 2404 435478
rect 37804 435476 38404 435478
rect 73804 435476 74404 435478
rect 109804 435476 110404 435478
rect 145804 435476 146404 435478
rect 469804 435476 470404 435478
rect 505804 435476 506404 435478
rect 541804 435476 542404 435478
rect 577804 435476 578404 435478
rect 585320 435476 585920 435478
rect -2936 435454 156000 435476
rect -2936 435218 -1814 435454
rect -1578 435218 1986 435454
rect 2222 435218 37986 435454
rect 38222 435218 73986 435454
rect 74222 435218 109986 435454
rect 110222 435218 145986 435454
rect 146222 435218 156000 435454
rect -2936 435134 156000 435218
rect -2936 434898 -1814 435134
rect -1578 434898 1986 435134
rect 2222 434898 37986 435134
rect 38222 434898 73986 435134
rect 74222 434898 109986 435134
rect 110222 434898 145986 435134
rect 146222 434898 156000 435134
rect -2936 434876 156000 434898
rect 440000 435454 586860 435476
rect 440000 435218 469986 435454
rect 470222 435218 505986 435454
rect 506222 435218 541986 435454
rect 542222 435218 577986 435454
rect 578222 435218 585502 435454
rect 585738 435218 586860 435454
rect 440000 435134 586860 435218
rect 440000 434898 469986 435134
rect 470222 434898 505986 435134
rect 506222 434898 541986 435134
rect 542222 434898 577986 435134
rect 578222 434898 585502 435134
rect 585738 434898 586860 435134
rect 440000 434876 586860 434898
rect -1996 434874 -1396 434876
rect 1804 434874 2404 434876
rect 37804 434874 38404 434876
rect 73804 434874 74404 434876
rect 109804 434874 110404 434876
rect 145804 434874 146404 434876
rect 469804 434874 470404 434876
rect 505804 434874 506404 434876
rect 541804 434874 542404 434876
rect 577804 434874 578404 434876
rect 585320 434874 585920 434876
rect -8576 428276 -7976 428278
rect 30604 428276 31204 428278
rect 66604 428276 67204 428278
rect 102604 428276 103204 428278
rect 138604 428276 139204 428278
rect 462604 428276 463204 428278
rect 498604 428276 499204 428278
rect 534604 428276 535204 428278
rect 570604 428276 571204 428278
rect 591900 428276 592500 428278
rect -8576 428254 156000 428276
rect -8576 428018 -8394 428254
rect -8158 428018 30786 428254
rect 31022 428018 66786 428254
rect 67022 428018 102786 428254
rect 103022 428018 138786 428254
rect 139022 428018 156000 428254
rect -8576 427934 156000 428018
rect -8576 427698 -8394 427934
rect -8158 427698 30786 427934
rect 31022 427698 66786 427934
rect 67022 427698 102786 427934
rect 103022 427698 138786 427934
rect 139022 427698 156000 427934
rect -8576 427676 156000 427698
rect 440000 428254 592500 428276
rect 440000 428018 462786 428254
rect 463022 428018 498786 428254
rect 499022 428018 534786 428254
rect 535022 428018 570786 428254
rect 571022 428018 592082 428254
rect 592318 428018 592500 428254
rect 440000 427934 592500 428018
rect 440000 427698 462786 427934
rect 463022 427698 498786 427934
rect 499022 427698 534786 427934
rect 535022 427698 570786 427934
rect 571022 427698 592082 427934
rect 592318 427698 592500 427934
rect 440000 427676 592500 427698
rect -8576 427674 -7976 427676
rect 30604 427674 31204 427676
rect 66604 427674 67204 427676
rect 102604 427674 103204 427676
rect 138604 427674 139204 427676
rect 462604 427674 463204 427676
rect 498604 427674 499204 427676
rect 534604 427674 535204 427676
rect 570604 427674 571204 427676
rect 591900 427674 592500 427676
rect -6696 424676 -6096 424678
rect 27004 424676 27604 424678
rect 63004 424676 63604 424678
rect 99004 424676 99604 424678
rect 135004 424676 135604 424678
rect 459004 424676 459604 424678
rect 495004 424676 495604 424678
rect 531004 424676 531604 424678
rect 567004 424676 567604 424678
rect 590020 424676 590620 424678
rect -6696 424654 156000 424676
rect -6696 424418 -6514 424654
rect -6278 424418 27186 424654
rect 27422 424418 63186 424654
rect 63422 424418 99186 424654
rect 99422 424418 135186 424654
rect 135422 424418 156000 424654
rect -6696 424334 156000 424418
rect -6696 424098 -6514 424334
rect -6278 424098 27186 424334
rect 27422 424098 63186 424334
rect 63422 424098 99186 424334
rect 99422 424098 135186 424334
rect 135422 424098 156000 424334
rect -6696 424076 156000 424098
rect 440000 424654 590620 424676
rect 440000 424418 459186 424654
rect 459422 424418 495186 424654
rect 495422 424418 531186 424654
rect 531422 424418 567186 424654
rect 567422 424418 590202 424654
rect 590438 424418 590620 424654
rect 440000 424334 590620 424418
rect 440000 424098 459186 424334
rect 459422 424098 495186 424334
rect 495422 424098 531186 424334
rect 531422 424098 567186 424334
rect 567422 424098 590202 424334
rect 590438 424098 590620 424334
rect 440000 424076 590620 424098
rect -6696 424074 -6096 424076
rect 27004 424074 27604 424076
rect 63004 424074 63604 424076
rect 99004 424074 99604 424076
rect 135004 424074 135604 424076
rect 459004 424074 459604 424076
rect 495004 424074 495604 424076
rect 531004 424074 531604 424076
rect 567004 424074 567604 424076
rect 590020 424074 590620 424076
rect -4816 421076 -4216 421078
rect 23404 421076 24004 421078
rect 59404 421076 60004 421078
rect 95404 421076 96004 421078
rect 131404 421076 132004 421078
rect 455404 421076 456004 421078
rect 491404 421076 492004 421078
rect 527404 421076 528004 421078
rect 563404 421076 564004 421078
rect 588140 421076 588740 421078
rect -4816 421054 156000 421076
rect -4816 420818 -4634 421054
rect -4398 420818 23586 421054
rect 23822 420818 59586 421054
rect 59822 420818 95586 421054
rect 95822 420818 131586 421054
rect 131822 420818 156000 421054
rect -4816 420734 156000 420818
rect -4816 420498 -4634 420734
rect -4398 420498 23586 420734
rect 23822 420498 59586 420734
rect 59822 420498 95586 420734
rect 95822 420498 131586 420734
rect 131822 420498 156000 420734
rect -4816 420476 156000 420498
rect 440000 421054 588740 421076
rect 440000 420818 455586 421054
rect 455822 420818 491586 421054
rect 491822 420818 527586 421054
rect 527822 420818 563586 421054
rect 563822 420818 588322 421054
rect 588558 420818 588740 421054
rect 440000 420734 588740 420818
rect 440000 420498 455586 420734
rect 455822 420498 491586 420734
rect 491822 420498 527586 420734
rect 527822 420498 563586 420734
rect 563822 420498 588322 420734
rect 588558 420498 588740 420734
rect 440000 420476 588740 420498
rect -4816 420474 -4216 420476
rect 23404 420474 24004 420476
rect 59404 420474 60004 420476
rect 95404 420474 96004 420476
rect 131404 420474 132004 420476
rect 455404 420474 456004 420476
rect 491404 420474 492004 420476
rect 527404 420474 528004 420476
rect 563404 420474 564004 420476
rect 588140 420474 588740 420476
rect -2936 417476 -2336 417478
rect 19804 417476 20404 417478
rect 55804 417476 56404 417478
rect 91804 417476 92404 417478
rect 127804 417476 128404 417478
rect 451804 417476 452404 417478
rect 487804 417476 488404 417478
rect 523804 417476 524404 417478
rect 559804 417476 560404 417478
rect 586260 417476 586860 417478
rect -2936 417454 156000 417476
rect -2936 417218 -2754 417454
rect -2518 417218 19986 417454
rect 20222 417218 55986 417454
rect 56222 417218 91986 417454
rect 92222 417218 127986 417454
rect 128222 417218 156000 417454
rect -2936 417134 156000 417218
rect -2936 416898 -2754 417134
rect -2518 416898 19986 417134
rect 20222 416898 55986 417134
rect 56222 416898 91986 417134
rect 92222 416898 127986 417134
rect 128222 416898 156000 417134
rect -2936 416876 156000 416898
rect 440000 417454 586860 417476
rect 440000 417218 451986 417454
rect 452222 417218 487986 417454
rect 488222 417218 523986 417454
rect 524222 417218 559986 417454
rect 560222 417218 586442 417454
rect 586678 417218 586860 417454
rect 440000 417134 586860 417218
rect 440000 416898 451986 417134
rect 452222 416898 487986 417134
rect 488222 416898 523986 417134
rect 524222 416898 559986 417134
rect 560222 416898 586442 417134
rect 586678 416898 586860 417134
rect 440000 416876 586860 416898
rect -2936 416874 -2336 416876
rect 19804 416874 20404 416876
rect 55804 416874 56404 416876
rect 91804 416874 92404 416876
rect 127804 416874 128404 416876
rect 451804 416874 452404 416876
rect 487804 416874 488404 416876
rect 523804 416874 524404 416876
rect 559804 416874 560404 416876
rect 586260 416874 586860 416876
rect -7636 410276 -7036 410278
rect 12604 410276 13204 410278
rect 48604 410276 49204 410278
rect 84604 410276 85204 410278
rect 120604 410276 121204 410278
rect 444604 410276 445204 410278
rect 480604 410276 481204 410278
rect 516604 410276 517204 410278
rect 552604 410276 553204 410278
rect 590960 410276 591560 410278
rect -8576 410254 156000 410276
rect -8576 410018 -7454 410254
rect -7218 410018 12786 410254
rect 13022 410018 48786 410254
rect 49022 410018 84786 410254
rect 85022 410018 120786 410254
rect 121022 410018 156000 410254
rect -8576 409934 156000 410018
rect -8576 409698 -7454 409934
rect -7218 409698 12786 409934
rect 13022 409698 48786 409934
rect 49022 409698 84786 409934
rect 85022 409698 120786 409934
rect 121022 409698 156000 409934
rect -8576 409676 156000 409698
rect 440000 410254 592500 410276
rect 440000 410018 444786 410254
rect 445022 410018 480786 410254
rect 481022 410018 516786 410254
rect 517022 410018 552786 410254
rect 553022 410018 591142 410254
rect 591378 410018 592500 410254
rect 440000 409934 592500 410018
rect 440000 409698 444786 409934
rect 445022 409698 480786 409934
rect 481022 409698 516786 409934
rect 517022 409698 552786 409934
rect 553022 409698 591142 409934
rect 591378 409698 592500 409934
rect 440000 409676 592500 409698
rect -7636 409674 -7036 409676
rect 12604 409674 13204 409676
rect 48604 409674 49204 409676
rect 84604 409674 85204 409676
rect 120604 409674 121204 409676
rect 444604 409674 445204 409676
rect 480604 409674 481204 409676
rect 516604 409674 517204 409676
rect 552604 409674 553204 409676
rect 590960 409674 591560 409676
rect -5756 406676 -5156 406678
rect 9004 406676 9604 406678
rect 45004 406676 45604 406678
rect 81004 406676 81604 406678
rect 117004 406676 117604 406678
rect 153004 406676 153604 406678
rect 441004 406676 441604 406678
rect 477004 406676 477604 406678
rect 513004 406676 513604 406678
rect 549004 406676 549604 406678
rect 589080 406676 589680 406678
rect -6696 406654 156000 406676
rect -6696 406418 -5574 406654
rect -5338 406418 9186 406654
rect 9422 406418 45186 406654
rect 45422 406418 81186 406654
rect 81422 406418 117186 406654
rect 117422 406418 153186 406654
rect 153422 406418 156000 406654
rect -6696 406334 156000 406418
rect -6696 406098 -5574 406334
rect -5338 406098 9186 406334
rect 9422 406098 45186 406334
rect 45422 406098 81186 406334
rect 81422 406098 117186 406334
rect 117422 406098 153186 406334
rect 153422 406098 156000 406334
rect -6696 406076 156000 406098
rect 440000 406654 590620 406676
rect 440000 406418 441186 406654
rect 441422 406418 477186 406654
rect 477422 406418 513186 406654
rect 513422 406418 549186 406654
rect 549422 406418 589262 406654
rect 589498 406418 590620 406654
rect 440000 406334 590620 406418
rect 440000 406098 441186 406334
rect 441422 406098 477186 406334
rect 477422 406098 513186 406334
rect 513422 406098 549186 406334
rect 549422 406098 589262 406334
rect 589498 406098 590620 406334
rect 440000 406076 590620 406098
rect -5756 406074 -5156 406076
rect 9004 406074 9604 406076
rect 45004 406074 45604 406076
rect 81004 406074 81604 406076
rect 117004 406074 117604 406076
rect 153004 406074 153604 406076
rect 441004 406074 441604 406076
rect 477004 406074 477604 406076
rect 513004 406074 513604 406076
rect 549004 406074 549604 406076
rect 589080 406074 589680 406076
rect -3876 403076 -3276 403078
rect 5404 403076 6004 403078
rect 41404 403076 42004 403078
rect 77404 403076 78004 403078
rect 113404 403076 114004 403078
rect 149404 403076 150004 403078
rect 473404 403076 474004 403078
rect 509404 403076 510004 403078
rect 545404 403076 546004 403078
rect 581404 403076 582004 403078
rect 587200 403076 587800 403078
rect -4816 403054 156000 403076
rect -4816 402818 -3694 403054
rect -3458 402818 5586 403054
rect 5822 402818 41586 403054
rect 41822 402818 77586 403054
rect 77822 402818 113586 403054
rect 113822 402818 149586 403054
rect 149822 402818 156000 403054
rect -4816 402734 156000 402818
rect -4816 402498 -3694 402734
rect -3458 402498 5586 402734
rect 5822 402498 41586 402734
rect 41822 402498 77586 402734
rect 77822 402498 113586 402734
rect 113822 402498 149586 402734
rect 149822 402498 156000 402734
rect -4816 402476 156000 402498
rect 440000 403054 588740 403076
rect 440000 402818 473586 403054
rect 473822 402818 509586 403054
rect 509822 402818 545586 403054
rect 545822 402818 581586 403054
rect 581822 402818 587382 403054
rect 587618 402818 588740 403054
rect 440000 402734 588740 402818
rect 440000 402498 473586 402734
rect 473822 402498 509586 402734
rect 509822 402498 545586 402734
rect 545822 402498 581586 402734
rect 581822 402498 587382 402734
rect 587618 402498 588740 402734
rect 440000 402476 588740 402498
rect -3876 402474 -3276 402476
rect 5404 402474 6004 402476
rect 41404 402474 42004 402476
rect 77404 402474 78004 402476
rect 113404 402474 114004 402476
rect 149404 402474 150004 402476
rect 473404 402474 474004 402476
rect 509404 402474 510004 402476
rect 545404 402474 546004 402476
rect 581404 402474 582004 402476
rect 587200 402474 587800 402476
rect -1996 399476 -1396 399478
rect 1804 399476 2404 399478
rect 37804 399476 38404 399478
rect 73804 399476 74404 399478
rect 109804 399476 110404 399478
rect 145804 399476 146404 399478
rect 469804 399476 470404 399478
rect 505804 399476 506404 399478
rect 541804 399476 542404 399478
rect 577804 399476 578404 399478
rect 585320 399476 585920 399478
rect -2936 399454 156000 399476
rect -2936 399218 -1814 399454
rect -1578 399218 1986 399454
rect 2222 399218 37986 399454
rect 38222 399218 73986 399454
rect 74222 399218 109986 399454
rect 110222 399218 145986 399454
rect 146222 399218 156000 399454
rect -2936 399134 156000 399218
rect -2936 398898 -1814 399134
rect -1578 398898 1986 399134
rect 2222 398898 37986 399134
rect 38222 398898 73986 399134
rect 74222 398898 109986 399134
rect 110222 398898 145986 399134
rect 146222 398898 156000 399134
rect -2936 398876 156000 398898
rect 440000 399454 586860 399476
rect 440000 399218 469986 399454
rect 470222 399218 505986 399454
rect 506222 399218 541986 399454
rect 542222 399218 577986 399454
rect 578222 399218 585502 399454
rect 585738 399218 586860 399454
rect 440000 399134 586860 399218
rect 440000 398898 469986 399134
rect 470222 398898 505986 399134
rect 506222 398898 541986 399134
rect 542222 398898 577986 399134
rect 578222 398898 585502 399134
rect 585738 398898 586860 399134
rect 440000 398876 586860 398898
rect -1996 398874 -1396 398876
rect 1804 398874 2404 398876
rect 37804 398874 38404 398876
rect 73804 398874 74404 398876
rect 109804 398874 110404 398876
rect 145804 398874 146404 398876
rect 469804 398874 470404 398876
rect 505804 398874 506404 398876
rect 541804 398874 542404 398876
rect 577804 398874 578404 398876
rect 585320 398874 585920 398876
rect -8576 392276 -7976 392278
rect 30604 392276 31204 392278
rect 66604 392276 67204 392278
rect 102604 392276 103204 392278
rect 138604 392276 139204 392278
rect 462604 392276 463204 392278
rect 498604 392276 499204 392278
rect 534604 392276 535204 392278
rect 570604 392276 571204 392278
rect 591900 392276 592500 392278
rect -8576 392254 156000 392276
rect -8576 392018 -8394 392254
rect -8158 392018 30786 392254
rect 31022 392018 66786 392254
rect 67022 392018 102786 392254
rect 103022 392018 138786 392254
rect 139022 392018 156000 392254
rect -8576 391934 156000 392018
rect -8576 391698 -8394 391934
rect -8158 391698 30786 391934
rect 31022 391698 66786 391934
rect 67022 391698 102786 391934
rect 103022 391698 138786 391934
rect 139022 391698 156000 391934
rect -8576 391676 156000 391698
rect 440000 392254 592500 392276
rect 440000 392018 462786 392254
rect 463022 392018 498786 392254
rect 499022 392018 534786 392254
rect 535022 392018 570786 392254
rect 571022 392018 592082 392254
rect 592318 392018 592500 392254
rect 440000 391934 592500 392018
rect 440000 391698 462786 391934
rect 463022 391698 498786 391934
rect 499022 391698 534786 391934
rect 535022 391698 570786 391934
rect 571022 391698 592082 391934
rect 592318 391698 592500 391934
rect 440000 391676 592500 391698
rect -8576 391674 -7976 391676
rect 30604 391674 31204 391676
rect 66604 391674 67204 391676
rect 102604 391674 103204 391676
rect 138604 391674 139204 391676
rect 462604 391674 463204 391676
rect 498604 391674 499204 391676
rect 534604 391674 535204 391676
rect 570604 391674 571204 391676
rect 591900 391674 592500 391676
rect -6696 388676 -6096 388678
rect 27004 388676 27604 388678
rect 63004 388676 63604 388678
rect 99004 388676 99604 388678
rect 135004 388676 135604 388678
rect 459004 388676 459604 388678
rect 495004 388676 495604 388678
rect 531004 388676 531604 388678
rect 567004 388676 567604 388678
rect 590020 388676 590620 388678
rect -6696 388654 156000 388676
rect -6696 388418 -6514 388654
rect -6278 388418 27186 388654
rect 27422 388418 63186 388654
rect 63422 388418 99186 388654
rect 99422 388418 135186 388654
rect 135422 388418 156000 388654
rect -6696 388334 156000 388418
rect -6696 388098 -6514 388334
rect -6278 388098 27186 388334
rect 27422 388098 63186 388334
rect 63422 388098 99186 388334
rect 99422 388098 135186 388334
rect 135422 388098 156000 388334
rect -6696 388076 156000 388098
rect 440000 388654 590620 388676
rect 440000 388418 459186 388654
rect 459422 388418 495186 388654
rect 495422 388418 531186 388654
rect 531422 388418 567186 388654
rect 567422 388418 590202 388654
rect 590438 388418 590620 388654
rect 440000 388334 590620 388418
rect 440000 388098 459186 388334
rect 459422 388098 495186 388334
rect 495422 388098 531186 388334
rect 531422 388098 567186 388334
rect 567422 388098 590202 388334
rect 590438 388098 590620 388334
rect 440000 388076 590620 388098
rect -6696 388074 -6096 388076
rect 27004 388074 27604 388076
rect 63004 388074 63604 388076
rect 99004 388074 99604 388076
rect 135004 388074 135604 388076
rect 459004 388074 459604 388076
rect 495004 388074 495604 388076
rect 531004 388074 531604 388076
rect 567004 388074 567604 388076
rect 590020 388074 590620 388076
rect -4816 385076 -4216 385078
rect 23404 385076 24004 385078
rect 59404 385076 60004 385078
rect 95404 385076 96004 385078
rect 131404 385076 132004 385078
rect 455404 385076 456004 385078
rect 491404 385076 492004 385078
rect 527404 385076 528004 385078
rect 563404 385076 564004 385078
rect 588140 385076 588740 385078
rect -4816 385054 156000 385076
rect -4816 384818 -4634 385054
rect -4398 384818 23586 385054
rect 23822 384818 59586 385054
rect 59822 384818 95586 385054
rect 95822 384818 131586 385054
rect 131822 384818 156000 385054
rect -4816 384734 156000 384818
rect -4816 384498 -4634 384734
rect -4398 384498 23586 384734
rect 23822 384498 59586 384734
rect 59822 384498 95586 384734
rect 95822 384498 131586 384734
rect 131822 384498 156000 384734
rect -4816 384476 156000 384498
rect 440000 385054 588740 385076
rect 440000 384818 455586 385054
rect 455822 384818 491586 385054
rect 491822 384818 527586 385054
rect 527822 384818 563586 385054
rect 563822 384818 588322 385054
rect 588558 384818 588740 385054
rect 440000 384734 588740 384818
rect 440000 384498 455586 384734
rect 455822 384498 491586 384734
rect 491822 384498 527586 384734
rect 527822 384498 563586 384734
rect 563822 384498 588322 384734
rect 588558 384498 588740 384734
rect 440000 384476 588740 384498
rect -4816 384474 -4216 384476
rect 23404 384474 24004 384476
rect 59404 384474 60004 384476
rect 95404 384474 96004 384476
rect 131404 384474 132004 384476
rect 455404 384474 456004 384476
rect 491404 384474 492004 384476
rect 527404 384474 528004 384476
rect 563404 384474 564004 384476
rect 588140 384474 588740 384476
rect -2936 381476 -2336 381478
rect 19804 381476 20404 381478
rect 55804 381476 56404 381478
rect 91804 381476 92404 381478
rect 127804 381476 128404 381478
rect 451804 381476 452404 381478
rect 487804 381476 488404 381478
rect 523804 381476 524404 381478
rect 559804 381476 560404 381478
rect 586260 381476 586860 381478
rect -2936 381454 156000 381476
rect -2936 381218 -2754 381454
rect -2518 381218 19986 381454
rect 20222 381218 55986 381454
rect 56222 381218 91986 381454
rect 92222 381218 127986 381454
rect 128222 381218 156000 381454
rect -2936 381134 156000 381218
rect -2936 380898 -2754 381134
rect -2518 380898 19986 381134
rect 20222 380898 55986 381134
rect 56222 380898 91986 381134
rect 92222 380898 127986 381134
rect 128222 380898 156000 381134
rect -2936 380876 156000 380898
rect 440000 381454 586860 381476
rect 440000 381218 451986 381454
rect 452222 381218 487986 381454
rect 488222 381218 523986 381454
rect 524222 381218 559986 381454
rect 560222 381218 586442 381454
rect 586678 381218 586860 381454
rect 440000 381134 586860 381218
rect 440000 380898 451986 381134
rect 452222 380898 487986 381134
rect 488222 380898 523986 381134
rect 524222 380898 559986 381134
rect 560222 380898 586442 381134
rect 586678 380898 586860 381134
rect 440000 380876 586860 380898
rect -2936 380874 -2336 380876
rect 19804 380874 20404 380876
rect 55804 380874 56404 380876
rect 91804 380874 92404 380876
rect 127804 380874 128404 380876
rect 451804 380874 452404 380876
rect 487804 380874 488404 380876
rect 523804 380874 524404 380876
rect 559804 380874 560404 380876
rect 586260 380874 586860 380876
rect -7636 374276 -7036 374278
rect 12604 374276 13204 374278
rect 48604 374276 49204 374278
rect 84604 374276 85204 374278
rect 120604 374276 121204 374278
rect 444604 374276 445204 374278
rect 480604 374276 481204 374278
rect 516604 374276 517204 374278
rect 552604 374276 553204 374278
rect 590960 374276 591560 374278
rect -8576 374254 156000 374276
rect -8576 374018 -7454 374254
rect -7218 374018 12786 374254
rect 13022 374018 48786 374254
rect 49022 374018 84786 374254
rect 85022 374018 120786 374254
rect 121022 374018 156000 374254
rect -8576 373934 156000 374018
rect -8576 373698 -7454 373934
rect -7218 373698 12786 373934
rect 13022 373698 48786 373934
rect 49022 373698 84786 373934
rect 85022 373698 120786 373934
rect 121022 373698 156000 373934
rect -8576 373676 156000 373698
rect 440000 374254 592500 374276
rect 440000 374018 444786 374254
rect 445022 374018 480786 374254
rect 481022 374018 516786 374254
rect 517022 374018 552786 374254
rect 553022 374018 591142 374254
rect 591378 374018 592500 374254
rect 440000 373934 592500 374018
rect 440000 373698 444786 373934
rect 445022 373698 480786 373934
rect 481022 373698 516786 373934
rect 517022 373698 552786 373934
rect 553022 373698 591142 373934
rect 591378 373698 592500 373934
rect 440000 373676 592500 373698
rect -7636 373674 -7036 373676
rect 12604 373674 13204 373676
rect 48604 373674 49204 373676
rect 84604 373674 85204 373676
rect 120604 373674 121204 373676
rect 444604 373674 445204 373676
rect 480604 373674 481204 373676
rect 516604 373674 517204 373676
rect 552604 373674 553204 373676
rect 590960 373674 591560 373676
rect -5756 370676 -5156 370678
rect 9004 370676 9604 370678
rect 45004 370676 45604 370678
rect 81004 370676 81604 370678
rect 117004 370676 117604 370678
rect 153004 370676 153604 370678
rect 441004 370676 441604 370678
rect 477004 370676 477604 370678
rect 513004 370676 513604 370678
rect 549004 370676 549604 370678
rect 589080 370676 589680 370678
rect -6696 370654 156000 370676
rect -6696 370418 -5574 370654
rect -5338 370418 9186 370654
rect 9422 370418 45186 370654
rect 45422 370418 81186 370654
rect 81422 370418 117186 370654
rect 117422 370418 153186 370654
rect 153422 370418 156000 370654
rect -6696 370334 156000 370418
rect -6696 370098 -5574 370334
rect -5338 370098 9186 370334
rect 9422 370098 45186 370334
rect 45422 370098 81186 370334
rect 81422 370098 117186 370334
rect 117422 370098 153186 370334
rect 153422 370098 156000 370334
rect -6696 370076 156000 370098
rect 440000 370654 590620 370676
rect 440000 370418 441186 370654
rect 441422 370418 477186 370654
rect 477422 370418 513186 370654
rect 513422 370418 549186 370654
rect 549422 370418 589262 370654
rect 589498 370418 590620 370654
rect 440000 370334 590620 370418
rect 440000 370098 441186 370334
rect 441422 370098 477186 370334
rect 477422 370098 513186 370334
rect 513422 370098 549186 370334
rect 549422 370098 589262 370334
rect 589498 370098 590620 370334
rect 440000 370076 590620 370098
rect -5756 370074 -5156 370076
rect 9004 370074 9604 370076
rect 45004 370074 45604 370076
rect 81004 370074 81604 370076
rect 117004 370074 117604 370076
rect 153004 370074 153604 370076
rect 441004 370074 441604 370076
rect 477004 370074 477604 370076
rect 513004 370074 513604 370076
rect 549004 370074 549604 370076
rect 589080 370074 589680 370076
rect -3876 367076 -3276 367078
rect 5404 367076 6004 367078
rect 41404 367076 42004 367078
rect 77404 367076 78004 367078
rect 113404 367076 114004 367078
rect 149404 367076 150004 367078
rect 473404 367076 474004 367078
rect 509404 367076 510004 367078
rect 545404 367076 546004 367078
rect 581404 367076 582004 367078
rect 587200 367076 587800 367078
rect -4816 367054 156000 367076
rect -4816 366818 -3694 367054
rect -3458 366818 5586 367054
rect 5822 366818 41586 367054
rect 41822 366818 77586 367054
rect 77822 366818 113586 367054
rect 113822 366818 149586 367054
rect 149822 366818 156000 367054
rect -4816 366734 156000 366818
rect -4816 366498 -3694 366734
rect -3458 366498 5586 366734
rect 5822 366498 41586 366734
rect 41822 366498 77586 366734
rect 77822 366498 113586 366734
rect 113822 366498 149586 366734
rect 149822 366498 156000 366734
rect -4816 366476 156000 366498
rect 440000 367054 588740 367076
rect 440000 366818 473586 367054
rect 473822 366818 509586 367054
rect 509822 366818 545586 367054
rect 545822 366818 581586 367054
rect 581822 366818 587382 367054
rect 587618 366818 588740 367054
rect 440000 366734 588740 366818
rect 440000 366498 473586 366734
rect 473822 366498 509586 366734
rect 509822 366498 545586 366734
rect 545822 366498 581586 366734
rect 581822 366498 587382 366734
rect 587618 366498 588740 366734
rect 440000 366476 588740 366498
rect -3876 366474 -3276 366476
rect 5404 366474 6004 366476
rect 41404 366474 42004 366476
rect 77404 366474 78004 366476
rect 113404 366474 114004 366476
rect 149404 366474 150004 366476
rect 473404 366474 474004 366476
rect 509404 366474 510004 366476
rect 545404 366474 546004 366476
rect 581404 366474 582004 366476
rect 587200 366474 587800 366476
rect -1996 363476 -1396 363478
rect 1804 363476 2404 363478
rect 37804 363476 38404 363478
rect 73804 363476 74404 363478
rect 109804 363476 110404 363478
rect 145804 363476 146404 363478
rect 469804 363476 470404 363478
rect 505804 363476 506404 363478
rect 541804 363476 542404 363478
rect 577804 363476 578404 363478
rect 585320 363476 585920 363478
rect -2936 363454 156000 363476
rect -2936 363218 -1814 363454
rect -1578 363218 1986 363454
rect 2222 363218 37986 363454
rect 38222 363218 73986 363454
rect 74222 363218 109986 363454
rect 110222 363218 145986 363454
rect 146222 363218 156000 363454
rect -2936 363134 156000 363218
rect -2936 362898 -1814 363134
rect -1578 362898 1986 363134
rect 2222 362898 37986 363134
rect 38222 362898 73986 363134
rect 74222 362898 109986 363134
rect 110222 362898 145986 363134
rect 146222 362898 156000 363134
rect -2936 362876 156000 362898
rect 440000 363454 586860 363476
rect 440000 363218 469986 363454
rect 470222 363218 505986 363454
rect 506222 363218 541986 363454
rect 542222 363218 577986 363454
rect 578222 363218 585502 363454
rect 585738 363218 586860 363454
rect 440000 363134 586860 363218
rect 440000 362898 469986 363134
rect 470222 362898 505986 363134
rect 506222 362898 541986 363134
rect 542222 362898 577986 363134
rect 578222 362898 585502 363134
rect 585738 362898 586860 363134
rect 440000 362876 586860 362898
rect -1996 362874 -1396 362876
rect 1804 362874 2404 362876
rect 37804 362874 38404 362876
rect 73804 362874 74404 362876
rect 109804 362874 110404 362876
rect 145804 362874 146404 362876
rect 469804 362874 470404 362876
rect 505804 362874 506404 362876
rect 541804 362874 542404 362876
rect 577804 362874 578404 362876
rect 585320 362874 585920 362876
rect -8576 356276 -7976 356278
rect 30604 356276 31204 356278
rect 66604 356276 67204 356278
rect 102604 356276 103204 356278
rect 138604 356276 139204 356278
rect 462604 356276 463204 356278
rect 498604 356276 499204 356278
rect 534604 356276 535204 356278
rect 570604 356276 571204 356278
rect 591900 356276 592500 356278
rect -8576 356254 156000 356276
rect -8576 356018 -8394 356254
rect -8158 356018 30786 356254
rect 31022 356018 66786 356254
rect 67022 356018 102786 356254
rect 103022 356018 138786 356254
rect 139022 356018 156000 356254
rect -8576 355934 156000 356018
rect -8576 355698 -8394 355934
rect -8158 355698 30786 355934
rect 31022 355698 66786 355934
rect 67022 355698 102786 355934
rect 103022 355698 138786 355934
rect 139022 355698 156000 355934
rect -8576 355676 156000 355698
rect 440000 356254 592500 356276
rect 440000 356018 462786 356254
rect 463022 356018 498786 356254
rect 499022 356018 534786 356254
rect 535022 356018 570786 356254
rect 571022 356018 592082 356254
rect 592318 356018 592500 356254
rect 440000 355934 592500 356018
rect 440000 355698 462786 355934
rect 463022 355698 498786 355934
rect 499022 355698 534786 355934
rect 535022 355698 570786 355934
rect 571022 355698 592082 355934
rect 592318 355698 592500 355934
rect 440000 355676 592500 355698
rect -8576 355674 -7976 355676
rect 30604 355674 31204 355676
rect 66604 355674 67204 355676
rect 102604 355674 103204 355676
rect 138604 355674 139204 355676
rect 462604 355674 463204 355676
rect 498604 355674 499204 355676
rect 534604 355674 535204 355676
rect 570604 355674 571204 355676
rect 591900 355674 592500 355676
rect -6696 352676 -6096 352678
rect 27004 352676 27604 352678
rect 63004 352676 63604 352678
rect 99004 352676 99604 352678
rect 135004 352676 135604 352678
rect 459004 352676 459604 352678
rect 495004 352676 495604 352678
rect 531004 352676 531604 352678
rect 567004 352676 567604 352678
rect 590020 352676 590620 352678
rect -6696 352654 156000 352676
rect -6696 352418 -6514 352654
rect -6278 352418 27186 352654
rect 27422 352418 63186 352654
rect 63422 352418 99186 352654
rect 99422 352418 135186 352654
rect 135422 352418 156000 352654
rect -6696 352334 156000 352418
rect -6696 352098 -6514 352334
rect -6278 352098 27186 352334
rect 27422 352098 63186 352334
rect 63422 352098 99186 352334
rect 99422 352098 135186 352334
rect 135422 352098 156000 352334
rect -6696 352076 156000 352098
rect 440000 352654 590620 352676
rect 440000 352418 459186 352654
rect 459422 352418 495186 352654
rect 495422 352418 531186 352654
rect 531422 352418 567186 352654
rect 567422 352418 590202 352654
rect 590438 352418 590620 352654
rect 440000 352334 590620 352418
rect 440000 352098 459186 352334
rect 459422 352098 495186 352334
rect 495422 352098 531186 352334
rect 531422 352098 567186 352334
rect 567422 352098 590202 352334
rect 590438 352098 590620 352334
rect 440000 352076 590620 352098
rect -6696 352074 -6096 352076
rect 27004 352074 27604 352076
rect 63004 352074 63604 352076
rect 99004 352074 99604 352076
rect 135004 352074 135604 352076
rect 459004 352074 459604 352076
rect 495004 352074 495604 352076
rect 531004 352074 531604 352076
rect 567004 352074 567604 352076
rect 590020 352074 590620 352076
rect -4816 349076 -4216 349078
rect 23404 349076 24004 349078
rect 59404 349076 60004 349078
rect 95404 349076 96004 349078
rect 131404 349076 132004 349078
rect 455404 349076 456004 349078
rect 491404 349076 492004 349078
rect 527404 349076 528004 349078
rect 563404 349076 564004 349078
rect 588140 349076 588740 349078
rect -4816 349054 156000 349076
rect -4816 348818 -4634 349054
rect -4398 348818 23586 349054
rect 23822 348818 59586 349054
rect 59822 348818 95586 349054
rect 95822 348818 131586 349054
rect 131822 348818 156000 349054
rect -4816 348734 156000 348818
rect -4816 348498 -4634 348734
rect -4398 348498 23586 348734
rect 23822 348498 59586 348734
rect 59822 348498 95586 348734
rect 95822 348498 131586 348734
rect 131822 348498 156000 348734
rect -4816 348476 156000 348498
rect 440000 349054 588740 349076
rect 440000 348818 455586 349054
rect 455822 348818 491586 349054
rect 491822 348818 527586 349054
rect 527822 348818 563586 349054
rect 563822 348818 588322 349054
rect 588558 348818 588740 349054
rect 440000 348734 588740 348818
rect 440000 348498 455586 348734
rect 455822 348498 491586 348734
rect 491822 348498 527586 348734
rect 527822 348498 563586 348734
rect 563822 348498 588322 348734
rect 588558 348498 588740 348734
rect 440000 348476 588740 348498
rect -4816 348474 -4216 348476
rect 23404 348474 24004 348476
rect 59404 348474 60004 348476
rect 95404 348474 96004 348476
rect 131404 348474 132004 348476
rect 455404 348474 456004 348476
rect 491404 348474 492004 348476
rect 527404 348474 528004 348476
rect 563404 348474 564004 348476
rect 588140 348474 588740 348476
rect -2936 345476 -2336 345478
rect 19804 345476 20404 345478
rect 55804 345476 56404 345478
rect 91804 345476 92404 345478
rect 127804 345476 128404 345478
rect 451804 345476 452404 345478
rect 487804 345476 488404 345478
rect 523804 345476 524404 345478
rect 559804 345476 560404 345478
rect 586260 345476 586860 345478
rect -2936 345454 156000 345476
rect -2936 345218 -2754 345454
rect -2518 345218 19986 345454
rect 20222 345218 55986 345454
rect 56222 345218 91986 345454
rect 92222 345218 127986 345454
rect 128222 345218 156000 345454
rect -2936 345134 156000 345218
rect -2936 344898 -2754 345134
rect -2518 344898 19986 345134
rect 20222 344898 55986 345134
rect 56222 344898 91986 345134
rect 92222 344898 127986 345134
rect 128222 344898 156000 345134
rect -2936 344876 156000 344898
rect 440000 345454 586860 345476
rect 440000 345218 451986 345454
rect 452222 345218 487986 345454
rect 488222 345218 523986 345454
rect 524222 345218 559986 345454
rect 560222 345218 586442 345454
rect 586678 345218 586860 345454
rect 440000 345134 586860 345218
rect 440000 344898 451986 345134
rect 452222 344898 487986 345134
rect 488222 344898 523986 345134
rect 524222 344898 559986 345134
rect 560222 344898 586442 345134
rect 586678 344898 586860 345134
rect 440000 344876 586860 344898
rect -2936 344874 -2336 344876
rect 19804 344874 20404 344876
rect 55804 344874 56404 344876
rect 91804 344874 92404 344876
rect 127804 344874 128404 344876
rect 451804 344874 452404 344876
rect 487804 344874 488404 344876
rect 523804 344874 524404 344876
rect 559804 344874 560404 344876
rect 586260 344874 586860 344876
rect -7636 338276 -7036 338278
rect 12604 338276 13204 338278
rect 48604 338276 49204 338278
rect 84604 338276 85204 338278
rect 120604 338276 121204 338278
rect 444604 338276 445204 338278
rect 480604 338276 481204 338278
rect 516604 338276 517204 338278
rect 552604 338276 553204 338278
rect 590960 338276 591560 338278
rect -8576 338254 156000 338276
rect -8576 338018 -7454 338254
rect -7218 338018 12786 338254
rect 13022 338018 48786 338254
rect 49022 338018 84786 338254
rect 85022 338018 120786 338254
rect 121022 338018 156000 338254
rect -8576 337934 156000 338018
rect -8576 337698 -7454 337934
rect -7218 337698 12786 337934
rect 13022 337698 48786 337934
rect 49022 337698 84786 337934
rect 85022 337698 120786 337934
rect 121022 337698 156000 337934
rect -8576 337676 156000 337698
rect 440000 338254 592500 338276
rect 440000 338018 444786 338254
rect 445022 338018 480786 338254
rect 481022 338018 516786 338254
rect 517022 338018 552786 338254
rect 553022 338018 591142 338254
rect 591378 338018 592500 338254
rect 440000 337934 592500 338018
rect 440000 337698 444786 337934
rect 445022 337698 480786 337934
rect 481022 337698 516786 337934
rect 517022 337698 552786 337934
rect 553022 337698 591142 337934
rect 591378 337698 592500 337934
rect 440000 337676 592500 337698
rect -7636 337674 -7036 337676
rect 12604 337674 13204 337676
rect 48604 337674 49204 337676
rect 84604 337674 85204 337676
rect 120604 337674 121204 337676
rect 444604 337674 445204 337676
rect 480604 337674 481204 337676
rect 516604 337674 517204 337676
rect 552604 337674 553204 337676
rect 590960 337674 591560 337676
rect -5756 334676 -5156 334678
rect 9004 334676 9604 334678
rect 45004 334676 45604 334678
rect 81004 334676 81604 334678
rect 117004 334676 117604 334678
rect 153004 334676 153604 334678
rect 441004 334676 441604 334678
rect 477004 334676 477604 334678
rect 513004 334676 513604 334678
rect 549004 334676 549604 334678
rect 589080 334676 589680 334678
rect -6696 334654 156000 334676
rect -6696 334418 -5574 334654
rect -5338 334418 9186 334654
rect 9422 334418 45186 334654
rect 45422 334418 81186 334654
rect 81422 334418 117186 334654
rect 117422 334418 153186 334654
rect 153422 334418 156000 334654
rect -6696 334334 156000 334418
rect -6696 334098 -5574 334334
rect -5338 334098 9186 334334
rect 9422 334098 45186 334334
rect 45422 334098 81186 334334
rect 81422 334098 117186 334334
rect 117422 334098 153186 334334
rect 153422 334098 156000 334334
rect -6696 334076 156000 334098
rect 440000 334654 590620 334676
rect 440000 334418 441186 334654
rect 441422 334418 477186 334654
rect 477422 334418 513186 334654
rect 513422 334418 549186 334654
rect 549422 334418 589262 334654
rect 589498 334418 590620 334654
rect 440000 334334 590620 334418
rect 440000 334098 441186 334334
rect 441422 334098 477186 334334
rect 477422 334098 513186 334334
rect 513422 334098 549186 334334
rect 549422 334098 589262 334334
rect 589498 334098 590620 334334
rect 440000 334076 590620 334098
rect -5756 334074 -5156 334076
rect 9004 334074 9604 334076
rect 45004 334074 45604 334076
rect 81004 334074 81604 334076
rect 117004 334074 117604 334076
rect 153004 334074 153604 334076
rect 441004 334074 441604 334076
rect 477004 334074 477604 334076
rect 513004 334074 513604 334076
rect 549004 334074 549604 334076
rect 589080 334074 589680 334076
rect -3876 331076 -3276 331078
rect 5404 331076 6004 331078
rect 41404 331076 42004 331078
rect 77404 331076 78004 331078
rect 113404 331076 114004 331078
rect 149404 331076 150004 331078
rect 473404 331076 474004 331078
rect 509404 331076 510004 331078
rect 545404 331076 546004 331078
rect 581404 331076 582004 331078
rect 587200 331076 587800 331078
rect -4816 331054 156000 331076
rect -4816 330818 -3694 331054
rect -3458 330818 5586 331054
rect 5822 330818 41586 331054
rect 41822 330818 77586 331054
rect 77822 330818 113586 331054
rect 113822 330818 149586 331054
rect 149822 330818 156000 331054
rect -4816 330734 156000 330818
rect -4816 330498 -3694 330734
rect -3458 330498 5586 330734
rect 5822 330498 41586 330734
rect 41822 330498 77586 330734
rect 77822 330498 113586 330734
rect 113822 330498 149586 330734
rect 149822 330498 156000 330734
rect -4816 330476 156000 330498
rect 440000 331054 588740 331076
rect 440000 330818 473586 331054
rect 473822 330818 509586 331054
rect 509822 330818 545586 331054
rect 545822 330818 581586 331054
rect 581822 330818 587382 331054
rect 587618 330818 588740 331054
rect 440000 330734 588740 330818
rect 440000 330498 473586 330734
rect 473822 330498 509586 330734
rect 509822 330498 545586 330734
rect 545822 330498 581586 330734
rect 581822 330498 587382 330734
rect 587618 330498 588740 330734
rect 440000 330476 588740 330498
rect -3876 330474 -3276 330476
rect 5404 330474 6004 330476
rect 41404 330474 42004 330476
rect 77404 330474 78004 330476
rect 113404 330474 114004 330476
rect 149404 330474 150004 330476
rect 473404 330474 474004 330476
rect 509404 330474 510004 330476
rect 545404 330474 546004 330476
rect 581404 330474 582004 330476
rect 587200 330474 587800 330476
rect -1996 327476 -1396 327478
rect 1804 327476 2404 327478
rect 37804 327476 38404 327478
rect 73804 327476 74404 327478
rect 109804 327476 110404 327478
rect 145804 327476 146404 327478
rect 469804 327476 470404 327478
rect 505804 327476 506404 327478
rect 541804 327476 542404 327478
rect 577804 327476 578404 327478
rect 585320 327476 585920 327478
rect -2936 327454 156000 327476
rect -2936 327218 -1814 327454
rect -1578 327218 1986 327454
rect 2222 327218 37986 327454
rect 38222 327218 73986 327454
rect 74222 327218 109986 327454
rect 110222 327218 145986 327454
rect 146222 327218 156000 327454
rect -2936 327134 156000 327218
rect -2936 326898 -1814 327134
rect -1578 326898 1986 327134
rect 2222 326898 37986 327134
rect 38222 326898 73986 327134
rect 74222 326898 109986 327134
rect 110222 326898 145986 327134
rect 146222 326898 156000 327134
rect -2936 326876 156000 326898
rect 440000 327454 586860 327476
rect 440000 327218 469986 327454
rect 470222 327218 505986 327454
rect 506222 327218 541986 327454
rect 542222 327218 577986 327454
rect 578222 327218 585502 327454
rect 585738 327218 586860 327454
rect 440000 327134 586860 327218
rect 440000 326898 469986 327134
rect 470222 326898 505986 327134
rect 506222 326898 541986 327134
rect 542222 326898 577986 327134
rect 578222 326898 585502 327134
rect 585738 326898 586860 327134
rect 440000 326876 586860 326898
rect -1996 326874 -1396 326876
rect 1804 326874 2404 326876
rect 37804 326874 38404 326876
rect 73804 326874 74404 326876
rect 109804 326874 110404 326876
rect 145804 326874 146404 326876
rect 469804 326874 470404 326876
rect 505804 326874 506404 326876
rect 541804 326874 542404 326876
rect 577804 326874 578404 326876
rect 585320 326874 585920 326876
rect -8576 320276 -7976 320278
rect 30604 320276 31204 320278
rect 66604 320276 67204 320278
rect 102604 320276 103204 320278
rect 138604 320276 139204 320278
rect 174604 320276 175204 320278
rect 210604 320276 211204 320278
rect 246604 320276 247204 320278
rect 282604 320276 283204 320278
rect 318604 320276 319204 320278
rect 354604 320276 355204 320278
rect 390604 320276 391204 320278
rect 426604 320276 427204 320278
rect 462604 320276 463204 320278
rect 498604 320276 499204 320278
rect 534604 320276 535204 320278
rect 570604 320276 571204 320278
rect 591900 320276 592500 320278
rect -8576 320254 592500 320276
rect -8576 320018 -8394 320254
rect -8158 320018 30786 320254
rect 31022 320018 66786 320254
rect 67022 320018 102786 320254
rect 103022 320018 138786 320254
rect 139022 320018 174786 320254
rect 175022 320018 210786 320254
rect 211022 320018 246786 320254
rect 247022 320018 282786 320254
rect 283022 320018 318786 320254
rect 319022 320018 354786 320254
rect 355022 320018 390786 320254
rect 391022 320018 426786 320254
rect 427022 320018 462786 320254
rect 463022 320018 498786 320254
rect 499022 320018 534786 320254
rect 535022 320018 570786 320254
rect 571022 320018 592082 320254
rect 592318 320018 592500 320254
rect -8576 319934 592500 320018
rect -8576 319698 -8394 319934
rect -8158 319698 30786 319934
rect 31022 319698 66786 319934
rect 67022 319698 102786 319934
rect 103022 319698 138786 319934
rect 139022 319698 174786 319934
rect 175022 319698 210786 319934
rect 211022 319698 246786 319934
rect 247022 319698 282786 319934
rect 283022 319698 318786 319934
rect 319022 319698 354786 319934
rect 355022 319698 390786 319934
rect 391022 319698 426786 319934
rect 427022 319698 462786 319934
rect 463022 319698 498786 319934
rect 499022 319698 534786 319934
rect 535022 319698 570786 319934
rect 571022 319698 592082 319934
rect 592318 319698 592500 319934
rect -8576 319676 592500 319698
rect -8576 319674 -7976 319676
rect 30604 319674 31204 319676
rect 66604 319674 67204 319676
rect 102604 319674 103204 319676
rect 138604 319674 139204 319676
rect 174604 319674 175204 319676
rect 210604 319674 211204 319676
rect 246604 319674 247204 319676
rect 282604 319674 283204 319676
rect 318604 319674 319204 319676
rect 354604 319674 355204 319676
rect 390604 319674 391204 319676
rect 426604 319674 427204 319676
rect 462604 319674 463204 319676
rect 498604 319674 499204 319676
rect 534604 319674 535204 319676
rect 570604 319674 571204 319676
rect 591900 319674 592500 319676
rect -6696 316676 -6096 316678
rect 27004 316676 27604 316678
rect 63004 316676 63604 316678
rect 99004 316676 99604 316678
rect 135004 316676 135604 316678
rect 171004 316676 171604 316678
rect 207004 316676 207604 316678
rect 243004 316676 243604 316678
rect 279004 316676 279604 316678
rect 315004 316676 315604 316678
rect 351004 316676 351604 316678
rect 387004 316676 387604 316678
rect 423004 316676 423604 316678
rect 459004 316676 459604 316678
rect 495004 316676 495604 316678
rect 531004 316676 531604 316678
rect 567004 316676 567604 316678
rect 590020 316676 590620 316678
rect -6696 316654 590620 316676
rect -6696 316418 -6514 316654
rect -6278 316418 27186 316654
rect 27422 316418 63186 316654
rect 63422 316418 99186 316654
rect 99422 316418 135186 316654
rect 135422 316418 171186 316654
rect 171422 316418 207186 316654
rect 207422 316418 243186 316654
rect 243422 316418 279186 316654
rect 279422 316418 315186 316654
rect 315422 316418 351186 316654
rect 351422 316418 387186 316654
rect 387422 316418 423186 316654
rect 423422 316418 459186 316654
rect 459422 316418 495186 316654
rect 495422 316418 531186 316654
rect 531422 316418 567186 316654
rect 567422 316418 590202 316654
rect 590438 316418 590620 316654
rect -6696 316334 590620 316418
rect -6696 316098 -6514 316334
rect -6278 316098 27186 316334
rect 27422 316098 63186 316334
rect 63422 316098 99186 316334
rect 99422 316098 135186 316334
rect 135422 316098 171186 316334
rect 171422 316098 207186 316334
rect 207422 316098 243186 316334
rect 243422 316098 279186 316334
rect 279422 316098 315186 316334
rect 315422 316098 351186 316334
rect 351422 316098 387186 316334
rect 387422 316098 423186 316334
rect 423422 316098 459186 316334
rect 459422 316098 495186 316334
rect 495422 316098 531186 316334
rect 531422 316098 567186 316334
rect 567422 316098 590202 316334
rect 590438 316098 590620 316334
rect -6696 316076 590620 316098
rect -6696 316074 -6096 316076
rect 27004 316074 27604 316076
rect 63004 316074 63604 316076
rect 99004 316074 99604 316076
rect 135004 316074 135604 316076
rect 171004 316074 171604 316076
rect 207004 316074 207604 316076
rect 243004 316074 243604 316076
rect 279004 316074 279604 316076
rect 315004 316074 315604 316076
rect 351004 316074 351604 316076
rect 387004 316074 387604 316076
rect 423004 316074 423604 316076
rect 459004 316074 459604 316076
rect 495004 316074 495604 316076
rect 531004 316074 531604 316076
rect 567004 316074 567604 316076
rect 590020 316074 590620 316076
rect -4816 313076 -4216 313078
rect 23404 313076 24004 313078
rect 59404 313076 60004 313078
rect 95404 313076 96004 313078
rect 131404 313076 132004 313078
rect 167404 313076 168004 313078
rect 203404 313076 204004 313078
rect 239404 313076 240004 313078
rect 275404 313076 276004 313078
rect 311404 313076 312004 313078
rect 347404 313076 348004 313078
rect 383404 313076 384004 313078
rect 419404 313076 420004 313078
rect 455404 313076 456004 313078
rect 491404 313076 492004 313078
rect 527404 313076 528004 313078
rect 563404 313076 564004 313078
rect 588140 313076 588740 313078
rect -4816 313054 588740 313076
rect -4816 312818 -4634 313054
rect -4398 312818 23586 313054
rect 23822 312818 59586 313054
rect 59822 312818 95586 313054
rect 95822 312818 131586 313054
rect 131822 312818 167586 313054
rect 167822 312818 203586 313054
rect 203822 312818 239586 313054
rect 239822 312818 275586 313054
rect 275822 312818 311586 313054
rect 311822 312818 347586 313054
rect 347822 312818 383586 313054
rect 383822 312818 419586 313054
rect 419822 312818 455586 313054
rect 455822 312818 491586 313054
rect 491822 312818 527586 313054
rect 527822 312818 563586 313054
rect 563822 312818 588322 313054
rect 588558 312818 588740 313054
rect -4816 312734 588740 312818
rect -4816 312498 -4634 312734
rect -4398 312498 23586 312734
rect 23822 312498 59586 312734
rect 59822 312498 95586 312734
rect 95822 312498 131586 312734
rect 131822 312498 167586 312734
rect 167822 312498 203586 312734
rect 203822 312498 239586 312734
rect 239822 312498 275586 312734
rect 275822 312498 311586 312734
rect 311822 312498 347586 312734
rect 347822 312498 383586 312734
rect 383822 312498 419586 312734
rect 419822 312498 455586 312734
rect 455822 312498 491586 312734
rect 491822 312498 527586 312734
rect 527822 312498 563586 312734
rect 563822 312498 588322 312734
rect 588558 312498 588740 312734
rect -4816 312476 588740 312498
rect -4816 312474 -4216 312476
rect 23404 312474 24004 312476
rect 59404 312474 60004 312476
rect 95404 312474 96004 312476
rect 131404 312474 132004 312476
rect 167404 312474 168004 312476
rect 203404 312474 204004 312476
rect 239404 312474 240004 312476
rect 275404 312474 276004 312476
rect 311404 312474 312004 312476
rect 347404 312474 348004 312476
rect 383404 312474 384004 312476
rect 419404 312474 420004 312476
rect 455404 312474 456004 312476
rect 491404 312474 492004 312476
rect 527404 312474 528004 312476
rect 563404 312474 564004 312476
rect 588140 312474 588740 312476
rect -2936 309476 -2336 309478
rect 19804 309476 20404 309478
rect 55804 309476 56404 309478
rect 91804 309476 92404 309478
rect 127804 309476 128404 309478
rect 163804 309476 164404 309478
rect 199804 309476 200404 309478
rect 235804 309476 236404 309478
rect 271804 309476 272404 309478
rect 307804 309476 308404 309478
rect 343804 309476 344404 309478
rect 379804 309476 380404 309478
rect 415804 309476 416404 309478
rect 451804 309476 452404 309478
rect 487804 309476 488404 309478
rect 523804 309476 524404 309478
rect 559804 309476 560404 309478
rect 586260 309476 586860 309478
rect -2936 309454 586860 309476
rect -2936 309218 -2754 309454
rect -2518 309218 19986 309454
rect 20222 309218 55986 309454
rect 56222 309218 91986 309454
rect 92222 309218 127986 309454
rect 128222 309218 163986 309454
rect 164222 309218 199986 309454
rect 200222 309218 235986 309454
rect 236222 309218 271986 309454
rect 272222 309218 307986 309454
rect 308222 309218 343986 309454
rect 344222 309218 379986 309454
rect 380222 309218 415986 309454
rect 416222 309218 451986 309454
rect 452222 309218 487986 309454
rect 488222 309218 523986 309454
rect 524222 309218 559986 309454
rect 560222 309218 586442 309454
rect 586678 309218 586860 309454
rect -2936 309134 586860 309218
rect -2936 308898 -2754 309134
rect -2518 308898 19986 309134
rect 20222 308898 55986 309134
rect 56222 308898 91986 309134
rect 92222 308898 127986 309134
rect 128222 308898 163986 309134
rect 164222 308898 199986 309134
rect 200222 308898 235986 309134
rect 236222 308898 271986 309134
rect 272222 308898 307986 309134
rect 308222 308898 343986 309134
rect 344222 308898 379986 309134
rect 380222 308898 415986 309134
rect 416222 308898 451986 309134
rect 452222 308898 487986 309134
rect 488222 308898 523986 309134
rect 524222 308898 559986 309134
rect 560222 308898 586442 309134
rect 586678 308898 586860 309134
rect -2936 308876 586860 308898
rect -2936 308874 -2336 308876
rect 19804 308874 20404 308876
rect 55804 308874 56404 308876
rect 91804 308874 92404 308876
rect 127804 308874 128404 308876
rect 163804 308874 164404 308876
rect 199804 308874 200404 308876
rect 235804 308874 236404 308876
rect 271804 308874 272404 308876
rect 307804 308874 308404 308876
rect 343804 308874 344404 308876
rect 379804 308874 380404 308876
rect 415804 308874 416404 308876
rect 451804 308874 452404 308876
rect 487804 308874 488404 308876
rect 523804 308874 524404 308876
rect 559804 308874 560404 308876
rect 586260 308874 586860 308876
rect -7636 302276 -7036 302278
rect 12604 302276 13204 302278
rect 48604 302276 49204 302278
rect 84604 302276 85204 302278
rect 120604 302276 121204 302278
rect 156604 302276 157204 302278
rect 192604 302276 193204 302278
rect 228604 302276 229204 302278
rect 264604 302276 265204 302278
rect 300604 302276 301204 302278
rect 336604 302276 337204 302278
rect 372604 302276 373204 302278
rect 408604 302276 409204 302278
rect 444604 302276 445204 302278
rect 480604 302276 481204 302278
rect 516604 302276 517204 302278
rect 552604 302276 553204 302278
rect 590960 302276 591560 302278
rect -8576 302254 592500 302276
rect -8576 302018 -7454 302254
rect -7218 302018 12786 302254
rect 13022 302018 48786 302254
rect 49022 302018 84786 302254
rect 85022 302018 120786 302254
rect 121022 302018 156786 302254
rect 157022 302018 192786 302254
rect 193022 302018 228786 302254
rect 229022 302018 264786 302254
rect 265022 302018 300786 302254
rect 301022 302018 336786 302254
rect 337022 302018 372786 302254
rect 373022 302018 408786 302254
rect 409022 302018 444786 302254
rect 445022 302018 480786 302254
rect 481022 302018 516786 302254
rect 517022 302018 552786 302254
rect 553022 302018 591142 302254
rect 591378 302018 592500 302254
rect -8576 301934 592500 302018
rect -8576 301698 -7454 301934
rect -7218 301698 12786 301934
rect 13022 301698 48786 301934
rect 49022 301698 84786 301934
rect 85022 301698 120786 301934
rect 121022 301698 156786 301934
rect 157022 301698 192786 301934
rect 193022 301698 228786 301934
rect 229022 301698 264786 301934
rect 265022 301698 300786 301934
rect 301022 301698 336786 301934
rect 337022 301698 372786 301934
rect 373022 301698 408786 301934
rect 409022 301698 444786 301934
rect 445022 301698 480786 301934
rect 481022 301698 516786 301934
rect 517022 301698 552786 301934
rect 553022 301698 591142 301934
rect 591378 301698 592500 301934
rect -8576 301676 592500 301698
rect -7636 301674 -7036 301676
rect 12604 301674 13204 301676
rect 48604 301674 49204 301676
rect 84604 301674 85204 301676
rect 120604 301674 121204 301676
rect 156604 301674 157204 301676
rect 192604 301674 193204 301676
rect 228604 301674 229204 301676
rect 264604 301674 265204 301676
rect 300604 301674 301204 301676
rect 336604 301674 337204 301676
rect 372604 301674 373204 301676
rect 408604 301674 409204 301676
rect 444604 301674 445204 301676
rect 480604 301674 481204 301676
rect 516604 301674 517204 301676
rect 552604 301674 553204 301676
rect 590960 301674 591560 301676
rect -5756 298676 -5156 298678
rect 9004 298676 9604 298678
rect 45004 298676 45604 298678
rect 81004 298676 81604 298678
rect 117004 298676 117604 298678
rect 153004 298676 153604 298678
rect 189004 298676 189604 298678
rect 225004 298676 225604 298678
rect 261004 298676 261604 298678
rect 297004 298676 297604 298678
rect 333004 298676 333604 298678
rect 369004 298676 369604 298678
rect 405004 298676 405604 298678
rect 441004 298676 441604 298678
rect 477004 298676 477604 298678
rect 513004 298676 513604 298678
rect 549004 298676 549604 298678
rect 589080 298676 589680 298678
rect -6696 298654 590620 298676
rect -6696 298418 -5574 298654
rect -5338 298418 9186 298654
rect 9422 298418 45186 298654
rect 45422 298418 81186 298654
rect 81422 298418 117186 298654
rect 117422 298418 153186 298654
rect 153422 298418 189186 298654
rect 189422 298418 225186 298654
rect 225422 298418 261186 298654
rect 261422 298418 297186 298654
rect 297422 298418 333186 298654
rect 333422 298418 369186 298654
rect 369422 298418 405186 298654
rect 405422 298418 441186 298654
rect 441422 298418 477186 298654
rect 477422 298418 513186 298654
rect 513422 298418 549186 298654
rect 549422 298418 589262 298654
rect 589498 298418 590620 298654
rect -6696 298334 590620 298418
rect -6696 298098 -5574 298334
rect -5338 298098 9186 298334
rect 9422 298098 45186 298334
rect 45422 298098 81186 298334
rect 81422 298098 117186 298334
rect 117422 298098 153186 298334
rect 153422 298098 189186 298334
rect 189422 298098 225186 298334
rect 225422 298098 261186 298334
rect 261422 298098 297186 298334
rect 297422 298098 333186 298334
rect 333422 298098 369186 298334
rect 369422 298098 405186 298334
rect 405422 298098 441186 298334
rect 441422 298098 477186 298334
rect 477422 298098 513186 298334
rect 513422 298098 549186 298334
rect 549422 298098 589262 298334
rect 589498 298098 590620 298334
rect -6696 298076 590620 298098
rect -5756 298074 -5156 298076
rect 9004 298074 9604 298076
rect 45004 298074 45604 298076
rect 81004 298074 81604 298076
rect 117004 298074 117604 298076
rect 153004 298074 153604 298076
rect 189004 298074 189604 298076
rect 225004 298074 225604 298076
rect 261004 298074 261604 298076
rect 297004 298074 297604 298076
rect 333004 298074 333604 298076
rect 369004 298074 369604 298076
rect 405004 298074 405604 298076
rect 441004 298074 441604 298076
rect 477004 298074 477604 298076
rect 513004 298074 513604 298076
rect 549004 298074 549604 298076
rect 589080 298074 589680 298076
rect -3876 295076 -3276 295078
rect 5404 295076 6004 295078
rect 41404 295076 42004 295078
rect 77404 295076 78004 295078
rect 113404 295076 114004 295078
rect 149404 295076 150004 295078
rect 185404 295076 186004 295078
rect 221404 295076 222004 295078
rect 257404 295076 258004 295078
rect 293404 295076 294004 295078
rect 329404 295076 330004 295078
rect 365404 295076 366004 295078
rect 401404 295076 402004 295078
rect 437404 295076 438004 295078
rect 473404 295076 474004 295078
rect 509404 295076 510004 295078
rect 545404 295076 546004 295078
rect 581404 295076 582004 295078
rect 587200 295076 587800 295078
rect -4816 295054 588740 295076
rect -4816 294818 -3694 295054
rect -3458 294818 5586 295054
rect 5822 294818 41586 295054
rect 41822 294818 77586 295054
rect 77822 294818 113586 295054
rect 113822 294818 149586 295054
rect 149822 294818 185586 295054
rect 185822 294818 221586 295054
rect 221822 294818 257586 295054
rect 257822 294818 293586 295054
rect 293822 294818 329586 295054
rect 329822 294818 365586 295054
rect 365822 294818 401586 295054
rect 401822 294818 437586 295054
rect 437822 294818 473586 295054
rect 473822 294818 509586 295054
rect 509822 294818 545586 295054
rect 545822 294818 581586 295054
rect 581822 294818 587382 295054
rect 587618 294818 588740 295054
rect -4816 294734 588740 294818
rect -4816 294498 -3694 294734
rect -3458 294498 5586 294734
rect 5822 294498 41586 294734
rect 41822 294498 77586 294734
rect 77822 294498 113586 294734
rect 113822 294498 149586 294734
rect 149822 294498 185586 294734
rect 185822 294498 221586 294734
rect 221822 294498 257586 294734
rect 257822 294498 293586 294734
rect 293822 294498 329586 294734
rect 329822 294498 365586 294734
rect 365822 294498 401586 294734
rect 401822 294498 437586 294734
rect 437822 294498 473586 294734
rect 473822 294498 509586 294734
rect 509822 294498 545586 294734
rect 545822 294498 581586 294734
rect 581822 294498 587382 294734
rect 587618 294498 588740 294734
rect -4816 294476 588740 294498
rect -3876 294474 -3276 294476
rect 5404 294474 6004 294476
rect 41404 294474 42004 294476
rect 77404 294474 78004 294476
rect 113404 294474 114004 294476
rect 149404 294474 150004 294476
rect 185404 294474 186004 294476
rect 221404 294474 222004 294476
rect 257404 294474 258004 294476
rect 293404 294474 294004 294476
rect 329404 294474 330004 294476
rect 365404 294474 366004 294476
rect 401404 294474 402004 294476
rect 437404 294474 438004 294476
rect 473404 294474 474004 294476
rect 509404 294474 510004 294476
rect 545404 294474 546004 294476
rect 581404 294474 582004 294476
rect 587200 294474 587800 294476
rect -1996 291476 -1396 291478
rect 1804 291476 2404 291478
rect 37804 291476 38404 291478
rect 73804 291476 74404 291478
rect 109804 291476 110404 291478
rect 145804 291476 146404 291478
rect 181804 291476 182404 291478
rect 217804 291476 218404 291478
rect 253804 291476 254404 291478
rect 289804 291476 290404 291478
rect 325804 291476 326404 291478
rect 361804 291476 362404 291478
rect 397804 291476 398404 291478
rect 433804 291476 434404 291478
rect 469804 291476 470404 291478
rect 505804 291476 506404 291478
rect 541804 291476 542404 291478
rect 577804 291476 578404 291478
rect 585320 291476 585920 291478
rect -2936 291454 586860 291476
rect -2936 291218 -1814 291454
rect -1578 291218 1986 291454
rect 2222 291218 37986 291454
rect 38222 291218 73986 291454
rect 74222 291218 109986 291454
rect 110222 291218 145986 291454
rect 146222 291218 181986 291454
rect 182222 291218 217986 291454
rect 218222 291218 253986 291454
rect 254222 291218 289986 291454
rect 290222 291218 325986 291454
rect 326222 291218 361986 291454
rect 362222 291218 397986 291454
rect 398222 291218 433986 291454
rect 434222 291218 469986 291454
rect 470222 291218 505986 291454
rect 506222 291218 541986 291454
rect 542222 291218 577986 291454
rect 578222 291218 585502 291454
rect 585738 291218 586860 291454
rect -2936 291134 586860 291218
rect -2936 290898 -1814 291134
rect -1578 290898 1986 291134
rect 2222 290898 37986 291134
rect 38222 290898 73986 291134
rect 74222 290898 109986 291134
rect 110222 290898 145986 291134
rect 146222 290898 181986 291134
rect 182222 290898 217986 291134
rect 218222 290898 253986 291134
rect 254222 290898 289986 291134
rect 290222 290898 325986 291134
rect 326222 290898 361986 291134
rect 362222 290898 397986 291134
rect 398222 290898 433986 291134
rect 434222 290898 469986 291134
rect 470222 290898 505986 291134
rect 506222 290898 541986 291134
rect 542222 290898 577986 291134
rect 578222 290898 585502 291134
rect 585738 290898 586860 291134
rect -2936 290876 586860 290898
rect -1996 290874 -1396 290876
rect 1804 290874 2404 290876
rect 37804 290874 38404 290876
rect 73804 290874 74404 290876
rect 109804 290874 110404 290876
rect 145804 290874 146404 290876
rect 181804 290874 182404 290876
rect 217804 290874 218404 290876
rect 253804 290874 254404 290876
rect 289804 290874 290404 290876
rect 325804 290874 326404 290876
rect 361804 290874 362404 290876
rect 397804 290874 398404 290876
rect 433804 290874 434404 290876
rect 469804 290874 470404 290876
rect 505804 290874 506404 290876
rect 541804 290874 542404 290876
rect 577804 290874 578404 290876
rect 585320 290874 585920 290876
rect -8576 284276 -7976 284278
rect 30604 284276 31204 284278
rect 66604 284276 67204 284278
rect 102604 284276 103204 284278
rect 138604 284276 139204 284278
rect 174604 284276 175204 284278
rect 210604 284276 211204 284278
rect 246604 284276 247204 284278
rect 282604 284276 283204 284278
rect 318604 284276 319204 284278
rect 354604 284276 355204 284278
rect 390604 284276 391204 284278
rect 426604 284276 427204 284278
rect 462604 284276 463204 284278
rect 498604 284276 499204 284278
rect 534604 284276 535204 284278
rect 570604 284276 571204 284278
rect 591900 284276 592500 284278
rect -8576 284254 592500 284276
rect -8576 284018 -8394 284254
rect -8158 284018 30786 284254
rect 31022 284018 66786 284254
rect 67022 284018 102786 284254
rect 103022 284018 138786 284254
rect 139022 284018 174786 284254
rect 175022 284018 210786 284254
rect 211022 284018 246786 284254
rect 247022 284018 282786 284254
rect 283022 284018 318786 284254
rect 319022 284018 354786 284254
rect 355022 284018 390786 284254
rect 391022 284018 426786 284254
rect 427022 284018 462786 284254
rect 463022 284018 498786 284254
rect 499022 284018 534786 284254
rect 535022 284018 570786 284254
rect 571022 284018 592082 284254
rect 592318 284018 592500 284254
rect -8576 283934 592500 284018
rect -8576 283698 -8394 283934
rect -8158 283698 30786 283934
rect 31022 283698 66786 283934
rect 67022 283698 102786 283934
rect 103022 283698 138786 283934
rect 139022 283698 174786 283934
rect 175022 283698 210786 283934
rect 211022 283698 246786 283934
rect 247022 283698 282786 283934
rect 283022 283698 318786 283934
rect 319022 283698 354786 283934
rect 355022 283698 390786 283934
rect 391022 283698 426786 283934
rect 427022 283698 462786 283934
rect 463022 283698 498786 283934
rect 499022 283698 534786 283934
rect 535022 283698 570786 283934
rect 571022 283698 592082 283934
rect 592318 283698 592500 283934
rect -8576 283676 592500 283698
rect -8576 283674 -7976 283676
rect 30604 283674 31204 283676
rect 66604 283674 67204 283676
rect 102604 283674 103204 283676
rect 138604 283674 139204 283676
rect 174604 283674 175204 283676
rect 210604 283674 211204 283676
rect 246604 283674 247204 283676
rect 282604 283674 283204 283676
rect 318604 283674 319204 283676
rect 354604 283674 355204 283676
rect 390604 283674 391204 283676
rect 426604 283674 427204 283676
rect 462604 283674 463204 283676
rect 498604 283674 499204 283676
rect 534604 283674 535204 283676
rect 570604 283674 571204 283676
rect 591900 283674 592500 283676
rect -6696 280676 -6096 280678
rect 27004 280676 27604 280678
rect 63004 280676 63604 280678
rect 99004 280676 99604 280678
rect 135004 280676 135604 280678
rect 171004 280676 171604 280678
rect 207004 280676 207604 280678
rect 243004 280676 243604 280678
rect 279004 280676 279604 280678
rect 315004 280676 315604 280678
rect 351004 280676 351604 280678
rect 387004 280676 387604 280678
rect 423004 280676 423604 280678
rect 459004 280676 459604 280678
rect 495004 280676 495604 280678
rect 531004 280676 531604 280678
rect 567004 280676 567604 280678
rect 590020 280676 590620 280678
rect -6696 280654 590620 280676
rect -6696 280418 -6514 280654
rect -6278 280418 27186 280654
rect 27422 280418 63186 280654
rect 63422 280418 99186 280654
rect 99422 280418 135186 280654
rect 135422 280418 171186 280654
rect 171422 280418 207186 280654
rect 207422 280418 243186 280654
rect 243422 280418 279186 280654
rect 279422 280418 315186 280654
rect 315422 280418 351186 280654
rect 351422 280418 387186 280654
rect 387422 280418 423186 280654
rect 423422 280418 459186 280654
rect 459422 280418 495186 280654
rect 495422 280418 531186 280654
rect 531422 280418 567186 280654
rect 567422 280418 590202 280654
rect 590438 280418 590620 280654
rect -6696 280334 590620 280418
rect -6696 280098 -6514 280334
rect -6278 280098 27186 280334
rect 27422 280098 63186 280334
rect 63422 280098 99186 280334
rect 99422 280098 135186 280334
rect 135422 280098 171186 280334
rect 171422 280098 207186 280334
rect 207422 280098 243186 280334
rect 243422 280098 279186 280334
rect 279422 280098 315186 280334
rect 315422 280098 351186 280334
rect 351422 280098 387186 280334
rect 387422 280098 423186 280334
rect 423422 280098 459186 280334
rect 459422 280098 495186 280334
rect 495422 280098 531186 280334
rect 531422 280098 567186 280334
rect 567422 280098 590202 280334
rect 590438 280098 590620 280334
rect -6696 280076 590620 280098
rect -6696 280074 -6096 280076
rect 27004 280074 27604 280076
rect 63004 280074 63604 280076
rect 99004 280074 99604 280076
rect 135004 280074 135604 280076
rect 171004 280074 171604 280076
rect 207004 280074 207604 280076
rect 243004 280074 243604 280076
rect 279004 280074 279604 280076
rect 315004 280074 315604 280076
rect 351004 280074 351604 280076
rect 387004 280074 387604 280076
rect 423004 280074 423604 280076
rect 459004 280074 459604 280076
rect 495004 280074 495604 280076
rect 531004 280074 531604 280076
rect 567004 280074 567604 280076
rect 590020 280074 590620 280076
rect -4816 277076 -4216 277078
rect 23404 277076 24004 277078
rect 59404 277076 60004 277078
rect 95404 277076 96004 277078
rect 131404 277076 132004 277078
rect 167404 277076 168004 277078
rect 203404 277076 204004 277078
rect 239404 277076 240004 277078
rect 275404 277076 276004 277078
rect 311404 277076 312004 277078
rect 347404 277076 348004 277078
rect 383404 277076 384004 277078
rect 419404 277076 420004 277078
rect 455404 277076 456004 277078
rect 491404 277076 492004 277078
rect 527404 277076 528004 277078
rect 563404 277076 564004 277078
rect 588140 277076 588740 277078
rect -4816 277054 588740 277076
rect -4816 276818 -4634 277054
rect -4398 276818 23586 277054
rect 23822 276818 59586 277054
rect 59822 276818 95586 277054
rect 95822 276818 131586 277054
rect 131822 276818 167586 277054
rect 167822 276818 203586 277054
rect 203822 276818 239586 277054
rect 239822 276818 275586 277054
rect 275822 276818 311586 277054
rect 311822 276818 347586 277054
rect 347822 276818 383586 277054
rect 383822 276818 419586 277054
rect 419822 276818 455586 277054
rect 455822 276818 491586 277054
rect 491822 276818 527586 277054
rect 527822 276818 563586 277054
rect 563822 276818 588322 277054
rect 588558 276818 588740 277054
rect -4816 276734 588740 276818
rect -4816 276498 -4634 276734
rect -4398 276498 23586 276734
rect 23822 276498 59586 276734
rect 59822 276498 95586 276734
rect 95822 276498 131586 276734
rect 131822 276498 167586 276734
rect 167822 276498 203586 276734
rect 203822 276498 239586 276734
rect 239822 276498 275586 276734
rect 275822 276498 311586 276734
rect 311822 276498 347586 276734
rect 347822 276498 383586 276734
rect 383822 276498 419586 276734
rect 419822 276498 455586 276734
rect 455822 276498 491586 276734
rect 491822 276498 527586 276734
rect 527822 276498 563586 276734
rect 563822 276498 588322 276734
rect 588558 276498 588740 276734
rect -4816 276476 588740 276498
rect -4816 276474 -4216 276476
rect 23404 276474 24004 276476
rect 59404 276474 60004 276476
rect 95404 276474 96004 276476
rect 131404 276474 132004 276476
rect 167404 276474 168004 276476
rect 203404 276474 204004 276476
rect 239404 276474 240004 276476
rect 275404 276474 276004 276476
rect 311404 276474 312004 276476
rect 347404 276474 348004 276476
rect 383404 276474 384004 276476
rect 419404 276474 420004 276476
rect 455404 276474 456004 276476
rect 491404 276474 492004 276476
rect 527404 276474 528004 276476
rect 563404 276474 564004 276476
rect 588140 276474 588740 276476
rect -2936 273476 -2336 273478
rect 19804 273476 20404 273478
rect 55804 273476 56404 273478
rect 91804 273476 92404 273478
rect 127804 273476 128404 273478
rect 163804 273476 164404 273478
rect 199804 273476 200404 273478
rect 235804 273476 236404 273478
rect 271804 273476 272404 273478
rect 307804 273476 308404 273478
rect 343804 273476 344404 273478
rect 379804 273476 380404 273478
rect 415804 273476 416404 273478
rect 451804 273476 452404 273478
rect 487804 273476 488404 273478
rect 523804 273476 524404 273478
rect 559804 273476 560404 273478
rect 586260 273476 586860 273478
rect -2936 273454 586860 273476
rect -2936 273218 -2754 273454
rect -2518 273218 19986 273454
rect 20222 273218 55986 273454
rect 56222 273218 91986 273454
rect 92222 273218 127986 273454
rect 128222 273218 163986 273454
rect 164222 273218 199986 273454
rect 200222 273218 235986 273454
rect 236222 273218 271986 273454
rect 272222 273218 307986 273454
rect 308222 273218 343986 273454
rect 344222 273218 379986 273454
rect 380222 273218 415986 273454
rect 416222 273218 451986 273454
rect 452222 273218 487986 273454
rect 488222 273218 523986 273454
rect 524222 273218 559986 273454
rect 560222 273218 586442 273454
rect 586678 273218 586860 273454
rect -2936 273134 586860 273218
rect -2936 272898 -2754 273134
rect -2518 272898 19986 273134
rect 20222 272898 55986 273134
rect 56222 272898 91986 273134
rect 92222 272898 127986 273134
rect 128222 272898 163986 273134
rect 164222 272898 199986 273134
rect 200222 272898 235986 273134
rect 236222 272898 271986 273134
rect 272222 272898 307986 273134
rect 308222 272898 343986 273134
rect 344222 272898 379986 273134
rect 380222 272898 415986 273134
rect 416222 272898 451986 273134
rect 452222 272898 487986 273134
rect 488222 272898 523986 273134
rect 524222 272898 559986 273134
rect 560222 272898 586442 273134
rect 586678 272898 586860 273134
rect -2936 272876 586860 272898
rect -2936 272874 -2336 272876
rect 19804 272874 20404 272876
rect 55804 272874 56404 272876
rect 91804 272874 92404 272876
rect 127804 272874 128404 272876
rect 163804 272874 164404 272876
rect 199804 272874 200404 272876
rect 235804 272874 236404 272876
rect 271804 272874 272404 272876
rect 307804 272874 308404 272876
rect 343804 272874 344404 272876
rect 379804 272874 380404 272876
rect 415804 272874 416404 272876
rect 451804 272874 452404 272876
rect 487804 272874 488404 272876
rect 523804 272874 524404 272876
rect 559804 272874 560404 272876
rect 586260 272874 586860 272876
rect -7636 266276 -7036 266278
rect 12604 266276 13204 266278
rect 48604 266276 49204 266278
rect 84604 266276 85204 266278
rect 120604 266276 121204 266278
rect 156604 266276 157204 266278
rect 192604 266276 193204 266278
rect 228604 266276 229204 266278
rect 264604 266276 265204 266278
rect 300604 266276 301204 266278
rect 336604 266276 337204 266278
rect 372604 266276 373204 266278
rect 408604 266276 409204 266278
rect 444604 266276 445204 266278
rect 480604 266276 481204 266278
rect 516604 266276 517204 266278
rect 552604 266276 553204 266278
rect 590960 266276 591560 266278
rect -8576 266254 592500 266276
rect -8576 266018 -7454 266254
rect -7218 266018 12786 266254
rect 13022 266018 48786 266254
rect 49022 266018 84786 266254
rect 85022 266018 120786 266254
rect 121022 266018 156786 266254
rect 157022 266018 192786 266254
rect 193022 266018 228786 266254
rect 229022 266018 264786 266254
rect 265022 266018 300786 266254
rect 301022 266018 336786 266254
rect 337022 266018 372786 266254
rect 373022 266018 408786 266254
rect 409022 266018 444786 266254
rect 445022 266018 480786 266254
rect 481022 266018 516786 266254
rect 517022 266018 552786 266254
rect 553022 266018 591142 266254
rect 591378 266018 592500 266254
rect -8576 265934 592500 266018
rect -8576 265698 -7454 265934
rect -7218 265698 12786 265934
rect 13022 265698 48786 265934
rect 49022 265698 84786 265934
rect 85022 265698 120786 265934
rect 121022 265698 156786 265934
rect 157022 265698 192786 265934
rect 193022 265698 228786 265934
rect 229022 265698 264786 265934
rect 265022 265698 300786 265934
rect 301022 265698 336786 265934
rect 337022 265698 372786 265934
rect 373022 265698 408786 265934
rect 409022 265698 444786 265934
rect 445022 265698 480786 265934
rect 481022 265698 516786 265934
rect 517022 265698 552786 265934
rect 553022 265698 591142 265934
rect 591378 265698 592500 265934
rect -8576 265676 592500 265698
rect -7636 265674 -7036 265676
rect 12604 265674 13204 265676
rect 48604 265674 49204 265676
rect 84604 265674 85204 265676
rect 120604 265674 121204 265676
rect 156604 265674 157204 265676
rect 192604 265674 193204 265676
rect 228604 265674 229204 265676
rect 264604 265674 265204 265676
rect 300604 265674 301204 265676
rect 336604 265674 337204 265676
rect 372604 265674 373204 265676
rect 408604 265674 409204 265676
rect 444604 265674 445204 265676
rect 480604 265674 481204 265676
rect 516604 265674 517204 265676
rect 552604 265674 553204 265676
rect 590960 265674 591560 265676
rect -5756 262676 -5156 262678
rect 9004 262676 9604 262678
rect 45004 262676 45604 262678
rect 81004 262676 81604 262678
rect 117004 262676 117604 262678
rect 153004 262676 153604 262678
rect 189004 262676 189604 262678
rect 225004 262676 225604 262678
rect 261004 262676 261604 262678
rect 297004 262676 297604 262678
rect 333004 262676 333604 262678
rect 369004 262676 369604 262678
rect 405004 262676 405604 262678
rect 441004 262676 441604 262678
rect 477004 262676 477604 262678
rect 513004 262676 513604 262678
rect 549004 262676 549604 262678
rect 589080 262676 589680 262678
rect -6696 262654 590620 262676
rect -6696 262418 -5574 262654
rect -5338 262418 9186 262654
rect 9422 262418 45186 262654
rect 45422 262418 81186 262654
rect 81422 262418 117186 262654
rect 117422 262418 153186 262654
rect 153422 262418 189186 262654
rect 189422 262418 225186 262654
rect 225422 262418 261186 262654
rect 261422 262418 297186 262654
rect 297422 262418 333186 262654
rect 333422 262418 369186 262654
rect 369422 262418 405186 262654
rect 405422 262418 441186 262654
rect 441422 262418 477186 262654
rect 477422 262418 513186 262654
rect 513422 262418 549186 262654
rect 549422 262418 589262 262654
rect 589498 262418 590620 262654
rect -6696 262334 590620 262418
rect -6696 262098 -5574 262334
rect -5338 262098 9186 262334
rect 9422 262098 45186 262334
rect 45422 262098 81186 262334
rect 81422 262098 117186 262334
rect 117422 262098 153186 262334
rect 153422 262098 189186 262334
rect 189422 262098 225186 262334
rect 225422 262098 261186 262334
rect 261422 262098 297186 262334
rect 297422 262098 333186 262334
rect 333422 262098 369186 262334
rect 369422 262098 405186 262334
rect 405422 262098 441186 262334
rect 441422 262098 477186 262334
rect 477422 262098 513186 262334
rect 513422 262098 549186 262334
rect 549422 262098 589262 262334
rect 589498 262098 590620 262334
rect -6696 262076 590620 262098
rect -5756 262074 -5156 262076
rect 9004 262074 9604 262076
rect 45004 262074 45604 262076
rect 81004 262074 81604 262076
rect 117004 262074 117604 262076
rect 153004 262074 153604 262076
rect 189004 262074 189604 262076
rect 225004 262074 225604 262076
rect 261004 262074 261604 262076
rect 297004 262074 297604 262076
rect 333004 262074 333604 262076
rect 369004 262074 369604 262076
rect 405004 262074 405604 262076
rect 441004 262074 441604 262076
rect 477004 262074 477604 262076
rect 513004 262074 513604 262076
rect 549004 262074 549604 262076
rect 589080 262074 589680 262076
rect -3876 259076 -3276 259078
rect 5404 259076 6004 259078
rect 41404 259076 42004 259078
rect 77404 259076 78004 259078
rect 113404 259076 114004 259078
rect 149404 259076 150004 259078
rect 185404 259076 186004 259078
rect 221404 259076 222004 259078
rect 257404 259076 258004 259078
rect 293404 259076 294004 259078
rect 329404 259076 330004 259078
rect 365404 259076 366004 259078
rect 401404 259076 402004 259078
rect 437404 259076 438004 259078
rect 473404 259076 474004 259078
rect 509404 259076 510004 259078
rect 545404 259076 546004 259078
rect 581404 259076 582004 259078
rect 587200 259076 587800 259078
rect -4816 259054 588740 259076
rect -4816 258818 -3694 259054
rect -3458 258818 5586 259054
rect 5822 258818 41586 259054
rect 41822 258818 77586 259054
rect 77822 258818 113586 259054
rect 113822 258818 149586 259054
rect 149822 258818 185586 259054
rect 185822 258818 221586 259054
rect 221822 258818 257586 259054
rect 257822 258818 293586 259054
rect 293822 258818 329586 259054
rect 329822 258818 365586 259054
rect 365822 258818 401586 259054
rect 401822 258818 437586 259054
rect 437822 258818 473586 259054
rect 473822 258818 509586 259054
rect 509822 258818 545586 259054
rect 545822 258818 581586 259054
rect 581822 258818 587382 259054
rect 587618 258818 588740 259054
rect -4816 258734 588740 258818
rect -4816 258498 -3694 258734
rect -3458 258498 5586 258734
rect 5822 258498 41586 258734
rect 41822 258498 77586 258734
rect 77822 258498 113586 258734
rect 113822 258498 149586 258734
rect 149822 258498 185586 258734
rect 185822 258498 221586 258734
rect 221822 258498 257586 258734
rect 257822 258498 293586 258734
rect 293822 258498 329586 258734
rect 329822 258498 365586 258734
rect 365822 258498 401586 258734
rect 401822 258498 437586 258734
rect 437822 258498 473586 258734
rect 473822 258498 509586 258734
rect 509822 258498 545586 258734
rect 545822 258498 581586 258734
rect 581822 258498 587382 258734
rect 587618 258498 588740 258734
rect -4816 258476 588740 258498
rect -3876 258474 -3276 258476
rect 5404 258474 6004 258476
rect 41404 258474 42004 258476
rect 77404 258474 78004 258476
rect 113404 258474 114004 258476
rect 149404 258474 150004 258476
rect 185404 258474 186004 258476
rect 221404 258474 222004 258476
rect 257404 258474 258004 258476
rect 293404 258474 294004 258476
rect 329404 258474 330004 258476
rect 365404 258474 366004 258476
rect 401404 258474 402004 258476
rect 437404 258474 438004 258476
rect 473404 258474 474004 258476
rect 509404 258474 510004 258476
rect 545404 258474 546004 258476
rect 581404 258474 582004 258476
rect 587200 258474 587800 258476
rect -1996 255476 -1396 255478
rect 1804 255476 2404 255478
rect 37804 255476 38404 255478
rect 73804 255476 74404 255478
rect 109804 255476 110404 255478
rect 145804 255476 146404 255478
rect 181804 255476 182404 255478
rect 217804 255476 218404 255478
rect 253804 255476 254404 255478
rect 289804 255476 290404 255478
rect 325804 255476 326404 255478
rect 361804 255476 362404 255478
rect 397804 255476 398404 255478
rect 433804 255476 434404 255478
rect 469804 255476 470404 255478
rect 505804 255476 506404 255478
rect 541804 255476 542404 255478
rect 577804 255476 578404 255478
rect 585320 255476 585920 255478
rect -2936 255454 586860 255476
rect -2936 255218 -1814 255454
rect -1578 255218 1986 255454
rect 2222 255218 37986 255454
rect 38222 255218 73986 255454
rect 74222 255218 109986 255454
rect 110222 255218 145986 255454
rect 146222 255218 181986 255454
rect 182222 255218 217986 255454
rect 218222 255218 253986 255454
rect 254222 255218 289986 255454
rect 290222 255218 325986 255454
rect 326222 255218 361986 255454
rect 362222 255218 397986 255454
rect 398222 255218 433986 255454
rect 434222 255218 469986 255454
rect 470222 255218 505986 255454
rect 506222 255218 541986 255454
rect 542222 255218 577986 255454
rect 578222 255218 585502 255454
rect 585738 255218 586860 255454
rect -2936 255134 586860 255218
rect -2936 254898 -1814 255134
rect -1578 254898 1986 255134
rect 2222 254898 37986 255134
rect 38222 254898 73986 255134
rect 74222 254898 109986 255134
rect 110222 254898 145986 255134
rect 146222 254898 181986 255134
rect 182222 254898 217986 255134
rect 218222 254898 253986 255134
rect 254222 254898 289986 255134
rect 290222 254898 325986 255134
rect 326222 254898 361986 255134
rect 362222 254898 397986 255134
rect 398222 254898 433986 255134
rect 434222 254898 469986 255134
rect 470222 254898 505986 255134
rect 506222 254898 541986 255134
rect 542222 254898 577986 255134
rect 578222 254898 585502 255134
rect 585738 254898 586860 255134
rect -2936 254876 586860 254898
rect -1996 254874 -1396 254876
rect 1804 254874 2404 254876
rect 37804 254874 38404 254876
rect 73804 254874 74404 254876
rect 109804 254874 110404 254876
rect 145804 254874 146404 254876
rect 181804 254874 182404 254876
rect 217804 254874 218404 254876
rect 253804 254874 254404 254876
rect 289804 254874 290404 254876
rect 325804 254874 326404 254876
rect 361804 254874 362404 254876
rect 397804 254874 398404 254876
rect 433804 254874 434404 254876
rect 469804 254874 470404 254876
rect 505804 254874 506404 254876
rect 541804 254874 542404 254876
rect 577804 254874 578404 254876
rect 585320 254874 585920 254876
rect -8576 248276 -7976 248278
rect 30604 248276 31204 248278
rect 66604 248276 67204 248278
rect 102604 248276 103204 248278
rect 138604 248276 139204 248278
rect 174604 248276 175204 248278
rect 210604 248276 211204 248278
rect 246604 248276 247204 248278
rect 282604 248276 283204 248278
rect 318604 248276 319204 248278
rect 354604 248276 355204 248278
rect 390604 248276 391204 248278
rect 426604 248276 427204 248278
rect 462604 248276 463204 248278
rect 498604 248276 499204 248278
rect 534604 248276 535204 248278
rect 570604 248276 571204 248278
rect 591900 248276 592500 248278
rect -8576 248254 592500 248276
rect -8576 248018 -8394 248254
rect -8158 248018 30786 248254
rect 31022 248018 66786 248254
rect 67022 248018 102786 248254
rect 103022 248018 138786 248254
rect 139022 248018 174786 248254
rect 175022 248018 210786 248254
rect 211022 248018 246786 248254
rect 247022 248018 282786 248254
rect 283022 248018 318786 248254
rect 319022 248018 354786 248254
rect 355022 248018 390786 248254
rect 391022 248018 426786 248254
rect 427022 248018 462786 248254
rect 463022 248018 498786 248254
rect 499022 248018 534786 248254
rect 535022 248018 570786 248254
rect 571022 248018 592082 248254
rect 592318 248018 592500 248254
rect -8576 247934 592500 248018
rect -8576 247698 -8394 247934
rect -8158 247698 30786 247934
rect 31022 247698 66786 247934
rect 67022 247698 102786 247934
rect 103022 247698 138786 247934
rect 139022 247698 174786 247934
rect 175022 247698 210786 247934
rect 211022 247698 246786 247934
rect 247022 247698 282786 247934
rect 283022 247698 318786 247934
rect 319022 247698 354786 247934
rect 355022 247698 390786 247934
rect 391022 247698 426786 247934
rect 427022 247698 462786 247934
rect 463022 247698 498786 247934
rect 499022 247698 534786 247934
rect 535022 247698 570786 247934
rect 571022 247698 592082 247934
rect 592318 247698 592500 247934
rect -8576 247676 592500 247698
rect -8576 247674 -7976 247676
rect 30604 247674 31204 247676
rect 66604 247674 67204 247676
rect 102604 247674 103204 247676
rect 138604 247674 139204 247676
rect 174604 247674 175204 247676
rect 210604 247674 211204 247676
rect 246604 247674 247204 247676
rect 282604 247674 283204 247676
rect 318604 247674 319204 247676
rect 354604 247674 355204 247676
rect 390604 247674 391204 247676
rect 426604 247674 427204 247676
rect 462604 247674 463204 247676
rect 498604 247674 499204 247676
rect 534604 247674 535204 247676
rect 570604 247674 571204 247676
rect 591900 247674 592500 247676
rect -6696 244676 -6096 244678
rect 27004 244676 27604 244678
rect 63004 244676 63604 244678
rect 99004 244676 99604 244678
rect 135004 244676 135604 244678
rect 171004 244676 171604 244678
rect 207004 244676 207604 244678
rect 243004 244676 243604 244678
rect 279004 244676 279604 244678
rect 315004 244676 315604 244678
rect 351004 244676 351604 244678
rect 387004 244676 387604 244678
rect 423004 244676 423604 244678
rect 459004 244676 459604 244678
rect 495004 244676 495604 244678
rect 531004 244676 531604 244678
rect 567004 244676 567604 244678
rect 590020 244676 590620 244678
rect -6696 244654 590620 244676
rect -6696 244418 -6514 244654
rect -6278 244418 27186 244654
rect 27422 244418 63186 244654
rect 63422 244418 99186 244654
rect 99422 244418 135186 244654
rect 135422 244418 171186 244654
rect 171422 244418 207186 244654
rect 207422 244418 243186 244654
rect 243422 244418 279186 244654
rect 279422 244418 315186 244654
rect 315422 244418 351186 244654
rect 351422 244418 387186 244654
rect 387422 244418 423186 244654
rect 423422 244418 459186 244654
rect 459422 244418 495186 244654
rect 495422 244418 531186 244654
rect 531422 244418 567186 244654
rect 567422 244418 590202 244654
rect 590438 244418 590620 244654
rect -6696 244334 590620 244418
rect -6696 244098 -6514 244334
rect -6278 244098 27186 244334
rect 27422 244098 63186 244334
rect 63422 244098 99186 244334
rect 99422 244098 135186 244334
rect 135422 244098 171186 244334
rect 171422 244098 207186 244334
rect 207422 244098 243186 244334
rect 243422 244098 279186 244334
rect 279422 244098 315186 244334
rect 315422 244098 351186 244334
rect 351422 244098 387186 244334
rect 387422 244098 423186 244334
rect 423422 244098 459186 244334
rect 459422 244098 495186 244334
rect 495422 244098 531186 244334
rect 531422 244098 567186 244334
rect 567422 244098 590202 244334
rect 590438 244098 590620 244334
rect -6696 244076 590620 244098
rect -6696 244074 -6096 244076
rect 27004 244074 27604 244076
rect 63004 244074 63604 244076
rect 99004 244074 99604 244076
rect 135004 244074 135604 244076
rect 171004 244074 171604 244076
rect 207004 244074 207604 244076
rect 243004 244074 243604 244076
rect 279004 244074 279604 244076
rect 315004 244074 315604 244076
rect 351004 244074 351604 244076
rect 387004 244074 387604 244076
rect 423004 244074 423604 244076
rect 459004 244074 459604 244076
rect 495004 244074 495604 244076
rect 531004 244074 531604 244076
rect 567004 244074 567604 244076
rect 590020 244074 590620 244076
rect -4816 241076 -4216 241078
rect 23404 241076 24004 241078
rect 59404 241076 60004 241078
rect 95404 241076 96004 241078
rect 131404 241076 132004 241078
rect 167404 241076 168004 241078
rect 203404 241076 204004 241078
rect 239404 241076 240004 241078
rect 275404 241076 276004 241078
rect 311404 241076 312004 241078
rect 347404 241076 348004 241078
rect 383404 241076 384004 241078
rect 419404 241076 420004 241078
rect 455404 241076 456004 241078
rect 491404 241076 492004 241078
rect 527404 241076 528004 241078
rect 563404 241076 564004 241078
rect 588140 241076 588740 241078
rect -4816 241054 588740 241076
rect -4816 240818 -4634 241054
rect -4398 240818 23586 241054
rect 23822 240818 59586 241054
rect 59822 240818 95586 241054
rect 95822 240818 131586 241054
rect 131822 240818 167586 241054
rect 167822 240818 203586 241054
rect 203822 240818 239586 241054
rect 239822 240818 275586 241054
rect 275822 240818 311586 241054
rect 311822 240818 347586 241054
rect 347822 240818 383586 241054
rect 383822 240818 419586 241054
rect 419822 240818 455586 241054
rect 455822 240818 491586 241054
rect 491822 240818 527586 241054
rect 527822 240818 563586 241054
rect 563822 240818 588322 241054
rect 588558 240818 588740 241054
rect -4816 240734 588740 240818
rect -4816 240498 -4634 240734
rect -4398 240498 23586 240734
rect 23822 240498 59586 240734
rect 59822 240498 95586 240734
rect 95822 240498 131586 240734
rect 131822 240498 167586 240734
rect 167822 240498 203586 240734
rect 203822 240498 239586 240734
rect 239822 240498 275586 240734
rect 275822 240498 311586 240734
rect 311822 240498 347586 240734
rect 347822 240498 383586 240734
rect 383822 240498 419586 240734
rect 419822 240498 455586 240734
rect 455822 240498 491586 240734
rect 491822 240498 527586 240734
rect 527822 240498 563586 240734
rect 563822 240498 588322 240734
rect 588558 240498 588740 240734
rect -4816 240476 588740 240498
rect -4816 240474 -4216 240476
rect 23404 240474 24004 240476
rect 59404 240474 60004 240476
rect 95404 240474 96004 240476
rect 131404 240474 132004 240476
rect 167404 240474 168004 240476
rect 203404 240474 204004 240476
rect 239404 240474 240004 240476
rect 275404 240474 276004 240476
rect 311404 240474 312004 240476
rect 347404 240474 348004 240476
rect 383404 240474 384004 240476
rect 419404 240474 420004 240476
rect 455404 240474 456004 240476
rect 491404 240474 492004 240476
rect 527404 240474 528004 240476
rect 563404 240474 564004 240476
rect 588140 240474 588740 240476
rect -2936 237476 -2336 237478
rect 19804 237476 20404 237478
rect 55804 237476 56404 237478
rect 91804 237476 92404 237478
rect 127804 237476 128404 237478
rect 163804 237476 164404 237478
rect 199804 237476 200404 237478
rect 235804 237476 236404 237478
rect 271804 237476 272404 237478
rect 307804 237476 308404 237478
rect 343804 237476 344404 237478
rect 379804 237476 380404 237478
rect 415804 237476 416404 237478
rect 451804 237476 452404 237478
rect 487804 237476 488404 237478
rect 523804 237476 524404 237478
rect 559804 237476 560404 237478
rect 586260 237476 586860 237478
rect -2936 237454 586860 237476
rect -2936 237218 -2754 237454
rect -2518 237218 19986 237454
rect 20222 237218 55986 237454
rect 56222 237218 91986 237454
rect 92222 237218 127986 237454
rect 128222 237218 163986 237454
rect 164222 237218 199986 237454
rect 200222 237218 235986 237454
rect 236222 237218 271986 237454
rect 272222 237218 307986 237454
rect 308222 237218 343986 237454
rect 344222 237218 379986 237454
rect 380222 237218 415986 237454
rect 416222 237218 451986 237454
rect 452222 237218 487986 237454
rect 488222 237218 523986 237454
rect 524222 237218 559986 237454
rect 560222 237218 586442 237454
rect 586678 237218 586860 237454
rect -2936 237134 586860 237218
rect -2936 236898 -2754 237134
rect -2518 236898 19986 237134
rect 20222 236898 55986 237134
rect 56222 236898 91986 237134
rect 92222 236898 127986 237134
rect 128222 236898 163986 237134
rect 164222 236898 199986 237134
rect 200222 236898 235986 237134
rect 236222 236898 271986 237134
rect 272222 236898 307986 237134
rect 308222 236898 343986 237134
rect 344222 236898 379986 237134
rect 380222 236898 415986 237134
rect 416222 236898 451986 237134
rect 452222 236898 487986 237134
rect 488222 236898 523986 237134
rect 524222 236898 559986 237134
rect 560222 236898 586442 237134
rect 586678 236898 586860 237134
rect -2936 236876 586860 236898
rect -2936 236874 -2336 236876
rect 19804 236874 20404 236876
rect 55804 236874 56404 236876
rect 91804 236874 92404 236876
rect 127804 236874 128404 236876
rect 163804 236874 164404 236876
rect 199804 236874 200404 236876
rect 235804 236874 236404 236876
rect 271804 236874 272404 236876
rect 307804 236874 308404 236876
rect 343804 236874 344404 236876
rect 379804 236874 380404 236876
rect 415804 236874 416404 236876
rect 451804 236874 452404 236876
rect 487804 236874 488404 236876
rect 523804 236874 524404 236876
rect 559804 236874 560404 236876
rect 586260 236874 586860 236876
rect -7636 230276 -7036 230278
rect 12604 230276 13204 230278
rect 48604 230276 49204 230278
rect 84604 230276 85204 230278
rect 120604 230276 121204 230278
rect 156604 230276 157204 230278
rect 192604 230276 193204 230278
rect 228604 230276 229204 230278
rect 264604 230276 265204 230278
rect 300604 230276 301204 230278
rect 336604 230276 337204 230278
rect 372604 230276 373204 230278
rect 408604 230276 409204 230278
rect 444604 230276 445204 230278
rect 480604 230276 481204 230278
rect 516604 230276 517204 230278
rect 552604 230276 553204 230278
rect 590960 230276 591560 230278
rect -8576 230254 592500 230276
rect -8576 230018 -7454 230254
rect -7218 230018 12786 230254
rect 13022 230018 48786 230254
rect 49022 230018 84786 230254
rect 85022 230018 120786 230254
rect 121022 230018 156786 230254
rect 157022 230018 192786 230254
rect 193022 230018 228786 230254
rect 229022 230018 264786 230254
rect 265022 230018 300786 230254
rect 301022 230018 336786 230254
rect 337022 230018 372786 230254
rect 373022 230018 408786 230254
rect 409022 230018 444786 230254
rect 445022 230018 480786 230254
rect 481022 230018 516786 230254
rect 517022 230018 552786 230254
rect 553022 230018 591142 230254
rect 591378 230018 592500 230254
rect -8576 229934 592500 230018
rect -8576 229698 -7454 229934
rect -7218 229698 12786 229934
rect 13022 229698 48786 229934
rect 49022 229698 84786 229934
rect 85022 229698 120786 229934
rect 121022 229698 156786 229934
rect 157022 229698 192786 229934
rect 193022 229698 228786 229934
rect 229022 229698 264786 229934
rect 265022 229698 300786 229934
rect 301022 229698 336786 229934
rect 337022 229698 372786 229934
rect 373022 229698 408786 229934
rect 409022 229698 444786 229934
rect 445022 229698 480786 229934
rect 481022 229698 516786 229934
rect 517022 229698 552786 229934
rect 553022 229698 591142 229934
rect 591378 229698 592500 229934
rect -8576 229676 592500 229698
rect -7636 229674 -7036 229676
rect 12604 229674 13204 229676
rect 48604 229674 49204 229676
rect 84604 229674 85204 229676
rect 120604 229674 121204 229676
rect 156604 229674 157204 229676
rect 192604 229674 193204 229676
rect 228604 229674 229204 229676
rect 264604 229674 265204 229676
rect 300604 229674 301204 229676
rect 336604 229674 337204 229676
rect 372604 229674 373204 229676
rect 408604 229674 409204 229676
rect 444604 229674 445204 229676
rect 480604 229674 481204 229676
rect 516604 229674 517204 229676
rect 552604 229674 553204 229676
rect 590960 229674 591560 229676
rect -5756 226676 -5156 226678
rect 9004 226676 9604 226678
rect 45004 226676 45604 226678
rect 81004 226676 81604 226678
rect 117004 226676 117604 226678
rect 153004 226676 153604 226678
rect 189004 226676 189604 226678
rect 225004 226676 225604 226678
rect 261004 226676 261604 226678
rect 297004 226676 297604 226678
rect 333004 226676 333604 226678
rect 369004 226676 369604 226678
rect 405004 226676 405604 226678
rect 441004 226676 441604 226678
rect 477004 226676 477604 226678
rect 513004 226676 513604 226678
rect 549004 226676 549604 226678
rect 589080 226676 589680 226678
rect -6696 226654 590620 226676
rect -6696 226418 -5574 226654
rect -5338 226418 9186 226654
rect 9422 226418 45186 226654
rect 45422 226418 81186 226654
rect 81422 226418 117186 226654
rect 117422 226418 153186 226654
rect 153422 226418 189186 226654
rect 189422 226418 225186 226654
rect 225422 226418 261186 226654
rect 261422 226418 297186 226654
rect 297422 226418 333186 226654
rect 333422 226418 369186 226654
rect 369422 226418 405186 226654
rect 405422 226418 441186 226654
rect 441422 226418 477186 226654
rect 477422 226418 513186 226654
rect 513422 226418 549186 226654
rect 549422 226418 589262 226654
rect 589498 226418 590620 226654
rect -6696 226334 590620 226418
rect -6696 226098 -5574 226334
rect -5338 226098 9186 226334
rect 9422 226098 45186 226334
rect 45422 226098 81186 226334
rect 81422 226098 117186 226334
rect 117422 226098 153186 226334
rect 153422 226098 189186 226334
rect 189422 226098 225186 226334
rect 225422 226098 261186 226334
rect 261422 226098 297186 226334
rect 297422 226098 333186 226334
rect 333422 226098 369186 226334
rect 369422 226098 405186 226334
rect 405422 226098 441186 226334
rect 441422 226098 477186 226334
rect 477422 226098 513186 226334
rect 513422 226098 549186 226334
rect 549422 226098 589262 226334
rect 589498 226098 590620 226334
rect -6696 226076 590620 226098
rect -5756 226074 -5156 226076
rect 9004 226074 9604 226076
rect 45004 226074 45604 226076
rect 81004 226074 81604 226076
rect 117004 226074 117604 226076
rect 153004 226074 153604 226076
rect 189004 226074 189604 226076
rect 225004 226074 225604 226076
rect 261004 226074 261604 226076
rect 297004 226074 297604 226076
rect 333004 226074 333604 226076
rect 369004 226074 369604 226076
rect 405004 226074 405604 226076
rect 441004 226074 441604 226076
rect 477004 226074 477604 226076
rect 513004 226074 513604 226076
rect 549004 226074 549604 226076
rect 589080 226074 589680 226076
rect -3876 223076 -3276 223078
rect 5404 223076 6004 223078
rect 41404 223076 42004 223078
rect 77404 223076 78004 223078
rect 113404 223076 114004 223078
rect 149404 223076 150004 223078
rect 185404 223076 186004 223078
rect 221404 223076 222004 223078
rect 257404 223076 258004 223078
rect 293404 223076 294004 223078
rect 329404 223076 330004 223078
rect 365404 223076 366004 223078
rect 401404 223076 402004 223078
rect 437404 223076 438004 223078
rect 473404 223076 474004 223078
rect 509404 223076 510004 223078
rect 545404 223076 546004 223078
rect 581404 223076 582004 223078
rect 587200 223076 587800 223078
rect -4816 223054 588740 223076
rect -4816 222818 -3694 223054
rect -3458 222818 5586 223054
rect 5822 222818 41586 223054
rect 41822 222818 77586 223054
rect 77822 222818 113586 223054
rect 113822 222818 149586 223054
rect 149822 222818 185586 223054
rect 185822 222818 221586 223054
rect 221822 222818 257586 223054
rect 257822 222818 293586 223054
rect 293822 222818 329586 223054
rect 329822 222818 365586 223054
rect 365822 222818 401586 223054
rect 401822 222818 437586 223054
rect 437822 222818 473586 223054
rect 473822 222818 509586 223054
rect 509822 222818 545586 223054
rect 545822 222818 581586 223054
rect 581822 222818 587382 223054
rect 587618 222818 588740 223054
rect -4816 222734 588740 222818
rect -4816 222498 -3694 222734
rect -3458 222498 5586 222734
rect 5822 222498 41586 222734
rect 41822 222498 77586 222734
rect 77822 222498 113586 222734
rect 113822 222498 149586 222734
rect 149822 222498 185586 222734
rect 185822 222498 221586 222734
rect 221822 222498 257586 222734
rect 257822 222498 293586 222734
rect 293822 222498 329586 222734
rect 329822 222498 365586 222734
rect 365822 222498 401586 222734
rect 401822 222498 437586 222734
rect 437822 222498 473586 222734
rect 473822 222498 509586 222734
rect 509822 222498 545586 222734
rect 545822 222498 581586 222734
rect 581822 222498 587382 222734
rect 587618 222498 588740 222734
rect -4816 222476 588740 222498
rect -3876 222474 -3276 222476
rect 5404 222474 6004 222476
rect 41404 222474 42004 222476
rect 77404 222474 78004 222476
rect 113404 222474 114004 222476
rect 149404 222474 150004 222476
rect 185404 222474 186004 222476
rect 221404 222474 222004 222476
rect 257404 222474 258004 222476
rect 293404 222474 294004 222476
rect 329404 222474 330004 222476
rect 365404 222474 366004 222476
rect 401404 222474 402004 222476
rect 437404 222474 438004 222476
rect 473404 222474 474004 222476
rect 509404 222474 510004 222476
rect 545404 222474 546004 222476
rect 581404 222474 582004 222476
rect 587200 222474 587800 222476
rect -1996 219476 -1396 219478
rect 1804 219476 2404 219478
rect 37804 219476 38404 219478
rect 73804 219476 74404 219478
rect 109804 219476 110404 219478
rect 145804 219476 146404 219478
rect 181804 219476 182404 219478
rect 217804 219476 218404 219478
rect 253804 219476 254404 219478
rect 289804 219476 290404 219478
rect 325804 219476 326404 219478
rect 361804 219476 362404 219478
rect 397804 219476 398404 219478
rect 433804 219476 434404 219478
rect 469804 219476 470404 219478
rect 505804 219476 506404 219478
rect 541804 219476 542404 219478
rect 577804 219476 578404 219478
rect 585320 219476 585920 219478
rect -2936 219454 586860 219476
rect -2936 219218 -1814 219454
rect -1578 219218 1986 219454
rect 2222 219218 37986 219454
rect 38222 219218 73986 219454
rect 74222 219218 109986 219454
rect 110222 219218 145986 219454
rect 146222 219218 181986 219454
rect 182222 219218 217986 219454
rect 218222 219218 253986 219454
rect 254222 219218 289986 219454
rect 290222 219218 325986 219454
rect 326222 219218 361986 219454
rect 362222 219218 397986 219454
rect 398222 219218 433986 219454
rect 434222 219218 469986 219454
rect 470222 219218 505986 219454
rect 506222 219218 541986 219454
rect 542222 219218 577986 219454
rect 578222 219218 585502 219454
rect 585738 219218 586860 219454
rect -2936 219134 586860 219218
rect -2936 218898 -1814 219134
rect -1578 218898 1986 219134
rect 2222 218898 37986 219134
rect 38222 218898 73986 219134
rect 74222 218898 109986 219134
rect 110222 218898 145986 219134
rect 146222 218898 181986 219134
rect 182222 218898 217986 219134
rect 218222 218898 253986 219134
rect 254222 218898 289986 219134
rect 290222 218898 325986 219134
rect 326222 218898 361986 219134
rect 362222 218898 397986 219134
rect 398222 218898 433986 219134
rect 434222 218898 469986 219134
rect 470222 218898 505986 219134
rect 506222 218898 541986 219134
rect 542222 218898 577986 219134
rect 578222 218898 585502 219134
rect 585738 218898 586860 219134
rect -2936 218876 586860 218898
rect -1996 218874 -1396 218876
rect 1804 218874 2404 218876
rect 37804 218874 38404 218876
rect 73804 218874 74404 218876
rect 109804 218874 110404 218876
rect 145804 218874 146404 218876
rect 181804 218874 182404 218876
rect 217804 218874 218404 218876
rect 253804 218874 254404 218876
rect 289804 218874 290404 218876
rect 325804 218874 326404 218876
rect 361804 218874 362404 218876
rect 397804 218874 398404 218876
rect 433804 218874 434404 218876
rect 469804 218874 470404 218876
rect 505804 218874 506404 218876
rect 541804 218874 542404 218876
rect 577804 218874 578404 218876
rect 585320 218874 585920 218876
rect -8576 212276 -7976 212278
rect 30604 212276 31204 212278
rect 66604 212276 67204 212278
rect 102604 212276 103204 212278
rect 138604 212276 139204 212278
rect 174604 212276 175204 212278
rect 210604 212276 211204 212278
rect 246604 212276 247204 212278
rect 282604 212276 283204 212278
rect 318604 212276 319204 212278
rect 354604 212276 355204 212278
rect 390604 212276 391204 212278
rect 426604 212276 427204 212278
rect 462604 212276 463204 212278
rect 498604 212276 499204 212278
rect 534604 212276 535204 212278
rect 570604 212276 571204 212278
rect 591900 212276 592500 212278
rect -8576 212254 592500 212276
rect -8576 212018 -8394 212254
rect -8158 212018 30786 212254
rect 31022 212018 66786 212254
rect 67022 212018 102786 212254
rect 103022 212018 138786 212254
rect 139022 212018 174786 212254
rect 175022 212018 210786 212254
rect 211022 212018 246786 212254
rect 247022 212018 282786 212254
rect 283022 212018 318786 212254
rect 319022 212018 354786 212254
rect 355022 212018 390786 212254
rect 391022 212018 426786 212254
rect 427022 212018 462786 212254
rect 463022 212018 498786 212254
rect 499022 212018 534786 212254
rect 535022 212018 570786 212254
rect 571022 212018 592082 212254
rect 592318 212018 592500 212254
rect -8576 211934 592500 212018
rect -8576 211698 -8394 211934
rect -8158 211698 30786 211934
rect 31022 211698 66786 211934
rect 67022 211698 102786 211934
rect 103022 211698 138786 211934
rect 139022 211698 174786 211934
rect 175022 211698 210786 211934
rect 211022 211698 246786 211934
rect 247022 211698 282786 211934
rect 283022 211698 318786 211934
rect 319022 211698 354786 211934
rect 355022 211698 390786 211934
rect 391022 211698 426786 211934
rect 427022 211698 462786 211934
rect 463022 211698 498786 211934
rect 499022 211698 534786 211934
rect 535022 211698 570786 211934
rect 571022 211698 592082 211934
rect 592318 211698 592500 211934
rect -8576 211676 592500 211698
rect -8576 211674 -7976 211676
rect 30604 211674 31204 211676
rect 66604 211674 67204 211676
rect 102604 211674 103204 211676
rect 138604 211674 139204 211676
rect 174604 211674 175204 211676
rect 210604 211674 211204 211676
rect 246604 211674 247204 211676
rect 282604 211674 283204 211676
rect 318604 211674 319204 211676
rect 354604 211674 355204 211676
rect 390604 211674 391204 211676
rect 426604 211674 427204 211676
rect 462604 211674 463204 211676
rect 498604 211674 499204 211676
rect 534604 211674 535204 211676
rect 570604 211674 571204 211676
rect 591900 211674 592500 211676
rect -6696 208676 -6096 208678
rect 27004 208676 27604 208678
rect 63004 208676 63604 208678
rect 99004 208676 99604 208678
rect 135004 208676 135604 208678
rect 171004 208676 171604 208678
rect 207004 208676 207604 208678
rect 243004 208676 243604 208678
rect 279004 208676 279604 208678
rect 315004 208676 315604 208678
rect 351004 208676 351604 208678
rect 387004 208676 387604 208678
rect 423004 208676 423604 208678
rect 459004 208676 459604 208678
rect 495004 208676 495604 208678
rect 531004 208676 531604 208678
rect 567004 208676 567604 208678
rect 590020 208676 590620 208678
rect -6696 208654 590620 208676
rect -6696 208418 -6514 208654
rect -6278 208418 27186 208654
rect 27422 208418 63186 208654
rect 63422 208418 99186 208654
rect 99422 208418 135186 208654
rect 135422 208418 171186 208654
rect 171422 208418 207186 208654
rect 207422 208418 243186 208654
rect 243422 208418 279186 208654
rect 279422 208418 315186 208654
rect 315422 208418 351186 208654
rect 351422 208418 387186 208654
rect 387422 208418 423186 208654
rect 423422 208418 459186 208654
rect 459422 208418 495186 208654
rect 495422 208418 531186 208654
rect 531422 208418 567186 208654
rect 567422 208418 590202 208654
rect 590438 208418 590620 208654
rect -6696 208334 590620 208418
rect -6696 208098 -6514 208334
rect -6278 208098 27186 208334
rect 27422 208098 63186 208334
rect 63422 208098 99186 208334
rect 99422 208098 135186 208334
rect 135422 208098 171186 208334
rect 171422 208098 207186 208334
rect 207422 208098 243186 208334
rect 243422 208098 279186 208334
rect 279422 208098 315186 208334
rect 315422 208098 351186 208334
rect 351422 208098 387186 208334
rect 387422 208098 423186 208334
rect 423422 208098 459186 208334
rect 459422 208098 495186 208334
rect 495422 208098 531186 208334
rect 531422 208098 567186 208334
rect 567422 208098 590202 208334
rect 590438 208098 590620 208334
rect -6696 208076 590620 208098
rect -6696 208074 -6096 208076
rect 27004 208074 27604 208076
rect 63004 208074 63604 208076
rect 99004 208074 99604 208076
rect 135004 208074 135604 208076
rect 171004 208074 171604 208076
rect 207004 208074 207604 208076
rect 243004 208074 243604 208076
rect 279004 208074 279604 208076
rect 315004 208074 315604 208076
rect 351004 208074 351604 208076
rect 387004 208074 387604 208076
rect 423004 208074 423604 208076
rect 459004 208074 459604 208076
rect 495004 208074 495604 208076
rect 531004 208074 531604 208076
rect 567004 208074 567604 208076
rect 590020 208074 590620 208076
rect -4816 205076 -4216 205078
rect 23404 205076 24004 205078
rect 59404 205076 60004 205078
rect 95404 205076 96004 205078
rect 131404 205076 132004 205078
rect 167404 205076 168004 205078
rect 203404 205076 204004 205078
rect 239404 205076 240004 205078
rect 275404 205076 276004 205078
rect 311404 205076 312004 205078
rect 347404 205076 348004 205078
rect 383404 205076 384004 205078
rect 419404 205076 420004 205078
rect 455404 205076 456004 205078
rect 491404 205076 492004 205078
rect 527404 205076 528004 205078
rect 563404 205076 564004 205078
rect 588140 205076 588740 205078
rect -4816 205054 588740 205076
rect -4816 204818 -4634 205054
rect -4398 204818 23586 205054
rect 23822 204818 59586 205054
rect 59822 204818 95586 205054
rect 95822 204818 131586 205054
rect 131822 204818 167586 205054
rect 167822 204818 203586 205054
rect 203822 204818 239586 205054
rect 239822 204818 275586 205054
rect 275822 204818 311586 205054
rect 311822 204818 347586 205054
rect 347822 204818 383586 205054
rect 383822 204818 419586 205054
rect 419822 204818 455586 205054
rect 455822 204818 491586 205054
rect 491822 204818 527586 205054
rect 527822 204818 563586 205054
rect 563822 204818 588322 205054
rect 588558 204818 588740 205054
rect -4816 204734 588740 204818
rect -4816 204498 -4634 204734
rect -4398 204498 23586 204734
rect 23822 204498 59586 204734
rect 59822 204498 95586 204734
rect 95822 204498 131586 204734
rect 131822 204498 167586 204734
rect 167822 204498 203586 204734
rect 203822 204498 239586 204734
rect 239822 204498 275586 204734
rect 275822 204498 311586 204734
rect 311822 204498 347586 204734
rect 347822 204498 383586 204734
rect 383822 204498 419586 204734
rect 419822 204498 455586 204734
rect 455822 204498 491586 204734
rect 491822 204498 527586 204734
rect 527822 204498 563586 204734
rect 563822 204498 588322 204734
rect 588558 204498 588740 204734
rect -4816 204476 588740 204498
rect -4816 204474 -4216 204476
rect 23404 204474 24004 204476
rect 59404 204474 60004 204476
rect 95404 204474 96004 204476
rect 131404 204474 132004 204476
rect 167404 204474 168004 204476
rect 203404 204474 204004 204476
rect 239404 204474 240004 204476
rect 275404 204474 276004 204476
rect 311404 204474 312004 204476
rect 347404 204474 348004 204476
rect 383404 204474 384004 204476
rect 419404 204474 420004 204476
rect 455404 204474 456004 204476
rect 491404 204474 492004 204476
rect 527404 204474 528004 204476
rect 563404 204474 564004 204476
rect 588140 204474 588740 204476
rect -2936 201476 -2336 201478
rect 19804 201476 20404 201478
rect 55804 201476 56404 201478
rect 91804 201476 92404 201478
rect 127804 201476 128404 201478
rect 163804 201476 164404 201478
rect 199804 201476 200404 201478
rect 235804 201476 236404 201478
rect 271804 201476 272404 201478
rect 307804 201476 308404 201478
rect 343804 201476 344404 201478
rect 379804 201476 380404 201478
rect 415804 201476 416404 201478
rect 451804 201476 452404 201478
rect 487804 201476 488404 201478
rect 523804 201476 524404 201478
rect 559804 201476 560404 201478
rect 586260 201476 586860 201478
rect -2936 201454 586860 201476
rect -2936 201218 -2754 201454
rect -2518 201218 19986 201454
rect 20222 201218 55986 201454
rect 56222 201218 91986 201454
rect 92222 201218 127986 201454
rect 128222 201218 163986 201454
rect 164222 201218 199986 201454
rect 200222 201218 235986 201454
rect 236222 201218 271986 201454
rect 272222 201218 307986 201454
rect 308222 201218 343986 201454
rect 344222 201218 379986 201454
rect 380222 201218 415986 201454
rect 416222 201218 451986 201454
rect 452222 201218 487986 201454
rect 488222 201218 523986 201454
rect 524222 201218 559986 201454
rect 560222 201218 586442 201454
rect 586678 201218 586860 201454
rect -2936 201134 586860 201218
rect -2936 200898 -2754 201134
rect -2518 200898 19986 201134
rect 20222 200898 55986 201134
rect 56222 200898 91986 201134
rect 92222 200898 127986 201134
rect 128222 200898 163986 201134
rect 164222 200898 199986 201134
rect 200222 200898 235986 201134
rect 236222 200898 271986 201134
rect 272222 200898 307986 201134
rect 308222 200898 343986 201134
rect 344222 200898 379986 201134
rect 380222 200898 415986 201134
rect 416222 200898 451986 201134
rect 452222 200898 487986 201134
rect 488222 200898 523986 201134
rect 524222 200898 559986 201134
rect 560222 200898 586442 201134
rect 586678 200898 586860 201134
rect -2936 200876 586860 200898
rect -2936 200874 -2336 200876
rect 19804 200874 20404 200876
rect 55804 200874 56404 200876
rect 91804 200874 92404 200876
rect 127804 200874 128404 200876
rect 163804 200874 164404 200876
rect 199804 200874 200404 200876
rect 235804 200874 236404 200876
rect 271804 200874 272404 200876
rect 307804 200874 308404 200876
rect 343804 200874 344404 200876
rect 379804 200874 380404 200876
rect 415804 200874 416404 200876
rect 451804 200874 452404 200876
rect 487804 200874 488404 200876
rect 523804 200874 524404 200876
rect 559804 200874 560404 200876
rect 586260 200874 586860 200876
rect -7636 194276 -7036 194278
rect 12604 194276 13204 194278
rect 48604 194276 49204 194278
rect 84604 194276 85204 194278
rect 120604 194276 121204 194278
rect 156604 194276 157204 194278
rect 192604 194276 193204 194278
rect 228604 194276 229204 194278
rect 264604 194276 265204 194278
rect 300604 194276 301204 194278
rect 336604 194276 337204 194278
rect 372604 194276 373204 194278
rect 408604 194276 409204 194278
rect 444604 194276 445204 194278
rect 480604 194276 481204 194278
rect 516604 194276 517204 194278
rect 552604 194276 553204 194278
rect 590960 194276 591560 194278
rect -8576 194254 592500 194276
rect -8576 194018 -7454 194254
rect -7218 194018 12786 194254
rect 13022 194018 48786 194254
rect 49022 194018 84786 194254
rect 85022 194018 120786 194254
rect 121022 194018 156786 194254
rect 157022 194018 192786 194254
rect 193022 194018 228786 194254
rect 229022 194018 264786 194254
rect 265022 194018 300786 194254
rect 301022 194018 336786 194254
rect 337022 194018 372786 194254
rect 373022 194018 408786 194254
rect 409022 194018 444786 194254
rect 445022 194018 480786 194254
rect 481022 194018 516786 194254
rect 517022 194018 552786 194254
rect 553022 194018 591142 194254
rect 591378 194018 592500 194254
rect -8576 193934 592500 194018
rect -8576 193698 -7454 193934
rect -7218 193698 12786 193934
rect 13022 193698 48786 193934
rect 49022 193698 84786 193934
rect 85022 193698 120786 193934
rect 121022 193698 156786 193934
rect 157022 193698 192786 193934
rect 193022 193698 228786 193934
rect 229022 193698 264786 193934
rect 265022 193698 300786 193934
rect 301022 193698 336786 193934
rect 337022 193698 372786 193934
rect 373022 193698 408786 193934
rect 409022 193698 444786 193934
rect 445022 193698 480786 193934
rect 481022 193698 516786 193934
rect 517022 193698 552786 193934
rect 553022 193698 591142 193934
rect 591378 193698 592500 193934
rect -8576 193676 592500 193698
rect -7636 193674 -7036 193676
rect 12604 193674 13204 193676
rect 48604 193674 49204 193676
rect 84604 193674 85204 193676
rect 120604 193674 121204 193676
rect 156604 193674 157204 193676
rect 192604 193674 193204 193676
rect 228604 193674 229204 193676
rect 264604 193674 265204 193676
rect 300604 193674 301204 193676
rect 336604 193674 337204 193676
rect 372604 193674 373204 193676
rect 408604 193674 409204 193676
rect 444604 193674 445204 193676
rect 480604 193674 481204 193676
rect 516604 193674 517204 193676
rect 552604 193674 553204 193676
rect 590960 193674 591560 193676
rect -5756 190676 -5156 190678
rect 9004 190676 9604 190678
rect 45004 190676 45604 190678
rect 81004 190676 81604 190678
rect 117004 190676 117604 190678
rect 153004 190676 153604 190678
rect 189004 190676 189604 190678
rect 225004 190676 225604 190678
rect 261004 190676 261604 190678
rect 297004 190676 297604 190678
rect 333004 190676 333604 190678
rect 369004 190676 369604 190678
rect 405004 190676 405604 190678
rect 441004 190676 441604 190678
rect 477004 190676 477604 190678
rect 513004 190676 513604 190678
rect 549004 190676 549604 190678
rect 589080 190676 589680 190678
rect -6696 190654 590620 190676
rect -6696 190418 -5574 190654
rect -5338 190418 9186 190654
rect 9422 190418 45186 190654
rect 45422 190418 81186 190654
rect 81422 190418 117186 190654
rect 117422 190418 153186 190654
rect 153422 190418 189186 190654
rect 189422 190418 225186 190654
rect 225422 190418 261186 190654
rect 261422 190418 297186 190654
rect 297422 190418 333186 190654
rect 333422 190418 369186 190654
rect 369422 190418 405186 190654
rect 405422 190418 441186 190654
rect 441422 190418 477186 190654
rect 477422 190418 513186 190654
rect 513422 190418 549186 190654
rect 549422 190418 589262 190654
rect 589498 190418 590620 190654
rect -6696 190334 590620 190418
rect -6696 190098 -5574 190334
rect -5338 190098 9186 190334
rect 9422 190098 45186 190334
rect 45422 190098 81186 190334
rect 81422 190098 117186 190334
rect 117422 190098 153186 190334
rect 153422 190098 189186 190334
rect 189422 190098 225186 190334
rect 225422 190098 261186 190334
rect 261422 190098 297186 190334
rect 297422 190098 333186 190334
rect 333422 190098 369186 190334
rect 369422 190098 405186 190334
rect 405422 190098 441186 190334
rect 441422 190098 477186 190334
rect 477422 190098 513186 190334
rect 513422 190098 549186 190334
rect 549422 190098 589262 190334
rect 589498 190098 590620 190334
rect -6696 190076 590620 190098
rect -5756 190074 -5156 190076
rect 9004 190074 9604 190076
rect 45004 190074 45604 190076
rect 81004 190074 81604 190076
rect 117004 190074 117604 190076
rect 153004 190074 153604 190076
rect 189004 190074 189604 190076
rect 225004 190074 225604 190076
rect 261004 190074 261604 190076
rect 297004 190074 297604 190076
rect 333004 190074 333604 190076
rect 369004 190074 369604 190076
rect 405004 190074 405604 190076
rect 441004 190074 441604 190076
rect 477004 190074 477604 190076
rect 513004 190074 513604 190076
rect 549004 190074 549604 190076
rect 589080 190074 589680 190076
rect -3876 187076 -3276 187078
rect 5404 187076 6004 187078
rect 41404 187076 42004 187078
rect 77404 187076 78004 187078
rect 113404 187076 114004 187078
rect 149404 187076 150004 187078
rect 185404 187076 186004 187078
rect 221404 187076 222004 187078
rect 257404 187076 258004 187078
rect 293404 187076 294004 187078
rect 329404 187076 330004 187078
rect 365404 187076 366004 187078
rect 401404 187076 402004 187078
rect 437404 187076 438004 187078
rect 473404 187076 474004 187078
rect 509404 187076 510004 187078
rect 545404 187076 546004 187078
rect 581404 187076 582004 187078
rect 587200 187076 587800 187078
rect -4816 187054 588740 187076
rect -4816 186818 -3694 187054
rect -3458 186818 5586 187054
rect 5822 186818 41586 187054
rect 41822 186818 77586 187054
rect 77822 186818 113586 187054
rect 113822 186818 149586 187054
rect 149822 186818 185586 187054
rect 185822 186818 221586 187054
rect 221822 186818 257586 187054
rect 257822 186818 293586 187054
rect 293822 186818 329586 187054
rect 329822 186818 365586 187054
rect 365822 186818 401586 187054
rect 401822 186818 437586 187054
rect 437822 186818 473586 187054
rect 473822 186818 509586 187054
rect 509822 186818 545586 187054
rect 545822 186818 581586 187054
rect 581822 186818 587382 187054
rect 587618 186818 588740 187054
rect -4816 186734 588740 186818
rect -4816 186498 -3694 186734
rect -3458 186498 5586 186734
rect 5822 186498 41586 186734
rect 41822 186498 77586 186734
rect 77822 186498 113586 186734
rect 113822 186498 149586 186734
rect 149822 186498 185586 186734
rect 185822 186498 221586 186734
rect 221822 186498 257586 186734
rect 257822 186498 293586 186734
rect 293822 186498 329586 186734
rect 329822 186498 365586 186734
rect 365822 186498 401586 186734
rect 401822 186498 437586 186734
rect 437822 186498 473586 186734
rect 473822 186498 509586 186734
rect 509822 186498 545586 186734
rect 545822 186498 581586 186734
rect 581822 186498 587382 186734
rect 587618 186498 588740 186734
rect -4816 186476 588740 186498
rect -3876 186474 -3276 186476
rect 5404 186474 6004 186476
rect 41404 186474 42004 186476
rect 77404 186474 78004 186476
rect 113404 186474 114004 186476
rect 149404 186474 150004 186476
rect 185404 186474 186004 186476
rect 221404 186474 222004 186476
rect 257404 186474 258004 186476
rect 293404 186474 294004 186476
rect 329404 186474 330004 186476
rect 365404 186474 366004 186476
rect 401404 186474 402004 186476
rect 437404 186474 438004 186476
rect 473404 186474 474004 186476
rect 509404 186474 510004 186476
rect 545404 186474 546004 186476
rect 581404 186474 582004 186476
rect 587200 186474 587800 186476
rect -1996 183476 -1396 183478
rect 1804 183476 2404 183478
rect 37804 183476 38404 183478
rect 73804 183476 74404 183478
rect 109804 183476 110404 183478
rect 145804 183476 146404 183478
rect 181804 183476 182404 183478
rect 217804 183476 218404 183478
rect 253804 183476 254404 183478
rect 289804 183476 290404 183478
rect 325804 183476 326404 183478
rect 361804 183476 362404 183478
rect 397804 183476 398404 183478
rect 433804 183476 434404 183478
rect 469804 183476 470404 183478
rect 505804 183476 506404 183478
rect 541804 183476 542404 183478
rect 577804 183476 578404 183478
rect 585320 183476 585920 183478
rect -2936 183454 586860 183476
rect -2936 183218 -1814 183454
rect -1578 183218 1986 183454
rect 2222 183218 37986 183454
rect 38222 183218 73986 183454
rect 74222 183218 109986 183454
rect 110222 183218 145986 183454
rect 146222 183218 181986 183454
rect 182222 183218 217986 183454
rect 218222 183218 253986 183454
rect 254222 183218 289986 183454
rect 290222 183218 325986 183454
rect 326222 183218 361986 183454
rect 362222 183218 397986 183454
rect 398222 183218 433986 183454
rect 434222 183218 469986 183454
rect 470222 183218 505986 183454
rect 506222 183218 541986 183454
rect 542222 183218 577986 183454
rect 578222 183218 585502 183454
rect 585738 183218 586860 183454
rect -2936 183134 586860 183218
rect -2936 182898 -1814 183134
rect -1578 182898 1986 183134
rect 2222 182898 37986 183134
rect 38222 182898 73986 183134
rect 74222 182898 109986 183134
rect 110222 182898 145986 183134
rect 146222 182898 181986 183134
rect 182222 182898 217986 183134
rect 218222 182898 253986 183134
rect 254222 182898 289986 183134
rect 290222 182898 325986 183134
rect 326222 182898 361986 183134
rect 362222 182898 397986 183134
rect 398222 182898 433986 183134
rect 434222 182898 469986 183134
rect 470222 182898 505986 183134
rect 506222 182898 541986 183134
rect 542222 182898 577986 183134
rect 578222 182898 585502 183134
rect 585738 182898 586860 183134
rect -2936 182876 586860 182898
rect -1996 182874 -1396 182876
rect 1804 182874 2404 182876
rect 37804 182874 38404 182876
rect 73804 182874 74404 182876
rect 109804 182874 110404 182876
rect 145804 182874 146404 182876
rect 181804 182874 182404 182876
rect 217804 182874 218404 182876
rect 253804 182874 254404 182876
rect 289804 182874 290404 182876
rect 325804 182874 326404 182876
rect 361804 182874 362404 182876
rect 397804 182874 398404 182876
rect 433804 182874 434404 182876
rect 469804 182874 470404 182876
rect 505804 182874 506404 182876
rect 541804 182874 542404 182876
rect 577804 182874 578404 182876
rect 585320 182874 585920 182876
rect -8576 176276 -7976 176278
rect 30604 176276 31204 176278
rect 66604 176276 67204 176278
rect 102604 176276 103204 176278
rect 138604 176276 139204 176278
rect 174604 176276 175204 176278
rect 210604 176276 211204 176278
rect 246604 176276 247204 176278
rect 282604 176276 283204 176278
rect 318604 176276 319204 176278
rect 354604 176276 355204 176278
rect 390604 176276 391204 176278
rect 426604 176276 427204 176278
rect 462604 176276 463204 176278
rect 498604 176276 499204 176278
rect 534604 176276 535204 176278
rect 570604 176276 571204 176278
rect 591900 176276 592500 176278
rect -8576 176254 592500 176276
rect -8576 176018 -8394 176254
rect -8158 176018 30786 176254
rect 31022 176018 66786 176254
rect 67022 176018 102786 176254
rect 103022 176018 138786 176254
rect 139022 176018 174786 176254
rect 175022 176018 210786 176254
rect 211022 176018 246786 176254
rect 247022 176018 282786 176254
rect 283022 176018 318786 176254
rect 319022 176018 354786 176254
rect 355022 176018 390786 176254
rect 391022 176018 426786 176254
rect 427022 176018 462786 176254
rect 463022 176018 498786 176254
rect 499022 176018 534786 176254
rect 535022 176018 570786 176254
rect 571022 176018 592082 176254
rect 592318 176018 592500 176254
rect -8576 175934 592500 176018
rect -8576 175698 -8394 175934
rect -8158 175698 30786 175934
rect 31022 175698 66786 175934
rect 67022 175698 102786 175934
rect 103022 175698 138786 175934
rect 139022 175698 174786 175934
rect 175022 175698 210786 175934
rect 211022 175698 246786 175934
rect 247022 175698 282786 175934
rect 283022 175698 318786 175934
rect 319022 175698 354786 175934
rect 355022 175698 390786 175934
rect 391022 175698 426786 175934
rect 427022 175698 462786 175934
rect 463022 175698 498786 175934
rect 499022 175698 534786 175934
rect 535022 175698 570786 175934
rect 571022 175698 592082 175934
rect 592318 175698 592500 175934
rect -8576 175676 592500 175698
rect -8576 175674 -7976 175676
rect 30604 175674 31204 175676
rect 66604 175674 67204 175676
rect 102604 175674 103204 175676
rect 138604 175674 139204 175676
rect 174604 175674 175204 175676
rect 210604 175674 211204 175676
rect 246604 175674 247204 175676
rect 282604 175674 283204 175676
rect 318604 175674 319204 175676
rect 354604 175674 355204 175676
rect 390604 175674 391204 175676
rect 426604 175674 427204 175676
rect 462604 175674 463204 175676
rect 498604 175674 499204 175676
rect 534604 175674 535204 175676
rect 570604 175674 571204 175676
rect 591900 175674 592500 175676
rect -6696 172676 -6096 172678
rect 27004 172676 27604 172678
rect 63004 172676 63604 172678
rect 99004 172676 99604 172678
rect 135004 172676 135604 172678
rect 171004 172676 171604 172678
rect 207004 172676 207604 172678
rect 243004 172676 243604 172678
rect 279004 172676 279604 172678
rect 315004 172676 315604 172678
rect 351004 172676 351604 172678
rect 387004 172676 387604 172678
rect 423004 172676 423604 172678
rect 459004 172676 459604 172678
rect 495004 172676 495604 172678
rect 531004 172676 531604 172678
rect 567004 172676 567604 172678
rect 590020 172676 590620 172678
rect -6696 172654 590620 172676
rect -6696 172418 -6514 172654
rect -6278 172418 27186 172654
rect 27422 172418 63186 172654
rect 63422 172418 99186 172654
rect 99422 172418 135186 172654
rect 135422 172418 171186 172654
rect 171422 172418 207186 172654
rect 207422 172418 243186 172654
rect 243422 172418 279186 172654
rect 279422 172418 315186 172654
rect 315422 172418 351186 172654
rect 351422 172418 387186 172654
rect 387422 172418 423186 172654
rect 423422 172418 459186 172654
rect 459422 172418 495186 172654
rect 495422 172418 531186 172654
rect 531422 172418 567186 172654
rect 567422 172418 590202 172654
rect 590438 172418 590620 172654
rect -6696 172334 590620 172418
rect -6696 172098 -6514 172334
rect -6278 172098 27186 172334
rect 27422 172098 63186 172334
rect 63422 172098 99186 172334
rect 99422 172098 135186 172334
rect 135422 172098 171186 172334
rect 171422 172098 207186 172334
rect 207422 172098 243186 172334
rect 243422 172098 279186 172334
rect 279422 172098 315186 172334
rect 315422 172098 351186 172334
rect 351422 172098 387186 172334
rect 387422 172098 423186 172334
rect 423422 172098 459186 172334
rect 459422 172098 495186 172334
rect 495422 172098 531186 172334
rect 531422 172098 567186 172334
rect 567422 172098 590202 172334
rect 590438 172098 590620 172334
rect -6696 172076 590620 172098
rect -6696 172074 -6096 172076
rect 27004 172074 27604 172076
rect 63004 172074 63604 172076
rect 99004 172074 99604 172076
rect 135004 172074 135604 172076
rect 171004 172074 171604 172076
rect 207004 172074 207604 172076
rect 243004 172074 243604 172076
rect 279004 172074 279604 172076
rect 315004 172074 315604 172076
rect 351004 172074 351604 172076
rect 387004 172074 387604 172076
rect 423004 172074 423604 172076
rect 459004 172074 459604 172076
rect 495004 172074 495604 172076
rect 531004 172074 531604 172076
rect 567004 172074 567604 172076
rect 590020 172074 590620 172076
rect -4816 169076 -4216 169078
rect 23404 169076 24004 169078
rect 59404 169076 60004 169078
rect 95404 169076 96004 169078
rect 131404 169076 132004 169078
rect 167404 169076 168004 169078
rect 203404 169076 204004 169078
rect 239404 169076 240004 169078
rect 275404 169076 276004 169078
rect 311404 169076 312004 169078
rect 347404 169076 348004 169078
rect 383404 169076 384004 169078
rect 419404 169076 420004 169078
rect 455404 169076 456004 169078
rect 491404 169076 492004 169078
rect 527404 169076 528004 169078
rect 563404 169076 564004 169078
rect 588140 169076 588740 169078
rect -4816 169054 588740 169076
rect -4816 168818 -4634 169054
rect -4398 168818 23586 169054
rect 23822 168818 59586 169054
rect 59822 168818 95586 169054
rect 95822 168818 131586 169054
rect 131822 168818 167586 169054
rect 167822 168818 203586 169054
rect 203822 168818 239586 169054
rect 239822 168818 275586 169054
rect 275822 168818 311586 169054
rect 311822 168818 347586 169054
rect 347822 168818 383586 169054
rect 383822 168818 419586 169054
rect 419822 168818 455586 169054
rect 455822 168818 491586 169054
rect 491822 168818 527586 169054
rect 527822 168818 563586 169054
rect 563822 168818 588322 169054
rect 588558 168818 588740 169054
rect -4816 168734 588740 168818
rect -4816 168498 -4634 168734
rect -4398 168498 23586 168734
rect 23822 168498 59586 168734
rect 59822 168498 95586 168734
rect 95822 168498 131586 168734
rect 131822 168498 167586 168734
rect 167822 168498 203586 168734
rect 203822 168498 239586 168734
rect 239822 168498 275586 168734
rect 275822 168498 311586 168734
rect 311822 168498 347586 168734
rect 347822 168498 383586 168734
rect 383822 168498 419586 168734
rect 419822 168498 455586 168734
rect 455822 168498 491586 168734
rect 491822 168498 527586 168734
rect 527822 168498 563586 168734
rect 563822 168498 588322 168734
rect 588558 168498 588740 168734
rect -4816 168476 588740 168498
rect -4816 168474 -4216 168476
rect 23404 168474 24004 168476
rect 59404 168474 60004 168476
rect 95404 168474 96004 168476
rect 131404 168474 132004 168476
rect 167404 168474 168004 168476
rect 203404 168474 204004 168476
rect 239404 168474 240004 168476
rect 275404 168474 276004 168476
rect 311404 168474 312004 168476
rect 347404 168474 348004 168476
rect 383404 168474 384004 168476
rect 419404 168474 420004 168476
rect 455404 168474 456004 168476
rect 491404 168474 492004 168476
rect 527404 168474 528004 168476
rect 563404 168474 564004 168476
rect 588140 168474 588740 168476
rect -2936 165476 -2336 165478
rect 19804 165476 20404 165478
rect 55804 165476 56404 165478
rect 91804 165476 92404 165478
rect 127804 165476 128404 165478
rect 163804 165476 164404 165478
rect 199804 165476 200404 165478
rect 235804 165476 236404 165478
rect 271804 165476 272404 165478
rect 307804 165476 308404 165478
rect 343804 165476 344404 165478
rect 379804 165476 380404 165478
rect 415804 165476 416404 165478
rect 451804 165476 452404 165478
rect 487804 165476 488404 165478
rect 523804 165476 524404 165478
rect 559804 165476 560404 165478
rect 586260 165476 586860 165478
rect -2936 165454 586860 165476
rect -2936 165218 -2754 165454
rect -2518 165218 19986 165454
rect 20222 165218 55986 165454
rect 56222 165218 91986 165454
rect 92222 165218 127986 165454
rect 128222 165218 163986 165454
rect 164222 165218 199986 165454
rect 200222 165218 235986 165454
rect 236222 165218 271986 165454
rect 272222 165218 307986 165454
rect 308222 165218 343986 165454
rect 344222 165218 379986 165454
rect 380222 165218 415986 165454
rect 416222 165218 451986 165454
rect 452222 165218 487986 165454
rect 488222 165218 523986 165454
rect 524222 165218 559986 165454
rect 560222 165218 586442 165454
rect 586678 165218 586860 165454
rect -2936 165134 586860 165218
rect -2936 164898 -2754 165134
rect -2518 164898 19986 165134
rect 20222 164898 55986 165134
rect 56222 164898 91986 165134
rect 92222 164898 127986 165134
rect 128222 164898 163986 165134
rect 164222 164898 199986 165134
rect 200222 164898 235986 165134
rect 236222 164898 271986 165134
rect 272222 164898 307986 165134
rect 308222 164898 343986 165134
rect 344222 164898 379986 165134
rect 380222 164898 415986 165134
rect 416222 164898 451986 165134
rect 452222 164898 487986 165134
rect 488222 164898 523986 165134
rect 524222 164898 559986 165134
rect 560222 164898 586442 165134
rect 586678 164898 586860 165134
rect -2936 164876 586860 164898
rect -2936 164874 -2336 164876
rect 19804 164874 20404 164876
rect 55804 164874 56404 164876
rect 91804 164874 92404 164876
rect 127804 164874 128404 164876
rect 163804 164874 164404 164876
rect 199804 164874 200404 164876
rect 235804 164874 236404 164876
rect 271804 164874 272404 164876
rect 307804 164874 308404 164876
rect 343804 164874 344404 164876
rect 379804 164874 380404 164876
rect 415804 164874 416404 164876
rect 451804 164874 452404 164876
rect 487804 164874 488404 164876
rect 523804 164874 524404 164876
rect 559804 164874 560404 164876
rect 586260 164874 586860 164876
rect -7636 158276 -7036 158278
rect 12604 158276 13204 158278
rect 48604 158276 49204 158278
rect 84604 158276 85204 158278
rect 120604 158276 121204 158278
rect 156604 158276 157204 158278
rect 192604 158276 193204 158278
rect 228604 158276 229204 158278
rect 264604 158276 265204 158278
rect 300604 158276 301204 158278
rect 336604 158276 337204 158278
rect 372604 158276 373204 158278
rect 408604 158276 409204 158278
rect 444604 158276 445204 158278
rect 480604 158276 481204 158278
rect 516604 158276 517204 158278
rect 552604 158276 553204 158278
rect 590960 158276 591560 158278
rect -8576 158254 592500 158276
rect -8576 158018 -7454 158254
rect -7218 158018 12786 158254
rect 13022 158018 48786 158254
rect 49022 158018 84786 158254
rect 85022 158018 120786 158254
rect 121022 158018 156786 158254
rect 157022 158018 192786 158254
rect 193022 158018 228786 158254
rect 229022 158018 264786 158254
rect 265022 158018 300786 158254
rect 301022 158018 336786 158254
rect 337022 158018 372786 158254
rect 373022 158018 408786 158254
rect 409022 158018 444786 158254
rect 445022 158018 480786 158254
rect 481022 158018 516786 158254
rect 517022 158018 552786 158254
rect 553022 158018 591142 158254
rect 591378 158018 592500 158254
rect -8576 157934 592500 158018
rect -8576 157698 -7454 157934
rect -7218 157698 12786 157934
rect 13022 157698 48786 157934
rect 49022 157698 84786 157934
rect 85022 157698 120786 157934
rect 121022 157698 156786 157934
rect 157022 157698 192786 157934
rect 193022 157698 228786 157934
rect 229022 157698 264786 157934
rect 265022 157698 300786 157934
rect 301022 157698 336786 157934
rect 337022 157698 372786 157934
rect 373022 157698 408786 157934
rect 409022 157698 444786 157934
rect 445022 157698 480786 157934
rect 481022 157698 516786 157934
rect 517022 157698 552786 157934
rect 553022 157698 591142 157934
rect 591378 157698 592500 157934
rect -8576 157676 592500 157698
rect -7636 157674 -7036 157676
rect 12604 157674 13204 157676
rect 48604 157674 49204 157676
rect 84604 157674 85204 157676
rect 120604 157674 121204 157676
rect 156604 157674 157204 157676
rect 192604 157674 193204 157676
rect 228604 157674 229204 157676
rect 264604 157674 265204 157676
rect 300604 157674 301204 157676
rect 336604 157674 337204 157676
rect 372604 157674 373204 157676
rect 408604 157674 409204 157676
rect 444604 157674 445204 157676
rect 480604 157674 481204 157676
rect 516604 157674 517204 157676
rect 552604 157674 553204 157676
rect 590960 157674 591560 157676
rect -5756 154676 -5156 154678
rect 9004 154676 9604 154678
rect 45004 154676 45604 154678
rect 81004 154676 81604 154678
rect 117004 154676 117604 154678
rect 153004 154676 153604 154678
rect 189004 154676 189604 154678
rect 225004 154676 225604 154678
rect 261004 154676 261604 154678
rect 297004 154676 297604 154678
rect 333004 154676 333604 154678
rect 369004 154676 369604 154678
rect 405004 154676 405604 154678
rect 441004 154676 441604 154678
rect 477004 154676 477604 154678
rect 513004 154676 513604 154678
rect 549004 154676 549604 154678
rect 589080 154676 589680 154678
rect -6696 154654 590620 154676
rect -6696 154418 -5574 154654
rect -5338 154418 9186 154654
rect 9422 154418 45186 154654
rect 45422 154418 81186 154654
rect 81422 154418 117186 154654
rect 117422 154418 153186 154654
rect 153422 154418 189186 154654
rect 189422 154418 225186 154654
rect 225422 154418 261186 154654
rect 261422 154418 297186 154654
rect 297422 154418 333186 154654
rect 333422 154418 369186 154654
rect 369422 154418 405186 154654
rect 405422 154418 441186 154654
rect 441422 154418 477186 154654
rect 477422 154418 513186 154654
rect 513422 154418 549186 154654
rect 549422 154418 589262 154654
rect 589498 154418 590620 154654
rect -6696 154334 590620 154418
rect -6696 154098 -5574 154334
rect -5338 154098 9186 154334
rect 9422 154098 45186 154334
rect 45422 154098 81186 154334
rect 81422 154098 117186 154334
rect 117422 154098 153186 154334
rect 153422 154098 189186 154334
rect 189422 154098 225186 154334
rect 225422 154098 261186 154334
rect 261422 154098 297186 154334
rect 297422 154098 333186 154334
rect 333422 154098 369186 154334
rect 369422 154098 405186 154334
rect 405422 154098 441186 154334
rect 441422 154098 477186 154334
rect 477422 154098 513186 154334
rect 513422 154098 549186 154334
rect 549422 154098 589262 154334
rect 589498 154098 590620 154334
rect -6696 154076 590620 154098
rect -5756 154074 -5156 154076
rect 9004 154074 9604 154076
rect 45004 154074 45604 154076
rect 81004 154074 81604 154076
rect 117004 154074 117604 154076
rect 153004 154074 153604 154076
rect 189004 154074 189604 154076
rect 225004 154074 225604 154076
rect 261004 154074 261604 154076
rect 297004 154074 297604 154076
rect 333004 154074 333604 154076
rect 369004 154074 369604 154076
rect 405004 154074 405604 154076
rect 441004 154074 441604 154076
rect 477004 154074 477604 154076
rect 513004 154074 513604 154076
rect 549004 154074 549604 154076
rect 589080 154074 589680 154076
rect -3876 151076 -3276 151078
rect 5404 151076 6004 151078
rect 41404 151076 42004 151078
rect 77404 151076 78004 151078
rect 113404 151076 114004 151078
rect 149404 151076 150004 151078
rect 185404 151076 186004 151078
rect 221404 151076 222004 151078
rect 257404 151076 258004 151078
rect 293404 151076 294004 151078
rect 329404 151076 330004 151078
rect 365404 151076 366004 151078
rect 401404 151076 402004 151078
rect 437404 151076 438004 151078
rect 473404 151076 474004 151078
rect 509404 151076 510004 151078
rect 545404 151076 546004 151078
rect 581404 151076 582004 151078
rect 587200 151076 587800 151078
rect -4816 151054 588740 151076
rect -4816 150818 -3694 151054
rect -3458 150818 5586 151054
rect 5822 150818 41586 151054
rect 41822 150818 77586 151054
rect 77822 150818 113586 151054
rect 113822 150818 149586 151054
rect 149822 150818 185586 151054
rect 185822 150818 221586 151054
rect 221822 150818 257586 151054
rect 257822 150818 293586 151054
rect 293822 150818 329586 151054
rect 329822 150818 365586 151054
rect 365822 150818 401586 151054
rect 401822 150818 437586 151054
rect 437822 150818 473586 151054
rect 473822 150818 509586 151054
rect 509822 150818 545586 151054
rect 545822 150818 581586 151054
rect 581822 150818 587382 151054
rect 587618 150818 588740 151054
rect -4816 150734 588740 150818
rect -4816 150498 -3694 150734
rect -3458 150498 5586 150734
rect 5822 150498 41586 150734
rect 41822 150498 77586 150734
rect 77822 150498 113586 150734
rect 113822 150498 149586 150734
rect 149822 150498 185586 150734
rect 185822 150498 221586 150734
rect 221822 150498 257586 150734
rect 257822 150498 293586 150734
rect 293822 150498 329586 150734
rect 329822 150498 365586 150734
rect 365822 150498 401586 150734
rect 401822 150498 437586 150734
rect 437822 150498 473586 150734
rect 473822 150498 509586 150734
rect 509822 150498 545586 150734
rect 545822 150498 581586 150734
rect 581822 150498 587382 150734
rect 587618 150498 588740 150734
rect -4816 150476 588740 150498
rect -3876 150474 -3276 150476
rect 5404 150474 6004 150476
rect 41404 150474 42004 150476
rect 77404 150474 78004 150476
rect 113404 150474 114004 150476
rect 149404 150474 150004 150476
rect 185404 150474 186004 150476
rect 221404 150474 222004 150476
rect 257404 150474 258004 150476
rect 293404 150474 294004 150476
rect 329404 150474 330004 150476
rect 365404 150474 366004 150476
rect 401404 150474 402004 150476
rect 437404 150474 438004 150476
rect 473404 150474 474004 150476
rect 509404 150474 510004 150476
rect 545404 150474 546004 150476
rect 581404 150474 582004 150476
rect 587200 150474 587800 150476
rect -1996 147476 -1396 147478
rect 1804 147476 2404 147478
rect 37804 147476 38404 147478
rect 73804 147476 74404 147478
rect 109804 147476 110404 147478
rect 145804 147476 146404 147478
rect 181804 147476 182404 147478
rect 217804 147476 218404 147478
rect 253804 147476 254404 147478
rect 289804 147476 290404 147478
rect 325804 147476 326404 147478
rect 361804 147476 362404 147478
rect 397804 147476 398404 147478
rect 433804 147476 434404 147478
rect 469804 147476 470404 147478
rect 505804 147476 506404 147478
rect 541804 147476 542404 147478
rect 577804 147476 578404 147478
rect 585320 147476 585920 147478
rect -2936 147454 586860 147476
rect -2936 147218 -1814 147454
rect -1578 147218 1986 147454
rect 2222 147218 37986 147454
rect 38222 147218 73986 147454
rect 74222 147218 109986 147454
rect 110222 147218 145986 147454
rect 146222 147218 181986 147454
rect 182222 147218 217986 147454
rect 218222 147218 253986 147454
rect 254222 147218 289986 147454
rect 290222 147218 325986 147454
rect 326222 147218 361986 147454
rect 362222 147218 397986 147454
rect 398222 147218 433986 147454
rect 434222 147218 469986 147454
rect 470222 147218 505986 147454
rect 506222 147218 541986 147454
rect 542222 147218 577986 147454
rect 578222 147218 585502 147454
rect 585738 147218 586860 147454
rect -2936 147134 586860 147218
rect -2936 146898 -1814 147134
rect -1578 146898 1986 147134
rect 2222 146898 37986 147134
rect 38222 146898 73986 147134
rect 74222 146898 109986 147134
rect 110222 146898 145986 147134
rect 146222 146898 181986 147134
rect 182222 146898 217986 147134
rect 218222 146898 253986 147134
rect 254222 146898 289986 147134
rect 290222 146898 325986 147134
rect 326222 146898 361986 147134
rect 362222 146898 397986 147134
rect 398222 146898 433986 147134
rect 434222 146898 469986 147134
rect 470222 146898 505986 147134
rect 506222 146898 541986 147134
rect 542222 146898 577986 147134
rect 578222 146898 585502 147134
rect 585738 146898 586860 147134
rect -2936 146876 586860 146898
rect -1996 146874 -1396 146876
rect 1804 146874 2404 146876
rect 37804 146874 38404 146876
rect 73804 146874 74404 146876
rect 109804 146874 110404 146876
rect 145804 146874 146404 146876
rect 181804 146874 182404 146876
rect 217804 146874 218404 146876
rect 253804 146874 254404 146876
rect 289804 146874 290404 146876
rect 325804 146874 326404 146876
rect 361804 146874 362404 146876
rect 397804 146874 398404 146876
rect 433804 146874 434404 146876
rect 469804 146874 470404 146876
rect 505804 146874 506404 146876
rect 541804 146874 542404 146876
rect 577804 146874 578404 146876
rect 585320 146874 585920 146876
rect -8576 140276 -7976 140278
rect 30604 140276 31204 140278
rect 66604 140276 67204 140278
rect 102604 140276 103204 140278
rect 138604 140276 139204 140278
rect 174604 140276 175204 140278
rect 210604 140276 211204 140278
rect 246604 140276 247204 140278
rect 282604 140276 283204 140278
rect 318604 140276 319204 140278
rect 354604 140276 355204 140278
rect 390604 140276 391204 140278
rect 426604 140276 427204 140278
rect 462604 140276 463204 140278
rect 498604 140276 499204 140278
rect 534604 140276 535204 140278
rect 570604 140276 571204 140278
rect 591900 140276 592500 140278
rect -8576 140254 592500 140276
rect -8576 140018 -8394 140254
rect -8158 140018 30786 140254
rect 31022 140018 66786 140254
rect 67022 140018 102786 140254
rect 103022 140018 138786 140254
rect 139022 140018 174786 140254
rect 175022 140018 210786 140254
rect 211022 140018 246786 140254
rect 247022 140018 282786 140254
rect 283022 140018 318786 140254
rect 319022 140018 354786 140254
rect 355022 140018 390786 140254
rect 391022 140018 426786 140254
rect 427022 140018 462786 140254
rect 463022 140018 498786 140254
rect 499022 140018 534786 140254
rect 535022 140018 570786 140254
rect 571022 140018 592082 140254
rect 592318 140018 592500 140254
rect -8576 139934 592500 140018
rect -8576 139698 -8394 139934
rect -8158 139698 30786 139934
rect 31022 139698 66786 139934
rect 67022 139698 102786 139934
rect 103022 139698 138786 139934
rect 139022 139698 174786 139934
rect 175022 139698 210786 139934
rect 211022 139698 246786 139934
rect 247022 139698 282786 139934
rect 283022 139698 318786 139934
rect 319022 139698 354786 139934
rect 355022 139698 390786 139934
rect 391022 139698 426786 139934
rect 427022 139698 462786 139934
rect 463022 139698 498786 139934
rect 499022 139698 534786 139934
rect 535022 139698 570786 139934
rect 571022 139698 592082 139934
rect 592318 139698 592500 139934
rect -8576 139676 592500 139698
rect -8576 139674 -7976 139676
rect 30604 139674 31204 139676
rect 66604 139674 67204 139676
rect 102604 139674 103204 139676
rect 138604 139674 139204 139676
rect 174604 139674 175204 139676
rect 210604 139674 211204 139676
rect 246604 139674 247204 139676
rect 282604 139674 283204 139676
rect 318604 139674 319204 139676
rect 354604 139674 355204 139676
rect 390604 139674 391204 139676
rect 426604 139674 427204 139676
rect 462604 139674 463204 139676
rect 498604 139674 499204 139676
rect 534604 139674 535204 139676
rect 570604 139674 571204 139676
rect 591900 139674 592500 139676
rect -6696 136676 -6096 136678
rect 27004 136676 27604 136678
rect 63004 136676 63604 136678
rect 99004 136676 99604 136678
rect 135004 136676 135604 136678
rect 171004 136676 171604 136678
rect 207004 136676 207604 136678
rect 243004 136676 243604 136678
rect 279004 136676 279604 136678
rect 315004 136676 315604 136678
rect 351004 136676 351604 136678
rect 387004 136676 387604 136678
rect 423004 136676 423604 136678
rect 459004 136676 459604 136678
rect 495004 136676 495604 136678
rect 531004 136676 531604 136678
rect 567004 136676 567604 136678
rect 590020 136676 590620 136678
rect -6696 136654 590620 136676
rect -6696 136418 -6514 136654
rect -6278 136418 27186 136654
rect 27422 136418 63186 136654
rect 63422 136418 99186 136654
rect 99422 136418 135186 136654
rect 135422 136418 171186 136654
rect 171422 136418 207186 136654
rect 207422 136418 243186 136654
rect 243422 136418 279186 136654
rect 279422 136418 315186 136654
rect 315422 136418 351186 136654
rect 351422 136418 387186 136654
rect 387422 136418 423186 136654
rect 423422 136418 459186 136654
rect 459422 136418 495186 136654
rect 495422 136418 531186 136654
rect 531422 136418 567186 136654
rect 567422 136418 590202 136654
rect 590438 136418 590620 136654
rect -6696 136334 590620 136418
rect -6696 136098 -6514 136334
rect -6278 136098 27186 136334
rect 27422 136098 63186 136334
rect 63422 136098 99186 136334
rect 99422 136098 135186 136334
rect 135422 136098 171186 136334
rect 171422 136098 207186 136334
rect 207422 136098 243186 136334
rect 243422 136098 279186 136334
rect 279422 136098 315186 136334
rect 315422 136098 351186 136334
rect 351422 136098 387186 136334
rect 387422 136098 423186 136334
rect 423422 136098 459186 136334
rect 459422 136098 495186 136334
rect 495422 136098 531186 136334
rect 531422 136098 567186 136334
rect 567422 136098 590202 136334
rect 590438 136098 590620 136334
rect -6696 136076 590620 136098
rect -6696 136074 -6096 136076
rect 27004 136074 27604 136076
rect 63004 136074 63604 136076
rect 99004 136074 99604 136076
rect 135004 136074 135604 136076
rect 171004 136074 171604 136076
rect 207004 136074 207604 136076
rect 243004 136074 243604 136076
rect 279004 136074 279604 136076
rect 315004 136074 315604 136076
rect 351004 136074 351604 136076
rect 387004 136074 387604 136076
rect 423004 136074 423604 136076
rect 459004 136074 459604 136076
rect 495004 136074 495604 136076
rect 531004 136074 531604 136076
rect 567004 136074 567604 136076
rect 590020 136074 590620 136076
rect -4816 133076 -4216 133078
rect 23404 133076 24004 133078
rect 59404 133076 60004 133078
rect 95404 133076 96004 133078
rect 131404 133076 132004 133078
rect 167404 133076 168004 133078
rect 203404 133076 204004 133078
rect 239404 133076 240004 133078
rect 275404 133076 276004 133078
rect 311404 133076 312004 133078
rect 347404 133076 348004 133078
rect 383404 133076 384004 133078
rect 419404 133076 420004 133078
rect 455404 133076 456004 133078
rect 491404 133076 492004 133078
rect 527404 133076 528004 133078
rect 563404 133076 564004 133078
rect 588140 133076 588740 133078
rect -4816 133054 588740 133076
rect -4816 132818 -4634 133054
rect -4398 132818 23586 133054
rect 23822 132818 59586 133054
rect 59822 132818 95586 133054
rect 95822 132818 131586 133054
rect 131822 132818 167586 133054
rect 167822 132818 203586 133054
rect 203822 132818 239586 133054
rect 239822 132818 275586 133054
rect 275822 132818 311586 133054
rect 311822 132818 347586 133054
rect 347822 132818 383586 133054
rect 383822 132818 419586 133054
rect 419822 132818 455586 133054
rect 455822 132818 491586 133054
rect 491822 132818 527586 133054
rect 527822 132818 563586 133054
rect 563822 132818 588322 133054
rect 588558 132818 588740 133054
rect -4816 132734 588740 132818
rect -4816 132498 -4634 132734
rect -4398 132498 23586 132734
rect 23822 132498 59586 132734
rect 59822 132498 95586 132734
rect 95822 132498 131586 132734
rect 131822 132498 167586 132734
rect 167822 132498 203586 132734
rect 203822 132498 239586 132734
rect 239822 132498 275586 132734
rect 275822 132498 311586 132734
rect 311822 132498 347586 132734
rect 347822 132498 383586 132734
rect 383822 132498 419586 132734
rect 419822 132498 455586 132734
rect 455822 132498 491586 132734
rect 491822 132498 527586 132734
rect 527822 132498 563586 132734
rect 563822 132498 588322 132734
rect 588558 132498 588740 132734
rect -4816 132476 588740 132498
rect -4816 132474 -4216 132476
rect 23404 132474 24004 132476
rect 59404 132474 60004 132476
rect 95404 132474 96004 132476
rect 131404 132474 132004 132476
rect 167404 132474 168004 132476
rect 203404 132474 204004 132476
rect 239404 132474 240004 132476
rect 275404 132474 276004 132476
rect 311404 132474 312004 132476
rect 347404 132474 348004 132476
rect 383404 132474 384004 132476
rect 419404 132474 420004 132476
rect 455404 132474 456004 132476
rect 491404 132474 492004 132476
rect 527404 132474 528004 132476
rect 563404 132474 564004 132476
rect 588140 132474 588740 132476
rect -2936 129476 -2336 129478
rect 19804 129476 20404 129478
rect 55804 129476 56404 129478
rect 91804 129476 92404 129478
rect 127804 129476 128404 129478
rect 163804 129476 164404 129478
rect 199804 129476 200404 129478
rect 235804 129476 236404 129478
rect 271804 129476 272404 129478
rect 307804 129476 308404 129478
rect 343804 129476 344404 129478
rect 379804 129476 380404 129478
rect 415804 129476 416404 129478
rect 451804 129476 452404 129478
rect 487804 129476 488404 129478
rect 523804 129476 524404 129478
rect 559804 129476 560404 129478
rect 586260 129476 586860 129478
rect -2936 129454 586860 129476
rect -2936 129218 -2754 129454
rect -2518 129218 19986 129454
rect 20222 129218 55986 129454
rect 56222 129218 91986 129454
rect 92222 129218 127986 129454
rect 128222 129218 163986 129454
rect 164222 129218 199986 129454
rect 200222 129218 235986 129454
rect 236222 129218 271986 129454
rect 272222 129218 307986 129454
rect 308222 129218 343986 129454
rect 344222 129218 379986 129454
rect 380222 129218 415986 129454
rect 416222 129218 451986 129454
rect 452222 129218 487986 129454
rect 488222 129218 523986 129454
rect 524222 129218 559986 129454
rect 560222 129218 586442 129454
rect 586678 129218 586860 129454
rect -2936 129134 586860 129218
rect -2936 128898 -2754 129134
rect -2518 128898 19986 129134
rect 20222 128898 55986 129134
rect 56222 128898 91986 129134
rect 92222 128898 127986 129134
rect 128222 128898 163986 129134
rect 164222 128898 199986 129134
rect 200222 128898 235986 129134
rect 236222 128898 271986 129134
rect 272222 128898 307986 129134
rect 308222 128898 343986 129134
rect 344222 128898 379986 129134
rect 380222 128898 415986 129134
rect 416222 128898 451986 129134
rect 452222 128898 487986 129134
rect 488222 128898 523986 129134
rect 524222 128898 559986 129134
rect 560222 128898 586442 129134
rect 586678 128898 586860 129134
rect -2936 128876 586860 128898
rect -2936 128874 -2336 128876
rect 19804 128874 20404 128876
rect 55804 128874 56404 128876
rect 91804 128874 92404 128876
rect 127804 128874 128404 128876
rect 163804 128874 164404 128876
rect 199804 128874 200404 128876
rect 235804 128874 236404 128876
rect 271804 128874 272404 128876
rect 307804 128874 308404 128876
rect 343804 128874 344404 128876
rect 379804 128874 380404 128876
rect 415804 128874 416404 128876
rect 451804 128874 452404 128876
rect 487804 128874 488404 128876
rect 523804 128874 524404 128876
rect 559804 128874 560404 128876
rect 586260 128874 586860 128876
rect -7636 122276 -7036 122278
rect 12604 122276 13204 122278
rect 48604 122276 49204 122278
rect 84604 122276 85204 122278
rect 120604 122276 121204 122278
rect 156604 122276 157204 122278
rect 192604 122276 193204 122278
rect 228604 122276 229204 122278
rect 264604 122276 265204 122278
rect 300604 122276 301204 122278
rect 336604 122276 337204 122278
rect 372604 122276 373204 122278
rect 408604 122276 409204 122278
rect 444604 122276 445204 122278
rect 480604 122276 481204 122278
rect 516604 122276 517204 122278
rect 552604 122276 553204 122278
rect 590960 122276 591560 122278
rect -8576 122254 592500 122276
rect -8576 122018 -7454 122254
rect -7218 122018 12786 122254
rect 13022 122018 48786 122254
rect 49022 122018 84786 122254
rect 85022 122018 120786 122254
rect 121022 122018 156786 122254
rect 157022 122018 192786 122254
rect 193022 122018 228786 122254
rect 229022 122018 264786 122254
rect 265022 122018 300786 122254
rect 301022 122018 336786 122254
rect 337022 122018 372786 122254
rect 373022 122018 408786 122254
rect 409022 122018 444786 122254
rect 445022 122018 480786 122254
rect 481022 122018 516786 122254
rect 517022 122018 552786 122254
rect 553022 122018 591142 122254
rect 591378 122018 592500 122254
rect -8576 121934 592500 122018
rect -8576 121698 -7454 121934
rect -7218 121698 12786 121934
rect 13022 121698 48786 121934
rect 49022 121698 84786 121934
rect 85022 121698 120786 121934
rect 121022 121698 156786 121934
rect 157022 121698 192786 121934
rect 193022 121698 228786 121934
rect 229022 121698 264786 121934
rect 265022 121698 300786 121934
rect 301022 121698 336786 121934
rect 337022 121698 372786 121934
rect 373022 121698 408786 121934
rect 409022 121698 444786 121934
rect 445022 121698 480786 121934
rect 481022 121698 516786 121934
rect 517022 121698 552786 121934
rect 553022 121698 591142 121934
rect 591378 121698 592500 121934
rect -8576 121676 592500 121698
rect -7636 121674 -7036 121676
rect 12604 121674 13204 121676
rect 48604 121674 49204 121676
rect 84604 121674 85204 121676
rect 120604 121674 121204 121676
rect 156604 121674 157204 121676
rect 192604 121674 193204 121676
rect 228604 121674 229204 121676
rect 264604 121674 265204 121676
rect 300604 121674 301204 121676
rect 336604 121674 337204 121676
rect 372604 121674 373204 121676
rect 408604 121674 409204 121676
rect 444604 121674 445204 121676
rect 480604 121674 481204 121676
rect 516604 121674 517204 121676
rect 552604 121674 553204 121676
rect 590960 121674 591560 121676
rect -5756 118676 -5156 118678
rect 9004 118676 9604 118678
rect 45004 118676 45604 118678
rect 81004 118676 81604 118678
rect 117004 118676 117604 118678
rect 153004 118676 153604 118678
rect 189004 118676 189604 118678
rect 225004 118676 225604 118678
rect 261004 118676 261604 118678
rect 297004 118676 297604 118678
rect 333004 118676 333604 118678
rect 369004 118676 369604 118678
rect 405004 118676 405604 118678
rect 441004 118676 441604 118678
rect 477004 118676 477604 118678
rect 513004 118676 513604 118678
rect 549004 118676 549604 118678
rect 589080 118676 589680 118678
rect -6696 118654 590620 118676
rect -6696 118418 -5574 118654
rect -5338 118418 9186 118654
rect 9422 118418 45186 118654
rect 45422 118418 81186 118654
rect 81422 118418 117186 118654
rect 117422 118418 153186 118654
rect 153422 118418 189186 118654
rect 189422 118418 225186 118654
rect 225422 118418 261186 118654
rect 261422 118418 297186 118654
rect 297422 118418 333186 118654
rect 333422 118418 369186 118654
rect 369422 118418 405186 118654
rect 405422 118418 441186 118654
rect 441422 118418 477186 118654
rect 477422 118418 513186 118654
rect 513422 118418 549186 118654
rect 549422 118418 589262 118654
rect 589498 118418 590620 118654
rect -6696 118334 590620 118418
rect -6696 118098 -5574 118334
rect -5338 118098 9186 118334
rect 9422 118098 45186 118334
rect 45422 118098 81186 118334
rect 81422 118098 117186 118334
rect 117422 118098 153186 118334
rect 153422 118098 189186 118334
rect 189422 118098 225186 118334
rect 225422 118098 261186 118334
rect 261422 118098 297186 118334
rect 297422 118098 333186 118334
rect 333422 118098 369186 118334
rect 369422 118098 405186 118334
rect 405422 118098 441186 118334
rect 441422 118098 477186 118334
rect 477422 118098 513186 118334
rect 513422 118098 549186 118334
rect 549422 118098 589262 118334
rect 589498 118098 590620 118334
rect -6696 118076 590620 118098
rect -5756 118074 -5156 118076
rect 9004 118074 9604 118076
rect 45004 118074 45604 118076
rect 81004 118074 81604 118076
rect 117004 118074 117604 118076
rect 153004 118074 153604 118076
rect 189004 118074 189604 118076
rect 225004 118074 225604 118076
rect 261004 118074 261604 118076
rect 297004 118074 297604 118076
rect 333004 118074 333604 118076
rect 369004 118074 369604 118076
rect 405004 118074 405604 118076
rect 441004 118074 441604 118076
rect 477004 118074 477604 118076
rect 513004 118074 513604 118076
rect 549004 118074 549604 118076
rect 589080 118074 589680 118076
rect -3876 115076 -3276 115078
rect 5404 115076 6004 115078
rect 41404 115076 42004 115078
rect 77404 115076 78004 115078
rect 113404 115076 114004 115078
rect 149404 115076 150004 115078
rect 185404 115076 186004 115078
rect 221404 115076 222004 115078
rect 257404 115076 258004 115078
rect 293404 115076 294004 115078
rect 329404 115076 330004 115078
rect 365404 115076 366004 115078
rect 401404 115076 402004 115078
rect 437404 115076 438004 115078
rect 473404 115076 474004 115078
rect 509404 115076 510004 115078
rect 545404 115076 546004 115078
rect 581404 115076 582004 115078
rect 587200 115076 587800 115078
rect -4816 115054 588740 115076
rect -4816 114818 -3694 115054
rect -3458 114818 5586 115054
rect 5822 114818 41586 115054
rect 41822 114818 77586 115054
rect 77822 114818 113586 115054
rect 113822 114818 149586 115054
rect 149822 114818 185586 115054
rect 185822 114818 221586 115054
rect 221822 114818 257586 115054
rect 257822 114818 293586 115054
rect 293822 114818 329586 115054
rect 329822 114818 365586 115054
rect 365822 114818 401586 115054
rect 401822 114818 437586 115054
rect 437822 114818 473586 115054
rect 473822 114818 509586 115054
rect 509822 114818 545586 115054
rect 545822 114818 581586 115054
rect 581822 114818 587382 115054
rect 587618 114818 588740 115054
rect -4816 114734 588740 114818
rect -4816 114498 -3694 114734
rect -3458 114498 5586 114734
rect 5822 114498 41586 114734
rect 41822 114498 77586 114734
rect 77822 114498 113586 114734
rect 113822 114498 149586 114734
rect 149822 114498 185586 114734
rect 185822 114498 221586 114734
rect 221822 114498 257586 114734
rect 257822 114498 293586 114734
rect 293822 114498 329586 114734
rect 329822 114498 365586 114734
rect 365822 114498 401586 114734
rect 401822 114498 437586 114734
rect 437822 114498 473586 114734
rect 473822 114498 509586 114734
rect 509822 114498 545586 114734
rect 545822 114498 581586 114734
rect 581822 114498 587382 114734
rect 587618 114498 588740 114734
rect -4816 114476 588740 114498
rect -3876 114474 -3276 114476
rect 5404 114474 6004 114476
rect 41404 114474 42004 114476
rect 77404 114474 78004 114476
rect 113404 114474 114004 114476
rect 149404 114474 150004 114476
rect 185404 114474 186004 114476
rect 221404 114474 222004 114476
rect 257404 114474 258004 114476
rect 293404 114474 294004 114476
rect 329404 114474 330004 114476
rect 365404 114474 366004 114476
rect 401404 114474 402004 114476
rect 437404 114474 438004 114476
rect 473404 114474 474004 114476
rect 509404 114474 510004 114476
rect 545404 114474 546004 114476
rect 581404 114474 582004 114476
rect 587200 114474 587800 114476
rect -1996 111476 -1396 111478
rect 1804 111476 2404 111478
rect 37804 111476 38404 111478
rect 73804 111476 74404 111478
rect 109804 111476 110404 111478
rect 145804 111476 146404 111478
rect 181804 111476 182404 111478
rect 217804 111476 218404 111478
rect 253804 111476 254404 111478
rect 289804 111476 290404 111478
rect 325804 111476 326404 111478
rect 361804 111476 362404 111478
rect 397804 111476 398404 111478
rect 433804 111476 434404 111478
rect 469804 111476 470404 111478
rect 505804 111476 506404 111478
rect 541804 111476 542404 111478
rect 577804 111476 578404 111478
rect 585320 111476 585920 111478
rect -2936 111454 586860 111476
rect -2936 111218 -1814 111454
rect -1578 111218 1986 111454
rect 2222 111218 37986 111454
rect 38222 111218 73986 111454
rect 74222 111218 109986 111454
rect 110222 111218 145986 111454
rect 146222 111218 181986 111454
rect 182222 111218 217986 111454
rect 218222 111218 253986 111454
rect 254222 111218 289986 111454
rect 290222 111218 325986 111454
rect 326222 111218 361986 111454
rect 362222 111218 397986 111454
rect 398222 111218 433986 111454
rect 434222 111218 469986 111454
rect 470222 111218 505986 111454
rect 506222 111218 541986 111454
rect 542222 111218 577986 111454
rect 578222 111218 585502 111454
rect 585738 111218 586860 111454
rect -2936 111134 586860 111218
rect -2936 110898 -1814 111134
rect -1578 110898 1986 111134
rect 2222 110898 37986 111134
rect 38222 110898 73986 111134
rect 74222 110898 109986 111134
rect 110222 110898 145986 111134
rect 146222 110898 181986 111134
rect 182222 110898 217986 111134
rect 218222 110898 253986 111134
rect 254222 110898 289986 111134
rect 290222 110898 325986 111134
rect 326222 110898 361986 111134
rect 362222 110898 397986 111134
rect 398222 110898 433986 111134
rect 434222 110898 469986 111134
rect 470222 110898 505986 111134
rect 506222 110898 541986 111134
rect 542222 110898 577986 111134
rect 578222 110898 585502 111134
rect 585738 110898 586860 111134
rect -2936 110876 586860 110898
rect -1996 110874 -1396 110876
rect 1804 110874 2404 110876
rect 37804 110874 38404 110876
rect 73804 110874 74404 110876
rect 109804 110874 110404 110876
rect 145804 110874 146404 110876
rect 181804 110874 182404 110876
rect 217804 110874 218404 110876
rect 253804 110874 254404 110876
rect 289804 110874 290404 110876
rect 325804 110874 326404 110876
rect 361804 110874 362404 110876
rect 397804 110874 398404 110876
rect 433804 110874 434404 110876
rect 469804 110874 470404 110876
rect 505804 110874 506404 110876
rect 541804 110874 542404 110876
rect 577804 110874 578404 110876
rect 585320 110874 585920 110876
rect -8576 104276 -7976 104278
rect 30604 104276 31204 104278
rect 66604 104276 67204 104278
rect 102604 104276 103204 104278
rect 138604 104276 139204 104278
rect 174604 104276 175204 104278
rect 210604 104276 211204 104278
rect 246604 104276 247204 104278
rect 282604 104276 283204 104278
rect 318604 104276 319204 104278
rect 354604 104276 355204 104278
rect 390604 104276 391204 104278
rect 426604 104276 427204 104278
rect 462604 104276 463204 104278
rect 498604 104276 499204 104278
rect 534604 104276 535204 104278
rect 570604 104276 571204 104278
rect 591900 104276 592500 104278
rect -8576 104254 592500 104276
rect -8576 104018 -8394 104254
rect -8158 104018 30786 104254
rect 31022 104018 66786 104254
rect 67022 104018 102786 104254
rect 103022 104018 138786 104254
rect 139022 104018 174786 104254
rect 175022 104018 210786 104254
rect 211022 104018 246786 104254
rect 247022 104018 282786 104254
rect 283022 104018 318786 104254
rect 319022 104018 354786 104254
rect 355022 104018 390786 104254
rect 391022 104018 426786 104254
rect 427022 104018 462786 104254
rect 463022 104018 498786 104254
rect 499022 104018 534786 104254
rect 535022 104018 570786 104254
rect 571022 104018 592082 104254
rect 592318 104018 592500 104254
rect -8576 103934 592500 104018
rect -8576 103698 -8394 103934
rect -8158 103698 30786 103934
rect 31022 103698 66786 103934
rect 67022 103698 102786 103934
rect 103022 103698 138786 103934
rect 139022 103698 174786 103934
rect 175022 103698 210786 103934
rect 211022 103698 246786 103934
rect 247022 103698 282786 103934
rect 283022 103698 318786 103934
rect 319022 103698 354786 103934
rect 355022 103698 390786 103934
rect 391022 103698 426786 103934
rect 427022 103698 462786 103934
rect 463022 103698 498786 103934
rect 499022 103698 534786 103934
rect 535022 103698 570786 103934
rect 571022 103698 592082 103934
rect 592318 103698 592500 103934
rect -8576 103676 592500 103698
rect -8576 103674 -7976 103676
rect 30604 103674 31204 103676
rect 66604 103674 67204 103676
rect 102604 103674 103204 103676
rect 138604 103674 139204 103676
rect 174604 103674 175204 103676
rect 210604 103674 211204 103676
rect 246604 103674 247204 103676
rect 282604 103674 283204 103676
rect 318604 103674 319204 103676
rect 354604 103674 355204 103676
rect 390604 103674 391204 103676
rect 426604 103674 427204 103676
rect 462604 103674 463204 103676
rect 498604 103674 499204 103676
rect 534604 103674 535204 103676
rect 570604 103674 571204 103676
rect 591900 103674 592500 103676
rect -6696 100676 -6096 100678
rect 27004 100676 27604 100678
rect 63004 100676 63604 100678
rect 99004 100676 99604 100678
rect 135004 100676 135604 100678
rect 171004 100676 171604 100678
rect 207004 100676 207604 100678
rect 243004 100676 243604 100678
rect 279004 100676 279604 100678
rect 315004 100676 315604 100678
rect 351004 100676 351604 100678
rect 387004 100676 387604 100678
rect 423004 100676 423604 100678
rect 459004 100676 459604 100678
rect 495004 100676 495604 100678
rect 531004 100676 531604 100678
rect 567004 100676 567604 100678
rect 590020 100676 590620 100678
rect -6696 100654 590620 100676
rect -6696 100418 -6514 100654
rect -6278 100418 27186 100654
rect 27422 100418 63186 100654
rect 63422 100418 99186 100654
rect 99422 100418 135186 100654
rect 135422 100418 171186 100654
rect 171422 100418 207186 100654
rect 207422 100418 243186 100654
rect 243422 100418 279186 100654
rect 279422 100418 315186 100654
rect 315422 100418 351186 100654
rect 351422 100418 387186 100654
rect 387422 100418 423186 100654
rect 423422 100418 459186 100654
rect 459422 100418 495186 100654
rect 495422 100418 531186 100654
rect 531422 100418 567186 100654
rect 567422 100418 590202 100654
rect 590438 100418 590620 100654
rect -6696 100334 590620 100418
rect -6696 100098 -6514 100334
rect -6278 100098 27186 100334
rect 27422 100098 63186 100334
rect 63422 100098 99186 100334
rect 99422 100098 135186 100334
rect 135422 100098 171186 100334
rect 171422 100098 207186 100334
rect 207422 100098 243186 100334
rect 243422 100098 279186 100334
rect 279422 100098 315186 100334
rect 315422 100098 351186 100334
rect 351422 100098 387186 100334
rect 387422 100098 423186 100334
rect 423422 100098 459186 100334
rect 459422 100098 495186 100334
rect 495422 100098 531186 100334
rect 531422 100098 567186 100334
rect 567422 100098 590202 100334
rect 590438 100098 590620 100334
rect -6696 100076 590620 100098
rect -6696 100074 -6096 100076
rect 27004 100074 27604 100076
rect 63004 100074 63604 100076
rect 99004 100074 99604 100076
rect 135004 100074 135604 100076
rect 171004 100074 171604 100076
rect 207004 100074 207604 100076
rect 243004 100074 243604 100076
rect 279004 100074 279604 100076
rect 315004 100074 315604 100076
rect 351004 100074 351604 100076
rect 387004 100074 387604 100076
rect 423004 100074 423604 100076
rect 459004 100074 459604 100076
rect 495004 100074 495604 100076
rect 531004 100074 531604 100076
rect 567004 100074 567604 100076
rect 590020 100074 590620 100076
rect -4816 97076 -4216 97078
rect 23404 97076 24004 97078
rect 59404 97076 60004 97078
rect 95404 97076 96004 97078
rect 131404 97076 132004 97078
rect 167404 97076 168004 97078
rect 203404 97076 204004 97078
rect 239404 97076 240004 97078
rect 275404 97076 276004 97078
rect 311404 97076 312004 97078
rect 347404 97076 348004 97078
rect 383404 97076 384004 97078
rect 419404 97076 420004 97078
rect 455404 97076 456004 97078
rect 491404 97076 492004 97078
rect 527404 97076 528004 97078
rect 563404 97076 564004 97078
rect 588140 97076 588740 97078
rect -4816 97054 588740 97076
rect -4816 96818 -4634 97054
rect -4398 96818 23586 97054
rect 23822 96818 59586 97054
rect 59822 96818 95586 97054
rect 95822 96818 131586 97054
rect 131822 96818 167586 97054
rect 167822 96818 203586 97054
rect 203822 96818 239586 97054
rect 239822 96818 275586 97054
rect 275822 96818 311586 97054
rect 311822 96818 347586 97054
rect 347822 96818 383586 97054
rect 383822 96818 419586 97054
rect 419822 96818 455586 97054
rect 455822 96818 491586 97054
rect 491822 96818 527586 97054
rect 527822 96818 563586 97054
rect 563822 96818 588322 97054
rect 588558 96818 588740 97054
rect -4816 96734 588740 96818
rect -4816 96498 -4634 96734
rect -4398 96498 23586 96734
rect 23822 96498 59586 96734
rect 59822 96498 95586 96734
rect 95822 96498 131586 96734
rect 131822 96498 167586 96734
rect 167822 96498 203586 96734
rect 203822 96498 239586 96734
rect 239822 96498 275586 96734
rect 275822 96498 311586 96734
rect 311822 96498 347586 96734
rect 347822 96498 383586 96734
rect 383822 96498 419586 96734
rect 419822 96498 455586 96734
rect 455822 96498 491586 96734
rect 491822 96498 527586 96734
rect 527822 96498 563586 96734
rect 563822 96498 588322 96734
rect 588558 96498 588740 96734
rect -4816 96476 588740 96498
rect -4816 96474 -4216 96476
rect 23404 96474 24004 96476
rect 59404 96474 60004 96476
rect 95404 96474 96004 96476
rect 131404 96474 132004 96476
rect 167404 96474 168004 96476
rect 203404 96474 204004 96476
rect 239404 96474 240004 96476
rect 275404 96474 276004 96476
rect 311404 96474 312004 96476
rect 347404 96474 348004 96476
rect 383404 96474 384004 96476
rect 419404 96474 420004 96476
rect 455404 96474 456004 96476
rect 491404 96474 492004 96476
rect 527404 96474 528004 96476
rect 563404 96474 564004 96476
rect 588140 96474 588740 96476
rect -2936 93476 -2336 93478
rect 19804 93476 20404 93478
rect 55804 93476 56404 93478
rect 91804 93476 92404 93478
rect 127804 93476 128404 93478
rect 163804 93476 164404 93478
rect 199804 93476 200404 93478
rect 235804 93476 236404 93478
rect 271804 93476 272404 93478
rect 307804 93476 308404 93478
rect 343804 93476 344404 93478
rect 379804 93476 380404 93478
rect 415804 93476 416404 93478
rect 451804 93476 452404 93478
rect 487804 93476 488404 93478
rect 523804 93476 524404 93478
rect 559804 93476 560404 93478
rect 586260 93476 586860 93478
rect -2936 93454 586860 93476
rect -2936 93218 -2754 93454
rect -2518 93218 19986 93454
rect 20222 93218 55986 93454
rect 56222 93218 91986 93454
rect 92222 93218 127986 93454
rect 128222 93218 163986 93454
rect 164222 93218 199986 93454
rect 200222 93218 235986 93454
rect 236222 93218 271986 93454
rect 272222 93218 307986 93454
rect 308222 93218 343986 93454
rect 344222 93218 379986 93454
rect 380222 93218 415986 93454
rect 416222 93218 451986 93454
rect 452222 93218 487986 93454
rect 488222 93218 523986 93454
rect 524222 93218 559986 93454
rect 560222 93218 586442 93454
rect 586678 93218 586860 93454
rect -2936 93134 586860 93218
rect -2936 92898 -2754 93134
rect -2518 92898 19986 93134
rect 20222 92898 55986 93134
rect 56222 92898 91986 93134
rect 92222 92898 127986 93134
rect 128222 92898 163986 93134
rect 164222 92898 199986 93134
rect 200222 92898 235986 93134
rect 236222 92898 271986 93134
rect 272222 92898 307986 93134
rect 308222 92898 343986 93134
rect 344222 92898 379986 93134
rect 380222 92898 415986 93134
rect 416222 92898 451986 93134
rect 452222 92898 487986 93134
rect 488222 92898 523986 93134
rect 524222 92898 559986 93134
rect 560222 92898 586442 93134
rect 586678 92898 586860 93134
rect -2936 92876 586860 92898
rect -2936 92874 -2336 92876
rect 19804 92874 20404 92876
rect 55804 92874 56404 92876
rect 91804 92874 92404 92876
rect 127804 92874 128404 92876
rect 163804 92874 164404 92876
rect 199804 92874 200404 92876
rect 235804 92874 236404 92876
rect 271804 92874 272404 92876
rect 307804 92874 308404 92876
rect 343804 92874 344404 92876
rect 379804 92874 380404 92876
rect 415804 92874 416404 92876
rect 451804 92874 452404 92876
rect 487804 92874 488404 92876
rect 523804 92874 524404 92876
rect 559804 92874 560404 92876
rect 586260 92874 586860 92876
rect -7636 86276 -7036 86278
rect 12604 86276 13204 86278
rect 48604 86276 49204 86278
rect 84604 86276 85204 86278
rect 120604 86276 121204 86278
rect 156604 86276 157204 86278
rect 192604 86276 193204 86278
rect 228604 86276 229204 86278
rect 264604 86276 265204 86278
rect 300604 86276 301204 86278
rect 336604 86276 337204 86278
rect 372604 86276 373204 86278
rect 408604 86276 409204 86278
rect 444604 86276 445204 86278
rect 480604 86276 481204 86278
rect 516604 86276 517204 86278
rect 552604 86276 553204 86278
rect 590960 86276 591560 86278
rect -8576 86254 592500 86276
rect -8576 86018 -7454 86254
rect -7218 86018 12786 86254
rect 13022 86018 48786 86254
rect 49022 86018 84786 86254
rect 85022 86018 120786 86254
rect 121022 86018 156786 86254
rect 157022 86018 192786 86254
rect 193022 86018 228786 86254
rect 229022 86018 264786 86254
rect 265022 86018 300786 86254
rect 301022 86018 336786 86254
rect 337022 86018 372786 86254
rect 373022 86018 408786 86254
rect 409022 86018 444786 86254
rect 445022 86018 480786 86254
rect 481022 86018 516786 86254
rect 517022 86018 552786 86254
rect 553022 86018 591142 86254
rect 591378 86018 592500 86254
rect -8576 85934 592500 86018
rect -8576 85698 -7454 85934
rect -7218 85698 12786 85934
rect 13022 85698 48786 85934
rect 49022 85698 84786 85934
rect 85022 85698 120786 85934
rect 121022 85698 156786 85934
rect 157022 85698 192786 85934
rect 193022 85698 228786 85934
rect 229022 85698 264786 85934
rect 265022 85698 300786 85934
rect 301022 85698 336786 85934
rect 337022 85698 372786 85934
rect 373022 85698 408786 85934
rect 409022 85698 444786 85934
rect 445022 85698 480786 85934
rect 481022 85698 516786 85934
rect 517022 85698 552786 85934
rect 553022 85698 591142 85934
rect 591378 85698 592500 85934
rect -8576 85676 592500 85698
rect -7636 85674 -7036 85676
rect 12604 85674 13204 85676
rect 48604 85674 49204 85676
rect 84604 85674 85204 85676
rect 120604 85674 121204 85676
rect 156604 85674 157204 85676
rect 192604 85674 193204 85676
rect 228604 85674 229204 85676
rect 264604 85674 265204 85676
rect 300604 85674 301204 85676
rect 336604 85674 337204 85676
rect 372604 85674 373204 85676
rect 408604 85674 409204 85676
rect 444604 85674 445204 85676
rect 480604 85674 481204 85676
rect 516604 85674 517204 85676
rect 552604 85674 553204 85676
rect 590960 85674 591560 85676
rect -5756 82676 -5156 82678
rect 9004 82676 9604 82678
rect 45004 82676 45604 82678
rect 81004 82676 81604 82678
rect 117004 82676 117604 82678
rect 153004 82676 153604 82678
rect 189004 82676 189604 82678
rect 225004 82676 225604 82678
rect 261004 82676 261604 82678
rect 297004 82676 297604 82678
rect 333004 82676 333604 82678
rect 369004 82676 369604 82678
rect 405004 82676 405604 82678
rect 441004 82676 441604 82678
rect 477004 82676 477604 82678
rect 513004 82676 513604 82678
rect 549004 82676 549604 82678
rect 589080 82676 589680 82678
rect -6696 82654 590620 82676
rect -6696 82418 -5574 82654
rect -5338 82418 9186 82654
rect 9422 82418 45186 82654
rect 45422 82418 81186 82654
rect 81422 82418 117186 82654
rect 117422 82418 153186 82654
rect 153422 82418 189186 82654
rect 189422 82418 225186 82654
rect 225422 82418 261186 82654
rect 261422 82418 297186 82654
rect 297422 82418 333186 82654
rect 333422 82418 369186 82654
rect 369422 82418 405186 82654
rect 405422 82418 441186 82654
rect 441422 82418 477186 82654
rect 477422 82418 513186 82654
rect 513422 82418 549186 82654
rect 549422 82418 589262 82654
rect 589498 82418 590620 82654
rect -6696 82334 590620 82418
rect -6696 82098 -5574 82334
rect -5338 82098 9186 82334
rect 9422 82098 45186 82334
rect 45422 82098 81186 82334
rect 81422 82098 117186 82334
rect 117422 82098 153186 82334
rect 153422 82098 189186 82334
rect 189422 82098 225186 82334
rect 225422 82098 261186 82334
rect 261422 82098 297186 82334
rect 297422 82098 333186 82334
rect 333422 82098 369186 82334
rect 369422 82098 405186 82334
rect 405422 82098 441186 82334
rect 441422 82098 477186 82334
rect 477422 82098 513186 82334
rect 513422 82098 549186 82334
rect 549422 82098 589262 82334
rect 589498 82098 590620 82334
rect -6696 82076 590620 82098
rect -5756 82074 -5156 82076
rect 9004 82074 9604 82076
rect 45004 82074 45604 82076
rect 81004 82074 81604 82076
rect 117004 82074 117604 82076
rect 153004 82074 153604 82076
rect 189004 82074 189604 82076
rect 225004 82074 225604 82076
rect 261004 82074 261604 82076
rect 297004 82074 297604 82076
rect 333004 82074 333604 82076
rect 369004 82074 369604 82076
rect 405004 82074 405604 82076
rect 441004 82074 441604 82076
rect 477004 82074 477604 82076
rect 513004 82074 513604 82076
rect 549004 82074 549604 82076
rect 589080 82074 589680 82076
rect -3876 79076 -3276 79078
rect 5404 79076 6004 79078
rect 41404 79076 42004 79078
rect 77404 79076 78004 79078
rect 113404 79076 114004 79078
rect 149404 79076 150004 79078
rect 185404 79076 186004 79078
rect 221404 79076 222004 79078
rect 257404 79076 258004 79078
rect 293404 79076 294004 79078
rect 329404 79076 330004 79078
rect 365404 79076 366004 79078
rect 401404 79076 402004 79078
rect 437404 79076 438004 79078
rect 473404 79076 474004 79078
rect 509404 79076 510004 79078
rect 545404 79076 546004 79078
rect 581404 79076 582004 79078
rect 587200 79076 587800 79078
rect -4816 79054 588740 79076
rect -4816 78818 -3694 79054
rect -3458 78818 5586 79054
rect 5822 78818 41586 79054
rect 41822 78818 77586 79054
rect 77822 78818 113586 79054
rect 113822 78818 149586 79054
rect 149822 78818 185586 79054
rect 185822 78818 221586 79054
rect 221822 78818 257586 79054
rect 257822 78818 293586 79054
rect 293822 78818 329586 79054
rect 329822 78818 365586 79054
rect 365822 78818 401586 79054
rect 401822 78818 437586 79054
rect 437822 78818 473586 79054
rect 473822 78818 509586 79054
rect 509822 78818 545586 79054
rect 545822 78818 581586 79054
rect 581822 78818 587382 79054
rect 587618 78818 588740 79054
rect -4816 78734 588740 78818
rect -4816 78498 -3694 78734
rect -3458 78498 5586 78734
rect 5822 78498 41586 78734
rect 41822 78498 77586 78734
rect 77822 78498 113586 78734
rect 113822 78498 149586 78734
rect 149822 78498 185586 78734
rect 185822 78498 221586 78734
rect 221822 78498 257586 78734
rect 257822 78498 293586 78734
rect 293822 78498 329586 78734
rect 329822 78498 365586 78734
rect 365822 78498 401586 78734
rect 401822 78498 437586 78734
rect 437822 78498 473586 78734
rect 473822 78498 509586 78734
rect 509822 78498 545586 78734
rect 545822 78498 581586 78734
rect 581822 78498 587382 78734
rect 587618 78498 588740 78734
rect -4816 78476 588740 78498
rect -3876 78474 -3276 78476
rect 5404 78474 6004 78476
rect 41404 78474 42004 78476
rect 77404 78474 78004 78476
rect 113404 78474 114004 78476
rect 149404 78474 150004 78476
rect 185404 78474 186004 78476
rect 221404 78474 222004 78476
rect 257404 78474 258004 78476
rect 293404 78474 294004 78476
rect 329404 78474 330004 78476
rect 365404 78474 366004 78476
rect 401404 78474 402004 78476
rect 437404 78474 438004 78476
rect 473404 78474 474004 78476
rect 509404 78474 510004 78476
rect 545404 78474 546004 78476
rect 581404 78474 582004 78476
rect 587200 78474 587800 78476
rect -1996 75476 -1396 75478
rect 1804 75476 2404 75478
rect 37804 75476 38404 75478
rect 73804 75476 74404 75478
rect 109804 75476 110404 75478
rect 145804 75476 146404 75478
rect 181804 75476 182404 75478
rect 217804 75476 218404 75478
rect 253804 75476 254404 75478
rect 289804 75476 290404 75478
rect 325804 75476 326404 75478
rect 361804 75476 362404 75478
rect 397804 75476 398404 75478
rect 433804 75476 434404 75478
rect 469804 75476 470404 75478
rect 505804 75476 506404 75478
rect 541804 75476 542404 75478
rect 577804 75476 578404 75478
rect 585320 75476 585920 75478
rect -2936 75454 586860 75476
rect -2936 75218 -1814 75454
rect -1578 75218 1986 75454
rect 2222 75218 37986 75454
rect 38222 75218 73986 75454
rect 74222 75218 109986 75454
rect 110222 75218 145986 75454
rect 146222 75218 181986 75454
rect 182222 75218 217986 75454
rect 218222 75218 253986 75454
rect 254222 75218 289986 75454
rect 290222 75218 325986 75454
rect 326222 75218 361986 75454
rect 362222 75218 397986 75454
rect 398222 75218 433986 75454
rect 434222 75218 469986 75454
rect 470222 75218 505986 75454
rect 506222 75218 541986 75454
rect 542222 75218 577986 75454
rect 578222 75218 585502 75454
rect 585738 75218 586860 75454
rect -2936 75134 586860 75218
rect -2936 74898 -1814 75134
rect -1578 74898 1986 75134
rect 2222 74898 37986 75134
rect 38222 74898 73986 75134
rect 74222 74898 109986 75134
rect 110222 74898 145986 75134
rect 146222 74898 181986 75134
rect 182222 74898 217986 75134
rect 218222 74898 253986 75134
rect 254222 74898 289986 75134
rect 290222 74898 325986 75134
rect 326222 74898 361986 75134
rect 362222 74898 397986 75134
rect 398222 74898 433986 75134
rect 434222 74898 469986 75134
rect 470222 74898 505986 75134
rect 506222 74898 541986 75134
rect 542222 74898 577986 75134
rect 578222 74898 585502 75134
rect 585738 74898 586860 75134
rect -2936 74876 586860 74898
rect -1996 74874 -1396 74876
rect 1804 74874 2404 74876
rect 37804 74874 38404 74876
rect 73804 74874 74404 74876
rect 109804 74874 110404 74876
rect 145804 74874 146404 74876
rect 181804 74874 182404 74876
rect 217804 74874 218404 74876
rect 253804 74874 254404 74876
rect 289804 74874 290404 74876
rect 325804 74874 326404 74876
rect 361804 74874 362404 74876
rect 397804 74874 398404 74876
rect 433804 74874 434404 74876
rect 469804 74874 470404 74876
rect 505804 74874 506404 74876
rect 541804 74874 542404 74876
rect 577804 74874 578404 74876
rect 585320 74874 585920 74876
rect -8576 68276 -7976 68278
rect 30604 68276 31204 68278
rect 66604 68276 67204 68278
rect 102604 68276 103204 68278
rect 138604 68276 139204 68278
rect 174604 68276 175204 68278
rect 210604 68276 211204 68278
rect 246604 68276 247204 68278
rect 282604 68276 283204 68278
rect 318604 68276 319204 68278
rect 354604 68276 355204 68278
rect 390604 68276 391204 68278
rect 426604 68276 427204 68278
rect 462604 68276 463204 68278
rect 498604 68276 499204 68278
rect 534604 68276 535204 68278
rect 570604 68276 571204 68278
rect 591900 68276 592500 68278
rect -8576 68254 592500 68276
rect -8576 68018 -8394 68254
rect -8158 68018 30786 68254
rect 31022 68018 66786 68254
rect 67022 68018 102786 68254
rect 103022 68018 138786 68254
rect 139022 68018 174786 68254
rect 175022 68018 210786 68254
rect 211022 68018 246786 68254
rect 247022 68018 282786 68254
rect 283022 68018 318786 68254
rect 319022 68018 354786 68254
rect 355022 68018 390786 68254
rect 391022 68018 426786 68254
rect 427022 68018 462786 68254
rect 463022 68018 498786 68254
rect 499022 68018 534786 68254
rect 535022 68018 570786 68254
rect 571022 68018 592082 68254
rect 592318 68018 592500 68254
rect -8576 67934 592500 68018
rect -8576 67698 -8394 67934
rect -8158 67698 30786 67934
rect 31022 67698 66786 67934
rect 67022 67698 102786 67934
rect 103022 67698 138786 67934
rect 139022 67698 174786 67934
rect 175022 67698 210786 67934
rect 211022 67698 246786 67934
rect 247022 67698 282786 67934
rect 283022 67698 318786 67934
rect 319022 67698 354786 67934
rect 355022 67698 390786 67934
rect 391022 67698 426786 67934
rect 427022 67698 462786 67934
rect 463022 67698 498786 67934
rect 499022 67698 534786 67934
rect 535022 67698 570786 67934
rect 571022 67698 592082 67934
rect 592318 67698 592500 67934
rect -8576 67676 592500 67698
rect -8576 67674 -7976 67676
rect 30604 67674 31204 67676
rect 66604 67674 67204 67676
rect 102604 67674 103204 67676
rect 138604 67674 139204 67676
rect 174604 67674 175204 67676
rect 210604 67674 211204 67676
rect 246604 67674 247204 67676
rect 282604 67674 283204 67676
rect 318604 67674 319204 67676
rect 354604 67674 355204 67676
rect 390604 67674 391204 67676
rect 426604 67674 427204 67676
rect 462604 67674 463204 67676
rect 498604 67674 499204 67676
rect 534604 67674 535204 67676
rect 570604 67674 571204 67676
rect 591900 67674 592500 67676
rect -6696 64676 -6096 64678
rect 27004 64676 27604 64678
rect 63004 64676 63604 64678
rect 99004 64676 99604 64678
rect 135004 64676 135604 64678
rect 171004 64676 171604 64678
rect 207004 64676 207604 64678
rect 243004 64676 243604 64678
rect 279004 64676 279604 64678
rect 315004 64676 315604 64678
rect 351004 64676 351604 64678
rect 387004 64676 387604 64678
rect 423004 64676 423604 64678
rect 459004 64676 459604 64678
rect 495004 64676 495604 64678
rect 531004 64676 531604 64678
rect 567004 64676 567604 64678
rect 590020 64676 590620 64678
rect -6696 64654 590620 64676
rect -6696 64418 -6514 64654
rect -6278 64418 27186 64654
rect 27422 64418 63186 64654
rect 63422 64418 99186 64654
rect 99422 64418 135186 64654
rect 135422 64418 171186 64654
rect 171422 64418 207186 64654
rect 207422 64418 243186 64654
rect 243422 64418 279186 64654
rect 279422 64418 315186 64654
rect 315422 64418 351186 64654
rect 351422 64418 387186 64654
rect 387422 64418 423186 64654
rect 423422 64418 459186 64654
rect 459422 64418 495186 64654
rect 495422 64418 531186 64654
rect 531422 64418 567186 64654
rect 567422 64418 590202 64654
rect 590438 64418 590620 64654
rect -6696 64334 590620 64418
rect -6696 64098 -6514 64334
rect -6278 64098 27186 64334
rect 27422 64098 63186 64334
rect 63422 64098 99186 64334
rect 99422 64098 135186 64334
rect 135422 64098 171186 64334
rect 171422 64098 207186 64334
rect 207422 64098 243186 64334
rect 243422 64098 279186 64334
rect 279422 64098 315186 64334
rect 315422 64098 351186 64334
rect 351422 64098 387186 64334
rect 387422 64098 423186 64334
rect 423422 64098 459186 64334
rect 459422 64098 495186 64334
rect 495422 64098 531186 64334
rect 531422 64098 567186 64334
rect 567422 64098 590202 64334
rect 590438 64098 590620 64334
rect -6696 64076 590620 64098
rect -6696 64074 -6096 64076
rect 27004 64074 27604 64076
rect 63004 64074 63604 64076
rect 99004 64074 99604 64076
rect 135004 64074 135604 64076
rect 171004 64074 171604 64076
rect 207004 64074 207604 64076
rect 243004 64074 243604 64076
rect 279004 64074 279604 64076
rect 315004 64074 315604 64076
rect 351004 64074 351604 64076
rect 387004 64074 387604 64076
rect 423004 64074 423604 64076
rect 459004 64074 459604 64076
rect 495004 64074 495604 64076
rect 531004 64074 531604 64076
rect 567004 64074 567604 64076
rect 590020 64074 590620 64076
rect -4816 61076 -4216 61078
rect 23404 61076 24004 61078
rect 59404 61076 60004 61078
rect 95404 61076 96004 61078
rect 131404 61076 132004 61078
rect 167404 61076 168004 61078
rect 203404 61076 204004 61078
rect 239404 61076 240004 61078
rect 275404 61076 276004 61078
rect 311404 61076 312004 61078
rect 347404 61076 348004 61078
rect 383404 61076 384004 61078
rect 419404 61076 420004 61078
rect 455404 61076 456004 61078
rect 491404 61076 492004 61078
rect 527404 61076 528004 61078
rect 563404 61076 564004 61078
rect 588140 61076 588740 61078
rect -4816 61054 588740 61076
rect -4816 60818 -4634 61054
rect -4398 60818 23586 61054
rect 23822 60818 59586 61054
rect 59822 60818 95586 61054
rect 95822 60818 131586 61054
rect 131822 60818 167586 61054
rect 167822 60818 203586 61054
rect 203822 60818 239586 61054
rect 239822 60818 275586 61054
rect 275822 60818 311586 61054
rect 311822 60818 347586 61054
rect 347822 60818 383586 61054
rect 383822 60818 419586 61054
rect 419822 60818 455586 61054
rect 455822 60818 491586 61054
rect 491822 60818 527586 61054
rect 527822 60818 563586 61054
rect 563822 60818 588322 61054
rect 588558 60818 588740 61054
rect -4816 60734 588740 60818
rect -4816 60498 -4634 60734
rect -4398 60498 23586 60734
rect 23822 60498 59586 60734
rect 59822 60498 95586 60734
rect 95822 60498 131586 60734
rect 131822 60498 167586 60734
rect 167822 60498 203586 60734
rect 203822 60498 239586 60734
rect 239822 60498 275586 60734
rect 275822 60498 311586 60734
rect 311822 60498 347586 60734
rect 347822 60498 383586 60734
rect 383822 60498 419586 60734
rect 419822 60498 455586 60734
rect 455822 60498 491586 60734
rect 491822 60498 527586 60734
rect 527822 60498 563586 60734
rect 563822 60498 588322 60734
rect 588558 60498 588740 60734
rect -4816 60476 588740 60498
rect -4816 60474 -4216 60476
rect 23404 60474 24004 60476
rect 59404 60474 60004 60476
rect 95404 60474 96004 60476
rect 131404 60474 132004 60476
rect 167404 60474 168004 60476
rect 203404 60474 204004 60476
rect 239404 60474 240004 60476
rect 275404 60474 276004 60476
rect 311404 60474 312004 60476
rect 347404 60474 348004 60476
rect 383404 60474 384004 60476
rect 419404 60474 420004 60476
rect 455404 60474 456004 60476
rect 491404 60474 492004 60476
rect 527404 60474 528004 60476
rect 563404 60474 564004 60476
rect 588140 60474 588740 60476
rect -2936 57476 -2336 57478
rect 19804 57476 20404 57478
rect 55804 57476 56404 57478
rect 91804 57476 92404 57478
rect 127804 57476 128404 57478
rect 163804 57476 164404 57478
rect 199804 57476 200404 57478
rect 235804 57476 236404 57478
rect 271804 57476 272404 57478
rect 307804 57476 308404 57478
rect 343804 57476 344404 57478
rect 379804 57476 380404 57478
rect 415804 57476 416404 57478
rect 451804 57476 452404 57478
rect 487804 57476 488404 57478
rect 523804 57476 524404 57478
rect 559804 57476 560404 57478
rect 586260 57476 586860 57478
rect -2936 57454 586860 57476
rect -2936 57218 -2754 57454
rect -2518 57218 19986 57454
rect 20222 57218 55986 57454
rect 56222 57218 91986 57454
rect 92222 57218 127986 57454
rect 128222 57218 163986 57454
rect 164222 57218 199986 57454
rect 200222 57218 235986 57454
rect 236222 57218 271986 57454
rect 272222 57218 307986 57454
rect 308222 57218 343986 57454
rect 344222 57218 379986 57454
rect 380222 57218 415986 57454
rect 416222 57218 451986 57454
rect 452222 57218 487986 57454
rect 488222 57218 523986 57454
rect 524222 57218 559986 57454
rect 560222 57218 586442 57454
rect 586678 57218 586860 57454
rect -2936 57134 586860 57218
rect -2936 56898 -2754 57134
rect -2518 56898 19986 57134
rect 20222 56898 55986 57134
rect 56222 56898 91986 57134
rect 92222 56898 127986 57134
rect 128222 56898 163986 57134
rect 164222 56898 199986 57134
rect 200222 56898 235986 57134
rect 236222 56898 271986 57134
rect 272222 56898 307986 57134
rect 308222 56898 343986 57134
rect 344222 56898 379986 57134
rect 380222 56898 415986 57134
rect 416222 56898 451986 57134
rect 452222 56898 487986 57134
rect 488222 56898 523986 57134
rect 524222 56898 559986 57134
rect 560222 56898 586442 57134
rect 586678 56898 586860 57134
rect -2936 56876 586860 56898
rect -2936 56874 -2336 56876
rect 19804 56874 20404 56876
rect 55804 56874 56404 56876
rect 91804 56874 92404 56876
rect 127804 56874 128404 56876
rect 163804 56874 164404 56876
rect 199804 56874 200404 56876
rect 235804 56874 236404 56876
rect 271804 56874 272404 56876
rect 307804 56874 308404 56876
rect 343804 56874 344404 56876
rect 379804 56874 380404 56876
rect 415804 56874 416404 56876
rect 451804 56874 452404 56876
rect 487804 56874 488404 56876
rect 523804 56874 524404 56876
rect 559804 56874 560404 56876
rect 586260 56874 586860 56876
rect -7636 50276 -7036 50278
rect 12604 50276 13204 50278
rect 48604 50276 49204 50278
rect 84604 50276 85204 50278
rect 120604 50276 121204 50278
rect 156604 50276 157204 50278
rect 192604 50276 193204 50278
rect 228604 50276 229204 50278
rect 264604 50276 265204 50278
rect 300604 50276 301204 50278
rect 336604 50276 337204 50278
rect 372604 50276 373204 50278
rect 408604 50276 409204 50278
rect 444604 50276 445204 50278
rect 480604 50276 481204 50278
rect 516604 50276 517204 50278
rect 552604 50276 553204 50278
rect 590960 50276 591560 50278
rect -8576 50254 592500 50276
rect -8576 50018 -7454 50254
rect -7218 50018 12786 50254
rect 13022 50018 48786 50254
rect 49022 50018 84786 50254
rect 85022 50018 120786 50254
rect 121022 50018 156786 50254
rect 157022 50018 192786 50254
rect 193022 50018 228786 50254
rect 229022 50018 264786 50254
rect 265022 50018 300786 50254
rect 301022 50018 336786 50254
rect 337022 50018 372786 50254
rect 373022 50018 408786 50254
rect 409022 50018 444786 50254
rect 445022 50018 480786 50254
rect 481022 50018 516786 50254
rect 517022 50018 552786 50254
rect 553022 50018 591142 50254
rect 591378 50018 592500 50254
rect -8576 49934 592500 50018
rect -8576 49698 -7454 49934
rect -7218 49698 12786 49934
rect 13022 49698 48786 49934
rect 49022 49698 84786 49934
rect 85022 49698 120786 49934
rect 121022 49698 156786 49934
rect 157022 49698 192786 49934
rect 193022 49698 228786 49934
rect 229022 49698 264786 49934
rect 265022 49698 300786 49934
rect 301022 49698 336786 49934
rect 337022 49698 372786 49934
rect 373022 49698 408786 49934
rect 409022 49698 444786 49934
rect 445022 49698 480786 49934
rect 481022 49698 516786 49934
rect 517022 49698 552786 49934
rect 553022 49698 591142 49934
rect 591378 49698 592500 49934
rect -8576 49676 592500 49698
rect -7636 49674 -7036 49676
rect 12604 49674 13204 49676
rect 48604 49674 49204 49676
rect 84604 49674 85204 49676
rect 120604 49674 121204 49676
rect 156604 49674 157204 49676
rect 192604 49674 193204 49676
rect 228604 49674 229204 49676
rect 264604 49674 265204 49676
rect 300604 49674 301204 49676
rect 336604 49674 337204 49676
rect 372604 49674 373204 49676
rect 408604 49674 409204 49676
rect 444604 49674 445204 49676
rect 480604 49674 481204 49676
rect 516604 49674 517204 49676
rect 552604 49674 553204 49676
rect 590960 49674 591560 49676
rect -5756 46676 -5156 46678
rect 9004 46676 9604 46678
rect 45004 46676 45604 46678
rect 81004 46676 81604 46678
rect 117004 46676 117604 46678
rect 153004 46676 153604 46678
rect 189004 46676 189604 46678
rect 225004 46676 225604 46678
rect 261004 46676 261604 46678
rect 297004 46676 297604 46678
rect 333004 46676 333604 46678
rect 369004 46676 369604 46678
rect 405004 46676 405604 46678
rect 441004 46676 441604 46678
rect 477004 46676 477604 46678
rect 513004 46676 513604 46678
rect 549004 46676 549604 46678
rect 589080 46676 589680 46678
rect -6696 46654 590620 46676
rect -6696 46418 -5574 46654
rect -5338 46418 9186 46654
rect 9422 46418 45186 46654
rect 45422 46418 81186 46654
rect 81422 46418 117186 46654
rect 117422 46418 153186 46654
rect 153422 46418 189186 46654
rect 189422 46418 225186 46654
rect 225422 46418 261186 46654
rect 261422 46418 297186 46654
rect 297422 46418 333186 46654
rect 333422 46418 369186 46654
rect 369422 46418 405186 46654
rect 405422 46418 441186 46654
rect 441422 46418 477186 46654
rect 477422 46418 513186 46654
rect 513422 46418 549186 46654
rect 549422 46418 589262 46654
rect 589498 46418 590620 46654
rect -6696 46334 590620 46418
rect -6696 46098 -5574 46334
rect -5338 46098 9186 46334
rect 9422 46098 45186 46334
rect 45422 46098 81186 46334
rect 81422 46098 117186 46334
rect 117422 46098 153186 46334
rect 153422 46098 189186 46334
rect 189422 46098 225186 46334
rect 225422 46098 261186 46334
rect 261422 46098 297186 46334
rect 297422 46098 333186 46334
rect 333422 46098 369186 46334
rect 369422 46098 405186 46334
rect 405422 46098 441186 46334
rect 441422 46098 477186 46334
rect 477422 46098 513186 46334
rect 513422 46098 549186 46334
rect 549422 46098 589262 46334
rect 589498 46098 590620 46334
rect -6696 46076 590620 46098
rect -5756 46074 -5156 46076
rect 9004 46074 9604 46076
rect 45004 46074 45604 46076
rect 81004 46074 81604 46076
rect 117004 46074 117604 46076
rect 153004 46074 153604 46076
rect 189004 46074 189604 46076
rect 225004 46074 225604 46076
rect 261004 46074 261604 46076
rect 297004 46074 297604 46076
rect 333004 46074 333604 46076
rect 369004 46074 369604 46076
rect 405004 46074 405604 46076
rect 441004 46074 441604 46076
rect 477004 46074 477604 46076
rect 513004 46074 513604 46076
rect 549004 46074 549604 46076
rect 589080 46074 589680 46076
rect -3876 43076 -3276 43078
rect 5404 43076 6004 43078
rect 41404 43076 42004 43078
rect 77404 43076 78004 43078
rect 113404 43076 114004 43078
rect 149404 43076 150004 43078
rect 185404 43076 186004 43078
rect 221404 43076 222004 43078
rect 257404 43076 258004 43078
rect 293404 43076 294004 43078
rect 329404 43076 330004 43078
rect 365404 43076 366004 43078
rect 401404 43076 402004 43078
rect 437404 43076 438004 43078
rect 473404 43076 474004 43078
rect 509404 43076 510004 43078
rect 545404 43076 546004 43078
rect 581404 43076 582004 43078
rect 587200 43076 587800 43078
rect -4816 43054 588740 43076
rect -4816 42818 -3694 43054
rect -3458 42818 5586 43054
rect 5822 42818 41586 43054
rect 41822 42818 77586 43054
rect 77822 42818 113586 43054
rect 113822 42818 149586 43054
rect 149822 42818 185586 43054
rect 185822 42818 221586 43054
rect 221822 42818 257586 43054
rect 257822 42818 293586 43054
rect 293822 42818 329586 43054
rect 329822 42818 365586 43054
rect 365822 42818 401586 43054
rect 401822 42818 437586 43054
rect 437822 42818 473586 43054
rect 473822 42818 509586 43054
rect 509822 42818 545586 43054
rect 545822 42818 581586 43054
rect 581822 42818 587382 43054
rect 587618 42818 588740 43054
rect -4816 42734 588740 42818
rect -4816 42498 -3694 42734
rect -3458 42498 5586 42734
rect 5822 42498 41586 42734
rect 41822 42498 77586 42734
rect 77822 42498 113586 42734
rect 113822 42498 149586 42734
rect 149822 42498 185586 42734
rect 185822 42498 221586 42734
rect 221822 42498 257586 42734
rect 257822 42498 293586 42734
rect 293822 42498 329586 42734
rect 329822 42498 365586 42734
rect 365822 42498 401586 42734
rect 401822 42498 437586 42734
rect 437822 42498 473586 42734
rect 473822 42498 509586 42734
rect 509822 42498 545586 42734
rect 545822 42498 581586 42734
rect 581822 42498 587382 42734
rect 587618 42498 588740 42734
rect -4816 42476 588740 42498
rect -3876 42474 -3276 42476
rect 5404 42474 6004 42476
rect 41404 42474 42004 42476
rect 77404 42474 78004 42476
rect 113404 42474 114004 42476
rect 149404 42474 150004 42476
rect 185404 42474 186004 42476
rect 221404 42474 222004 42476
rect 257404 42474 258004 42476
rect 293404 42474 294004 42476
rect 329404 42474 330004 42476
rect 365404 42474 366004 42476
rect 401404 42474 402004 42476
rect 437404 42474 438004 42476
rect 473404 42474 474004 42476
rect 509404 42474 510004 42476
rect 545404 42474 546004 42476
rect 581404 42474 582004 42476
rect 587200 42474 587800 42476
rect -1996 39476 -1396 39478
rect 1804 39476 2404 39478
rect 37804 39476 38404 39478
rect 73804 39476 74404 39478
rect 109804 39476 110404 39478
rect 145804 39476 146404 39478
rect 181804 39476 182404 39478
rect 217804 39476 218404 39478
rect 253804 39476 254404 39478
rect 289804 39476 290404 39478
rect 325804 39476 326404 39478
rect 361804 39476 362404 39478
rect 397804 39476 398404 39478
rect 433804 39476 434404 39478
rect 469804 39476 470404 39478
rect 505804 39476 506404 39478
rect 541804 39476 542404 39478
rect 577804 39476 578404 39478
rect 585320 39476 585920 39478
rect -2936 39454 586860 39476
rect -2936 39218 -1814 39454
rect -1578 39218 1986 39454
rect 2222 39218 37986 39454
rect 38222 39218 73986 39454
rect 74222 39218 109986 39454
rect 110222 39218 145986 39454
rect 146222 39218 181986 39454
rect 182222 39218 217986 39454
rect 218222 39218 253986 39454
rect 254222 39218 289986 39454
rect 290222 39218 325986 39454
rect 326222 39218 361986 39454
rect 362222 39218 397986 39454
rect 398222 39218 433986 39454
rect 434222 39218 469986 39454
rect 470222 39218 505986 39454
rect 506222 39218 541986 39454
rect 542222 39218 577986 39454
rect 578222 39218 585502 39454
rect 585738 39218 586860 39454
rect -2936 39134 586860 39218
rect -2936 38898 -1814 39134
rect -1578 38898 1986 39134
rect 2222 38898 37986 39134
rect 38222 38898 73986 39134
rect 74222 38898 109986 39134
rect 110222 38898 145986 39134
rect 146222 38898 181986 39134
rect 182222 38898 217986 39134
rect 218222 38898 253986 39134
rect 254222 38898 289986 39134
rect 290222 38898 325986 39134
rect 326222 38898 361986 39134
rect 362222 38898 397986 39134
rect 398222 38898 433986 39134
rect 434222 38898 469986 39134
rect 470222 38898 505986 39134
rect 506222 38898 541986 39134
rect 542222 38898 577986 39134
rect 578222 38898 585502 39134
rect 585738 38898 586860 39134
rect -2936 38876 586860 38898
rect -1996 38874 -1396 38876
rect 1804 38874 2404 38876
rect 37804 38874 38404 38876
rect 73804 38874 74404 38876
rect 109804 38874 110404 38876
rect 145804 38874 146404 38876
rect 181804 38874 182404 38876
rect 217804 38874 218404 38876
rect 253804 38874 254404 38876
rect 289804 38874 290404 38876
rect 325804 38874 326404 38876
rect 361804 38874 362404 38876
rect 397804 38874 398404 38876
rect 433804 38874 434404 38876
rect 469804 38874 470404 38876
rect 505804 38874 506404 38876
rect 541804 38874 542404 38876
rect 577804 38874 578404 38876
rect 585320 38874 585920 38876
rect -8576 32276 -7976 32278
rect 30604 32276 31204 32278
rect 66604 32276 67204 32278
rect 102604 32276 103204 32278
rect 138604 32276 139204 32278
rect 174604 32276 175204 32278
rect 210604 32276 211204 32278
rect 246604 32276 247204 32278
rect 282604 32276 283204 32278
rect 318604 32276 319204 32278
rect 354604 32276 355204 32278
rect 390604 32276 391204 32278
rect 426604 32276 427204 32278
rect 462604 32276 463204 32278
rect 498604 32276 499204 32278
rect 534604 32276 535204 32278
rect 570604 32276 571204 32278
rect 591900 32276 592500 32278
rect -8576 32254 592500 32276
rect -8576 32018 -8394 32254
rect -8158 32018 30786 32254
rect 31022 32018 66786 32254
rect 67022 32018 102786 32254
rect 103022 32018 138786 32254
rect 139022 32018 174786 32254
rect 175022 32018 210786 32254
rect 211022 32018 246786 32254
rect 247022 32018 282786 32254
rect 283022 32018 318786 32254
rect 319022 32018 354786 32254
rect 355022 32018 390786 32254
rect 391022 32018 426786 32254
rect 427022 32018 462786 32254
rect 463022 32018 498786 32254
rect 499022 32018 534786 32254
rect 535022 32018 570786 32254
rect 571022 32018 592082 32254
rect 592318 32018 592500 32254
rect -8576 31934 592500 32018
rect -8576 31698 -8394 31934
rect -8158 31698 30786 31934
rect 31022 31698 66786 31934
rect 67022 31698 102786 31934
rect 103022 31698 138786 31934
rect 139022 31698 174786 31934
rect 175022 31698 210786 31934
rect 211022 31698 246786 31934
rect 247022 31698 282786 31934
rect 283022 31698 318786 31934
rect 319022 31698 354786 31934
rect 355022 31698 390786 31934
rect 391022 31698 426786 31934
rect 427022 31698 462786 31934
rect 463022 31698 498786 31934
rect 499022 31698 534786 31934
rect 535022 31698 570786 31934
rect 571022 31698 592082 31934
rect 592318 31698 592500 31934
rect -8576 31676 592500 31698
rect -8576 31674 -7976 31676
rect 30604 31674 31204 31676
rect 66604 31674 67204 31676
rect 102604 31674 103204 31676
rect 138604 31674 139204 31676
rect 174604 31674 175204 31676
rect 210604 31674 211204 31676
rect 246604 31674 247204 31676
rect 282604 31674 283204 31676
rect 318604 31674 319204 31676
rect 354604 31674 355204 31676
rect 390604 31674 391204 31676
rect 426604 31674 427204 31676
rect 462604 31674 463204 31676
rect 498604 31674 499204 31676
rect 534604 31674 535204 31676
rect 570604 31674 571204 31676
rect 591900 31674 592500 31676
rect -6696 28676 -6096 28678
rect 27004 28676 27604 28678
rect 63004 28676 63604 28678
rect 99004 28676 99604 28678
rect 135004 28676 135604 28678
rect 171004 28676 171604 28678
rect 207004 28676 207604 28678
rect 243004 28676 243604 28678
rect 279004 28676 279604 28678
rect 315004 28676 315604 28678
rect 351004 28676 351604 28678
rect 387004 28676 387604 28678
rect 423004 28676 423604 28678
rect 459004 28676 459604 28678
rect 495004 28676 495604 28678
rect 531004 28676 531604 28678
rect 567004 28676 567604 28678
rect 590020 28676 590620 28678
rect -6696 28654 590620 28676
rect -6696 28418 -6514 28654
rect -6278 28418 27186 28654
rect 27422 28418 63186 28654
rect 63422 28418 99186 28654
rect 99422 28418 135186 28654
rect 135422 28418 171186 28654
rect 171422 28418 207186 28654
rect 207422 28418 243186 28654
rect 243422 28418 279186 28654
rect 279422 28418 315186 28654
rect 315422 28418 351186 28654
rect 351422 28418 387186 28654
rect 387422 28418 423186 28654
rect 423422 28418 459186 28654
rect 459422 28418 495186 28654
rect 495422 28418 531186 28654
rect 531422 28418 567186 28654
rect 567422 28418 590202 28654
rect 590438 28418 590620 28654
rect -6696 28334 590620 28418
rect -6696 28098 -6514 28334
rect -6278 28098 27186 28334
rect 27422 28098 63186 28334
rect 63422 28098 99186 28334
rect 99422 28098 135186 28334
rect 135422 28098 171186 28334
rect 171422 28098 207186 28334
rect 207422 28098 243186 28334
rect 243422 28098 279186 28334
rect 279422 28098 315186 28334
rect 315422 28098 351186 28334
rect 351422 28098 387186 28334
rect 387422 28098 423186 28334
rect 423422 28098 459186 28334
rect 459422 28098 495186 28334
rect 495422 28098 531186 28334
rect 531422 28098 567186 28334
rect 567422 28098 590202 28334
rect 590438 28098 590620 28334
rect -6696 28076 590620 28098
rect -6696 28074 -6096 28076
rect 27004 28074 27604 28076
rect 63004 28074 63604 28076
rect 99004 28074 99604 28076
rect 135004 28074 135604 28076
rect 171004 28074 171604 28076
rect 207004 28074 207604 28076
rect 243004 28074 243604 28076
rect 279004 28074 279604 28076
rect 315004 28074 315604 28076
rect 351004 28074 351604 28076
rect 387004 28074 387604 28076
rect 423004 28074 423604 28076
rect 459004 28074 459604 28076
rect 495004 28074 495604 28076
rect 531004 28074 531604 28076
rect 567004 28074 567604 28076
rect 590020 28074 590620 28076
rect -4816 25076 -4216 25078
rect 23404 25076 24004 25078
rect 59404 25076 60004 25078
rect 95404 25076 96004 25078
rect 131404 25076 132004 25078
rect 167404 25076 168004 25078
rect 203404 25076 204004 25078
rect 239404 25076 240004 25078
rect 275404 25076 276004 25078
rect 311404 25076 312004 25078
rect 347404 25076 348004 25078
rect 383404 25076 384004 25078
rect 419404 25076 420004 25078
rect 455404 25076 456004 25078
rect 491404 25076 492004 25078
rect 527404 25076 528004 25078
rect 563404 25076 564004 25078
rect 588140 25076 588740 25078
rect -4816 25054 588740 25076
rect -4816 24818 -4634 25054
rect -4398 24818 23586 25054
rect 23822 24818 59586 25054
rect 59822 24818 95586 25054
rect 95822 24818 131586 25054
rect 131822 24818 167586 25054
rect 167822 24818 203586 25054
rect 203822 24818 239586 25054
rect 239822 24818 275586 25054
rect 275822 24818 311586 25054
rect 311822 24818 347586 25054
rect 347822 24818 383586 25054
rect 383822 24818 419586 25054
rect 419822 24818 455586 25054
rect 455822 24818 491586 25054
rect 491822 24818 527586 25054
rect 527822 24818 563586 25054
rect 563822 24818 588322 25054
rect 588558 24818 588740 25054
rect -4816 24734 588740 24818
rect -4816 24498 -4634 24734
rect -4398 24498 23586 24734
rect 23822 24498 59586 24734
rect 59822 24498 95586 24734
rect 95822 24498 131586 24734
rect 131822 24498 167586 24734
rect 167822 24498 203586 24734
rect 203822 24498 239586 24734
rect 239822 24498 275586 24734
rect 275822 24498 311586 24734
rect 311822 24498 347586 24734
rect 347822 24498 383586 24734
rect 383822 24498 419586 24734
rect 419822 24498 455586 24734
rect 455822 24498 491586 24734
rect 491822 24498 527586 24734
rect 527822 24498 563586 24734
rect 563822 24498 588322 24734
rect 588558 24498 588740 24734
rect -4816 24476 588740 24498
rect -4816 24474 -4216 24476
rect 23404 24474 24004 24476
rect 59404 24474 60004 24476
rect 95404 24474 96004 24476
rect 131404 24474 132004 24476
rect 167404 24474 168004 24476
rect 203404 24474 204004 24476
rect 239404 24474 240004 24476
rect 275404 24474 276004 24476
rect 311404 24474 312004 24476
rect 347404 24474 348004 24476
rect 383404 24474 384004 24476
rect 419404 24474 420004 24476
rect 455404 24474 456004 24476
rect 491404 24474 492004 24476
rect 527404 24474 528004 24476
rect 563404 24474 564004 24476
rect 588140 24474 588740 24476
rect -2936 21476 -2336 21478
rect 19804 21476 20404 21478
rect 55804 21476 56404 21478
rect 91804 21476 92404 21478
rect 127804 21476 128404 21478
rect 163804 21476 164404 21478
rect 199804 21476 200404 21478
rect 235804 21476 236404 21478
rect 271804 21476 272404 21478
rect 307804 21476 308404 21478
rect 343804 21476 344404 21478
rect 379804 21476 380404 21478
rect 415804 21476 416404 21478
rect 451804 21476 452404 21478
rect 487804 21476 488404 21478
rect 523804 21476 524404 21478
rect 559804 21476 560404 21478
rect 586260 21476 586860 21478
rect -2936 21454 586860 21476
rect -2936 21218 -2754 21454
rect -2518 21218 19986 21454
rect 20222 21218 55986 21454
rect 56222 21218 91986 21454
rect 92222 21218 127986 21454
rect 128222 21218 163986 21454
rect 164222 21218 199986 21454
rect 200222 21218 235986 21454
rect 236222 21218 271986 21454
rect 272222 21218 307986 21454
rect 308222 21218 343986 21454
rect 344222 21218 379986 21454
rect 380222 21218 415986 21454
rect 416222 21218 451986 21454
rect 452222 21218 487986 21454
rect 488222 21218 523986 21454
rect 524222 21218 559986 21454
rect 560222 21218 586442 21454
rect 586678 21218 586860 21454
rect -2936 21134 586860 21218
rect -2936 20898 -2754 21134
rect -2518 20898 19986 21134
rect 20222 20898 55986 21134
rect 56222 20898 91986 21134
rect 92222 20898 127986 21134
rect 128222 20898 163986 21134
rect 164222 20898 199986 21134
rect 200222 20898 235986 21134
rect 236222 20898 271986 21134
rect 272222 20898 307986 21134
rect 308222 20898 343986 21134
rect 344222 20898 379986 21134
rect 380222 20898 415986 21134
rect 416222 20898 451986 21134
rect 452222 20898 487986 21134
rect 488222 20898 523986 21134
rect 524222 20898 559986 21134
rect 560222 20898 586442 21134
rect 586678 20898 586860 21134
rect -2936 20876 586860 20898
rect -2936 20874 -2336 20876
rect 19804 20874 20404 20876
rect 55804 20874 56404 20876
rect 91804 20874 92404 20876
rect 127804 20874 128404 20876
rect 163804 20874 164404 20876
rect 199804 20874 200404 20876
rect 235804 20874 236404 20876
rect 271804 20874 272404 20876
rect 307804 20874 308404 20876
rect 343804 20874 344404 20876
rect 379804 20874 380404 20876
rect 415804 20874 416404 20876
rect 451804 20874 452404 20876
rect 487804 20874 488404 20876
rect 523804 20874 524404 20876
rect 559804 20874 560404 20876
rect 586260 20874 586860 20876
rect -7636 14276 -7036 14278
rect 12604 14276 13204 14278
rect 48604 14276 49204 14278
rect 84604 14276 85204 14278
rect 120604 14276 121204 14278
rect 156604 14276 157204 14278
rect 192604 14276 193204 14278
rect 228604 14276 229204 14278
rect 264604 14276 265204 14278
rect 300604 14276 301204 14278
rect 336604 14276 337204 14278
rect 372604 14276 373204 14278
rect 408604 14276 409204 14278
rect 444604 14276 445204 14278
rect 480604 14276 481204 14278
rect 516604 14276 517204 14278
rect 552604 14276 553204 14278
rect 590960 14276 591560 14278
rect -8576 14254 592500 14276
rect -8576 14018 -7454 14254
rect -7218 14018 12786 14254
rect 13022 14018 48786 14254
rect 49022 14018 84786 14254
rect 85022 14018 120786 14254
rect 121022 14018 156786 14254
rect 157022 14018 192786 14254
rect 193022 14018 228786 14254
rect 229022 14018 264786 14254
rect 265022 14018 300786 14254
rect 301022 14018 336786 14254
rect 337022 14018 372786 14254
rect 373022 14018 408786 14254
rect 409022 14018 444786 14254
rect 445022 14018 480786 14254
rect 481022 14018 516786 14254
rect 517022 14018 552786 14254
rect 553022 14018 591142 14254
rect 591378 14018 592500 14254
rect -8576 13934 592500 14018
rect -8576 13698 -7454 13934
rect -7218 13698 12786 13934
rect 13022 13698 48786 13934
rect 49022 13698 84786 13934
rect 85022 13698 120786 13934
rect 121022 13698 156786 13934
rect 157022 13698 192786 13934
rect 193022 13698 228786 13934
rect 229022 13698 264786 13934
rect 265022 13698 300786 13934
rect 301022 13698 336786 13934
rect 337022 13698 372786 13934
rect 373022 13698 408786 13934
rect 409022 13698 444786 13934
rect 445022 13698 480786 13934
rect 481022 13698 516786 13934
rect 517022 13698 552786 13934
rect 553022 13698 591142 13934
rect 591378 13698 592500 13934
rect -8576 13676 592500 13698
rect -7636 13674 -7036 13676
rect 12604 13674 13204 13676
rect 48604 13674 49204 13676
rect 84604 13674 85204 13676
rect 120604 13674 121204 13676
rect 156604 13674 157204 13676
rect 192604 13674 193204 13676
rect 228604 13674 229204 13676
rect 264604 13674 265204 13676
rect 300604 13674 301204 13676
rect 336604 13674 337204 13676
rect 372604 13674 373204 13676
rect 408604 13674 409204 13676
rect 444604 13674 445204 13676
rect 480604 13674 481204 13676
rect 516604 13674 517204 13676
rect 552604 13674 553204 13676
rect 590960 13674 591560 13676
rect -5756 10676 -5156 10678
rect 9004 10676 9604 10678
rect 45004 10676 45604 10678
rect 81004 10676 81604 10678
rect 117004 10676 117604 10678
rect 153004 10676 153604 10678
rect 189004 10676 189604 10678
rect 225004 10676 225604 10678
rect 261004 10676 261604 10678
rect 297004 10676 297604 10678
rect 333004 10676 333604 10678
rect 369004 10676 369604 10678
rect 405004 10676 405604 10678
rect 441004 10676 441604 10678
rect 477004 10676 477604 10678
rect 513004 10676 513604 10678
rect 549004 10676 549604 10678
rect 589080 10676 589680 10678
rect -6696 10654 590620 10676
rect -6696 10418 -5574 10654
rect -5338 10418 9186 10654
rect 9422 10418 45186 10654
rect 45422 10418 81186 10654
rect 81422 10418 117186 10654
rect 117422 10418 153186 10654
rect 153422 10418 189186 10654
rect 189422 10418 225186 10654
rect 225422 10418 261186 10654
rect 261422 10418 297186 10654
rect 297422 10418 333186 10654
rect 333422 10418 369186 10654
rect 369422 10418 405186 10654
rect 405422 10418 441186 10654
rect 441422 10418 477186 10654
rect 477422 10418 513186 10654
rect 513422 10418 549186 10654
rect 549422 10418 589262 10654
rect 589498 10418 590620 10654
rect -6696 10334 590620 10418
rect -6696 10098 -5574 10334
rect -5338 10098 9186 10334
rect 9422 10098 45186 10334
rect 45422 10098 81186 10334
rect 81422 10098 117186 10334
rect 117422 10098 153186 10334
rect 153422 10098 189186 10334
rect 189422 10098 225186 10334
rect 225422 10098 261186 10334
rect 261422 10098 297186 10334
rect 297422 10098 333186 10334
rect 333422 10098 369186 10334
rect 369422 10098 405186 10334
rect 405422 10098 441186 10334
rect 441422 10098 477186 10334
rect 477422 10098 513186 10334
rect 513422 10098 549186 10334
rect 549422 10098 589262 10334
rect 589498 10098 590620 10334
rect -6696 10076 590620 10098
rect -5756 10074 -5156 10076
rect 9004 10074 9604 10076
rect 45004 10074 45604 10076
rect 81004 10074 81604 10076
rect 117004 10074 117604 10076
rect 153004 10074 153604 10076
rect 189004 10074 189604 10076
rect 225004 10074 225604 10076
rect 261004 10074 261604 10076
rect 297004 10074 297604 10076
rect 333004 10074 333604 10076
rect 369004 10074 369604 10076
rect 405004 10074 405604 10076
rect 441004 10074 441604 10076
rect 477004 10074 477604 10076
rect 513004 10074 513604 10076
rect 549004 10074 549604 10076
rect 589080 10074 589680 10076
rect -3876 7076 -3276 7078
rect 5404 7076 6004 7078
rect 41404 7076 42004 7078
rect 77404 7076 78004 7078
rect 113404 7076 114004 7078
rect 149404 7076 150004 7078
rect 185404 7076 186004 7078
rect 221404 7076 222004 7078
rect 257404 7076 258004 7078
rect 293404 7076 294004 7078
rect 329404 7076 330004 7078
rect 365404 7076 366004 7078
rect 401404 7076 402004 7078
rect 437404 7076 438004 7078
rect 473404 7076 474004 7078
rect 509404 7076 510004 7078
rect 545404 7076 546004 7078
rect 581404 7076 582004 7078
rect 587200 7076 587800 7078
rect -4816 7054 588740 7076
rect -4816 6818 -3694 7054
rect -3458 6818 5586 7054
rect 5822 6818 41586 7054
rect 41822 6818 77586 7054
rect 77822 6818 113586 7054
rect 113822 6818 149586 7054
rect 149822 6818 185586 7054
rect 185822 6818 221586 7054
rect 221822 6818 257586 7054
rect 257822 6818 293586 7054
rect 293822 6818 329586 7054
rect 329822 6818 365586 7054
rect 365822 6818 401586 7054
rect 401822 6818 437586 7054
rect 437822 6818 473586 7054
rect 473822 6818 509586 7054
rect 509822 6818 545586 7054
rect 545822 6818 581586 7054
rect 581822 6818 587382 7054
rect 587618 6818 588740 7054
rect -4816 6734 588740 6818
rect -4816 6498 -3694 6734
rect -3458 6498 5586 6734
rect 5822 6498 41586 6734
rect 41822 6498 77586 6734
rect 77822 6498 113586 6734
rect 113822 6498 149586 6734
rect 149822 6498 185586 6734
rect 185822 6498 221586 6734
rect 221822 6498 257586 6734
rect 257822 6498 293586 6734
rect 293822 6498 329586 6734
rect 329822 6498 365586 6734
rect 365822 6498 401586 6734
rect 401822 6498 437586 6734
rect 437822 6498 473586 6734
rect 473822 6498 509586 6734
rect 509822 6498 545586 6734
rect 545822 6498 581586 6734
rect 581822 6498 587382 6734
rect 587618 6498 588740 6734
rect -4816 6476 588740 6498
rect -3876 6474 -3276 6476
rect 5404 6474 6004 6476
rect 41404 6474 42004 6476
rect 77404 6474 78004 6476
rect 113404 6474 114004 6476
rect 149404 6474 150004 6476
rect 185404 6474 186004 6476
rect 221404 6474 222004 6476
rect 257404 6474 258004 6476
rect 293404 6474 294004 6476
rect 329404 6474 330004 6476
rect 365404 6474 366004 6476
rect 401404 6474 402004 6476
rect 437404 6474 438004 6476
rect 473404 6474 474004 6476
rect 509404 6474 510004 6476
rect 545404 6474 546004 6476
rect 581404 6474 582004 6476
rect 587200 6474 587800 6476
rect -1996 3476 -1396 3478
rect 1804 3476 2404 3478
rect 37804 3476 38404 3478
rect 73804 3476 74404 3478
rect 109804 3476 110404 3478
rect 145804 3476 146404 3478
rect 181804 3476 182404 3478
rect 217804 3476 218404 3478
rect 253804 3476 254404 3478
rect 289804 3476 290404 3478
rect 325804 3476 326404 3478
rect 361804 3476 362404 3478
rect 397804 3476 398404 3478
rect 433804 3476 434404 3478
rect 469804 3476 470404 3478
rect 505804 3476 506404 3478
rect 541804 3476 542404 3478
rect 577804 3476 578404 3478
rect 585320 3476 585920 3478
rect -2936 3454 586860 3476
rect -2936 3218 -1814 3454
rect -1578 3218 1986 3454
rect 2222 3218 37986 3454
rect 38222 3218 73986 3454
rect 74222 3218 109986 3454
rect 110222 3218 145986 3454
rect 146222 3218 181986 3454
rect 182222 3218 217986 3454
rect 218222 3218 253986 3454
rect 254222 3218 289986 3454
rect 290222 3218 325986 3454
rect 326222 3218 361986 3454
rect 362222 3218 397986 3454
rect 398222 3218 433986 3454
rect 434222 3218 469986 3454
rect 470222 3218 505986 3454
rect 506222 3218 541986 3454
rect 542222 3218 577986 3454
rect 578222 3218 585502 3454
rect 585738 3218 586860 3454
rect -2936 3134 586860 3218
rect -2936 2898 -1814 3134
rect -1578 2898 1986 3134
rect 2222 2898 37986 3134
rect 38222 2898 73986 3134
rect 74222 2898 109986 3134
rect 110222 2898 145986 3134
rect 146222 2898 181986 3134
rect 182222 2898 217986 3134
rect 218222 2898 253986 3134
rect 254222 2898 289986 3134
rect 290222 2898 325986 3134
rect 326222 2898 361986 3134
rect 362222 2898 397986 3134
rect 398222 2898 433986 3134
rect 434222 2898 469986 3134
rect 470222 2898 505986 3134
rect 506222 2898 541986 3134
rect 542222 2898 577986 3134
rect 578222 2898 585502 3134
rect 585738 2898 586860 3134
rect -2936 2876 586860 2898
rect -1996 2874 -1396 2876
rect 1804 2874 2404 2876
rect 37804 2874 38404 2876
rect 73804 2874 74404 2876
rect 109804 2874 110404 2876
rect 145804 2874 146404 2876
rect 181804 2874 182404 2876
rect 217804 2874 218404 2876
rect 253804 2874 254404 2876
rect 289804 2874 290404 2876
rect 325804 2874 326404 2876
rect 361804 2874 362404 2876
rect 397804 2874 398404 2876
rect 433804 2874 434404 2876
rect 469804 2874 470404 2876
rect 505804 2874 506404 2876
rect 541804 2874 542404 2876
rect 577804 2874 578404 2876
rect 585320 2874 585920 2876
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 1986 -346
rect 2222 -582 37986 -346
rect 38222 -582 73986 -346
rect 74222 -582 109986 -346
rect 110222 -582 145986 -346
rect 146222 -582 181986 -346
rect 182222 -582 217986 -346
rect 218222 -582 253986 -346
rect 254222 -582 289986 -346
rect 290222 -582 325986 -346
rect 326222 -582 361986 -346
rect 362222 -582 397986 -346
rect 398222 -582 433986 -346
rect 434222 -582 469986 -346
rect 470222 -582 505986 -346
rect 506222 -582 541986 -346
rect 542222 -582 577986 -346
rect 578222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 1986 -666
rect 2222 -902 37986 -666
rect 38222 -902 73986 -666
rect 74222 -902 109986 -666
rect 110222 -902 145986 -666
rect 146222 -902 181986 -666
rect 182222 -902 217986 -666
rect 218222 -902 253986 -666
rect 254222 -902 289986 -666
rect 290222 -902 325986 -666
rect 326222 -902 361986 -666
rect 362222 -902 397986 -666
rect 398222 -902 433986 -666
rect 434222 -902 469986 -666
rect 470222 -902 505986 -666
rect 506222 -902 541986 -666
rect 542222 -902 577986 -666
rect 578222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 19986 -1286
rect 20222 -1522 55986 -1286
rect 56222 -1522 91986 -1286
rect 92222 -1522 127986 -1286
rect 128222 -1522 163986 -1286
rect 164222 -1522 199986 -1286
rect 200222 -1522 235986 -1286
rect 236222 -1522 271986 -1286
rect 272222 -1522 307986 -1286
rect 308222 -1522 343986 -1286
rect 344222 -1522 379986 -1286
rect 380222 -1522 415986 -1286
rect 416222 -1522 451986 -1286
rect 452222 -1522 487986 -1286
rect 488222 -1522 523986 -1286
rect 524222 -1522 559986 -1286
rect 560222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 19986 -1606
rect 20222 -1842 55986 -1606
rect 56222 -1842 91986 -1606
rect 92222 -1842 127986 -1606
rect 128222 -1842 163986 -1606
rect 164222 -1842 199986 -1606
rect 200222 -1842 235986 -1606
rect 236222 -1842 271986 -1606
rect 272222 -1842 307986 -1606
rect 308222 -1842 343986 -1606
rect 344222 -1842 379986 -1606
rect 380222 -1842 415986 -1606
rect 416222 -1842 451986 -1606
rect 452222 -1842 487986 -1606
rect 488222 -1842 523986 -1606
rect 524222 -1842 559986 -1606
rect 560222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 5586 -2226
rect 5822 -2462 41586 -2226
rect 41822 -2462 77586 -2226
rect 77822 -2462 113586 -2226
rect 113822 -2462 149586 -2226
rect 149822 -2462 185586 -2226
rect 185822 -2462 221586 -2226
rect 221822 -2462 257586 -2226
rect 257822 -2462 293586 -2226
rect 293822 -2462 329586 -2226
rect 329822 -2462 365586 -2226
rect 365822 -2462 401586 -2226
rect 401822 -2462 437586 -2226
rect 437822 -2462 473586 -2226
rect 473822 -2462 509586 -2226
rect 509822 -2462 545586 -2226
rect 545822 -2462 581586 -2226
rect 581822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 5586 -2546
rect 5822 -2782 41586 -2546
rect 41822 -2782 77586 -2546
rect 77822 -2782 113586 -2546
rect 113822 -2782 149586 -2546
rect 149822 -2782 185586 -2546
rect 185822 -2782 221586 -2546
rect 221822 -2782 257586 -2546
rect 257822 -2782 293586 -2546
rect 293822 -2782 329586 -2546
rect 329822 -2782 365586 -2546
rect 365822 -2782 401586 -2546
rect 401822 -2782 437586 -2546
rect 437822 -2782 473586 -2546
rect 473822 -2782 509586 -2546
rect 509822 -2782 545586 -2546
rect 545822 -2782 581586 -2546
rect 581822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 23586 -3166
rect 23822 -3402 59586 -3166
rect 59822 -3402 95586 -3166
rect 95822 -3402 131586 -3166
rect 131822 -3402 167586 -3166
rect 167822 -3402 203586 -3166
rect 203822 -3402 239586 -3166
rect 239822 -3402 275586 -3166
rect 275822 -3402 311586 -3166
rect 311822 -3402 347586 -3166
rect 347822 -3402 383586 -3166
rect 383822 -3402 419586 -3166
rect 419822 -3402 455586 -3166
rect 455822 -3402 491586 -3166
rect 491822 -3402 527586 -3166
rect 527822 -3402 563586 -3166
rect 563822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 23586 -3486
rect 23822 -3722 59586 -3486
rect 59822 -3722 95586 -3486
rect 95822 -3722 131586 -3486
rect 131822 -3722 167586 -3486
rect 167822 -3722 203586 -3486
rect 203822 -3722 239586 -3486
rect 239822 -3722 275586 -3486
rect 275822 -3722 311586 -3486
rect 311822 -3722 347586 -3486
rect 347822 -3722 383586 -3486
rect 383822 -3722 419586 -3486
rect 419822 -3722 455586 -3486
rect 455822 -3722 491586 -3486
rect 491822 -3722 527586 -3486
rect 527822 -3722 563586 -3486
rect 563822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 9186 -4106
rect 9422 -4342 45186 -4106
rect 45422 -4342 81186 -4106
rect 81422 -4342 117186 -4106
rect 117422 -4342 153186 -4106
rect 153422 -4342 189186 -4106
rect 189422 -4342 225186 -4106
rect 225422 -4342 261186 -4106
rect 261422 -4342 297186 -4106
rect 297422 -4342 333186 -4106
rect 333422 -4342 369186 -4106
rect 369422 -4342 405186 -4106
rect 405422 -4342 441186 -4106
rect 441422 -4342 477186 -4106
rect 477422 -4342 513186 -4106
rect 513422 -4342 549186 -4106
rect 549422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 9186 -4426
rect 9422 -4662 45186 -4426
rect 45422 -4662 81186 -4426
rect 81422 -4662 117186 -4426
rect 117422 -4662 153186 -4426
rect 153422 -4662 189186 -4426
rect 189422 -4662 225186 -4426
rect 225422 -4662 261186 -4426
rect 261422 -4662 297186 -4426
rect 297422 -4662 333186 -4426
rect 333422 -4662 369186 -4426
rect 369422 -4662 405186 -4426
rect 405422 -4662 441186 -4426
rect 441422 -4662 477186 -4426
rect 477422 -4662 513186 -4426
rect 513422 -4662 549186 -4426
rect 549422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 27186 -5046
rect 27422 -5282 63186 -5046
rect 63422 -5282 99186 -5046
rect 99422 -5282 135186 -5046
rect 135422 -5282 171186 -5046
rect 171422 -5282 207186 -5046
rect 207422 -5282 243186 -5046
rect 243422 -5282 279186 -5046
rect 279422 -5282 315186 -5046
rect 315422 -5282 351186 -5046
rect 351422 -5282 387186 -5046
rect 387422 -5282 423186 -5046
rect 423422 -5282 459186 -5046
rect 459422 -5282 495186 -5046
rect 495422 -5282 531186 -5046
rect 531422 -5282 567186 -5046
rect 567422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 27186 -5366
rect 27422 -5602 63186 -5366
rect 63422 -5602 99186 -5366
rect 99422 -5602 135186 -5366
rect 135422 -5602 171186 -5366
rect 171422 -5602 207186 -5366
rect 207422 -5602 243186 -5366
rect 243422 -5602 279186 -5366
rect 279422 -5602 315186 -5366
rect 315422 -5602 351186 -5366
rect 351422 -5602 387186 -5366
rect 387422 -5602 423186 -5366
rect 423422 -5602 459186 -5366
rect 459422 -5602 495186 -5366
rect 495422 -5602 531186 -5366
rect 531422 -5602 567186 -5366
rect 567422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 12786 -5986
rect 13022 -6222 48786 -5986
rect 49022 -6222 84786 -5986
rect 85022 -6222 120786 -5986
rect 121022 -6222 156786 -5986
rect 157022 -6222 192786 -5986
rect 193022 -6222 228786 -5986
rect 229022 -6222 264786 -5986
rect 265022 -6222 300786 -5986
rect 301022 -6222 336786 -5986
rect 337022 -6222 372786 -5986
rect 373022 -6222 408786 -5986
rect 409022 -6222 444786 -5986
rect 445022 -6222 480786 -5986
rect 481022 -6222 516786 -5986
rect 517022 -6222 552786 -5986
rect 553022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 12786 -6306
rect 13022 -6542 48786 -6306
rect 49022 -6542 84786 -6306
rect 85022 -6542 120786 -6306
rect 121022 -6542 156786 -6306
rect 157022 -6542 192786 -6306
rect 193022 -6542 228786 -6306
rect 229022 -6542 264786 -6306
rect 265022 -6542 300786 -6306
rect 301022 -6542 336786 -6306
rect 337022 -6542 372786 -6306
rect 373022 -6542 408786 -6306
rect 409022 -6542 444786 -6306
rect 445022 -6542 480786 -6306
rect 481022 -6542 516786 -6306
rect 517022 -6542 552786 -6306
rect 553022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 30786 -6926
rect 31022 -7162 66786 -6926
rect 67022 -7162 102786 -6926
rect 103022 -7162 138786 -6926
rect 139022 -7162 174786 -6926
rect 175022 -7162 210786 -6926
rect 211022 -7162 246786 -6926
rect 247022 -7162 282786 -6926
rect 283022 -7162 318786 -6926
rect 319022 -7162 354786 -6926
rect 355022 -7162 390786 -6926
rect 391022 -7162 426786 -6926
rect 427022 -7162 462786 -6926
rect 463022 -7162 498786 -6926
rect 499022 -7162 534786 -6926
rect 535022 -7162 570786 -6926
rect 571022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 30786 -7246
rect 31022 -7482 66786 -7246
rect 67022 -7482 102786 -7246
rect 103022 -7482 138786 -7246
rect 139022 -7482 174786 -7246
rect 175022 -7482 210786 -7246
rect 211022 -7482 246786 -7246
rect 247022 -7482 282786 -7246
rect 283022 -7482 318786 -7246
rect 319022 -7482 354786 -7246
rect 355022 -7482 390786 -7246
rect 391022 -7482 426786 -7246
rect 427022 -7482 462786 -7246
rect 463022 -7482 498786 -7246
rect 499022 -7482 534786 -7246
rect 535022 -7482 570786 -7246
rect 571022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
use adc_wrapper  mprj
timestamp 1626434083
transform 1 0 168000 0 1 338000
box 0 0 260000 160000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 533 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 599 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 600 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 601 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 602 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 603 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 604 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 605 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 606 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 607 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 608 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 609 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 610 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 611 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 612 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 613 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 614 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 615 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 616 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 617 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 618 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 619 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 620 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 621 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 622 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 623 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 624 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 625 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 626 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 627 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 628 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 629 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 630 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 577804 -1864 578404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 541804 -1864 542404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 505804 -1864 506404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 469804 -1864 470404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 433804 510000 434404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 397804 510000 398404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 361804 510000 362404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 325804 510000 326404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 289804 510000 290404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 253804 510000 254404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 217804 510000 218404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 181804 510000 182404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 145804 -1864 146404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 109804 -1864 110404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 73804 -1864 74404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 37804 -1864 38404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 1804 -1864 2404 705800 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 433804 -1864 434404 326000 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 397804 -1864 398404 326000 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 361804 -1864 362404 326000 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 325804 -1864 326404 326000 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 289804 -1864 290404 326000 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 253804 -1864 254404 326000 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 217804 -1864 218404 326000 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 181804 -1864 182404 326000 6 vccd1
port 663 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 664 nsew power bidirectional
rlabel metal5 s -2936 686876 586860 687476 6 vccd1
port 665 nsew power bidirectional
rlabel metal5 s -2936 650876 586860 651476 6 vccd1
port 666 nsew power bidirectional
rlabel metal5 s -2936 614876 586860 615476 6 vccd1
port 667 nsew power bidirectional
rlabel metal5 s -2936 578876 586860 579476 6 vccd1
port 668 nsew power bidirectional
rlabel metal5 s -2936 542876 586860 543476 6 vccd1
port 669 nsew power bidirectional
rlabel metal5 s 440000 506876 586860 507476 6 vccd1
port 670 nsew power bidirectional
rlabel metal5 s -2936 506876 156000 507476 6 vccd1
port 671 nsew power bidirectional
rlabel metal5 s 440000 470876 586860 471476 6 vccd1
port 672 nsew power bidirectional
rlabel metal5 s -2936 470876 156000 471476 6 vccd1
port 673 nsew power bidirectional
rlabel metal5 s 440000 434876 586860 435476 6 vccd1
port 674 nsew power bidirectional
rlabel metal5 s -2936 434876 156000 435476 6 vccd1
port 675 nsew power bidirectional
rlabel metal5 s 440000 398876 586860 399476 6 vccd1
port 676 nsew power bidirectional
rlabel metal5 s -2936 398876 156000 399476 6 vccd1
port 677 nsew power bidirectional
rlabel metal5 s 440000 362876 586860 363476 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s -2936 362876 156000 363476 6 vccd1
port 679 nsew power bidirectional
rlabel metal5 s 440000 326876 586860 327476 6 vccd1
port 680 nsew power bidirectional
rlabel metal5 s -2936 326876 156000 327476 6 vccd1
port 681 nsew power bidirectional
rlabel metal5 s -2936 290876 586860 291476 6 vccd1
port 682 nsew power bidirectional
rlabel metal5 s -2936 254876 586860 255476 6 vccd1
port 683 nsew power bidirectional
rlabel metal5 s -2936 218876 586860 219476 6 vccd1
port 684 nsew power bidirectional
rlabel metal5 s -2936 182876 586860 183476 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s -2936 146876 586860 147476 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s -2936 110876 586860 111476 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s -2936 74876 586860 75476 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s -2936 38876 586860 39476 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s -2936 2876 586860 3476 6 vccd1
port 690 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 691 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 692 nsew ground bidirectional
rlabel metal4 s 559804 -1864 560404 705800 6 vssd1
port 693 nsew ground bidirectional
rlabel metal4 s 523804 -1864 524404 705800 6 vssd1
port 694 nsew ground bidirectional
rlabel metal4 s 487804 -1864 488404 705800 6 vssd1
port 695 nsew ground bidirectional
rlabel metal4 s 451804 -1864 452404 705800 6 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s 415804 510000 416404 705800 6 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 379804 510000 380404 705800 6 vssd1
port 698 nsew ground bidirectional
rlabel metal4 s 343804 510000 344404 705800 6 vssd1
port 699 nsew ground bidirectional
rlabel metal4 s 307804 510000 308404 705800 6 vssd1
port 700 nsew ground bidirectional
rlabel metal4 s 271804 510000 272404 705800 6 vssd1
port 701 nsew ground bidirectional
rlabel metal4 s 235804 510000 236404 705800 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 199804 510000 200404 705800 6 vssd1
port 703 nsew ground bidirectional
rlabel metal4 s 163804 510000 164404 705800 6 vssd1
port 704 nsew ground bidirectional
rlabel metal4 s 127804 -1864 128404 705800 6 vssd1
port 705 nsew ground bidirectional
rlabel metal4 s 91804 -1864 92404 705800 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 55804 -1864 56404 705800 6 vssd1
port 707 nsew ground bidirectional
rlabel metal4 s 19804 -1864 20404 705800 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s 415804 -1864 416404 326000 6 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 379804 -1864 380404 326000 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 343804 -1864 344404 326000 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 307804 -1864 308404 326000 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 271804 -1864 272404 326000 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 235804 -1864 236404 326000 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 199804 -1864 200404 326000 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 163804 -1864 164404 326000 6 vssd1
port 717 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 718 nsew ground bidirectional
rlabel metal5 s -2936 668876 586860 669476 6 vssd1
port 719 nsew ground bidirectional
rlabel metal5 s -2936 632876 586860 633476 6 vssd1
port 720 nsew ground bidirectional
rlabel metal5 s -2936 596876 586860 597476 6 vssd1
port 721 nsew ground bidirectional
rlabel metal5 s -2936 560876 586860 561476 6 vssd1
port 722 nsew ground bidirectional
rlabel metal5 s -2936 524876 586860 525476 6 vssd1
port 723 nsew ground bidirectional
rlabel metal5 s 440000 488876 586860 489476 6 vssd1
port 724 nsew ground bidirectional
rlabel metal5 s -2936 488876 156000 489476 6 vssd1
port 725 nsew ground bidirectional
rlabel metal5 s 440000 452876 586860 453476 6 vssd1
port 726 nsew ground bidirectional
rlabel metal5 s -2936 452876 156000 453476 6 vssd1
port 727 nsew ground bidirectional
rlabel metal5 s 440000 416876 586860 417476 6 vssd1
port 728 nsew ground bidirectional
rlabel metal5 s -2936 416876 156000 417476 6 vssd1
port 729 nsew ground bidirectional
rlabel metal5 s 440000 380876 586860 381476 6 vssd1
port 730 nsew ground bidirectional
rlabel metal5 s -2936 380876 156000 381476 6 vssd1
port 731 nsew ground bidirectional
rlabel metal5 s 440000 344876 586860 345476 6 vssd1
port 732 nsew ground bidirectional
rlabel metal5 s -2936 344876 156000 345476 6 vssd1
port 733 nsew ground bidirectional
rlabel metal5 s -2936 308876 586860 309476 6 vssd1
port 734 nsew ground bidirectional
rlabel metal5 s -2936 272876 586860 273476 6 vssd1
port 735 nsew ground bidirectional
rlabel metal5 s -2936 236876 586860 237476 6 vssd1
port 736 nsew ground bidirectional
rlabel metal5 s -2936 200876 586860 201476 6 vssd1
port 737 nsew ground bidirectional
rlabel metal5 s -2936 164876 586860 165476 6 vssd1
port 738 nsew ground bidirectional
rlabel metal5 s -2936 128876 586860 129476 6 vssd1
port 739 nsew ground bidirectional
rlabel metal5 s -2936 92876 586860 93476 6 vssd1
port 740 nsew ground bidirectional
rlabel metal5 s -2936 56876 586860 57476 6 vssd1
port 741 nsew ground bidirectional
rlabel metal5 s -2936 20876 586860 21476 6 vssd1
port 742 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 743 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 744 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 707680 6 vccd2
port 745 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 707680 6 vccd2
port 746 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 707680 6 vccd2
port 747 nsew power bidirectional
rlabel metal4 s 437404 510000 438004 707680 6 vccd2
port 748 nsew power bidirectional
rlabel metal4 s 401404 510000 402004 707680 6 vccd2
port 749 nsew power bidirectional
rlabel metal4 s 365404 510000 366004 707680 6 vccd2
port 750 nsew power bidirectional
rlabel metal4 s 329404 510000 330004 707680 6 vccd2
port 751 nsew power bidirectional
rlabel metal4 s 293404 510000 294004 707680 6 vccd2
port 752 nsew power bidirectional
rlabel metal4 s 257404 510000 258004 707680 6 vccd2
port 753 nsew power bidirectional
rlabel metal4 s 221404 510000 222004 707680 6 vccd2
port 754 nsew power bidirectional
rlabel metal4 s 185404 510000 186004 707680 6 vccd2
port 755 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 707680 6 vccd2
port 756 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 707680 6 vccd2
port 757 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 707680 6 vccd2
port 758 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 707680 6 vccd2
port 759 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2
port 760 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 761 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 326000 6 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 326000 6 vccd2
port 764 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 326000 6 vccd2
port 765 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 326000 6 vccd2
port 766 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 326000 6 vccd2
port 767 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 326000 6 vccd2
port 768 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 326000 6 vccd2
port 769 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 326000 6 vccd2
port 770 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 771 nsew power bidirectional
rlabel metal5 s -4816 690476 588740 691076 6 vccd2
port 772 nsew power bidirectional
rlabel metal5 s -4816 654476 588740 655076 6 vccd2
port 773 nsew power bidirectional
rlabel metal5 s -4816 618476 588740 619076 6 vccd2
port 774 nsew power bidirectional
rlabel metal5 s -4816 582476 588740 583076 6 vccd2
port 775 nsew power bidirectional
rlabel metal5 s -4816 546476 588740 547076 6 vccd2
port 776 nsew power bidirectional
rlabel metal5 s -4816 510476 588740 511076 6 vccd2
port 777 nsew power bidirectional
rlabel metal5 s 440000 474476 588740 475076 6 vccd2
port 778 nsew power bidirectional
rlabel metal5 s -4816 474476 156000 475076 6 vccd2
port 779 nsew power bidirectional
rlabel metal5 s 440000 438476 588740 439076 6 vccd2
port 780 nsew power bidirectional
rlabel metal5 s -4816 438476 156000 439076 6 vccd2
port 781 nsew power bidirectional
rlabel metal5 s 440000 402476 588740 403076 6 vccd2
port 782 nsew power bidirectional
rlabel metal5 s -4816 402476 156000 403076 6 vccd2
port 783 nsew power bidirectional
rlabel metal5 s 440000 366476 588740 367076 6 vccd2
port 784 nsew power bidirectional
rlabel metal5 s -4816 366476 156000 367076 6 vccd2
port 785 nsew power bidirectional
rlabel metal5 s 440000 330476 588740 331076 6 vccd2
port 786 nsew power bidirectional
rlabel metal5 s -4816 330476 156000 331076 6 vccd2
port 787 nsew power bidirectional
rlabel metal5 s -4816 294476 588740 295076 6 vccd2
port 788 nsew power bidirectional
rlabel metal5 s -4816 258476 588740 259076 6 vccd2
port 789 nsew power bidirectional
rlabel metal5 s -4816 222476 588740 223076 6 vccd2
port 790 nsew power bidirectional
rlabel metal5 s -4816 186476 588740 187076 6 vccd2
port 791 nsew power bidirectional
rlabel metal5 s -4816 150476 588740 151076 6 vccd2
port 792 nsew power bidirectional
rlabel metal5 s -4816 114476 588740 115076 6 vccd2
port 793 nsew power bidirectional
rlabel metal5 s -4816 78476 588740 79076 6 vccd2
port 794 nsew power bidirectional
rlabel metal5 s -4816 42476 588740 43076 6 vccd2
port 795 nsew power bidirectional
rlabel metal5 s -4816 6476 588740 7076 6 vccd2
port 796 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 797 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 798 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 707680 6 vssd2
port 799 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 707680 6 vssd2
port 800 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 707680 6 vssd2
port 801 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 707680 6 vssd2
port 802 nsew ground bidirectional
rlabel metal4 s 419404 510000 420004 707680 6 vssd2
port 803 nsew ground bidirectional
rlabel metal4 s 383404 510000 384004 707680 6 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 347404 510000 348004 707680 6 vssd2
port 805 nsew ground bidirectional
rlabel metal4 s 311404 510000 312004 707680 6 vssd2
port 806 nsew ground bidirectional
rlabel metal4 s 275404 510000 276004 707680 6 vssd2
port 807 nsew ground bidirectional
rlabel metal4 s 239404 510000 240004 707680 6 vssd2
port 808 nsew ground bidirectional
rlabel metal4 s 203404 510000 204004 707680 6 vssd2
port 809 nsew ground bidirectional
rlabel metal4 s 167404 510000 168004 707680 6 vssd2
port 810 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 707680 6 vssd2
port 811 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 707680 6 vssd2
port 812 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 707680 6 vssd2
port 813 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 707680 6 vssd2
port 814 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 815 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 326000 6 vssd2
port 816 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 326000 6 vssd2
port 817 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 326000 6 vssd2
port 818 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 326000 6 vssd2
port 819 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 326000 6 vssd2
port 820 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 326000 6 vssd2
port 821 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 326000 6 vssd2
port 822 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 326000 6 vssd2
port 823 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 824 nsew ground bidirectional
rlabel metal5 s -4816 672476 588740 673076 6 vssd2
port 825 nsew ground bidirectional
rlabel metal5 s -4816 636476 588740 637076 6 vssd2
port 826 nsew ground bidirectional
rlabel metal5 s -4816 600476 588740 601076 6 vssd2
port 827 nsew ground bidirectional
rlabel metal5 s -4816 564476 588740 565076 6 vssd2
port 828 nsew ground bidirectional
rlabel metal5 s -4816 528476 588740 529076 6 vssd2
port 829 nsew ground bidirectional
rlabel metal5 s 440000 492476 588740 493076 6 vssd2
port 830 nsew ground bidirectional
rlabel metal5 s -4816 492476 156000 493076 6 vssd2
port 831 nsew ground bidirectional
rlabel metal5 s 440000 456476 588740 457076 6 vssd2
port 832 nsew ground bidirectional
rlabel metal5 s -4816 456476 156000 457076 6 vssd2
port 833 nsew ground bidirectional
rlabel metal5 s 440000 420476 588740 421076 6 vssd2
port 834 nsew ground bidirectional
rlabel metal5 s -4816 420476 156000 421076 6 vssd2
port 835 nsew ground bidirectional
rlabel metal5 s 440000 384476 588740 385076 6 vssd2
port 836 nsew ground bidirectional
rlabel metal5 s -4816 384476 156000 385076 6 vssd2
port 837 nsew ground bidirectional
rlabel metal5 s 440000 348476 588740 349076 6 vssd2
port 838 nsew ground bidirectional
rlabel metal5 s -4816 348476 156000 349076 6 vssd2
port 839 nsew ground bidirectional
rlabel metal5 s -4816 312476 588740 313076 6 vssd2
port 840 nsew ground bidirectional
rlabel metal5 s -4816 276476 588740 277076 6 vssd2
port 841 nsew ground bidirectional
rlabel metal5 s -4816 240476 588740 241076 6 vssd2
port 842 nsew ground bidirectional
rlabel metal5 s -4816 204476 588740 205076 6 vssd2
port 843 nsew ground bidirectional
rlabel metal5 s -4816 168476 588740 169076 6 vssd2
port 844 nsew ground bidirectional
rlabel metal5 s -4816 132476 588740 133076 6 vssd2
port 845 nsew ground bidirectional
rlabel metal5 s -4816 96476 588740 97076 6 vssd2
port 846 nsew ground bidirectional
rlabel metal5 s -4816 60476 588740 61076 6 vssd2
port 847 nsew ground bidirectional
rlabel metal5 s -4816 24476 588740 25076 6 vssd2
port 848 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 849 nsew ground bidirectional
rlabel metal4 s 549004 -5624 549604 709560 6 vdda1
port 850 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 709560 6 vdda1
port 851 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 709560 6 vdda1
port 852 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 709560 6 vdda1
port 853 nsew power bidirectional
rlabel metal4 s 405004 510000 405604 709560 6 vdda1
port 854 nsew power bidirectional
rlabel metal4 s 369004 510000 369604 709560 6 vdda1
port 855 nsew power bidirectional
rlabel metal4 s 333004 510000 333604 709560 6 vdda1
port 856 nsew power bidirectional
rlabel metal4 s 297004 510000 297604 709560 6 vdda1
port 857 nsew power bidirectional
rlabel metal4 s 261004 510000 261604 709560 6 vdda1
port 858 nsew power bidirectional
rlabel metal4 s 225004 510000 225604 709560 6 vdda1
port 859 nsew power bidirectional
rlabel metal4 s 189004 510000 189604 709560 6 vdda1
port 860 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 709560 6 vdda1
port 861 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 709560 6 vdda1
port 862 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 709560 6 vdda1
port 863 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 709560 6 vdda1
port 864 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1
port 865 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 866 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 867 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 326000 6 vdda1
port 868 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 326000 6 vdda1
port 869 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 326000 6 vdda1
port 870 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 326000 6 vdda1
port 871 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 326000 6 vdda1
port 872 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 326000 6 vdda1
port 873 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 326000 6 vdda1
port 874 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 875 nsew power bidirectional
rlabel metal5 s -6696 694076 590620 694676 6 vdda1
port 876 nsew power bidirectional
rlabel metal5 s -6696 658076 590620 658676 6 vdda1
port 877 nsew power bidirectional
rlabel metal5 s -6696 622076 590620 622676 6 vdda1
port 878 nsew power bidirectional
rlabel metal5 s -6696 586076 590620 586676 6 vdda1
port 879 nsew power bidirectional
rlabel metal5 s -6696 550076 590620 550676 6 vdda1
port 880 nsew power bidirectional
rlabel metal5 s -6696 514076 590620 514676 6 vdda1
port 881 nsew power bidirectional
rlabel metal5 s 440000 478076 590620 478676 6 vdda1
port 882 nsew power bidirectional
rlabel metal5 s -6696 478076 156000 478676 6 vdda1
port 883 nsew power bidirectional
rlabel metal5 s 440000 442076 590620 442676 6 vdda1
port 884 nsew power bidirectional
rlabel metal5 s -6696 442076 156000 442676 6 vdda1
port 885 nsew power bidirectional
rlabel metal5 s 440000 406076 590620 406676 6 vdda1
port 886 nsew power bidirectional
rlabel metal5 s -6696 406076 156000 406676 6 vdda1
port 887 nsew power bidirectional
rlabel metal5 s 440000 370076 590620 370676 6 vdda1
port 888 nsew power bidirectional
rlabel metal5 s -6696 370076 156000 370676 6 vdda1
port 889 nsew power bidirectional
rlabel metal5 s 440000 334076 590620 334676 6 vdda1
port 890 nsew power bidirectional
rlabel metal5 s -6696 334076 156000 334676 6 vdda1
port 891 nsew power bidirectional
rlabel metal5 s -6696 298076 590620 298676 6 vdda1
port 892 nsew power bidirectional
rlabel metal5 s -6696 262076 590620 262676 6 vdda1
port 893 nsew power bidirectional
rlabel metal5 s -6696 226076 590620 226676 6 vdda1
port 894 nsew power bidirectional
rlabel metal5 s -6696 190076 590620 190676 6 vdda1
port 895 nsew power bidirectional
rlabel metal5 s -6696 154076 590620 154676 6 vdda1
port 896 nsew power bidirectional
rlabel metal5 s -6696 118076 590620 118676 6 vdda1
port 897 nsew power bidirectional
rlabel metal5 s -6696 82076 590620 82676 6 vdda1
port 898 nsew power bidirectional
rlabel metal5 s -6696 46076 590620 46676 6 vdda1
port 899 nsew power bidirectional
rlabel metal5 s -6696 10076 590620 10676 6 vdda1
port 900 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 901 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 902 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 709560 6 vssa1
port 903 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 709560 6 vssa1
port 904 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 709560 6 vssa1
port 905 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 709560 6 vssa1
port 906 nsew ground bidirectional
rlabel metal4 s 423004 510000 423604 709560 6 vssa1
port 907 nsew ground bidirectional
rlabel metal4 s 387004 510000 387604 709560 6 vssa1
port 908 nsew ground bidirectional
rlabel metal4 s 351004 510000 351604 709560 6 vssa1
port 909 nsew ground bidirectional
rlabel metal4 s 315004 510000 315604 709560 6 vssa1
port 910 nsew ground bidirectional
rlabel metal4 s 279004 510000 279604 709560 6 vssa1
port 911 nsew ground bidirectional
rlabel metal4 s 243004 510000 243604 709560 6 vssa1
port 912 nsew ground bidirectional
rlabel metal4 s 207004 510000 207604 709560 6 vssa1
port 913 nsew ground bidirectional
rlabel metal4 s 171004 510000 171604 709560 6 vssa1
port 914 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 709560 6 vssa1
port 915 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 709560 6 vssa1
port 916 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 709560 6 vssa1
port 917 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 709560 6 vssa1
port 918 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 919 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 326000 6 vssa1
port 920 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 326000 6 vssa1
port 921 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 326000 6 vssa1
port 922 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 326000 6 vssa1
port 923 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 326000 6 vssa1
port 924 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 326000 6 vssa1
port 925 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 326000 6 vssa1
port 926 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 326000 6 vssa1
port 927 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 928 nsew ground bidirectional
rlabel metal5 s -6696 676076 590620 676676 6 vssa1
port 929 nsew ground bidirectional
rlabel metal5 s -6696 640076 590620 640676 6 vssa1
port 930 nsew ground bidirectional
rlabel metal5 s -6696 604076 590620 604676 6 vssa1
port 931 nsew ground bidirectional
rlabel metal5 s -6696 568076 590620 568676 6 vssa1
port 932 nsew ground bidirectional
rlabel metal5 s -6696 532076 590620 532676 6 vssa1
port 933 nsew ground bidirectional
rlabel metal5 s 440000 496076 590620 496676 6 vssa1
port 934 nsew ground bidirectional
rlabel metal5 s -6696 496076 156000 496676 6 vssa1
port 935 nsew ground bidirectional
rlabel metal5 s 440000 460076 590620 460676 6 vssa1
port 936 nsew ground bidirectional
rlabel metal5 s -6696 460076 156000 460676 6 vssa1
port 937 nsew ground bidirectional
rlabel metal5 s 440000 424076 590620 424676 6 vssa1
port 938 nsew ground bidirectional
rlabel metal5 s -6696 424076 156000 424676 6 vssa1
port 939 nsew ground bidirectional
rlabel metal5 s 440000 388076 590620 388676 6 vssa1
port 940 nsew ground bidirectional
rlabel metal5 s -6696 388076 156000 388676 6 vssa1
port 941 nsew ground bidirectional
rlabel metal5 s 440000 352076 590620 352676 6 vssa1
port 942 nsew ground bidirectional
rlabel metal5 s -6696 352076 156000 352676 6 vssa1
port 943 nsew ground bidirectional
rlabel metal5 s -6696 316076 590620 316676 6 vssa1
port 944 nsew ground bidirectional
rlabel metal5 s -6696 280076 590620 280676 6 vssa1
port 945 nsew ground bidirectional
rlabel metal5 s -6696 244076 590620 244676 6 vssa1
port 946 nsew ground bidirectional
rlabel metal5 s -6696 208076 590620 208676 6 vssa1
port 947 nsew ground bidirectional
rlabel metal5 s -6696 172076 590620 172676 6 vssa1
port 948 nsew ground bidirectional
rlabel metal5 s -6696 136076 590620 136676 6 vssa1
port 949 nsew ground bidirectional
rlabel metal5 s -6696 100076 590620 100676 6 vssa1
port 950 nsew ground bidirectional
rlabel metal5 s -6696 64076 590620 64676 6 vssa1
port 951 nsew ground bidirectional
rlabel metal5 s -6696 28076 590620 28676 6 vssa1
port 952 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 953 nsew ground bidirectional
rlabel metal4 s 552604 -7504 553204 711440 6 vdda2
port 954 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 711440 6 vdda2
port 955 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 711440 6 vdda2
port 956 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 711440 6 vdda2
port 957 nsew power bidirectional
rlabel metal4 s 408604 510000 409204 711440 6 vdda2
port 958 nsew power bidirectional
rlabel metal4 s 372604 510000 373204 711440 6 vdda2
port 959 nsew power bidirectional
rlabel metal4 s 336604 510000 337204 711440 6 vdda2
port 960 nsew power bidirectional
rlabel metal4 s 300604 510000 301204 711440 6 vdda2
port 961 nsew power bidirectional
rlabel metal4 s 264604 510000 265204 711440 6 vdda2
port 962 nsew power bidirectional
rlabel metal4 s 228604 510000 229204 711440 6 vdda2
port 963 nsew power bidirectional
rlabel metal4 s 192604 510000 193204 711440 6 vdda2
port 964 nsew power bidirectional
rlabel metal4 s 156604 510000 157204 711440 6 vdda2
port 965 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 711440 6 vdda2
port 966 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 711440 6 vdda2
port 967 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 711440 6 vdda2
port 968 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2
port 969 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 970 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 971 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 326000 6 vdda2
port 972 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 326000 6 vdda2
port 973 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 326000 6 vdda2
port 974 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 326000 6 vdda2
port 975 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 326000 6 vdda2
port 976 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 326000 6 vdda2
port 977 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 326000 6 vdda2
port 978 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 326000 6 vdda2
port 979 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 980 nsew power bidirectional
rlabel metal5 s -8576 697676 592500 698276 6 vdda2
port 981 nsew power bidirectional
rlabel metal5 s -8576 661676 592500 662276 6 vdda2
port 982 nsew power bidirectional
rlabel metal5 s -8576 625676 592500 626276 6 vdda2
port 983 nsew power bidirectional
rlabel metal5 s -8576 589676 592500 590276 6 vdda2
port 984 nsew power bidirectional
rlabel metal5 s -8576 553676 592500 554276 6 vdda2
port 985 nsew power bidirectional
rlabel metal5 s -8576 517676 592500 518276 6 vdda2
port 986 nsew power bidirectional
rlabel metal5 s 440000 481676 592500 482276 6 vdda2
port 987 nsew power bidirectional
rlabel metal5 s -8576 481676 156000 482276 6 vdda2
port 988 nsew power bidirectional
rlabel metal5 s 440000 445676 592500 446276 6 vdda2
port 989 nsew power bidirectional
rlabel metal5 s -8576 445676 156000 446276 6 vdda2
port 990 nsew power bidirectional
rlabel metal5 s 440000 409676 592500 410276 6 vdda2
port 991 nsew power bidirectional
rlabel metal5 s -8576 409676 156000 410276 6 vdda2
port 992 nsew power bidirectional
rlabel metal5 s 440000 373676 592500 374276 6 vdda2
port 993 nsew power bidirectional
rlabel metal5 s -8576 373676 156000 374276 6 vdda2
port 994 nsew power bidirectional
rlabel metal5 s 440000 337676 592500 338276 6 vdda2
port 995 nsew power bidirectional
rlabel metal5 s -8576 337676 156000 338276 6 vdda2
port 996 nsew power bidirectional
rlabel metal5 s -8576 301676 592500 302276 6 vdda2
port 997 nsew power bidirectional
rlabel metal5 s -8576 265676 592500 266276 6 vdda2
port 998 nsew power bidirectional
rlabel metal5 s -8576 229676 592500 230276 6 vdda2
port 999 nsew power bidirectional
rlabel metal5 s -8576 193676 592500 194276 6 vdda2
port 1000 nsew power bidirectional
rlabel metal5 s -8576 157676 592500 158276 6 vdda2
port 1001 nsew power bidirectional
rlabel metal5 s -8576 121676 592500 122276 6 vdda2
port 1002 nsew power bidirectional
rlabel metal5 s -8576 85676 592500 86276 6 vdda2
port 1003 nsew power bidirectional
rlabel metal5 s -8576 49676 592500 50276 6 vdda2
port 1004 nsew power bidirectional
rlabel metal5 s -8576 13676 592500 14276 6 vdda2
port 1005 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1006 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1007 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 711440 6 vssa2
port 1008 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 711440 6 vssa2
port 1009 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 711440 6 vssa2
port 1010 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 711440 6 vssa2
port 1011 nsew ground bidirectional
rlabel metal4 s 426604 510000 427204 711440 6 vssa2
port 1012 nsew ground bidirectional
rlabel metal4 s 390604 510000 391204 711440 6 vssa2
port 1013 nsew ground bidirectional
rlabel metal4 s 354604 510000 355204 711440 6 vssa2
port 1014 nsew ground bidirectional
rlabel metal4 s 318604 510000 319204 711440 6 vssa2
port 1015 nsew ground bidirectional
rlabel metal4 s 282604 510000 283204 711440 6 vssa2
port 1016 nsew ground bidirectional
rlabel metal4 s 246604 510000 247204 711440 6 vssa2
port 1017 nsew ground bidirectional
rlabel metal4 s 210604 510000 211204 711440 6 vssa2
port 1018 nsew ground bidirectional
rlabel metal4 s 174604 510000 175204 711440 6 vssa2
port 1019 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 711440 6 vssa2
port 1020 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 711440 6 vssa2
port 1021 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 711440 6 vssa2
port 1022 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 711440 6 vssa2
port 1023 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1024 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 326000 6 vssa2
port 1025 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 326000 6 vssa2
port 1026 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 326000 6 vssa2
port 1027 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 326000 6 vssa2
port 1028 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 326000 6 vssa2
port 1029 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 326000 6 vssa2
port 1030 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 326000 6 vssa2
port 1031 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 326000 6 vssa2
port 1032 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1033 nsew ground bidirectional
rlabel metal5 s -8576 679676 592500 680276 6 vssa2
port 1034 nsew ground bidirectional
rlabel metal5 s -8576 643676 592500 644276 6 vssa2
port 1035 nsew ground bidirectional
rlabel metal5 s -8576 607676 592500 608276 6 vssa2
port 1036 nsew ground bidirectional
rlabel metal5 s -8576 571676 592500 572276 6 vssa2
port 1037 nsew ground bidirectional
rlabel metal5 s -8576 535676 592500 536276 6 vssa2
port 1038 nsew ground bidirectional
rlabel metal5 s 440000 499676 592500 500276 6 vssa2
port 1039 nsew ground bidirectional
rlabel metal5 s -8576 499676 156000 500276 6 vssa2
port 1040 nsew ground bidirectional
rlabel metal5 s 440000 463676 592500 464276 6 vssa2
port 1041 nsew ground bidirectional
rlabel metal5 s -8576 463676 156000 464276 6 vssa2
port 1042 nsew ground bidirectional
rlabel metal5 s 440000 427676 592500 428276 6 vssa2
port 1043 nsew ground bidirectional
rlabel metal5 s -8576 427676 156000 428276 6 vssa2
port 1044 nsew ground bidirectional
rlabel metal5 s 440000 391676 592500 392276 6 vssa2
port 1045 nsew ground bidirectional
rlabel metal5 s -8576 391676 156000 392276 6 vssa2
port 1046 nsew ground bidirectional
rlabel metal5 s 440000 355676 592500 356276 6 vssa2
port 1047 nsew ground bidirectional
rlabel metal5 s -8576 355676 156000 356276 6 vssa2
port 1048 nsew ground bidirectional
rlabel metal5 s -8576 319676 592500 320276 6 vssa2
port 1049 nsew ground bidirectional
rlabel metal5 s -8576 283676 592500 284276 6 vssa2
port 1050 nsew ground bidirectional
rlabel metal5 s -8576 247676 592500 248276 6 vssa2
port 1051 nsew ground bidirectional
rlabel metal5 s -8576 211676 592500 212276 6 vssa2
port 1052 nsew ground bidirectional
rlabel metal5 s -8576 175676 592500 176276 6 vssa2
port 1053 nsew ground bidirectional
rlabel metal5 s -8576 139676 592500 140276 6 vssa2
port 1054 nsew ground bidirectional
rlabel metal5 s -8576 103676 592500 104276 6 vssa2
port 1055 nsew ground bidirectional
rlabel metal5 s -8576 67676 592500 68276 6 vssa2
port 1056 nsew ground bidirectional
rlabel metal5 s -8576 31676 592500 32276 6 vssa2
port 1057 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1058 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
