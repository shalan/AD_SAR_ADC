VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ACMP
  CLASS BLOCK ;
  FOREIGN ACMP ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.920 BY 100.400 ;
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.680 49.610 50.680 50.730 ;
    END
  END INN
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.680 19.710 50.680 20.830 ;
    END
  END INP
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.680 79.510 50.680 80.630 ;
    END
  END Q
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.680 79.510 14.680 80.630 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.680 49.610 14.680 50.730 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.680 19.710 14.680 20.830 ;
    END
  END clk
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.700 90.700 55.220 94.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.700 5.700 55.220 9.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 39.285 0.000 41.385 100.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.630 0.000 31.730 100.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.975 0.000 22.075 100.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 51.220 5.700 55.220 94.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.700 5.700 9.700 94.700 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.400 60.920 100.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 60.920 4.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 56.920 0.000 60.920 100.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.455 0.000 36.555 100.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.805 0.000 26.905 100.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 4.000 100.400 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 16.200 16.115 44.720 84.285 ;
      LAYER met1 ;
        RECT 15.810 15.960 46.030 84.440 ;
      LAYER met2 ;
        RECT 14.680 80.910 46.680 84.440 ;
        RECT 14.960 79.230 46.400 80.910 ;
        RECT 14.680 51.010 46.680 79.230 ;
        RECT 14.960 49.330 46.400 51.010 ;
        RECT 14.680 21.110 46.680 49.330 ;
        RECT 14.960 19.430 46.400 21.110 ;
        RECT 14.680 15.960 46.680 19.430 ;
      LAYER met3 ;
        RECT 19.975 16.035 41.380 84.365 ;
      LAYER met4 ;
        RECT 27.305 0.000 29.230 100.400 ;
        RECT 32.130 0.000 34.055 100.400 ;
        RECT 36.955 0.000 38.885 100.400 ;
  END
END ACMP
END LIBRARY

