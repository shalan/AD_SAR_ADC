magic
tech sky130A
magscale 1 2
timestamp 1626378704
<< obsli1 >>
rect 3240 3223 8944 6521
<< obsm1 >>
rect 3162 3192 9206 6552
<< metal2 >>
rect 2136 7622 2936 7846
rect 9336 7622 10136 7846
rect 2136 4954 2936 5178
rect 9336 4954 10136 5178
rect 2136 2286 2936 2510
rect 9336 2286 10136 2510
<< obsm2 >>
rect 2992 7566 9280 7748
rect 2936 5234 9336 7566
rect 2992 4898 9280 5234
rect 2936 2566 9336 4898
rect 2992 2384 9280 2566
<< metal3 >>
rect 0 8944 12184 9744
rect 1140 7804 11044 8604
rect 1140 1140 11044 1940
rect 0 0 12184 800
<< obsm3 >>
rect 3995 3207 8276 6537
<< metal4 >>
rect 0 0 800 9744
rect 1140 1140 1940 8604
rect 3995 0 4415 9744
rect 4961 0 5381 9744
rect 5926 0 6346 9744
rect 6891 0 7311 9744
rect 7857 0 8277 9744
rect 10244 1140 11044 8604
rect 11384 0 12184 9744
<< obsm4 >>
rect 5461 0 5846 9744
rect 6426 0 6811 9744
rect 7391 0 7777 9744
<< labels >>
rlabel metal2 s 9336 4954 10136 5178 6 INN
port 1 nsew signal input
rlabel metal2 s 9336 2286 10136 2510 6 INP
port 2 nsew signal input
rlabel metal2 s 9336 7622 10136 7846 6 Q
port 3 nsew signal output
rlabel metal2 s 2136 7622 2936 7846 6 VDD
port 4 nsew signal input
rlabel metal2 s 2136 4954 2936 5178 6 VSS
port 5 nsew signal input
rlabel metal2 s 2136 2286 2936 2510 6 clk
port 6 nsew signal input
rlabel metal3 s 1140 7804 11044 8604 6 vccd2
port 7 nsew power bidirectional
rlabel metal3 s 1140 1140 11044 1940 6 vccd2
port 8 nsew power bidirectional
rlabel metal4 s 7857 0 8277 9744 6 vccd2
port 9 nsew power bidirectional
rlabel metal4 s 5926 0 6346 9744 6 vccd2
port 10 nsew power bidirectional
rlabel metal4 s 3995 0 4415 9744 6 vccd2
port 11 nsew power bidirectional
rlabel metal4 s 10244 1140 11044 8604 6 vccd2
port 12 nsew power bidirectional
rlabel metal4 s 1140 1140 1940 8604 6 vccd2
port 13 nsew power bidirectional
rlabel metal3 s 0 8944 12184 9744 6 vssd2
port 14 nsew ground bidirectional
rlabel metal3 s 0 0 12184 800 6 vssd2
port 15 nsew ground bidirectional
rlabel metal4 s 11384 0 12184 9744 6 vssd2
port 16 nsew ground bidirectional
rlabel metal4 s 6891 0 7311 9744 6 vssd2
port 17 nsew ground bidirectional
rlabel metal4 s 4961 0 5381 9744 6 vssd2
port 18 nsew ground bidirectional
rlabel metal4 s 0 0 800 9744 6 vssd2
port 19 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 12184 9744
string LEFview TRUE
string GDS_FILE /project/openlane/ACMP/runs/ACMP/results/magic/ACMP.gds
string GDS_END 199476
string GDS_START 52858
<< end >>

