magic
tech sky130A
magscale 1 2
timestamp 1626642735
<< viali >>
rect 8053 16109 8087 16143
rect 3545 15973 3579 16007
rect 4189 15973 4223 16007
rect 7869 15973 7903 16007
rect 3729 15837 3763 15871
rect 7501 11689 7535 11723
rect 7685 11689 7719 11723
rect 7409 11621 7443 11655
rect 7409 11485 7443 11519
rect 7869 11281 7903 11315
rect 6857 11145 6891 11179
rect 7041 11145 7075 11179
rect 7133 11145 7167 11179
rect 7409 11145 7443 11179
rect 7869 11145 7903 11179
rect 8145 11077 8179 11111
rect 7961 11009 7995 11043
rect 6397 10941 6431 10975
rect 7225 10941 7259 10975
rect 7317 10941 7351 10975
rect 7133 10737 7167 10771
rect 7133 10533 7167 10567
rect 7225 10533 7259 10567
rect 7593 10533 7627 10567
rect 7409 10465 7443 10499
rect 7501 10465 7535 10499
rect 6627 10193 6661 10227
rect 7317 10193 7351 10227
rect 7501 10125 7535 10159
rect 3545 10057 3579 10091
rect 4189 10057 4223 10091
rect 6556 10057 6590 10091
rect 7133 10057 7167 10091
rect 7225 10057 7259 10091
rect 7409 10057 7443 10091
rect 7593 10057 7627 10091
rect 3729 9853 3763 9887
rect 6857 9649 6891 9683
rect 8007 9649 8041 9683
rect 7317 9513 7351 9547
rect 6857 9445 6891 9479
rect 7041 9445 7075 9479
rect 7133 9445 7167 9479
rect 7409 9445 7443 9479
rect 7904 9445 7938 9479
rect 6397 9309 6431 9343
rect 6995 9105 7029 9139
rect 6892 8969 6926 9003
rect 7593 8969 7627 9003
rect 8237 8969 8271 9003
rect 8053 8833 8087 8867
rect 6397 8765 6431 8799
rect 8053 4753 8087 4787
rect 7593 4617 7627 4651
rect 8237 4617 8271 4651
<< metal1 >>
rect 3240 16866 8944 16888
rect 3240 16814 4984 16866
rect 5036 16814 5048 16866
rect 5100 16814 5112 16866
rect 5164 16814 5176 16866
rect 5228 16814 5240 16866
rect 5292 16814 5304 16866
rect 5356 16814 6915 16866
rect 6967 16814 6979 16866
rect 7031 16814 7043 16866
rect 7095 16814 7107 16866
rect 7159 16814 7171 16866
rect 7223 16814 7235 16866
rect 7287 16814 8944 16866
rect 3240 16792 8944 16814
rect 3240 16322 8944 16344
rect 3240 16270 4019 16322
rect 4071 16270 4083 16322
rect 4135 16270 4147 16322
rect 4199 16270 4211 16322
rect 4263 16270 4275 16322
rect 4327 16270 4339 16322
rect 4391 16270 5950 16322
rect 6002 16270 6014 16322
rect 6066 16270 6078 16322
rect 6130 16270 6142 16322
rect 6194 16270 6206 16322
rect 6258 16270 6270 16322
rect 6322 16270 7880 16322
rect 7932 16270 7944 16322
rect 7996 16270 8008 16322
rect 8060 16270 8072 16322
rect 8124 16270 8136 16322
rect 8188 16270 8200 16322
rect 8252 16270 8944 16322
rect 3240 16248 8944 16270
rect 8041 16143 8099 16149
rect 8041 16109 8053 16143
rect 8087 16140 8099 16143
rect 9142 16140 9148 16152
rect 8087 16112 9148 16140
rect 8087 16109 8099 16112
rect 8041 16103 8099 16109
rect 9142 16100 9148 16112
rect 9200 16100 9206 16152
rect 3162 15964 3168 16016
rect 3220 16004 3226 16016
rect 3533 16007 3591 16013
rect 3533 16004 3545 16007
rect 3220 15976 3545 16004
rect 3220 15964 3226 15976
rect 3533 15973 3545 15976
rect 3579 16004 3591 16007
rect 4177 16007 4235 16013
rect 4177 16004 4189 16007
rect 3579 15976 4189 16004
rect 3579 15973 3591 15976
rect 3533 15967 3591 15973
rect 4177 15973 4189 15976
rect 4223 15973 4235 16007
rect 4177 15967 4235 15973
rect 7670 15964 7676 16016
rect 7728 16004 7734 16016
rect 7857 16007 7915 16013
rect 7857 16004 7869 16007
rect 7728 15976 7869 16004
rect 7728 15964 7734 15976
rect 7857 15973 7869 15976
rect 7903 15973 7915 16007
rect 7857 15967 7915 15973
rect 3717 15871 3775 15877
rect 3717 15837 3729 15871
rect 3763 15868 3775 15871
rect 6750 15868 6756 15880
rect 3763 15840 6756 15868
rect 3763 15837 3775 15840
rect 3717 15831 3775 15837
rect 6750 15828 6756 15840
rect 6808 15828 6814 15880
rect 3240 15778 8944 15800
rect 3240 15726 4984 15778
rect 5036 15726 5048 15778
rect 5100 15726 5112 15778
rect 5164 15726 5176 15778
rect 5228 15726 5240 15778
rect 5292 15726 5304 15778
rect 5356 15726 6915 15778
rect 6967 15726 6979 15778
rect 7031 15726 7043 15778
rect 7095 15726 7107 15778
rect 7159 15726 7171 15778
rect 7223 15726 7235 15778
rect 7287 15726 8944 15778
rect 3240 15704 8944 15726
rect 3240 15234 8944 15256
rect 3240 15182 4019 15234
rect 4071 15182 4083 15234
rect 4135 15182 4147 15234
rect 4199 15182 4211 15234
rect 4263 15182 4275 15234
rect 4327 15182 4339 15234
rect 4391 15182 5950 15234
rect 6002 15182 6014 15234
rect 6066 15182 6078 15234
rect 6130 15182 6142 15234
rect 6194 15182 6206 15234
rect 6258 15182 6270 15234
rect 6322 15182 7880 15234
rect 7932 15182 7944 15234
rect 7996 15182 8008 15234
rect 8060 15182 8072 15234
rect 8124 15182 8136 15234
rect 8188 15182 8200 15234
rect 8252 15182 8944 15234
rect 3240 15160 8944 15182
rect 3240 14690 8944 14712
rect 3240 14638 4984 14690
rect 5036 14638 5048 14690
rect 5100 14638 5112 14690
rect 5164 14638 5176 14690
rect 5228 14638 5240 14690
rect 5292 14638 5304 14690
rect 5356 14638 6915 14690
rect 6967 14638 6979 14690
rect 7031 14638 7043 14690
rect 7095 14638 7107 14690
rect 7159 14638 7171 14690
rect 7223 14638 7235 14690
rect 7287 14638 8944 14690
rect 3240 14616 8944 14638
rect 3240 14146 8944 14168
rect 3240 14094 4019 14146
rect 4071 14094 4083 14146
rect 4135 14094 4147 14146
rect 4199 14094 4211 14146
rect 4263 14094 4275 14146
rect 4327 14094 4339 14146
rect 4391 14094 5950 14146
rect 6002 14094 6014 14146
rect 6066 14094 6078 14146
rect 6130 14094 6142 14146
rect 6194 14094 6206 14146
rect 6258 14094 6270 14146
rect 6322 14094 7880 14146
rect 7932 14094 7944 14146
rect 7996 14094 8008 14146
rect 8060 14094 8072 14146
rect 8124 14094 8136 14146
rect 8188 14094 8200 14146
rect 8252 14094 8944 14146
rect 3240 14072 8944 14094
rect 3240 13602 8944 13624
rect 3240 13550 4984 13602
rect 5036 13550 5048 13602
rect 5100 13550 5112 13602
rect 5164 13550 5176 13602
rect 5228 13550 5240 13602
rect 5292 13550 5304 13602
rect 5356 13550 6915 13602
rect 6967 13550 6979 13602
rect 7031 13550 7043 13602
rect 7095 13550 7107 13602
rect 7159 13550 7171 13602
rect 7223 13550 7235 13602
rect 7287 13550 8944 13602
rect 3240 13528 8944 13550
rect 3240 13058 8944 13080
rect 3240 13006 4019 13058
rect 4071 13006 4083 13058
rect 4135 13006 4147 13058
rect 4199 13006 4211 13058
rect 4263 13006 4275 13058
rect 4327 13006 4339 13058
rect 4391 13006 5950 13058
rect 6002 13006 6014 13058
rect 6066 13006 6078 13058
rect 6130 13006 6142 13058
rect 6194 13006 6206 13058
rect 6258 13006 6270 13058
rect 6322 13006 7880 13058
rect 7932 13006 7944 13058
rect 7996 13006 8008 13058
rect 8060 13006 8072 13058
rect 8124 13006 8136 13058
rect 8188 13006 8200 13058
rect 8252 13006 8944 13058
rect 3240 12984 8944 13006
rect 3240 12514 8944 12536
rect 3240 12462 4984 12514
rect 5036 12462 5048 12514
rect 5100 12462 5112 12514
rect 5164 12462 5176 12514
rect 5228 12462 5240 12514
rect 5292 12462 5304 12514
rect 5356 12462 6915 12514
rect 6967 12462 6979 12514
rect 7031 12462 7043 12514
rect 7095 12462 7107 12514
rect 7159 12462 7171 12514
rect 7223 12462 7235 12514
rect 7287 12462 8944 12514
rect 3240 12440 8944 12462
rect 3240 11970 8944 11992
rect 3240 11918 4019 11970
rect 4071 11918 4083 11970
rect 4135 11918 4147 11970
rect 4199 11918 4211 11970
rect 4263 11918 4275 11970
rect 4327 11918 4339 11970
rect 4391 11918 5950 11970
rect 6002 11918 6014 11970
rect 6066 11918 6078 11970
rect 6130 11918 6142 11970
rect 6194 11918 6206 11970
rect 6258 11918 6270 11970
rect 6322 11918 7880 11970
rect 7932 11918 7944 11970
rect 7996 11918 8008 11970
rect 8060 11918 8072 11970
rect 8124 11918 8136 11970
rect 8188 11918 8200 11970
rect 8252 11918 8944 11970
rect 3240 11896 8944 11918
rect 6658 11680 6664 11732
rect 6716 11720 6722 11732
rect 7489 11723 7547 11729
rect 7489 11720 7501 11723
rect 6716 11692 7501 11720
rect 6716 11680 6722 11692
rect 7489 11689 7501 11692
rect 7535 11689 7547 11723
rect 7670 11720 7676 11732
rect 7631 11692 7676 11720
rect 7489 11683 7547 11689
rect 7670 11680 7676 11692
rect 7728 11680 7734 11732
rect 7394 11652 7400 11664
rect 7355 11624 7400 11652
rect 7394 11612 7400 11624
rect 7452 11612 7458 11664
rect 7397 11519 7455 11525
rect 7397 11485 7409 11519
rect 7443 11516 7455 11519
rect 7854 11516 7860 11528
rect 7443 11488 7860 11516
rect 7443 11485 7455 11488
rect 7397 11479 7455 11485
rect 7854 11476 7860 11488
rect 7912 11476 7918 11528
rect 3240 11426 8944 11448
rect 3240 11374 4984 11426
rect 5036 11374 5048 11426
rect 5100 11374 5112 11426
rect 5164 11374 5176 11426
rect 5228 11374 5240 11426
rect 5292 11374 5304 11426
rect 5356 11374 6915 11426
rect 6967 11374 6979 11426
rect 7031 11374 7043 11426
rect 7095 11374 7107 11426
rect 7159 11374 7171 11426
rect 7223 11374 7235 11426
rect 7287 11374 8944 11426
rect 3240 11352 8944 11374
rect 7670 11272 7676 11324
rect 7728 11312 7734 11324
rect 7857 11315 7915 11321
rect 7857 11312 7869 11315
rect 7728 11284 7869 11312
rect 7728 11272 7734 11284
rect 7857 11281 7869 11284
rect 7903 11281 7915 11315
rect 7857 11275 7915 11281
rect 6382 11204 6388 11256
rect 6440 11244 6446 11256
rect 6440 11216 7072 11244
rect 6440 11204 6446 11216
rect 6566 11136 6572 11188
rect 6624 11176 6630 11188
rect 7044 11185 7072 11216
rect 6845 11179 6903 11185
rect 6845 11176 6857 11179
rect 6624 11148 6857 11176
rect 6624 11136 6630 11148
rect 6845 11145 6857 11148
rect 6891 11145 6903 11179
rect 6845 11139 6903 11145
rect 7029 11179 7087 11185
rect 7029 11145 7041 11179
rect 7075 11145 7087 11179
rect 7029 11139 7087 11145
rect 7121 11179 7179 11185
rect 7121 11145 7133 11179
rect 7167 11145 7179 11179
rect 7121 11139 7179 11145
rect 6474 11068 6480 11120
rect 6532 11108 6538 11120
rect 7136 11108 7164 11139
rect 7302 11136 7308 11188
rect 7360 11176 7366 11188
rect 7397 11179 7455 11185
rect 7397 11176 7409 11179
rect 7360 11148 7409 11176
rect 7360 11136 7366 11148
rect 7397 11145 7409 11148
rect 7443 11145 7455 11179
rect 7854 11176 7860 11188
rect 7815 11148 7860 11176
rect 7397 11139 7455 11145
rect 7854 11136 7860 11148
rect 7912 11136 7918 11188
rect 6532 11080 7164 11108
rect 8133 11111 8191 11117
rect 6532 11068 6538 11080
rect 8133 11077 8145 11111
rect 8179 11108 8191 11111
rect 8314 11108 8320 11120
rect 8179 11080 8320 11108
rect 8179 11077 8191 11080
rect 8133 11071 8191 11077
rect 8314 11068 8320 11080
rect 8372 11068 8378 11120
rect 7118 11000 7124 11052
rect 7176 11040 7182 11052
rect 7578 11040 7584 11052
rect 7176 11012 7584 11040
rect 7176 11000 7182 11012
rect 7578 11000 7584 11012
rect 7636 11040 7642 11052
rect 7949 11043 8007 11049
rect 7949 11040 7961 11043
rect 7636 11012 7961 11040
rect 7636 11000 7642 11012
rect 7949 11009 7961 11012
rect 7995 11009 8007 11043
rect 7949 11003 8007 11009
rect 6382 10972 6388 10984
rect 6343 10944 6388 10972
rect 6382 10932 6388 10944
rect 6440 10932 6446 10984
rect 7026 10932 7032 10984
rect 7084 10972 7090 10984
rect 7213 10975 7271 10981
rect 7213 10972 7225 10975
rect 7084 10944 7225 10972
rect 7084 10932 7090 10944
rect 7213 10941 7225 10944
rect 7259 10941 7271 10975
rect 7213 10935 7271 10941
rect 7302 10932 7308 10984
rect 7360 10972 7366 10984
rect 7360 10944 7405 10972
rect 7360 10932 7366 10944
rect 3240 10882 8944 10904
rect 3240 10830 4019 10882
rect 4071 10830 4083 10882
rect 4135 10830 4147 10882
rect 4199 10830 4211 10882
rect 4263 10830 4275 10882
rect 4327 10830 4339 10882
rect 4391 10830 5950 10882
rect 6002 10830 6014 10882
rect 6066 10830 6078 10882
rect 6130 10830 6142 10882
rect 6194 10830 6206 10882
rect 6258 10830 6270 10882
rect 6322 10830 7880 10882
rect 7932 10830 7944 10882
rect 7996 10830 8008 10882
rect 8060 10830 8072 10882
rect 8124 10830 8136 10882
rect 8188 10830 8200 10882
rect 8252 10830 8944 10882
rect 3240 10808 8944 10830
rect 7121 10771 7179 10777
rect 7121 10737 7133 10771
rect 7167 10768 7179 10771
rect 7394 10768 7400 10780
rect 7167 10740 7400 10768
rect 7167 10737 7179 10740
rect 7121 10731 7179 10737
rect 7394 10728 7400 10740
rect 7452 10728 7458 10780
rect 7302 10660 7308 10712
rect 7360 10700 7366 10712
rect 7360 10672 7624 10700
rect 7360 10660 7366 10672
rect 6750 10592 6756 10644
rect 6808 10632 6814 10644
rect 6808 10604 7256 10632
rect 6808 10592 6814 10604
rect 7118 10564 7124 10576
rect 7079 10536 7124 10564
rect 7118 10524 7124 10536
rect 7176 10524 7182 10576
rect 7228 10573 7256 10604
rect 7213 10567 7271 10573
rect 7213 10533 7225 10567
rect 7259 10564 7271 10567
rect 7302 10564 7308 10576
rect 7259 10536 7308 10564
rect 7259 10533 7271 10536
rect 7213 10527 7271 10533
rect 7302 10524 7308 10536
rect 7360 10524 7366 10576
rect 7596 10573 7624 10672
rect 7581 10567 7639 10573
rect 7581 10533 7593 10567
rect 7627 10533 7639 10567
rect 7581 10527 7639 10533
rect 7394 10496 7400 10508
rect 7355 10468 7400 10496
rect 7394 10456 7400 10468
rect 7452 10456 7458 10508
rect 7489 10499 7547 10505
rect 7489 10465 7501 10499
rect 7535 10496 7547 10499
rect 7596 10496 7624 10527
rect 7535 10468 7624 10496
rect 7535 10465 7547 10468
rect 7489 10459 7547 10465
rect 6750 10388 6756 10440
rect 6808 10428 6814 10440
rect 7504 10428 7532 10459
rect 6808 10400 7532 10428
rect 6808 10388 6814 10400
rect 3240 10338 8944 10360
rect 3240 10286 4984 10338
rect 5036 10286 5048 10338
rect 5100 10286 5112 10338
rect 5164 10286 5176 10338
rect 5228 10286 5240 10338
rect 5292 10286 5304 10338
rect 5356 10286 6915 10338
rect 6967 10286 6979 10338
rect 7031 10286 7043 10338
rect 7095 10286 7107 10338
rect 7159 10286 7171 10338
rect 7223 10286 7235 10338
rect 7287 10286 8944 10338
rect 3240 10264 8944 10286
rect 6658 10233 6664 10236
rect 6615 10227 6664 10233
rect 6615 10193 6627 10227
rect 6661 10193 6664 10227
rect 6615 10187 6664 10193
rect 6658 10184 6664 10187
rect 6716 10184 6722 10236
rect 7305 10227 7363 10233
rect 7305 10193 7317 10227
rect 7351 10224 7363 10227
rect 7578 10224 7584 10236
rect 7351 10196 7584 10224
rect 7351 10193 7363 10196
rect 7305 10187 7363 10193
rect 7578 10184 7584 10196
rect 7636 10184 7642 10236
rect 7489 10159 7547 10165
rect 7489 10125 7501 10159
rect 7535 10156 7547 10159
rect 7535 10128 7624 10156
rect 7535 10125 7547 10128
rect 7489 10119 7547 10125
rect 3162 10048 3168 10100
rect 3220 10088 3226 10100
rect 6566 10097 6572 10100
rect 3533 10091 3591 10097
rect 3533 10088 3545 10091
rect 3220 10060 3545 10088
rect 3220 10048 3226 10060
rect 3533 10057 3545 10060
rect 3579 10088 3591 10091
rect 4177 10091 4235 10097
rect 4177 10088 4189 10091
rect 3579 10060 4189 10088
rect 3579 10057 3591 10060
rect 3533 10051 3591 10057
rect 4177 10057 4189 10060
rect 4223 10057 4235 10091
rect 4177 10051 4235 10057
rect 6544 10091 6572 10097
rect 6544 10057 6556 10091
rect 6544 10051 6572 10057
rect 6566 10048 6572 10051
rect 6624 10048 6630 10100
rect 7121 10091 7179 10097
rect 7121 10057 7133 10091
rect 7167 10057 7179 10091
rect 7121 10051 7179 10057
rect 7213 10091 7271 10097
rect 7213 10057 7225 10091
rect 7259 10088 7271 10091
rect 7302 10088 7308 10100
rect 7259 10060 7308 10088
rect 7259 10057 7271 10060
rect 7213 10051 7271 10057
rect 7136 10020 7164 10051
rect 7302 10048 7308 10060
rect 7360 10048 7366 10100
rect 7394 10048 7400 10100
rect 7452 10088 7458 10100
rect 7596 10097 7624 10128
rect 7581 10091 7639 10097
rect 7452 10060 7497 10088
rect 7452 10048 7458 10060
rect 7581 10057 7593 10091
rect 7627 10088 7639 10091
rect 7670 10088 7676 10100
rect 7627 10060 7676 10088
rect 7627 10057 7639 10060
rect 7581 10051 7639 10057
rect 7670 10048 7676 10060
rect 7728 10048 7734 10100
rect 7486 10020 7492 10032
rect 7136 9992 7492 10020
rect 7486 9980 7492 9992
rect 7544 9980 7550 10032
rect 3717 9887 3775 9893
rect 3717 9853 3729 9887
rect 3763 9884 3775 9887
rect 6474 9884 6480 9896
rect 3763 9856 6480 9884
rect 3763 9853 3775 9856
rect 3717 9847 3775 9853
rect 6474 9844 6480 9856
rect 6532 9844 6538 9896
rect 3240 9794 8944 9816
rect 3240 9742 4019 9794
rect 4071 9742 4083 9794
rect 4135 9742 4147 9794
rect 4199 9742 4211 9794
rect 4263 9742 4275 9794
rect 4327 9742 4339 9794
rect 4391 9742 5950 9794
rect 6002 9742 6014 9794
rect 6066 9742 6078 9794
rect 6130 9742 6142 9794
rect 6194 9742 6206 9794
rect 6258 9742 6270 9794
rect 6322 9742 7880 9794
rect 7932 9742 7944 9794
rect 7996 9742 8008 9794
rect 8060 9742 8072 9794
rect 8124 9742 8136 9794
rect 8188 9742 8200 9794
rect 8252 9742 8944 9794
rect 3240 9720 8944 9742
rect 6566 9640 6572 9692
rect 6624 9680 6630 9692
rect 6845 9683 6903 9689
rect 6845 9680 6857 9683
rect 6624 9652 6857 9680
rect 6624 9640 6630 9652
rect 6845 9649 6857 9652
rect 6891 9649 6903 9683
rect 6845 9643 6903 9649
rect 7995 9683 8053 9689
rect 7995 9649 8007 9683
rect 8041 9680 8053 9683
rect 8314 9680 8320 9692
rect 8041 9652 8320 9680
rect 8041 9649 8053 9652
rect 7995 9643 8053 9649
rect 8314 9640 8320 9652
rect 8372 9640 8378 9692
rect 6934 9572 6940 9624
rect 6992 9612 6998 9624
rect 6992 9584 7808 9612
rect 6992 9572 6998 9584
rect 6474 9504 6480 9556
rect 6532 9544 6538 9556
rect 7305 9547 7363 9553
rect 6532 9516 7164 9544
rect 6532 9504 6538 9516
rect 6842 9476 6848 9488
rect 6803 9448 6848 9476
rect 6842 9436 6848 9448
rect 6900 9436 6906 9488
rect 7136 9485 7164 9516
rect 7305 9513 7317 9547
rect 7351 9513 7363 9547
rect 7305 9507 7363 9513
rect 7029 9479 7087 9485
rect 7029 9445 7041 9479
rect 7075 9445 7087 9479
rect 7029 9439 7087 9445
rect 7121 9479 7179 9485
rect 7121 9445 7133 9479
rect 7167 9445 7179 9479
rect 7320 9476 7348 9507
rect 7397 9479 7455 9485
rect 7397 9476 7409 9479
rect 7320 9448 7409 9476
rect 7121 9439 7179 9445
rect 7397 9445 7409 9448
rect 7443 9476 7455 9479
rect 7670 9476 7676 9488
rect 7443 9448 7676 9476
rect 7443 9445 7455 9448
rect 7397 9439 7455 9445
rect 7044 9408 7072 9439
rect 7670 9436 7676 9448
rect 7728 9436 7734 9488
rect 7780 9476 7808 9584
rect 7892 9479 7950 9485
rect 7892 9476 7904 9479
rect 7780 9448 7904 9476
rect 7892 9445 7904 9448
rect 7938 9445 7950 9479
rect 7892 9439 7950 9445
rect 6400 9380 7072 9408
rect 6400 9352 6428 9380
rect 6382 9340 6388 9352
rect 6343 9312 6388 9340
rect 6382 9300 6388 9312
rect 6440 9300 6446 9352
rect 3240 9250 8944 9272
rect 3240 9198 4984 9250
rect 5036 9198 5048 9250
rect 5100 9198 5112 9250
rect 5164 9198 5176 9250
rect 5228 9198 5240 9250
rect 5292 9198 5304 9250
rect 5356 9198 6915 9250
rect 6967 9198 6979 9250
rect 7031 9198 7043 9250
rect 7095 9198 7107 9250
rect 7159 9198 7171 9250
rect 7223 9198 7235 9250
rect 7287 9198 8944 9250
rect 3240 9176 8944 9198
rect 6983 9139 7041 9145
rect 6983 9105 6995 9139
rect 7029 9136 7041 9139
rect 7394 9136 7400 9148
rect 7029 9108 7400 9136
rect 7029 9105 7041 9108
rect 6983 9099 7041 9105
rect 7394 9096 7400 9108
rect 7452 9096 7458 9148
rect 6382 8960 6388 9012
rect 6440 9000 6446 9012
rect 6880 9003 6938 9009
rect 6880 9000 6892 9003
rect 6440 8972 6892 9000
rect 6440 8960 6446 8972
rect 6880 8969 6892 8972
rect 6926 8969 6938 9003
rect 6880 8963 6938 8969
rect 7581 9003 7639 9009
rect 7581 8969 7593 9003
rect 7627 9000 7639 9003
rect 8225 9003 8283 9009
rect 8225 9000 8237 9003
rect 7627 8972 8237 9000
rect 7627 8969 7639 8972
rect 7581 8963 7639 8969
rect 8225 8969 8237 8972
rect 8271 9000 8283 9003
rect 9142 9000 9148 9012
rect 8271 8972 9148 9000
rect 8271 8969 8283 8972
rect 8225 8963 8283 8969
rect 9142 8960 9148 8972
rect 9200 8960 9206 9012
rect 6750 8824 6756 8876
rect 6808 8864 6814 8876
rect 8041 8867 8099 8873
rect 8041 8864 8053 8867
rect 6808 8836 8053 8864
rect 6808 8824 6814 8836
rect 8041 8833 8053 8836
rect 8087 8833 8099 8867
rect 8041 8827 8099 8833
rect 6382 8796 6388 8808
rect 6343 8768 6388 8796
rect 6382 8756 6388 8768
rect 6440 8756 6446 8808
rect 3240 8706 8944 8728
rect 3240 8654 4019 8706
rect 4071 8654 4083 8706
rect 4135 8654 4147 8706
rect 4199 8654 4211 8706
rect 4263 8654 4275 8706
rect 4327 8654 4339 8706
rect 4391 8654 5950 8706
rect 6002 8654 6014 8706
rect 6066 8654 6078 8706
rect 6130 8654 6142 8706
rect 6194 8654 6206 8706
rect 6258 8654 6270 8706
rect 6322 8654 7880 8706
rect 7932 8654 7944 8706
rect 7996 8654 8008 8706
rect 8060 8654 8072 8706
rect 8124 8654 8136 8706
rect 8188 8654 8200 8706
rect 8252 8654 8944 8706
rect 3240 8632 8944 8654
rect 3240 8162 8944 8184
rect 3240 8110 4984 8162
rect 5036 8110 5048 8162
rect 5100 8110 5112 8162
rect 5164 8110 5176 8162
rect 5228 8110 5240 8162
rect 5292 8110 5304 8162
rect 5356 8110 6915 8162
rect 6967 8110 6979 8162
rect 7031 8110 7043 8162
rect 7095 8110 7107 8162
rect 7159 8110 7171 8162
rect 7223 8110 7235 8162
rect 7287 8110 8944 8162
rect 3240 8088 8944 8110
rect 3240 7618 8944 7640
rect 3240 7566 4019 7618
rect 4071 7566 4083 7618
rect 4135 7566 4147 7618
rect 4199 7566 4211 7618
rect 4263 7566 4275 7618
rect 4327 7566 4339 7618
rect 4391 7566 5950 7618
rect 6002 7566 6014 7618
rect 6066 7566 6078 7618
rect 6130 7566 6142 7618
rect 6194 7566 6206 7618
rect 6258 7566 6270 7618
rect 6322 7566 7880 7618
rect 7932 7566 7944 7618
rect 7996 7566 8008 7618
rect 8060 7566 8072 7618
rect 8124 7566 8136 7618
rect 8188 7566 8200 7618
rect 8252 7566 8944 7618
rect 3240 7544 8944 7566
rect 3240 7074 8944 7096
rect 3240 7022 4984 7074
rect 5036 7022 5048 7074
rect 5100 7022 5112 7074
rect 5164 7022 5176 7074
rect 5228 7022 5240 7074
rect 5292 7022 5304 7074
rect 5356 7022 6915 7074
rect 6967 7022 6979 7074
rect 7031 7022 7043 7074
rect 7095 7022 7107 7074
rect 7159 7022 7171 7074
rect 7223 7022 7235 7074
rect 7287 7022 8944 7074
rect 3240 7000 8944 7022
rect 3162 6580 3168 6632
rect 3220 6620 3226 6632
rect 6382 6620 6388 6632
rect 3220 6592 6388 6620
rect 3220 6580 3226 6592
rect 6382 6580 6388 6592
rect 6440 6580 6446 6632
rect 3240 6530 8944 6552
rect 3240 6478 4019 6530
rect 4071 6478 4083 6530
rect 4135 6478 4147 6530
rect 4199 6478 4211 6530
rect 4263 6478 4275 6530
rect 4327 6478 4339 6530
rect 4391 6478 5950 6530
rect 6002 6478 6014 6530
rect 6066 6478 6078 6530
rect 6130 6478 6142 6530
rect 6194 6478 6206 6530
rect 6258 6478 6270 6530
rect 6322 6478 7880 6530
rect 7932 6478 7944 6530
rect 7996 6478 8008 6530
rect 8060 6478 8072 6530
rect 8124 6478 8136 6530
rect 8188 6478 8200 6530
rect 8252 6478 8944 6530
rect 3240 6456 8944 6478
rect 3240 5986 8944 6008
rect 3240 5934 4984 5986
rect 5036 5934 5048 5986
rect 5100 5934 5112 5986
rect 5164 5934 5176 5986
rect 5228 5934 5240 5986
rect 5292 5934 5304 5986
rect 5356 5934 6915 5986
rect 6967 5934 6979 5986
rect 7031 5934 7043 5986
rect 7095 5934 7107 5986
rect 7159 5934 7171 5986
rect 7223 5934 7235 5986
rect 7287 5934 8944 5986
rect 3240 5912 8944 5934
rect 3240 5442 8944 5464
rect 3240 5390 4019 5442
rect 4071 5390 4083 5442
rect 4135 5390 4147 5442
rect 4199 5390 4211 5442
rect 4263 5390 4275 5442
rect 4327 5390 4339 5442
rect 4391 5390 5950 5442
rect 6002 5390 6014 5442
rect 6066 5390 6078 5442
rect 6130 5390 6142 5442
rect 6194 5390 6206 5442
rect 6258 5390 6270 5442
rect 6322 5390 7880 5442
rect 7932 5390 7944 5442
rect 7996 5390 8008 5442
rect 8060 5390 8072 5442
rect 8124 5390 8136 5442
rect 8188 5390 8200 5442
rect 8252 5390 8944 5442
rect 3240 5368 8944 5390
rect 3240 4898 8944 4920
rect 3240 4846 4984 4898
rect 5036 4846 5048 4898
rect 5100 4846 5112 4898
rect 5164 4846 5176 4898
rect 5228 4846 5240 4898
rect 5292 4846 5304 4898
rect 5356 4846 6915 4898
rect 6967 4846 6979 4898
rect 7031 4846 7043 4898
rect 7095 4846 7107 4898
rect 7159 4846 7171 4898
rect 7223 4846 7235 4898
rect 7287 4846 8944 4898
rect 3240 4824 8944 4846
rect 7670 4744 7676 4796
rect 7728 4784 7734 4796
rect 8041 4787 8099 4793
rect 8041 4784 8053 4787
rect 7728 4756 8053 4784
rect 7728 4744 7734 4756
rect 8041 4753 8053 4756
rect 8087 4753 8099 4787
rect 8041 4747 8099 4753
rect 7581 4651 7639 4657
rect 7581 4617 7593 4651
rect 7627 4648 7639 4651
rect 8225 4651 8283 4657
rect 8225 4648 8237 4651
rect 7627 4620 8237 4648
rect 7627 4617 7639 4620
rect 7581 4611 7639 4617
rect 8225 4617 8237 4620
rect 8271 4648 8283 4651
rect 9142 4648 9148 4660
rect 8271 4620 9148 4648
rect 8271 4617 8283 4620
rect 8225 4611 8283 4617
rect 9142 4608 9148 4620
rect 9200 4608 9206 4660
rect 3240 4354 8944 4376
rect 3240 4302 4019 4354
rect 4071 4302 4083 4354
rect 4135 4302 4147 4354
rect 4199 4302 4211 4354
rect 4263 4302 4275 4354
rect 4327 4302 4339 4354
rect 4391 4302 5950 4354
rect 6002 4302 6014 4354
rect 6066 4302 6078 4354
rect 6130 4302 6142 4354
rect 6194 4302 6206 4354
rect 6258 4302 6270 4354
rect 6322 4302 7880 4354
rect 7932 4302 7944 4354
rect 7996 4302 8008 4354
rect 8060 4302 8072 4354
rect 8124 4302 8136 4354
rect 8188 4302 8200 4354
rect 8252 4302 8944 4354
rect 3240 4280 8944 4302
rect 3240 3810 8944 3832
rect 3240 3758 4984 3810
rect 5036 3758 5048 3810
rect 5100 3758 5112 3810
rect 5164 3758 5176 3810
rect 5228 3758 5240 3810
rect 5292 3758 5304 3810
rect 5356 3758 6915 3810
rect 6967 3758 6979 3810
rect 7031 3758 7043 3810
rect 7095 3758 7107 3810
rect 7159 3758 7171 3810
rect 7223 3758 7235 3810
rect 7287 3758 8944 3810
rect 3240 3736 8944 3758
rect 3240 3266 8944 3288
rect 3240 3214 4019 3266
rect 4071 3214 4083 3266
rect 4135 3214 4147 3266
rect 4199 3214 4211 3266
rect 4263 3214 4275 3266
rect 4327 3214 4339 3266
rect 4391 3214 5950 3266
rect 6002 3214 6014 3266
rect 6066 3214 6078 3266
rect 6130 3214 6142 3266
rect 6194 3214 6206 3266
rect 6258 3214 6270 3266
rect 6322 3214 7880 3266
rect 7932 3214 7944 3266
rect 7996 3214 8008 3266
rect 8060 3214 8072 3266
rect 8124 3214 8136 3266
rect 8188 3214 8200 3266
rect 8252 3214 8944 3266
rect 3240 3192 8944 3214
<< via1 >>
rect 4984 16814 5036 16866
rect 5048 16814 5100 16866
rect 5112 16814 5164 16866
rect 5176 16814 5228 16866
rect 5240 16814 5292 16866
rect 5304 16814 5356 16866
rect 6915 16814 6967 16866
rect 6979 16814 7031 16866
rect 7043 16814 7095 16866
rect 7107 16814 7159 16866
rect 7171 16814 7223 16866
rect 7235 16814 7287 16866
rect 4019 16270 4071 16322
rect 4083 16270 4135 16322
rect 4147 16270 4199 16322
rect 4211 16270 4263 16322
rect 4275 16270 4327 16322
rect 4339 16270 4391 16322
rect 5950 16270 6002 16322
rect 6014 16270 6066 16322
rect 6078 16270 6130 16322
rect 6142 16270 6194 16322
rect 6206 16270 6258 16322
rect 6270 16270 6322 16322
rect 7880 16270 7932 16322
rect 7944 16270 7996 16322
rect 8008 16270 8060 16322
rect 8072 16270 8124 16322
rect 8136 16270 8188 16322
rect 8200 16270 8252 16322
rect 9148 16100 9200 16152
rect 3168 15964 3220 16016
rect 7676 15964 7728 16016
rect 6756 15828 6808 15880
rect 4984 15726 5036 15778
rect 5048 15726 5100 15778
rect 5112 15726 5164 15778
rect 5176 15726 5228 15778
rect 5240 15726 5292 15778
rect 5304 15726 5356 15778
rect 6915 15726 6967 15778
rect 6979 15726 7031 15778
rect 7043 15726 7095 15778
rect 7107 15726 7159 15778
rect 7171 15726 7223 15778
rect 7235 15726 7287 15778
rect 4019 15182 4071 15234
rect 4083 15182 4135 15234
rect 4147 15182 4199 15234
rect 4211 15182 4263 15234
rect 4275 15182 4327 15234
rect 4339 15182 4391 15234
rect 5950 15182 6002 15234
rect 6014 15182 6066 15234
rect 6078 15182 6130 15234
rect 6142 15182 6194 15234
rect 6206 15182 6258 15234
rect 6270 15182 6322 15234
rect 7880 15182 7932 15234
rect 7944 15182 7996 15234
rect 8008 15182 8060 15234
rect 8072 15182 8124 15234
rect 8136 15182 8188 15234
rect 8200 15182 8252 15234
rect 4984 14638 5036 14690
rect 5048 14638 5100 14690
rect 5112 14638 5164 14690
rect 5176 14638 5228 14690
rect 5240 14638 5292 14690
rect 5304 14638 5356 14690
rect 6915 14638 6967 14690
rect 6979 14638 7031 14690
rect 7043 14638 7095 14690
rect 7107 14638 7159 14690
rect 7171 14638 7223 14690
rect 7235 14638 7287 14690
rect 4019 14094 4071 14146
rect 4083 14094 4135 14146
rect 4147 14094 4199 14146
rect 4211 14094 4263 14146
rect 4275 14094 4327 14146
rect 4339 14094 4391 14146
rect 5950 14094 6002 14146
rect 6014 14094 6066 14146
rect 6078 14094 6130 14146
rect 6142 14094 6194 14146
rect 6206 14094 6258 14146
rect 6270 14094 6322 14146
rect 7880 14094 7932 14146
rect 7944 14094 7996 14146
rect 8008 14094 8060 14146
rect 8072 14094 8124 14146
rect 8136 14094 8188 14146
rect 8200 14094 8252 14146
rect 4984 13550 5036 13602
rect 5048 13550 5100 13602
rect 5112 13550 5164 13602
rect 5176 13550 5228 13602
rect 5240 13550 5292 13602
rect 5304 13550 5356 13602
rect 6915 13550 6967 13602
rect 6979 13550 7031 13602
rect 7043 13550 7095 13602
rect 7107 13550 7159 13602
rect 7171 13550 7223 13602
rect 7235 13550 7287 13602
rect 4019 13006 4071 13058
rect 4083 13006 4135 13058
rect 4147 13006 4199 13058
rect 4211 13006 4263 13058
rect 4275 13006 4327 13058
rect 4339 13006 4391 13058
rect 5950 13006 6002 13058
rect 6014 13006 6066 13058
rect 6078 13006 6130 13058
rect 6142 13006 6194 13058
rect 6206 13006 6258 13058
rect 6270 13006 6322 13058
rect 7880 13006 7932 13058
rect 7944 13006 7996 13058
rect 8008 13006 8060 13058
rect 8072 13006 8124 13058
rect 8136 13006 8188 13058
rect 8200 13006 8252 13058
rect 4984 12462 5036 12514
rect 5048 12462 5100 12514
rect 5112 12462 5164 12514
rect 5176 12462 5228 12514
rect 5240 12462 5292 12514
rect 5304 12462 5356 12514
rect 6915 12462 6967 12514
rect 6979 12462 7031 12514
rect 7043 12462 7095 12514
rect 7107 12462 7159 12514
rect 7171 12462 7223 12514
rect 7235 12462 7287 12514
rect 4019 11918 4071 11970
rect 4083 11918 4135 11970
rect 4147 11918 4199 11970
rect 4211 11918 4263 11970
rect 4275 11918 4327 11970
rect 4339 11918 4391 11970
rect 5950 11918 6002 11970
rect 6014 11918 6066 11970
rect 6078 11918 6130 11970
rect 6142 11918 6194 11970
rect 6206 11918 6258 11970
rect 6270 11918 6322 11970
rect 7880 11918 7932 11970
rect 7944 11918 7996 11970
rect 8008 11918 8060 11970
rect 8072 11918 8124 11970
rect 8136 11918 8188 11970
rect 8200 11918 8252 11970
rect 6664 11680 6716 11732
rect 7676 11723 7728 11732
rect 7676 11689 7685 11723
rect 7685 11689 7719 11723
rect 7719 11689 7728 11723
rect 7676 11680 7728 11689
rect 7400 11655 7452 11664
rect 7400 11621 7409 11655
rect 7409 11621 7443 11655
rect 7443 11621 7452 11655
rect 7400 11612 7452 11621
rect 7860 11476 7912 11528
rect 4984 11374 5036 11426
rect 5048 11374 5100 11426
rect 5112 11374 5164 11426
rect 5176 11374 5228 11426
rect 5240 11374 5292 11426
rect 5304 11374 5356 11426
rect 6915 11374 6967 11426
rect 6979 11374 7031 11426
rect 7043 11374 7095 11426
rect 7107 11374 7159 11426
rect 7171 11374 7223 11426
rect 7235 11374 7287 11426
rect 7676 11272 7728 11324
rect 6388 11204 6440 11256
rect 6572 11136 6624 11188
rect 6480 11068 6532 11120
rect 7308 11136 7360 11188
rect 7860 11179 7912 11188
rect 7860 11145 7869 11179
rect 7869 11145 7903 11179
rect 7903 11145 7912 11179
rect 7860 11136 7912 11145
rect 8320 11068 8372 11120
rect 7124 11000 7176 11052
rect 7584 11000 7636 11052
rect 6388 10975 6440 10984
rect 6388 10941 6397 10975
rect 6397 10941 6431 10975
rect 6431 10941 6440 10975
rect 6388 10932 6440 10941
rect 7032 10932 7084 10984
rect 7308 10975 7360 10984
rect 7308 10941 7317 10975
rect 7317 10941 7351 10975
rect 7351 10941 7360 10975
rect 7308 10932 7360 10941
rect 4019 10830 4071 10882
rect 4083 10830 4135 10882
rect 4147 10830 4199 10882
rect 4211 10830 4263 10882
rect 4275 10830 4327 10882
rect 4339 10830 4391 10882
rect 5950 10830 6002 10882
rect 6014 10830 6066 10882
rect 6078 10830 6130 10882
rect 6142 10830 6194 10882
rect 6206 10830 6258 10882
rect 6270 10830 6322 10882
rect 7880 10830 7932 10882
rect 7944 10830 7996 10882
rect 8008 10830 8060 10882
rect 8072 10830 8124 10882
rect 8136 10830 8188 10882
rect 8200 10830 8252 10882
rect 7400 10728 7452 10780
rect 7308 10660 7360 10712
rect 6756 10592 6808 10644
rect 7124 10567 7176 10576
rect 7124 10533 7133 10567
rect 7133 10533 7167 10567
rect 7167 10533 7176 10567
rect 7124 10524 7176 10533
rect 7308 10524 7360 10576
rect 7400 10499 7452 10508
rect 7400 10465 7409 10499
rect 7409 10465 7443 10499
rect 7443 10465 7452 10499
rect 7400 10456 7452 10465
rect 6756 10388 6808 10440
rect 4984 10286 5036 10338
rect 5048 10286 5100 10338
rect 5112 10286 5164 10338
rect 5176 10286 5228 10338
rect 5240 10286 5292 10338
rect 5304 10286 5356 10338
rect 6915 10286 6967 10338
rect 6979 10286 7031 10338
rect 7043 10286 7095 10338
rect 7107 10286 7159 10338
rect 7171 10286 7223 10338
rect 7235 10286 7287 10338
rect 6664 10184 6716 10236
rect 7584 10184 7636 10236
rect 3168 10048 3220 10100
rect 6572 10091 6624 10100
rect 6572 10057 6590 10091
rect 6590 10057 6624 10091
rect 6572 10048 6624 10057
rect 7308 10048 7360 10100
rect 7400 10091 7452 10100
rect 7400 10057 7409 10091
rect 7409 10057 7443 10091
rect 7443 10057 7452 10091
rect 7400 10048 7452 10057
rect 7676 10048 7728 10100
rect 7492 9980 7544 10032
rect 6480 9844 6532 9896
rect 4019 9742 4071 9794
rect 4083 9742 4135 9794
rect 4147 9742 4199 9794
rect 4211 9742 4263 9794
rect 4275 9742 4327 9794
rect 4339 9742 4391 9794
rect 5950 9742 6002 9794
rect 6014 9742 6066 9794
rect 6078 9742 6130 9794
rect 6142 9742 6194 9794
rect 6206 9742 6258 9794
rect 6270 9742 6322 9794
rect 7880 9742 7932 9794
rect 7944 9742 7996 9794
rect 8008 9742 8060 9794
rect 8072 9742 8124 9794
rect 8136 9742 8188 9794
rect 8200 9742 8252 9794
rect 6572 9640 6624 9692
rect 8320 9640 8372 9692
rect 6940 9572 6992 9624
rect 6480 9504 6532 9556
rect 6848 9479 6900 9488
rect 6848 9445 6857 9479
rect 6857 9445 6891 9479
rect 6891 9445 6900 9479
rect 6848 9436 6900 9445
rect 7676 9436 7728 9488
rect 6388 9343 6440 9352
rect 6388 9309 6397 9343
rect 6397 9309 6431 9343
rect 6431 9309 6440 9343
rect 6388 9300 6440 9309
rect 4984 9198 5036 9250
rect 5048 9198 5100 9250
rect 5112 9198 5164 9250
rect 5176 9198 5228 9250
rect 5240 9198 5292 9250
rect 5304 9198 5356 9250
rect 6915 9198 6967 9250
rect 6979 9198 7031 9250
rect 7043 9198 7095 9250
rect 7107 9198 7159 9250
rect 7171 9198 7223 9250
rect 7235 9198 7287 9250
rect 7400 9096 7452 9148
rect 6388 8960 6440 9012
rect 9148 8960 9200 9012
rect 6756 8824 6808 8876
rect 6388 8799 6440 8808
rect 6388 8765 6397 8799
rect 6397 8765 6431 8799
rect 6431 8765 6440 8799
rect 6388 8756 6440 8765
rect 4019 8654 4071 8706
rect 4083 8654 4135 8706
rect 4147 8654 4199 8706
rect 4211 8654 4263 8706
rect 4275 8654 4327 8706
rect 4339 8654 4391 8706
rect 5950 8654 6002 8706
rect 6014 8654 6066 8706
rect 6078 8654 6130 8706
rect 6142 8654 6194 8706
rect 6206 8654 6258 8706
rect 6270 8654 6322 8706
rect 7880 8654 7932 8706
rect 7944 8654 7996 8706
rect 8008 8654 8060 8706
rect 8072 8654 8124 8706
rect 8136 8654 8188 8706
rect 8200 8654 8252 8706
rect 4984 8110 5036 8162
rect 5048 8110 5100 8162
rect 5112 8110 5164 8162
rect 5176 8110 5228 8162
rect 5240 8110 5292 8162
rect 5304 8110 5356 8162
rect 6915 8110 6967 8162
rect 6979 8110 7031 8162
rect 7043 8110 7095 8162
rect 7107 8110 7159 8162
rect 7171 8110 7223 8162
rect 7235 8110 7287 8162
rect 4019 7566 4071 7618
rect 4083 7566 4135 7618
rect 4147 7566 4199 7618
rect 4211 7566 4263 7618
rect 4275 7566 4327 7618
rect 4339 7566 4391 7618
rect 5950 7566 6002 7618
rect 6014 7566 6066 7618
rect 6078 7566 6130 7618
rect 6142 7566 6194 7618
rect 6206 7566 6258 7618
rect 6270 7566 6322 7618
rect 7880 7566 7932 7618
rect 7944 7566 7996 7618
rect 8008 7566 8060 7618
rect 8072 7566 8124 7618
rect 8136 7566 8188 7618
rect 8200 7566 8252 7618
rect 4984 7022 5036 7074
rect 5048 7022 5100 7074
rect 5112 7022 5164 7074
rect 5176 7022 5228 7074
rect 5240 7022 5292 7074
rect 5304 7022 5356 7074
rect 6915 7022 6967 7074
rect 6979 7022 7031 7074
rect 7043 7022 7095 7074
rect 7107 7022 7159 7074
rect 7171 7022 7223 7074
rect 7235 7022 7287 7074
rect 3168 6580 3220 6632
rect 6388 6580 6440 6632
rect 4019 6478 4071 6530
rect 4083 6478 4135 6530
rect 4147 6478 4199 6530
rect 4211 6478 4263 6530
rect 4275 6478 4327 6530
rect 4339 6478 4391 6530
rect 5950 6478 6002 6530
rect 6014 6478 6066 6530
rect 6078 6478 6130 6530
rect 6142 6478 6194 6530
rect 6206 6478 6258 6530
rect 6270 6478 6322 6530
rect 7880 6478 7932 6530
rect 7944 6478 7996 6530
rect 8008 6478 8060 6530
rect 8072 6478 8124 6530
rect 8136 6478 8188 6530
rect 8200 6478 8252 6530
rect 4984 5934 5036 5986
rect 5048 5934 5100 5986
rect 5112 5934 5164 5986
rect 5176 5934 5228 5986
rect 5240 5934 5292 5986
rect 5304 5934 5356 5986
rect 6915 5934 6967 5986
rect 6979 5934 7031 5986
rect 7043 5934 7095 5986
rect 7107 5934 7159 5986
rect 7171 5934 7223 5986
rect 7235 5934 7287 5986
rect 4019 5390 4071 5442
rect 4083 5390 4135 5442
rect 4147 5390 4199 5442
rect 4211 5390 4263 5442
rect 4275 5390 4327 5442
rect 4339 5390 4391 5442
rect 5950 5390 6002 5442
rect 6014 5390 6066 5442
rect 6078 5390 6130 5442
rect 6142 5390 6194 5442
rect 6206 5390 6258 5442
rect 6270 5390 6322 5442
rect 7880 5390 7932 5442
rect 7944 5390 7996 5442
rect 8008 5390 8060 5442
rect 8072 5390 8124 5442
rect 8136 5390 8188 5442
rect 8200 5390 8252 5442
rect 4984 4846 5036 4898
rect 5048 4846 5100 4898
rect 5112 4846 5164 4898
rect 5176 4846 5228 4898
rect 5240 4846 5292 4898
rect 5304 4846 5356 4898
rect 6915 4846 6967 4898
rect 6979 4846 7031 4898
rect 7043 4846 7095 4898
rect 7107 4846 7159 4898
rect 7171 4846 7223 4898
rect 7235 4846 7287 4898
rect 7676 4744 7728 4796
rect 9148 4608 9200 4660
rect 4019 4302 4071 4354
rect 4083 4302 4135 4354
rect 4147 4302 4199 4354
rect 4211 4302 4263 4354
rect 4275 4302 4327 4354
rect 4339 4302 4391 4354
rect 5950 4302 6002 4354
rect 6014 4302 6066 4354
rect 6078 4302 6130 4354
rect 6142 4302 6194 4354
rect 6206 4302 6258 4354
rect 6270 4302 6322 4354
rect 7880 4302 7932 4354
rect 7944 4302 7996 4354
rect 8008 4302 8060 4354
rect 8072 4302 8124 4354
rect 8136 4302 8188 4354
rect 8200 4302 8252 4354
rect 4984 3758 5036 3810
rect 5048 3758 5100 3810
rect 5112 3758 5164 3810
rect 5176 3758 5228 3810
rect 5240 3758 5292 3810
rect 5304 3758 5356 3810
rect 6915 3758 6967 3810
rect 6979 3758 7031 3810
rect 7043 3758 7095 3810
rect 7107 3758 7159 3810
rect 7171 3758 7223 3810
rect 7235 3758 7287 3810
rect 4019 3214 4071 3266
rect 4083 3214 4135 3266
rect 4147 3214 4199 3266
rect 4211 3214 4263 3266
rect 4275 3214 4327 3266
rect 4339 3214 4391 3266
rect 5950 3214 6002 3266
rect 6014 3214 6066 3266
rect 6078 3214 6130 3266
rect 6142 3214 6194 3266
rect 6206 3214 6258 3266
rect 6270 3214 6322 3266
rect 7880 3214 7932 3266
rect 7944 3214 7996 3266
rect 8008 3214 8060 3266
rect 8072 3214 8124 3266
rect 8136 3214 8188 3266
rect 8200 3214 8252 3266
<< metal2 >>
rect 4982 16868 5358 16888
rect 5038 16866 5062 16868
rect 5118 16866 5142 16868
rect 5198 16866 5222 16868
rect 5278 16866 5302 16868
rect 5038 16814 5048 16866
rect 5292 16814 5302 16866
rect 5038 16812 5062 16814
rect 5118 16812 5142 16814
rect 5198 16812 5222 16814
rect 5278 16812 5302 16814
rect 4982 16792 5358 16812
rect 6913 16868 7289 16888
rect 6969 16866 6993 16868
rect 7049 16866 7073 16868
rect 7129 16866 7153 16868
rect 7209 16866 7233 16868
rect 6969 16814 6979 16866
rect 7223 16814 7233 16866
rect 6969 16812 6993 16814
rect 7049 16812 7073 16814
rect 7129 16812 7153 16814
rect 7209 16812 7233 16814
rect 6913 16792 7289 16812
rect 4017 16324 4393 16344
rect 4073 16322 4097 16324
rect 4153 16322 4177 16324
rect 4233 16322 4257 16324
rect 4313 16322 4337 16324
rect 4073 16270 4083 16322
rect 4327 16270 4337 16322
rect 4073 16268 4097 16270
rect 4153 16268 4177 16270
rect 4233 16268 4257 16270
rect 4313 16268 4337 16270
rect 4017 16248 4393 16268
rect 5948 16324 6324 16344
rect 6004 16322 6028 16324
rect 6084 16322 6108 16324
rect 6164 16322 6188 16324
rect 6244 16322 6268 16324
rect 6004 16270 6014 16322
rect 6258 16270 6268 16322
rect 6004 16268 6028 16270
rect 6084 16268 6108 16270
rect 6164 16268 6188 16270
rect 6244 16268 6268 16270
rect 5948 16248 6324 16268
rect 7878 16324 8254 16344
rect 7934 16322 7958 16324
rect 8014 16322 8038 16324
rect 8094 16322 8118 16324
rect 8174 16322 8198 16324
rect 7934 16270 7944 16322
rect 8188 16270 8198 16322
rect 7934 16268 7958 16270
rect 8014 16268 8038 16270
rect 8094 16268 8118 16270
rect 8174 16268 8198 16270
rect 7878 16248 8254 16268
rect 9148 16152 9200 16158
rect 2136 16028 2936 16126
rect 9148 16094 9200 16100
rect 9160 16028 9188 16094
rect 9336 16028 10136 16126
rect 2136 16022 3208 16028
rect 2136 16016 3220 16022
rect 2136 16000 3168 16016
rect 2136 15902 2936 16000
rect 3168 15958 3220 15964
rect 7676 16016 7728 16022
rect 9160 16000 10136 16028
rect 7676 15958 7728 15964
rect 6756 15880 6808 15886
rect 6756 15822 6808 15828
rect 4982 15780 5358 15800
rect 5038 15778 5062 15780
rect 5118 15778 5142 15780
rect 5198 15778 5222 15780
rect 5278 15778 5302 15780
rect 5038 15726 5048 15778
rect 5292 15726 5302 15778
rect 5038 15724 5062 15726
rect 5118 15724 5142 15726
rect 5198 15724 5222 15726
rect 5278 15724 5302 15726
rect 4982 15704 5358 15724
rect 4017 15236 4393 15256
rect 4073 15234 4097 15236
rect 4153 15234 4177 15236
rect 4233 15234 4257 15236
rect 4313 15234 4337 15236
rect 4073 15182 4083 15234
rect 4327 15182 4337 15234
rect 4073 15180 4097 15182
rect 4153 15180 4177 15182
rect 4233 15180 4257 15182
rect 4313 15180 4337 15182
rect 4017 15160 4393 15180
rect 5948 15236 6324 15256
rect 6004 15234 6028 15236
rect 6084 15234 6108 15236
rect 6164 15234 6188 15236
rect 6244 15234 6268 15236
rect 6004 15182 6014 15234
rect 6258 15182 6268 15234
rect 6004 15180 6028 15182
rect 6084 15180 6108 15182
rect 6164 15180 6188 15182
rect 6244 15180 6268 15182
rect 5948 15160 6324 15180
rect 4982 14692 5358 14712
rect 5038 14690 5062 14692
rect 5118 14690 5142 14692
rect 5198 14690 5222 14692
rect 5278 14690 5302 14692
rect 5038 14638 5048 14690
rect 5292 14638 5302 14690
rect 5038 14636 5062 14638
rect 5118 14636 5142 14638
rect 5198 14636 5222 14638
rect 5278 14636 5302 14638
rect 4982 14616 5358 14636
rect 4017 14148 4393 14168
rect 4073 14146 4097 14148
rect 4153 14146 4177 14148
rect 4233 14146 4257 14148
rect 4313 14146 4337 14148
rect 4073 14094 4083 14146
rect 4327 14094 4337 14146
rect 4073 14092 4097 14094
rect 4153 14092 4177 14094
rect 4233 14092 4257 14094
rect 4313 14092 4337 14094
rect 4017 14072 4393 14092
rect 5948 14148 6324 14168
rect 6004 14146 6028 14148
rect 6084 14146 6108 14148
rect 6164 14146 6188 14148
rect 6244 14146 6268 14148
rect 6004 14094 6014 14146
rect 6258 14094 6268 14146
rect 6004 14092 6028 14094
rect 6084 14092 6108 14094
rect 6164 14092 6188 14094
rect 6244 14092 6268 14094
rect 5948 14072 6324 14092
rect 4982 13604 5358 13624
rect 5038 13602 5062 13604
rect 5118 13602 5142 13604
rect 5198 13602 5222 13604
rect 5278 13602 5302 13604
rect 5038 13550 5048 13602
rect 5292 13550 5302 13602
rect 5038 13548 5062 13550
rect 5118 13548 5142 13550
rect 5198 13548 5222 13550
rect 5278 13548 5302 13550
rect 4982 13528 5358 13548
rect 4017 13060 4393 13080
rect 4073 13058 4097 13060
rect 4153 13058 4177 13060
rect 4233 13058 4257 13060
rect 4313 13058 4337 13060
rect 4073 13006 4083 13058
rect 4327 13006 4337 13058
rect 4073 13004 4097 13006
rect 4153 13004 4177 13006
rect 4233 13004 4257 13006
rect 4313 13004 4337 13006
rect 4017 12984 4393 13004
rect 5948 13060 6324 13080
rect 6004 13058 6028 13060
rect 6084 13058 6108 13060
rect 6164 13058 6188 13060
rect 6244 13058 6268 13060
rect 6004 13006 6014 13058
rect 6258 13006 6268 13058
rect 6004 13004 6028 13006
rect 6084 13004 6108 13006
rect 6164 13004 6188 13006
rect 6244 13004 6268 13006
rect 5948 12984 6324 13004
rect 4982 12516 5358 12536
rect 5038 12514 5062 12516
rect 5118 12514 5142 12516
rect 5198 12514 5222 12516
rect 5278 12514 5302 12516
rect 5038 12462 5048 12514
rect 5292 12462 5302 12514
rect 5038 12460 5062 12462
rect 5118 12460 5142 12462
rect 5198 12460 5222 12462
rect 5278 12460 5302 12462
rect 4982 12440 5358 12460
rect 4017 11972 4393 11992
rect 4073 11970 4097 11972
rect 4153 11970 4177 11972
rect 4233 11970 4257 11972
rect 4313 11970 4337 11972
rect 4073 11918 4083 11970
rect 4327 11918 4337 11970
rect 4073 11916 4097 11918
rect 4153 11916 4177 11918
rect 4233 11916 4257 11918
rect 4313 11916 4337 11918
rect 4017 11896 4393 11916
rect 5948 11972 6324 11992
rect 6004 11970 6028 11972
rect 6084 11970 6108 11972
rect 6164 11970 6188 11972
rect 6244 11970 6268 11972
rect 6004 11918 6014 11970
rect 6258 11918 6268 11970
rect 6004 11916 6028 11918
rect 6084 11916 6108 11918
rect 6164 11916 6188 11918
rect 6244 11916 6268 11918
rect 5948 11896 6324 11916
rect 6664 11732 6716 11738
rect 6664 11674 6716 11680
rect 4982 11428 5358 11448
rect 5038 11426 5062 11428
rect 5118 11426 5142 11428
rect 5198 11426 5222 11428
rect 5278 11426 5302 11428
rect 5038 11374 5048 11426
rect 5292 11374 5302 11426
rect 5038 11372 5062 11374
rect 5118 11372 5142 11374
rect 5198 11372 5222 11374
rect 5278 11372 5302 11374
rect 4982 11352 5358 11372
rect 6388 11256 6440 11262
rect 6388 11198 6440 11204
rect 6400 10990 6428 11198
rect 6572 11188 6624 11194
rect 6572 11130 6624 11136
rect 6480 11120 6532 11126
rect 6480 11062 6532 11068
rect 6388 10984 6440 10990
rect 6388 10926 6440 10932
rect 4017 10884 4393 10904
rect 4073 10882 4097 10884
rect 4153 10882 4177 10884
rect 4233 10882 4257 10884
rect 4313 10882 4337 10884
rect 4073 10830 4083 10882
rect 4327 10830 4337 10882
rect 4073 10828 4097 10830
rect 4153 10828 4177 10830
rect 4233 10828 4257 10830
rect 4313 10828 4337 10830
rect 4017 10808 4393 10828
rect 5948 10884 6324 10904
rect 6004 10882 6028 10884
rect 6084 10882 6108 10884
rect 6164 10882 6188 10884
rect 6244 10882 6268 10884
rect 6004 10830 6014 10882
rect 6258 10830 6268 10882
rect 6004 10828 6028 10830
rect 6084 10828 6108 10830
rect 6164 10828 6188 10830
rect 6244 10828 6268 10830
rect 5948 10808 6324 10828
rect 4982 10340 5358 10360
rect 5038 10338 5062 10340
rect 5118 10338 5142 10340
rect 5198 10338 5222 10340
rect 5278 10338 5302 10340
rect 5038 10286 5048 10338
rect 5292 10286 5302 10338
rect 5038 10284 5062 10286
rect 5118 10284 5142 10286
rect 5198 10284 5222 10286
rect 5278 10284 5302 10286
rect 4982 10264 5358 10284
rect 2136 10048 2936 10146
rect 3168 10100 3220 10106
rect 2136 10042 3220 10048
rect 2136 10020 3208 10042
rect 2136 9922 2936 10020
rect 4017 9796 4393 9816
rect 4073 9794 4097 9796
rect 4153 9794 4177 9796
rect 4233 9794 4257 9796
rect 4313 9794 4337 9796
rect 4073 9742 4083 9794
rect 4327 9742 4337 9794
rect 4073 9740 4097 9742
rect 4153 9740 4177 9742
rect 4233 9740 4257 9742
rect 4313 9740 4337 9742
rect 4017 9720 4393 9740
rect 5948 9796 6324 9816
rect 6004 9794 6028 9796
rect 6084 9794 6108 9796
rect 6164 9794 6188 9796
rect 6244 9794 6268 9796
rect 6004 9742 6014 9794
rect 6258 9742 6268 9794
rect 6004 9740 6028 9742
rect 6084 9740 6108 9742
rect 6164 9740 6188 9742
rect 6244 9740 6268 9742
rect 5948 9720 6324 9740
rect 6400 9358 6428 10926
rect 6492 9902 6520 11062
rect 6584 10106 6612 11130
rect 6676 10242 6704 11674
rect 6768 10650 6796 15822
rect 6913 15780 7289 15800
rect 6969 15778 6993 15780
rect 7049 15778 7073 15780
rect 7129 15778 7153 15780
rect 7209 15778 7233 15780
rect 6969 15726 6979 15778
rect 7223 15726 7233 15778
rect 6969 15724 6993 15726
rect 7049 15724 7073 15726
rect 7129 15724 7153 15726
rect 7209 15724 7233 15726
rect 6913 15704 7289 15724
rect 6913 14692 7289 14712
rect 6969 14690 6993 14692
rect 7049 14690 7073 14692
rect 7129 14690 7153 14692
rect 7209 14690 7233 14692
rect 6969 14638 6979 14690
rect 7223 14638 7233 14690
rect 6969 14636 6993 14638
rect 7049 14636 7073 14638
rect 7129 14636 7153 14638
rect 7209 14636 7233 14638
rect 6913 14616 7289 14636
rect 6913 13604 7289 13624
rect 6969 13602 6993 13604
rect 7049 13602 7073 13604
rect 7129 13602 7153 13604
rect 7209 13602 7233 13604
rect 6969 13550 6979 13602
rect 7223 13550 7233 13602
rect 6969 13548 6993 13550
rect 7049 13548 7073 13550
rect 7129 13548 7153 13550
rect 7209 13548 7233 13550
rect 6913 13528 7289 13548
rect 6913 12516 7289 12536
rect 6969 12514 6993 12516
rect 7049 12514 7073 12516
rect 7129 12514 7153 12516
rect 7209 12514 7233 12516
rect 6969 12462 6979 12514
rect 7223 12462 7233 12514
rect 6969 12460 6993 12462
rect 7049 12460 7073 12462
rect 7129 12460 7153 12462
rect 7209 12460 7233 12462
rect 6913 12440 7289 12460
rect 7688 11738 7716 15958
rect 9336 15902 10136 16000
rect 7878 15236 8254 15256
rect 7934 15234 7958 15236
rect 8014 15234 8038 15236
rect 8094 15234 8118 15236
rect 8174 15234 8198 15236
rect 7934 15182 7944 15234
rect 8188 15182 8198 15234
rect 7934 15180 7958 15182
rect 8014 15180 8038 15182
rect 8094 15180 8118 15182
rect 8174 15180 8198 15182
rect 7878 15160 8254 15180
rect 7878 14148 8254 14168
rect 7934 14146 7958 14148
rect 8014 14146 8038 14148
rect 8094 14146 8118 14148
rect 8174 14146 8198 14148
rect 7934 14094 7944 14146
rect 8188 14094 8198 14146
rect 7934 14092 7958 14094
rect 8014 14092 8038 14094
rect 8094 14092 8118 14094
rect 8174 14092 8198 14094
rect 7878 14072 8254 14092
rect 7878 13060 8254 13080
rect 7934 13058 7958 13060
rect 8014 13058 8038 13060
rect 8094 13058 8118 13060
rect 8174 13058 8198 13060
rect 7934 13006 7944 13058
rect 8188 13006 8198 13058
rect 7934 13004 7958 13006
rect 8014 13004 8038 13006
rect 8094 13004 8118 13006
rect 8174 13004 8198 13006
rect 7878 12984 8254 13004
rect 7878 11972 8254 11992
rect 7934 11970 7958 11972
rect 8014 11970 8038 11972
rect 8094 11970 8118 11972
rect 8174 11970 8198 11972
rect 7934 11918 7944 11970
rect 8188 11918 8198 11970
rect 7934 11916 7958 11918
rect 8014 11916 8038 11918
rect 8094 11916 8118 11918
rect 8174 11916 8198 11918
rect 7878 11896 8254 11916
rect 7676 11732 7728 11738
rect 7676 11674 7728 11680
rect 7400 11664 7452 11670
rect 7400 11606 7452 11612
rect 6913 11428 7289 11448
rect 6969 11426 6993 11428
rect 7049 11426 7073 11428
rect 7129 11426 7153 11428
rect 7209 11426 7233 11428
rect 6969 11374 6979 11426
rect 7223 11374 7233 11426
rect 6969 11372 6993 11374
rect 7049 11372 7073 11374
rect 7129 11372 7153 11374
rect 7209 11372 7233 11374
rect 6913 11352 7289 11372
rect 7308 11188 7360 11194
rect 7308 11130 7360 11136
rect 7124 11052 7176 11058
rect 7124 10994 7176 11000
rect 7032 10984 7084 10990
rect 7032 10926 7084 10932
rect 6756 10644 6808 10650
rect 6756 10586 6808 10592
rect 7044 10553 7072 10926
rect 7136 10582 7164 10994
rect 7320 10990 7348 11130
rect 7308 10984 7360 10990
rect 7308 10926 7360 10932
rect 7320 10718 7348 10926
rect 7412 10786 7440 11606
rect 7688 11330 7716 11674
rect 7860 11528 7912 11534
rect 7860 11470 7912 11476
rect 7676 11324 7728 11330
rect 7676 11266 7728 11272
rect 7872 11194 7900 11470
rect 7860 11188 7912 11194
rect 7860 11130 7912 11136
rect 8320 11120 8372 11126
rect 8320 11062 8372 11068
rect 7584 11052 7636 11058
rect 7584 10994 7636 11000
rect 7400 10780 7452 10786
rect 7400 10722 7452 10728
rect 7308 10712 7360 10718
rect 7308 10654 7360 10660
rect 7412 10666 7440 10722
rect 7412 10638 7532 10666
rect 7124 10576 7176 10582
rect 7030 10544 7086 10553
rect 7124 10518 7176 10524
rect 7308 10576 7360 10582
rect 7308 10518 7360 10524
rect 7030 10479 7086 10488
rect 6756 10440 6808 10446
rect 6756 10382 6808 10388
rect 6664 10236 6716 10242
rect 6664 10178 6716 10184
rect 6572 10100 6624 10106
rect 6572 10042 6624 10048
rect 6480 9896 6532 9902
rect 6480 9838 6532 9844
rect 6492 9562 6520 9838
rect 6584 9698 6612 10042
rect 6572 9692 6624 9698
rect 6572 9634 6624 9640
rect 6480 9556 6532 9562
rect 6480 9498 6532 9504
rect 6388 9352 6440 9358
rect 6388 9294 6440 9300
rect 4982 9252 5358 9272
rect 5038 9250 5062 9252
rect 5118 9250 5142 9252
rect 5198 9250 5222 9252
rect 5278 9250 5302 9252
rect 5038 9198 5048 9250
rect 5292 9198 5302 9250
rect 5038 9196 5062 9198
rect 5118 9196 5142 9198
rect 5198 9196 5222 9198
rect 5278 9196 5302 9198
rect 4982 9176 5358 9196
rect 6400 9018 6428 9294
rect 6388 9012 6440 9018
rect 6388 8954 6440 8960
rect 6400 8814 6428 8954
rect 6768 8882 6796 10382
rect 6913 10340 7289 10360
rect 6969 10338 6993 10340
rect 7049 10338 7073 10340
rect 7129 10338 7153 10340
rect 7209 10338 7233 10340
rect 6969 10286 6979 10338
rect 7223 10286 7233 10338
rect 6969 10284 6993 10286
rect 7049 10284 7073 10286
rect 7129 10284 7153 10286
rect 7209 10284 7233 10286
rect 6913 10264 7289 10284
rect 6846 10136 6902 10145
rect 7320 10106 7348 10518
rect 7400 10508 7452 10514
rect 7400 10450 7452 10456
rect 7412 10106 7440 10450
rect 6846 10071 6902 10080
rect 7308 10100 7360 10106
rect 6860 9578 6888 10071
rect 7308 10042 7360 10048
rect 7400 10100 7452 10106
rect 7400 10042 7452 10048
rect 6940 9624 6992 9630
rect 6860 9572 6940 9578
rect 6860 9566 6992 9572
rect 6860 9550 6980 9566
rect 6860 9494 6888 9550
rect 6848 9488 6900 9494
rect 6848 9430 6900 9436
rect 6913 9252 7289 9272
rect 6969 9250 6993 9252
rect 7049 9250 7073 9252
rect 7129 9250 7153 9252
rect 7209 9250 7233 9252
rect 6969 9198 6979 9250
rect 7223 9198 7233 9250
rect 6969 9196 6993 9198
rect 7049 9196 7073 9198
rect 7129 9196 7153 9198
rect 7209 9196 7233 9198
rect 6913 9176 7289 9196
rect 7412 9154 7440 10042
rect 7504 10038 7532 10638
rect 7596 10242 7624 10994
rect 7878 10884 8254 10904
rect 7934 10882 7958 10884
rect 8014 10882 8038 10884
rect 8094 10882 8118 10884
rect 8174 10882 8198 10884
rect 7934 10830 7944 10882
rect 8188 10830 8198 10882
rect 7934 10828 7958 10830
rect 8014 10828 8038 10830
rect 8094 10828 8118 10830
rect 8174 10828 8198 10830
rect 7878 10808 8254 10828
rect 7584 10236 7636 10242
rect 7584 10178 7636 10184
rect 7676 10100 7728 10106
rect 7676 10042 7728 10048
rect 7492 10032 7544 10038
rect 7492 9974 7544 9980
rect 7688 9494 7716 10042
rect 7878 9796 8254 9816
rect 7934 9794 7958 9796
rect 8014 9794 8038 9796
rect 8094 9794 8118 9796
rect 8174 9794 8198 9796
rect 7934 9742 7944 9794
rect 8188 9742 8198 9794
rect 7934 9740 7958 9742
rect 8014 9740 8038 9742
rect 8094 9740 8118 9742
rect 8174 9740 8198 9742
rect 7878 9720 8254 9740
rect 8332 9698 8360 11062
rect 9336 10048 10136 10146
rect 9160 10020 10136 10048
rect 8320 9692 8372 9698
rect 8320 9634 8372 9640
rect 7676 9488 7728 9494
rect 7676 9430 7728 9436
rect 7400 9148 7452 9154
rect 7400 9090 7452 9096
rect 6756 8876 6808 8882
rect 6756 8818 6808 8824
rect 6388 8808 6440 8814
rect 6388 8750 6440 8756
rect 4017 8708 4393 8728
rect 4073 8706 4097 8708
rect 4153 8706 4177 8708
rect 4233 8706 4257 8708
rect 4313 8706 4337 8708
rect 4073 8654 4083 8706
rect 4327 8654 4337 8706
rect 4073 8652 4097 8654
rect 4153 8652 4177 8654
rect 4233 8652 4257 8654
rect 4313 8652 4337 8654
rect 4017 8632 4393 8652
rect 5948 8708 6324 8728
rect 6004 8706 6028 8708
rect 6084 8706 6108 8708
rect 6164 8706 6188 8708
rect 6244 8706 6268 8708
rect 6004 8654 6014 8706
rect 6258 8654 6268 8706
rect 6004 8652 6028 8654
rect 6084 8652 6108 8654
rect 6164 8652 6188 8654
rect 6244 8652 6268 8654
rect 5948 8632 6324 8652
rect 4982 8164 5358 8184
rect 5038 8162 5062 8164
rect 5118 8162 5142 8164
rect 5198 8162 5222 8164
rect 5278 8162 5302 8164
rect 5038 8110 5048 8162
rect 5292 8110 5302 8162
rect 5038 8108 5062 8110
rect 5118 8108 5142 8110
rect 5198 8108 5222 8110
rect 5278 8108 5302 8110
rect 4982 8088 5358 8108
rect 4017 7620 4393 7640
rect 4073 7618 4097 7620
rect 4153 7618 4177 7620
rect 4233 7618 4257 7620
rect 4313 7618 4337 7620
rect 4073 7566 4083 7618
rect 4327 7566 4337 7618
rect 4073 7564 4097 7566
rect 4153 7564 4177 7566
rect 4233 7564 4257 7566
rect 4313 7564 4337 7566
rect 4017 7544 4393 7564
rect 5948 7620 6324 7640
rect 6004 7618 6028 7620
rect 6084 7618 6108 7620
rect 6164 7618 6188 7620
rect 6244 7618 6268 7620
rect 6004 7566 6014 7618
rect 6258 7566 6268 7618
rect 6004 7564 6028 7566
rect 6084 7564 6108 7566
rect 6164 7564 6188 7566
rect 6244 7564 6268 7566
rect 5948 7544 6324 7564
rect 4982 7076 5358 7096
rect 5038 7074 5062 7076
rect 5118 7074 5142 7076
rect 5198 7074 5222 7076
rect 5278 7074 5302 7076
rect 5038 7022 5048 7074
rect 5292 7022 5302 7074
rect 5038 7020 5062 7022
rect 5118 7020 5142 7022
rect 5198 7020 5222 7022
rect 5278 7020 5302 7022
rect 4982 7000 5358 7020
rect 6400 6638 6428 8750
rect 6913 8164 7289 8184
rect 6969 8162 6993 8164
rect 7049 8162 7073 8164
rect 7129 8162 7153 8164
rect 7209 8162 7233 8164
rect 6969 8110 6979 8162
rect 7223 8110 7233 8162
rect 6969 8108 6993 8110
rect 7049 8108 7073 8110
rect 7129 8108 7153 8110
rect 7209 8108 7233 8110
rect 6913 8088 7289 8108
rect 6913 7076 7289 7096
rect 6969 7074 6993 7076
rect 7049 7074 7073 7076
rect 7129 7074 7153 7076
rect 7209 7074 7233 7076
rect 6969 7022 6979 7074
rect 7223 7022 7233 7074
rect 6969 7020 6993 7022
rect 7049 7020 7073 7022
rect 7129 7020 7153 7022
rect 7209 7020 7233 7022
rect 6913 7000 7289 7020
rect 3168 6632 3220 6638
rect 3168 6574 3220 6580
rect 6388 6632 6440 6638
rect 6388 6574 6440 6580
rect 2136 4068 2936 4166
rect 3180 4068 3208 6574
rect 4017 6532 4393 6552
rect 4073 6530 4097 6532
rect 4153 6530 4177 6532
rect 4233 6530 4257 6532
rect 4313 6530 4337 6532
rect 4073 6478 4083 6530
rect 4327 6478 4337 6530
rect 4073 6476 4097 6478
rect 4153 6476 4177 6478
rect 4233 6476 4257 6478
rect 4313 6476 4337 6478
rect 4017 6456 4393 6476
rect 5948 6532 6324 6552
rect 6004 6530 6028 6532
rect 6084 6530 6108 6532
rect 6164 6530 6188 6532
rect 6244 6530 6268 6532
rect 6004 6478 6014 6530
rect 6258 6478 6268 6530
rect 6004 6476 6028 6478
rect 6084 6476 6108 6478
rect 6164 6476 6188 6478
rect 6244 6476 6268 6478
rect 5948 6456 6324 6476
rect 4982 5988 5358 6008
rect 5038 5986 5062 5988
rect 5118 5986 5142 5988
rect 5198 5986 5222 5988
rect 5278 5986 5302 5988
rect 5038 5934 5048 5986
rect 5292 5934 5302 5986
rect 5038 5932 5062 5934
rect 5118 5932 5142 5934
rect 5198 5932 5222 5934
rect 5278 5932 5302 5934
rect 4982 5912 5358 5932
rect 6913 5988 7289 6008
rect 6969 5986 6993 5988
rect 7049 5986 7073 5988
rect 7129 5986 7153 5988
rect 7209 5986 7233 5988
rect 6969 5934 6979 5986
rect 7223 5934 7233 5986
rect 6969 5932 6993 5934
rect 7049 5932 7073 5934
rect 7129 5932 7153 5934
rect 7209 5932 7233 5934
rect 6913 5912 7289 5932
rect 4017 5444 4393 5464
rect 4073 5442 4097 5444
rect 4153 5442 4177 5444
rect 4233 5442 4257 5444
rect 4313 5442 4337 5444
rect 4073 5390 4083 5442
rect 4327 5390 4337 5442
rect 4073 5388 4097 5390
rect 4153 5388 4177 5390
rect 4233 5388 4257 5390
rect 4313 5388 4337 5390
rect 4017 5368 4393 5388
rect 5948 5444 6324 5464
rect 6004 5442 6028 5444
rect 6084 5442 6108 5444
rect 6164 5442 6188 5444
rect 6244 5442 6268 5444
rect 6004 5390 6014 5442
rect 6258 5390 6268 5442
rect 6004 5388 6028 5390
rect 6084 5388 6108 5390
rect 6164 5388 6188 5390
rect 6244 5388 6268 5390
rect 5948 5368 6324 5388
rect 4982 4900 5358 4920
rect 5038 4898 5062 4900
rect 5118 4898 5142 4900
rect 5198 4898 5222 4900
rect 5278 4898 5302 4900
rect 5038 4846 5048 4898
rect 5292 4846 5302 4898
rect 5038 4844 5062 4846
rect 5118 4844 5142 4846
rect 5198 4844 5222 4846
rect 5278 4844 5302 4846
rect 4982 4824 5358 4844
rect 6913 4900 7289 4920
rect 6969 4898 6993 4900
rect 7049 4898 7073 4900
rect 7129 4898 7153 4900
rect 7209 4898 7233 4900
rect 6969 4846 6979 4898
rect 7223 4846 7233 4898
rect 6969 4844 6993 4846
rect 7049 4844 7073 4846
rect 7129 4844 7153 4846
rect 7209 4844 7233 4846
rect 6913 4824 7289 4844
rect 7688 4802 7716 9430
rect 9160 9018 9188 10020
rect 9336 9922 10136 10020
rect 9148 9012 9200 9018
rect 9148 8954 9200 8960
rect 7878 8708 8254 8728
rect 7934 8706 7958 8708
rect 8014 8706 8038 8708
rect 8094 8706 8118 8708
rect 8174 8706 8198 8708
rect 7934 8654 7944 8706
rect 8188 8654 8198 8706
rect 7934 8652 7958 8654
rect 8014 8652 8038 8654
rect 8094 8652 8118 8654
rect 8174 8652 8198 8654
rect 7878 8632 8254 8652
rect 7878 7620 8254 7640
rect 7934 7618 7958 7620
rect 8014 7618 8038 7620
rect 8094 7618 8118 7620
rect 8174 7618 8198 7620
rect 7934 7566 7944 7618
rect 8188 7566 8198 7618
rect 7934 7564 7958 7566
rect 8014 7564 8038 7566
rect 8094 7564 8118 7566
rect 8174 7564 8198 7566
rect 7878 7544 8254 7564
rect 7878 6532 8254 6552
rect 7934 6530 7958 6532
rect 8014 6530 8038 6532
rect 8094 6530 8118 6532
rect 8174 6530 8198 6532
rect 7934 6478 7944 6530
rect 8188 6478 8198 6530
rect 7934 6476 7958 6478
rect 8014 6476 8038 6478
rect 8094 6476 8118 6478
rect 8174 6476 8198 6478
rect 7878 6456 8254 6476
rect 7878 5444 8254 5464
rect 7934 5442 7958 5444
rect 8014 5442 8038 5444
rect 8094 5442 8118 5444
rect 8174 5442 8198 5444
rect 7934 5390 7944 5442
rect 8188 5390 8198 5442
rect 7934 5388 7958 5390
rect 8014 5388 8038 5390
rect 8094 5388 8118 5390
rect 8174 5388 8198 5390
rect 7878 5368 8254 5388
rect 7676 4796 7728 4802
rect 7676 4738 7728 4744
rect 9148 4660 9200 4666
rect 9148 4602 9200 4608
rect 4017 4356 4393 4376
rect 4073 4354 4097 4356
rect 4153 4354 4177 4356
rect 4233 4354 4257 4356
rect 4313 4354 4337 4356
rect 4073 4302 4083 4354
rect 4327 4302 4337 4354
rect 4073 4300 4097 4302
rect 4153 4300 4177 4302
rect 4233 4300 4257 4302
rect 4313 4300 4337 4302
rect 4017 4280 4393 4300
rect 5948 4356 6324 4376
rect 6004 4354 6028 4356
rect 6084 4354 6108 4356
rect 6164 4354 6188 4356
rect 6244 4354 6268 4356
rect 6004 4302 6014 4354
rect 6258 4302 6268 4354
rect 6004 4300 6028 4302
rect 6084 4300 6108 4302
rect 6164 4300 6188 4302
rect 6244 4300 6268 4302
rect 5948 4280 6324 4300
rect 7878 4356 8254 4376
rect 7934 4354 7958 4356
rect 8014 4354 8038 4356
rect 8094 4354 8118 4356
rect 8174 4354 8198 4356
rect 7934 4302 7944 4354
rect 8188 4302 8198 4354
rect 7934 4300 7958 4302
rect 8014 4300 8038 4302
rect 8094 4300 8118 4302
rect 8174 4300 8198 4302
rect 7878 4280 8254 4300
rect 2136 4040 3208 4068
rect 9160 4068 9188 4602
rect 9336 4068 10136 4166
rect 9160 4040 10136 4068
rect 2136 3942 2936 4040
rect 9336 3942 10136 4040
rect 4982 3812 5358 3832
rect 5038 3810 5062 3812
rect 5118 3810 5142 3812
rect 5198 3810 5222 3812
rect 5278 3810 5302 3812
rect 5038 3758 5048 3810
rect 5292 3758 5302 3810
rect 5038 3756 5062 3758
rect 5118 3756 5142 3758
rect 5198 3756 5222 3758
rect 5278 3756 5302 3758
rect 4982 3736 5358 3756
rect 6913 3812 7289 3832
rect 6969 3810 6993 3812
rect 7049 3810 7073 3812
rect 7129 3810 7153 3812
rect 7209 3810 7233 3812
rect 6969 3758 6979 3810
rect 7223 3758 7233 3810
rect 6969 3756 6993 3758
rect 7049 3756 7073 3758
rect 7129 3756 7153 3758
rect 7209 3756 7233 3758
rect 6913 3736 7289 3756
rect 4017 3268 4393 3288
rect 4073 3266 4097 3268
rect 4153 3266 4177 3268
rect 4233 3266 4257 3268
rect 4313 3266 4337 3268
rect 4073 3214 4083 3266
rect 4327 3214 4337 3266
rect 4073 3212 4097 3214
rect 4153 3212 4177 3214
rect 4233 3212 4257 3214
rect 4313 3212 4337 3214
rect 4017 3192 4393 3212
rect 5948 3268 6324 3288
rect 6004 3266 6028 3268
rect 6084 3266 6108 3268
rect 6164 3266 6188 3268
rect 6244 3266 6268 3268
rect 6004 3214 6014 3266
rect 6258 3214 6268 3266
rect 6004 3212 6028 3214
rect 6084 3212 6108 3214
rect 6164 3212 6188 3214
rect 6244 3212 6268 3214
rect 5948 3192 6324 3212
rect 7878 3268 8254 3288
rect 7934 3266 7958 3268
rect 8014 3266 8038 3268
rect 8094 3266 8118 3268
rect 8174 3266 8198 3268
rect 7934 3214 7944 3266
rect 8188 3214 8198 3266
rect 7934 3212 7958 3214
rect 8014 3212 8038 3214
rect 8094 3212 8118 3214
rect 8174 3212 8198 3214
rect 7878 3192 8254 3212
<< via2 >>
rect 4982 16866 5038 16868
rect 5062 16866 5118 16868
rect 5142 16866 5198 16868
rect 5222 16866 5278 16868
rect 5302 16866 5358 16868
rect 4982 16814 4984 16866
rect 4984 16814 5036 16866
rect 5036 16814 5038 16866
rect 5062 16814 5100 16866
rect 5100 16814 5112 16866
rect 5112 16814 5118 16866
rect 5142 16814 5164 16866
rect 5164 16814 5176 16866
rect 5176 16814 5198 16866
rect 5222 16814 5228 16866
rect 5228 16814 5240 16866
rect 5240 16814 5278 16866
rect 5302 16814 5304 16866
rect 5304 16814 5356 16866
rect 5356 16814 5358 16866
rect 4982 16812 5038 16814
rect 5062 16812 5118 16814
rect 5142 16812 5198 16814
rect 5222 16812 5278 16814
rect 5302 16812 5358 16814
rect 6913 16866 6969 16868
rect 6993 16866 7049 16868
rect 7073 16866 7129 16868
rect 7153 16866 7209 16868
rect 7233 16866 7289 16868
rect 6913 16814 6915 16866
rect 6915 16814 6967 16866
rect 6967 16814 6969 16866
rect 6993 16814 7031 16866
rect 7031 16814 7043 16866
rect 7043 16814 7049 16866
rect 7073 16814 7095 16866
rect 7095 16814 7107 16866
rect 7107 16814 7129 16866
rect 7153 16814 7159 16866
rect 7159 16814 7171 16866
rect 7171 16814 7209 16866
rect 7233 16814 7235 16866
rect 7235 16814 7287 16866
rect 7287 16814 7289 16866
rect 6913 16812 6969 16814
rect 6993 16812 7049 16814
rect 7073 16812 7129 16814
rect 7153 16812 7209 16814
rect 7233 16812 7289 16814
rect 4017 16322 4073 16324
rect 4097 16322 4153 16324
rect 4177 16322 4233 16324
rect 4257 16322 4313 16324
rect 4337 16322 4393 16324
rect 4017 16270 4019 16322
rect 4019 16270 4071 16322
rect 4071 16270 4073 16322
rect 4097 16270 4135 16322
rect 4135 16270 4147 16322
rect 4147 16270 4153 16322
rect 4177 16270 4199 16322
rect 4199 16270 4211 16322
rect 4211 16270 4233 16322
rect 4257 16270 4263 16322
rect 4263 16270 4275 16322
rect 4275 16270 4313 16322
rect 4337 16270 4339 16322
rect 4339 16270 4391 16322
rect 4391 16270 4393 16322
rect 4017 16268 4073 16270
rect 4097 16268 4153 16270
rect 4177 16268 4233 16270
rect 4257 16268 4313 16270
rect 4337 16268 4393 16270
rect 5948 16322 6004 16324
rect 6028 16322 6084 16324
rect 6108 16322 6164 16324
rect 6188 16322 6244 16324
rect 6268 16322 6324 16324
rect 5948 16270 5950 16322
rect 5950 16270 6002 16322
rect 6002 16270 6004 16322
rect 6028 16270 6066 16322
rect 6066 16270 6078 16322
rect 6078 16270 6084 16322
rect 6108 16270 6130 16322
rect 6130 16270 6142 16322
rect 6142 16270 6164 16322
rect 6188 16270 6194 16322
rect 6194 16270 6206 16322
rect 6206 16270 6244 16322
rect 6268 16270 6270 16322
rect 6270 16270 6322 16322
rect 6322 16270 6324 16322
rect 5948 16268 6004 16270
rect 6028 16268 6084 16270
rect 6108 16268 6164 16270
rect 6188 16268 6244 16270
rect 6268 16268 6324 16270
rect 7878 16322 7934 16324
rect 7958 16322 8014 16324
rect 8038 16322 8094 16324
rect 8118 16322 8174 16324
rect 8198 16322 8254 16324
rect 7878 16270 7880 16322
rect 7880 16270 7932 16322
rect 7932 16270 7934 16322
rect 7958 16270 7996 16322
rect 7996 16270 8008 16322
rect 8008 16270 8014 16322
rect 8038 16270 8060 16322
rect 8060 16270 8072 16322
rect 8072 16270 8094 16322
rect 8118 16270 8124 16322
rect 8124 16270 8136 16322
rect 8136 16270 8174 16322
rect 8198 16270 8200 16322
rect 8200 16270 8252 16322
rect 8252 16270 8254 16322
rect 7878 16268 7934 16270
rect 7958 16268 8014 16270
rect 8038 16268 8094 16270
rect 8118 16268 8174 16270
rect 8198 16268 8254 16270
rect 4982 15778 5038 15780
rect 5062 15778 5118 15780
rect 5142 15778 5198 15780
rect 5222 15778 5278 15780
rect 5302 15778 5358 15780
rect 4982 15726 4984 15778
rect 4984 15726 5036 15778
rect 5036 15726 5038 15778
rect 5062 15726 5100 15778
rect 5100 15726 5112 15778
rect 5112 15726 5118 15778
rect 5142 15726 5164 15778
rect 5164 15726 5176 15778
rect 5176 15726 5198 15778
rect 5222 15726 5228 15778
rect 5228 15726 5240 15778
rect 5240 15726 5278 15778
rect 5302 15726 5304 15778
rect 5304 15726 5356 15778
rect 5356 15726 5358 15778
rect 4982 15724 5038 15726
rect 5062 15724 5118 15726
rect 5142 15724 5198 15726
rect 5222 15724 5278 15726
rect 5302 15724 5358 15726
rect 4017 15234 4073 15236
rect 4097 15234 4153 15236
rect 4177 15234 4233 15236
rect 4257 15234 4313 15236
rect 4337 15234 4393 15236
rect 4017 15182 4019 15234
rect 4019 15182 4071 15234
rect 4071 15182 4073 15234
rect 4097 15182 4135 15234
rect 4135 15182 4147 15234
rect 4147 15182 4153 15234
rect 4177 15182 4199 15234
rect 4199 15182 4211 15234
rect 4211 15182 4233 15234
rect 4257 15182 4263 15234
rect 4263 15182 4275 15234
rect 4275 15182 4313 15234
rect 4337 15182 4339 15234
rect 4339 15182 4391 15234
rect 4391 15182 4393 15234
rect 4017 15180 4073 15182
rect 4097 15180 4153 15182
rect 4177 15180 4233 15182
rect 4257 15180 4313 15182
rect 4337 15180 4393 15182
rect 5948 15234 6004 15236
rect 6028 15234 6084 15236
rect 6108 15234 6164 15236
rect 6188 15234 6244 15236
rect 6268 15234 6324 15236
rect 5948 15182 5950 15234
rect 5950 15182 6002 15234
rect 6002 15182 6004 15234
rect 6028 15182 6066 15234
rect 6066 15182 6078 15234
rect 6078 15182 6084 15234
rect 6108 15182 6130 15234
rect 6130 15182 6142 15234
rect 6142 15182 6164 15234
rect 6188 15182 6194 15234
rect 6194 15182 6206 15234
rect 6206 15182 6244 15234
rect 6268 15182 6270 15234
rect 6270 15182 6322 15234
rect 6322 15182 6324 15234
rect 5948 15180 6004 15182
rect 6028 15180 6084 15182
rect 6108 15180 6164 15182
rect 6188 15180 6244 15182
rect 6268 15180 6324 15182
rect 4982 14690 5038 14692
rect 5062 14690 5118 14692
rect 5142 14690 5198 14692
rect 5222 14690 5278 14692
rect 5302 14690 5358 14692
rect 4982 14638 4984 14690
rect 4984 14638 5036 14690
rect 5036 14638 5038 14690
rect 5062 14638 5100 14690
rect 5100 14638 5112 14690
rect 5112 14638 5118 14690
rect 5142 14638 5164 14690
rect 5164 14638 5176 14690
rect 5176 14638 5198 14690
rect 5222 14638 5228 14690
rect 5228 14638 5240 14690
rect 5240 14638 5278 14690
rect 5302 14638 5304 14690
rect 5304 14638 5356 14690
rect 5356 14638 5358 14690
rect 4982 14636 5038 14638
rect 5062 14636 5118 14638
rect 5142 14636 5198 14638
rect 5222 14636 5278 14638
rect 5302 14636 5358 14638
rect 4017 14146 4073 14148
rect 4097 14146 4153 14148
rect 4177 14146 4233 14148
rect 4257 14146 4313 14148
rect 4337 14146 4393 14148
rect 4017 14094 4019 14146
rect 4019 14094 4071 14146
rect 4071 14094 4073 14146
rect 4097 14094 4135 14146
rect 4135 14094 4147 14146
rect 4147 14094 4153 14146
rect 4177 14094 4199 14146
rect 4199 14094 4211 14146
rect 4211 14094 4233 14146
rect 4257 14094 4263 14146
rect 4263 14094 4275 14146
rect 4275 14094 4313 14146
rect 4337 14094 4339 14146
rect 4339 14094 4391 14146
rect 4391 14094 4393 14146
rect 4017 14092 4073 14094
rect 4097 14092 4153 14094
rect 4177 14092 4233 14094
rect 4257 14092 4313 14094
rect 4337 14092 4393 14094
rect 5948 14146 6004 14148
rect 6028 14146 6084 14148
rect 6108 14146 6164 14148
rect 6188 14146 6244 14148
rect 6268 14146 6324 14148
rect 5948 14094 5950 14146
rect 5950 14094 6002 14146
rect 6002 14094 6004 14146
rect 6028 14094 6066 14146
rect 6066 14094 6078 14146
rect 6078 14094 6084 14146
rect 6108 14094 6130 14146
rect 6130 14094 6142 14146
rect 6142 14094 6164 14146
rect 6188 14094 6194 14146
rect 6194 14094 6206 14146
rect 6206 14094 6244 14146
rect 6268 14094 6270 14146
rect 6270 14094 6322 14146
rect 6322 14094 6324 14146
rect 5948 14092 6004 14094
rect 6028 14092 6084 14094
rect 6108 14092 6164 14094
rect 6188 14092 6244 14094
rect 6268 14092 6324 14094
rect 4982 13602 5038 13604
rect 5062 13602 5118 13604
rect 5142 13602 5198 13604
rect 5222 13602 5278 13604
rect 5302 13602 5358 13604
rect 4982 13550 4984 13602
rect 4984 13550 5036 13602
rect 5036 13550 5038 13602
rect 5062 13550 5100 13602
rect 5100 13550 5112 13602
rect 5112 13550 5118 13602
rect 5142 13550 5164 13602
rect 5164 13550 5176 13602
rect 5176 13550 5198 13602
rect 5222 13550 5228 13602
rect 5228 13550 5240 13602
rect 5240 13550 5278 13602
rect 5302 13550 5304 13602
rect 5304 13550 5356 13602
rect 5356 13550 5358 13602
rect 4982 13548 5038 13550
rect 5062 13548 5118 13550
rect 5142 13548 5198 13550
rect 5222 13548 5278 13550
rect 5302 13548 5358 13550
rect 4017 13058 4073 13060
rect 4097 13058 4153 13060
rect 4177 13058 4233 13060
rect 4257 13058 4313 13060
rect 4337 13058 4393 13060
rect 4017 13006 4019 13058
rect 4019 13006 4071 13058
rect 4071 13006 4073 13058
rect 4097 13006 4135 13058
rect 4135 13006 4147 13058
rect 4147 13006 4153 13058
rect 4177 13006 4199 13058
rect 4199 13006 4211 13058
rect 4211 13006 4233 13058
rect 4257 13006 4263 13058
rect 4263 13006 4275 13058
rect 4275 13006 4313 13058
rect 4337 13006 4339 13058
rect 4339 13006 4391 13058
rect 4391 13006 4393 13058
rect 4017 13004 4073 13006
rect 4097 13004 4153 13006
rect 4177 13004 4233 13006
rect 4257 13004 4313 13006
rect 4337 13004 4393 13006
rect 5948 13058 6004 13060
rect 6028 13058 6084 13060
rect 6108 13058 6164 13060
rect 6188 13058 6244 13060
rect 6268 13058 6324 13060
rect 5948 13006 5950 13058
rect 5950 13006 6002 13058
rect 6002 13006 6004 13058
rect 6028 13006 6066 13058
rect 6066 13006 6078 13058
rect 6078 13006 6084 13058
rect 6108 13006 6130 13058
rect 6130 13006 6142 13058
rect 6142 13006 6164 13058
rect 6188 13006 6194 13058
rect 6194 13006 6206 13058
rect 6206 13006 6244 13058
rect 6268 13006 6270 13058
rect 6270 13006 6322 13058
rect 6322 13006 6324 13058
rect 5948 13004 6004 13006
rect 6028 13004 6084 13006
rect 6108 13004 6164 13006
rect 6188 13004 6244 13006
rect 6268 13004 6324 13006
rect 4982 12514 5038 12516
rect 5062 12514 5118 12516
rect 5142 12514 5198 12516
rect 5222 12514 5278 12516
rect 5302 12514 5358 12516
rect 4982 12462 4984 12514
rect 4984 12462 5036 12514
rect 5036 12462 5038 12514
rect 5062 12462 5100 12514
rect 5100 12462 5112 12514
rect 5112 12462 5118 12514
rect 5142 12462 5164 12514
rect 5164 12462 5176 12514
rect 5176 12462 5198 12514
rect 5222 12462 5228 12514
rect 5228 12462 5240 12514
rect 5240 12462 5278 12514
rect 5302 12462 5304 12514
rect 5304 12462 5356 12514
rect 5356 12462 5358 12514
rect 4982 12460 5038 12462
rect 5062 12460 5118 12462
rect 5142 12460 5198 12462
rect 5222 12460 5278 12462
rect 5302 12460 5358 12462
rect 4017 11970 4073 11972
rect 4097 11970 4153 11972
rect 4177 11970 4233 11972
rect 4257 11970 4313 11972
rect 4337 11970 4393 11972
rect 4017 11918 4019 11970
rect 4019 11918 4071 11970
rect 4071 11918 4073 11970
rect 4097 11918 4135 11970
rect 4135 11918 4147 11970
rect 4147 11918 4153 11970
rect 4177 11918 4199 11970
rect 4199 11918 4211 11970
rect 4211 11918 4233 11970
rect 4257 11918 4263 11970
rect 4263 11918 4275 11970
rect 4275 11918 4313 11970
rect 4337 11918 4339 11970
rect 4339 11918 4391 11970
rect 4391 11918 4393 11970
rect 4017 11916 4073 11918
rect 4097 11916 4153 11918
rect 4177 11916 4233 11918
rect 4257 11916 4313 11918
rect 4337 11916 4393 11918
rect 5948 11970 6004 11972
rect 6028 11970 6084 11972
rect 6108 11970 6164 11972
rect 6188 11970 6244 11972
rect 6268 11970 6324 11972
rect 5948 11918 5950 11970
rect 5950 11918 6002 11970
rect 6002 11918 6004 11970
rect 6028 11918 6066 11970
rect 6066 11918 6078 11970
rect 6078 11918 6084 11970
rect 6108 11918 6130 11970
rect 6130 11918 6142 11970
rect 6142 11918 6164 11970
rect 6188 11918 6194 11970
rect 6194 11918 6206 11970
rect 6206 11918 6244 11970
rect 6268 11918 6270 11970
rect 6270 11918 6322 11970
rect 6322 11918 6324 11970
rect 5948 11916 6004 11918
rect 6028 11916 6084 11918
rect 6108 11916 6164 11918
rect 6188 11916 6244 11918
rect 6268 11916 6324 11918
rect 4982 11426 5038 11428
rect 5062 11426 5118 11428
rect 5142 11426 5198 11428
rect 5222 11426 5278 11428
rect 5302 11426 5358 11428
rect 4982 11374 4984 11426
rect 4984 11374 5036 11426
rect 5036 11374 5038 11426
rect 5062 11374 5100 11426
rect 5100 11374 5112 11426
rect 5112 11374 5118 11426
rect 5142 11374 5164 11426
rect 5164 11374 5176 11426
rect 5176 11374 5198 11426
rect 5222 11374 5228 11426
rect 5228 11374 5240 11426
rect 5240 11374 5278 11426
rect 5302 11374 5304 11426
rect 5304 11374 5356 11426
rect 5356 11374 5358 11426
rect 4982 11372 5038 11374
rect 5062 11372 5118 11374
rect 5142 11372 5198 11374
rect 5222 11372 5278 11374
rect 5302 11372 5358 11374
rect 4017 10882 4073 10884
rect 4097 10882 4153 10884
rect 4177 10882 4233 10884
rect 4257 10882 4313 10884
rect 4337 10882 4393 10884
rect 4017 10830 4019 10882
rect 4019 10830 4071 10882
rect 4071 10830 4073 10882
rect 4097 10830 4135 10882
rect 4135 10830 4147 10882
rect 4147 10830 4153 10882
rect 4177 10830 4199 10882
rect 4199 10830 4211 10882
rect 4211 10830 4233 10882
rect 4257 10830 4263 10882
rect 4263 10830 4275 10882
rect 4275 10830 4313 10882
rect 4337 10830 4339 10882
rect 4339 10830 4391 10882
rect 4391 10830 4393 10882
rect 4017 10828 4073 10830
rect 4097 10828 4153 10830
rect 4177 10828 4233 10830
rect 4257 10828 4313 10830
rect 4337 10828 4393 10830
rect 5948 10882 6004 10884
rect 6028 10882 6084 10884
rect 6108 10882 6164 10884
rect 6188 10882 6244 10884
rect 6268 10882 6324 10884
rect 5948 10830 5950 10882
rect 5950 10830 6002 10882
rect 6002 10830 6004 10882
rect 6028 10830 6066 10882
rect 6066 10830 6078 10882
rect 6078 10830 6084 10882
rect 6108 10830 6130 10882
rect 6130 10830 6142 10882
rect 6142 10830 6164 10882
rect 6188 10830 6194 10882
rect 6194 10830 6206 10882
rect 6206 10830 6244 10882
rect 6268 10830 6270 10882
rect 6270 10830 6322 10882
rect 6322 10830 6324 10882
rect 5948 10828 6004 10830
rect 6028 10828 6084 10830
rect 6108 10828 6164 10830
rect 6188 10828 6244 10830
rect 6268 10828 6324 10830
rect 4982 10338 5038 10340
rect 5062 10338 5118 10340
rect 5142 10338 5198 10340
rect 5222 10338 5278 10340
rect 5302 10338 5358 10340
rect 4982 10286 4984 10338
rect 4984 10286 5036 10338
rect 5036 10286 5038 10338
rect 5062 10286 5100 10338
rect 5100 10286 5112 10338
rect 5112 10286 5118 10338
rect 5142 10286 5164 10338
rect 5164 10286 5176 10338
rect 5176 10286 5198 10338
rect 5222 10286 5228 10338
rect 5228 10286 5240 10338
rect 5240 10286 5278 10338
rect 5302 10286 5304 10338
rect 5304 10286 5356 10338
rect 5356 10286 5358 10338
rect 4982 10284 5038 10286
rect 5062 10284 5118 10286
rect 5142 10284 5198 10286
rect 5222 10284 5278 10286
rect 5302 10284 5358 10286
rect 4017 9794 4073 9796
rect 4097 9794 4153 9796
rect 4177 9794 4233 9796
rect 4257 9794 4313 9796
rect 4337 9794 4393 9796
rect 4017 9742 4019 9794
rect 4019 9742 4071 9794
rect 4071 9742 4073 9794
rect 4097 9742 4135 9794
rect 4135 9742 4147 9794
rect 4147 9742 4153 9794
rect 4177 9742 4199 9794
rect 4199 9742 4211 9794
rect 4211 9742 4233 9794
rect 4257 9742 4263 9794
rect 4263 9742 4275 9794
rect 4275 9742 4313 9794
rect 4337 9742 4339 9794
rect 4339 9742 4391 9794
rect 4391 9742 4393 9794
rect 4017 9740 4073 9742
rect 4097 9740 4153 9742
rect 4177 9740 4233 9742
rect 4257 9740 4313 9742
rect 4337 9740 4393 9742
rect 5948 9794 6004 9796
rect 6028 9794 6084 9796
rect 6108 9794 6164 9796
rect 6188 9794 6244 9796
rect 6268 9794 6324 9796
rect 5948 9742 5950 9794
rect 5950 9742 6002 9794
rect 6002 9742 6004 9794
rect 6028 9742 6066 9794
rect 6066 9742 6078 9794
rect 6078 9742 6084 9794
rect 6108 9742 6130 9794
rect 6130 9742 6142 9794
rect 6142 9742 6164 9794
rect 6188 9742 6194 9794
rect 6194 9742 6206 9794
rect 6206 9742 6244 9794
rect 6268 9742 6270 9794
rect 6270 9742 6322 9794
rect 6322 9742 6324 9794
rect 5948 9740 6004 9742
rect 6028 9740 6084 9742
rect 6108 9740 6164 9742
rect 6188 9740 6244 9742
rect 6268 9740 6324 9742
rect 6913 15778 6969 15780
rect 6993 15778 7049 15780
rect 7073 15778 7129 15780
rect 7153 15778 7209 15780
rect 7233 15778 7289 15780
rect 6913 15726 6915 15778
rect 6915 15726 6967 15778
rect 6967 15726 6969 15778
rect 6993 15726 7031 15778
rect 7031 15726 7043 15778
rect 7043 15726 7049 15778
rect 7073 15726 7095 15778
rect 7095 15726 7107 15778
rect 7107 15726 7129 15778
rect 7153 15726 7159 15778
rect 7159 15726 7171 15778
rect 7171 15726 7209 15778
rect 7233 15726 7235 15778
rect 7235 15726 7287 15778
rect 7287 15726 7289 15778
rect 6913 15724 6969 15726
rect 6993 15724 7049 15726
rect 7073 15724 7129 15726
rect 7153 15724 7209 15726
rect 7233 15724 7289 15726
rect 6913 14690 6969 14692
rect 6993 14690 7049 14692
rect 7073 14690 7129 14692
rect 7153 14690 7209 14692
rect 7233 14690 7289 14692
rect 6913 14638 6915 14690
rect 6915 14638 6967 14690
rect 6967 14638 6969 14690
rect 6993 14638 7031 14690
rect 7031 14638 7043 14690
rect 7043 14638 7049 14690
rect 7073 14638 7095 14690
rect 7095 14638 7107 14690
rect 7107 14638 7129 14690
rect 7153 14638 7159 14690
rect 7159 14638 7171 14690
rect 7171 14638 7209 14690
rect 7233 14638 7235 14690
rect 7235 14638 7287 14690
rect 7287 14638 7289 14690
rect 6913 14636 6969 14638
rect 6993 14636 7049 14638
rect 7073 14636 7129 14638
rect 7153 14636 7209 14638
rect 7233 14636 7289 14638
rect 6913 13602 6969 13604
rect 6993 13602 7049 13604
rect 7073 13602 7129 13604
rect 7153 13602 7209 13604
rect 7233 13602 7289 13604
rect 6913 13550 6915 13602
rect 6915 13550 6967 13602
rect 6967 13550 6969 13602
rect 6993 13550 7031 13602
rect 7031 13550 7043 13602
rect 7043 13550 7049 13602
rect 7073 13550 7095 13602
rect 7095 13550 7107 13602
rect 7107 13550 7129 13602
rect 7153 13550 7159 13602
rect 7159 13550 7171 13602
rect 7171 13550 7209 13602
rect 7233 13550 7235 13602
rect 7235 13550 7287 13602
rect 7287 13550 7289 13602
rect 6913 13548 6969 13550
rect 6993 13548 7049 13550
rect 7073 13548 7129 13550
rect 7153 13548 7209 13550
rect 7233 13548 7289 13550
rect 6913 12514 6969 12516
rect 6993 12514 7049 12516
rect 7073 12514 7129 12516
rect 7153 12514 7209 12516
rect 7233 12514 7289 12516
rect 6913 12462 6915 12514
rect 6915 12462 6967 12514
rect 6967 12462 6969 12514
rect 6993 12462 7031 12514
rect 7031 12462 7043 12514
rect 7043 12462 7049 12514
rect 7073 12462 7095 12514
rect 7095 12462 7107 12514
rect 7107 12462 7129 12514
rect 7153 12462 7159 12514
rect 7159 12462 7171 12514
rect 7171 12462 7209 12514
rect 7233 12462 7235 12514
rect 7235 12462 7287 12514
rect 7287 12462 7289 12514
rect 6913 12460 6969 12462
rect 6993 12460 7049 12462
rect 7073 12460 7129 12462
rect 7153 12460 7209 12462
rect 7233 12460 7289 12462
rect 7878 15234 7934 15236
rect 7958 15234 8014 15236
rect 8038 15234 8094 15236
rect 8118 15234 8174 15236
rect 8198 15234 8254 15236
rect 7878 15182 7880 15234
rect 7880 15182 7932 15234
rect 7932 15182 7934 15234
rect 7958 15182 7996 15234
rect 7996 15182 8008 15234
rect 8008 15182 8014 15234
rect 8038 15182 8060 15234
rect 8060 15182 8072 15234
rect 8072 15182 8094 15234
rect 8118 15182 8124 15234
rect 8124 15182 8136 15234
rect 8136 15182 8174 15234
rect 8198 15182 8200 15234
rect 8200 15182 8252 15234
rect 8252 15182 8254 15234
rect 7878 15180 7934 15182
rect 7958 15180 8014 15182
rect 8038 15180 8094 15182
rect 8118 15180 8174 15182
rect 8198 15180 8254 15182
rect 7878 14146 7934 14148
rect 7958 14146 8014 14148
rect 8038 14146 8094 14148
rect 8118 14146 8174 14148
rect 8198 14146 8254 14148
rect 7878 14094 7880 14146
rect 7880 14094 7932 14146
rect 7932 14094 7934 14146
rect 7958 14094 7996 14146
rect 7996 14094 8008 14146
rect 8008 14094 8014 14146
rect 8038 14094 8060 14146
rect 8060 14094 8072 14146
rect 8072 14094 8094 14146
rect 8118 14094 8124 14146
rect 8124 14094 8136 14146
rect 8136 14094 8174 14146
rect 8198 14094 8200 14146
rect 8200 14094 8252 14146
rect 8252 14094 8254 14146
rect 7878 14092 7934 14094
rect 7958 14092 8014 14094
rect 8038 14092 8094 14094
rect 8118 14092 8174 14094
rect 8198 14092 8254 14094
rect 7878 13058 7934 13060
rect 7958 13058 8014 13060
rect 8038 13058 8094 13060
rect 8118 13058 8174 13060
rect 8198 13058 8254 13060
rect 7878 13006 7880 13058
rect 7880 13006 7932 13058
rect 7932 13006 7934 13058
rect 7958 13006 7996 13058
rect 7996 13006 8008 13058
rect 8008 13006 8014 13058
rect 8038 13006 8060 13058
rect 8060 13006 8072 13058
rect 8072 13006 8094 13058
rect 8118 13006 8124 13058
rect 8124 13006 8136 13058
rect 8136 13006 8174 13058
rect 8198 13006 8200 13058
rect 8200 13006 8252 13058
rect 8252 13006 8254 13058
rect 7878 13004 7934 13006
rect 7958 13004 8014 13006
rect 8038 13004 8094 13006
rect 8118 13004 8174 13006
rect 8198 13004 8254 13006
rect 7878 11970 7934 11972
rect 7958 11970 8014 11972
rect 8038 11970 8094 11972
rect 8118 11970 8174 11972
rect 8198 11970 8254 11972
rect 7878 11918 7880 11970
rect 7880 11918 7932 11970
rect 7932 11918 7934 11970
rect 7958 11918 7996 11970
rect 7996 11918 8008 11970
rect 8008 11918 8014 11970
rect 8038 11918 8060 11970
rect 8060 11918 8072 11970
rect 8072 11918 8094 11970
rect 8118 11918 8124 11970
rect 8124 11918 8136 11970
rect 8136 11918 8174 11970
rect 8198 11918 8200 11970
rect 8200 11918 8252 11970
rect 8252 11918 8254 11970
rect 7878 11916 7934 11918
rect 7958 11916 8014 11918
rect 8038 11916 8094 11918
rect 8118 11916 8174 11918
rect 8198 11916 8254 11918
rect 6913 11426 6969 11428
rect 6993 11426 7049 11428
rect 7073 11426 7129 11428
rect 7153 11426 7209 11428
rect 7233 11426 7289 11428
rect 6913 11374 6915 11426
rect 6915 11374 6967 11426
rect 6967 11374 6969 11426
rect 6993 11374 7031 11426
rect 7031 11374 7043 11426
rect 7043 11374 7049 11426
rect 7073 11374 7095 11426
rect 7095 11374 7107 11426
rect 7107 11374 7129 11426
rect 7153 11374 7159 11426
rect 7159 11374 7171 11426
rect 7171 11374 7209 11426
rect 7233 11374 7235 11426
rect 7235 11374 7287 11426
rect 7287 11374 7289 11426
rect 6913 11372 6969 11374
rect 6993 11372 7049 11374
rect 7073 11372 7129 11374
rect 7153 11372 7209 11374
rect 7233 11372 7289 11374
rect 7030 10488 7086 10544
rect 4982 9250 5038 9252
rect 5062 9250 5118 9252
rect 5142 9250 5198 9252
rect 5222 9250 5278 9252
rect 5302 9250 5358 9252
rect 4982 9198 4984 9250
rect 4984 9198 5036 9250
rect 5036 9198 5038 9250
rect 5062 9198 5100 9250
rect 5100 9198 5112 9250
rect 5112 9198 5118 9250
rect 5142 9198 5164 9250
rect 5164 9198 5176 9250
rect 5176 9198 5198 9250
rect 5222 9198 5228 9250
rect 5228 9198 5240 9250
rect 5240 9198 5278 9250
rect 5302 9198 5304 9250
rect 5304 9198 5356 9250
rect 5356 9198 5358 9250
rect 4982 9196 5038 9198
rect 5062 9196 5118 9198
rect 5142 9196 5198 9198
rect 5222 9196 5278 9198
rect 5302 9196 5358 9198
rect 6913 10338 6969 10340
rect 6993 10338 7049 10340
rect 7073 10338 7129 10340
rect 7153 10338 7209 10340
rect 7233 10338 7289 10340
rect 6913 10286 6915 10338
rect 6915 10286 6967 10338
rect 6967 10286 6969 10338
rect 6993 10286 7031 10338
rect 7031 10286 7043 10338
rect 7043 10286 7049 10338
rect 7073 10286 7095 10338
rect 7095 10286 7107 10338
rect 7107 10286 7129 10338
rect 7153 10286 7159 10338
rect 7159 10286 7171 10338
rect 7171 10286 7209 10338
rect 7233 10286 7235 10338
rect 7235 10286 7287 10338
rect 7287 10286 7289 10338
rect 6913 10284 6969 10286
rect 6993 10284 7049 10286
rect 7073 10284 7129 10286
rect 7153 10284 7209 10286
rect 7233 10284 7289 10286
rect 6846 10080 6902 10136
rect 6913 9250 6969 9252
rect 6993 9250 7049 9252
rect 7073 9250 7129 9252
rect 7153 9250 7209 9252
rect 7233 9250 7289 9252
rect 6913 9198 6915 9250
rect 6915 9198 6967 9250
rect 6967 9198 6969 9250
rect 6993 9198 7031 9250
rect 7031 9198 7043 9250
rect 7043 9198 7049 9250
rect 7073 9198 7095 9250
rect 7095 9198 7107 9250
rect 7107 9198 7129 9250
rect 7153 9198 7159 9250
rect 7159 9198 7171 9250
rect 7171 9198 7209 9250
rect 7233 9198 7235 9250
rect 7235 9198 7287 9250
rect 7287 9198 7289 9250
rect 6913 9196 6969 9198
rect 6993 9196 7049 9198
rect 7073 9196 7129 9198
rect 7153 9196 7209 9198
rect 7233 9196 7289 9198
rect 7878 10882 7934 10884
rect 7958 10882 8014 10884
rect 8038 10882 8094 10884
rect 8118 10882 8174 10884
rect 8198 10882 8254 10884
rect 7878 10830 7880 10882
rect 7880 10830 7932 10882
rect 7932 10830 7934 10882
rect 7958 10830 7996 10882
rect 7996 10830 8008 10882
rect 8008 10830 8014 10882
rect 8038 10830 8060 10882
rect 8060 10830 8072 10882
rect 8072 10830 8094 10882
rect 8118 10830 8124 10882
rect 8124 10830 8136 10882
rect 8136 10830 8174 10882
rect 8198 10830 8200 10882
rect 8200 10830 8252 10882
rect 8252 10830 8254 10882
rect 7878 10828 7934 10830
rect 7958 10828 8014 10830
rect 8038 10828 8094 10830
rect 8118 10828 8174 10830
rect 8198 10828 8254 10830
rect 7878 9794 7934 9796
rect 7958 9794 8014 9796
rect 8038 9794 8094 9796
rect 8118 9794 8174 9796
rect 8198 9794 8254 9796
rect 7878 9742 7880 9794
rect 7880 9742 7932 9794
rect 7932 9742 7934 9794
rect 7958 9742 7996 9794
rect 7996 9742 8008 9794
rect 8008 9742 8014 9794
rect 8038 9742 8060 9794
rect 8060 9742 8072 9794
rect 8072 9742 8094 9794
rect 8118 9742 8124 9794
rect 8124 9742 8136 9794
rect 8136 9742 8174 9794
rect 8198 9742 8200 9794
rect 8200 9742 8252 9794
rect 8252 9742 8254 9794
rect 7878 9740 7934 9742
rect 7958 9740 8014 9742
rect 8038 9740 8094 9742
rect 8118 9740 8174 9742
rect 8198 9740 8254 9742
rect 4017 8706 4073 8708
rect 4097 8706 4153 8708
rect 4177 8706 4233 8708
rect 4257 8706 4313 8708
rect 4337 8706 4393 8708
rect 4017 8654 4019 8706
rect 4019 8654 4071 8706
rect 4071 8654 4073 8706
rect 4097 8654 4135 8706
rect 4135 8654 4147 8706
rect 4147 8654 4153 8706
rect 4177 8654 4199 8706
rect 4199 8654 4211 8706
rect 4211 8654 4233 8706
rect 4257 8654 4263 8706
rect 4263 8654 4275 8706
rect 4275 8654 4313 8706
rect 4337 8654 4339 8706
rect 4339 8654 4391 8706
rect 4391 8654 4393 8706
rect 4017 8652 4073 8654
rect 4097 8652 4153 8654
rect 4177 8652 4233 8654
rect 4257 8652 4313 8654
rect 4337 8652 4393 8654
rect 5948 8706 6004 8708
rect 6028 8706 6084 8708
rect 6108 8706 6164 8708
rect 6188 8706 6244 8708
rect 6268 8706 6324 8708
rect 5948 8654 5950 8706
rect 5950 8654 6002 8706
rect 6002 8654 6004 8706
rect 6028 8654 6066 8706
rect 6066 8654 6078 8706
rect 6078 8654 6084 8706
rect 6108 8654 6130 8706
rect 6130 8654 6142 8706
rect 6142 8654 6164 8706
rect 6188 8654 6194 8706
rect 6194 8654 6206 8706
rect 6206 8654 6244 8706
rect 6268 8654 6270 8706
rect 6270 8654 6322 8706
rect 6322 8654 6324 8706
rect 5948 8652 6004 8654
rect 6028 8652 6084 8654
rect 6108 8652 6164 8654
rect 6188 8652 6244 8654
rect 6268 8652 6324 8654
rect 4982 8162 5038 8164
rect 5062 8162 5118 8164
rect 5142 8162 5198 8164
rect 5222 8162 5278 8164
rect 5302 8162 5358 8164
rect 4982 8110 4984 8162
rect 4984 8110 5036 8162
rect 5036 8110 5038 8162
rect 5062 8110 5100 8162
rect 5100 8110 5112 8162
rect 5112 8110 5118 8162
rect 5142 8110 5164 8162
rect 5164 8110 5176 8162
rect 5176 8110 5198 8162
rect 5222 8110 5228 8162
rect 5228 8110 5240 8162
rect 5240 8110 5278 8162
rect 5302 8110 5304 8162
rect 5304 8110 5356 8162
rect 5356 8110 5358 8162
rect 4982 8108 5038 8110
rect 5062 8108 5118 8110
rect 5142 8108 5198 8110
rect 5222 8108 5278 8110
rect 5302 8108 5358 8110
rect 4017 7618 4073 7620
rect 4097 7618 4153 7620
rect 4177 7618 4233 7620
rect 4257 7618 4313 7620
rect 4337 7618 4393 7620
rect 4017 7566 4019 7618
rect 4019 7566 4071 7618
rect 4071 7566 4073 7618
rect 4097 7566 4135 7618
rect 4135 7566 4147 7618
rect 4147 7566 4153 7618
rect 4177 7566 4199 7618
rect 4199 7566 4211 7618
rect 4211 7566 4233 7618
rect 4257 7566 4263 7618
rect 4263 7566 4275 7618
rect 4275 7566 4313 7618
rect 4337 7566 4339 7618
rect 4339 7566 4391 7618
rect 4391 7566 4393 7618
rect 4017 7564 4073 7566
rect 4097 7564 4153 7566
rect 4177 7564 4233 7566
rect 4257 7564 4313 7566
rect 4337 7564 4393 7566
rect 5948 7618 6004 7620
rect 6028 7618 6084 7620
rect 6108 7618 6164 7620
rect 6188 7618 6244 7620
rect 6268 7618 6324 7620
rect 5948 7566 5950 7618
rect 5950 7566 6002 7618
rect 6002 7566 6004 7618
rect 6028 7566 6066 7618
rect 6066 7566 6078 7618
rect 6078 7566 6084 7618
rect 6108 7566 6130 7618
rect 6130 7566 6142 7618
rect 6142 7566 6164 7618
rect 6188 7566 6194 7618
rect 6194 7566 6206 7618
rect 6206 7566 6244 7618
rect 6268 7566 6270 7618
rect 6270 7566 6322 7618
rect 6322 7566 6324 7618
rect 5948 7564 6004 7566
rect 6028 7564 6084 7566
rect 6108 7564 6164 7566
rect 6188 7564 6244 7566
rect 6268 7564 6324 7566
rect 4982 7074 5038 7076
rect 5062 7074 5118 7076
rect 5142 7074 5198 7076
rect 5222 7074 5278 7076
rect 5302 7074 5358 7076
rect 4982 7022 4984 7074
rect 4984 7022 5036 7074
rect 5036 7022 5038 7074
rect 5062 7022 5100 7074
rect 5100 7022 5112 7074
rect 5112 7022 5118 7074
rect 5142 7022 5164 7074
rect 5164 7022 5176 7074
rect 5176 7022 5198 7074
rect 5222 7022 5228 7074
rect 5228 7022 5240 7074
rect 5240 7022 5278 7074
rect 5302 7022 5304 7074
rect 5304 7022 5356 7074
rect 5356 7022 5358 7074
rect 4982 7020 5038 7022
rect 5062 7020 5118 7022
rect 5142 7020 5198 7022
rect 5222 7020 5278 7022
rect 5302 7020 5358 7022
rect 6913 8162 6969 8164
rect 6993 8162 7049 8164
rect 7073 8162 7129 8164
rect 7153 8162 7209 8164
rect 7233 8162 7289 8164
rect 6913 8110 6915 8162
rect 6915 8110 6967 8162
rect 6967 8110 6969 8162
rect 6993 8110 7031 8162
rect 7031 8110 7043 8162
rect 7043 8110 7049 8162
rect 7073 8110 7095 8162
rect 7095 8110 7107 8162
rect 7107 8110 7129 8162
rect 7153 8110 7159 8162
rect 7159 8110 7171 8162
rect 7171 8110 7209 8162
rect 7233 8110 7235 8162
rect 7235 8110 7287 8162
rect 7287 8110 7289 8162
rect 6913 8108 6969 8110
rect 6993 8108 7049 8110
rect 7073 8108 7129 8110
rect 7153 8108 7209 8110
rect 7233 8108 7289 8110
rect 6913 7074 6969 7076
rect 6993 7074 7049 7076
rect 7073 7074 7129 7076
rect 7153 7074 7209 7076
rect 7233 7074 7289 7076
rect 6913 7022 6915 7074
rect 6915 7022 6967 7074
rect 6967 7022 6969 7074
rect 6993 7022 7031 7074
rect 7031 7022 7043 7074
rect 7043 7022 7049 7074
rect 7073 7022 7095 7074
rect 7095 7022 7107 7074
rect 7107 7022 7129 7074
rect 7153 7022 7159 7074
rect 7159 7022 7171 7074
rect 7171 7022 7209 7074
rect 7233 7022 7235 7074
rect 7235 7022 7287 7074
rect 7287 7022 7289 7074
rect 6913 7020 6969 7022
rect 6993 7020 7049 7022
rect 7073 7020 7129 7022
rect 7153 7020 7209 7022
rect 7233 7020 7289 7022
rect 4017 6530 4073 6532
rect 4097 6530 4153 6532
rect 4177 6530 4233 6532
rect 4257 6530 4313 6532
rect 4337 6530 4393 6532
rect 4017 6478 4019 6530
rect 4019 6478 4071 6530
rect 4071 6478 4073 6530
rect 4097 6478 4135 6530
rect 4135 6478 4147 6530
rect 4147 6478 4153 6530
rect 4177 6478 4199 6530
rect 4199 6478 4211 6530
rect 4211 6478 4233 6530
rect 4257 6478 4263 6530
rect 4263 6478 4275 6530
rect 4275 6478 4313 6530
rect 4337 6478 4339 6530
rect 4339 6478 4391 6530
rect 4391 6478 4393 6530
rect 4017 6476 4073 6478
rect 4097 6476 4153 6478
rect 4177 6476 4233 6478
rect 4257 6476 4313 6478
rect 4337 6476 4393 6478
rect 5948 6530 6004 6532
rect 6028 6530 6084 6532
rect 6108 6530 6164 6532
rect 6188 6530 6244 6532
rect 6268 6530 6324 6532
rect 5948 6478 5950 6530
rect 5950 6478 6002 6530
rect 6002 6478 6004 6530
rect 6028 6478 6066 6530
rect 6066 6478 6078 6530
rect 6078 6478 6084 6530
rect 6108 6478 6130 6530
rect 6130 6478 6142 6530
rect 6142 6478 6164 6530
rect 6188 6478 6194 6530
rect 6194 6478 6206 6530
rect 6206 6478 6244 6530
rect 6268 6478 6270 6530
rect 6270 6478 6322 6530
rect 6322 6478 6324 6530
rect 5948 6476 6004 6478
rect 6028 6476 6084 6478
rect 6108 6476 6164 6478
rect 6188 6476 6244 6478
rect 6268 6476 6324 6478
rect 4982 5986 5038 5988
rect 5062 5986 5118 5988
rect 5142 5986 5198 5988
rect 5222 5986 5278 5988
rect 5302 5986 5358 5988
rect 4982 5934 4984 5986
rect 4984 5934 5036 5986
rect 5036 5934 5038 5986
rect 5062 5934 5100 5986
rect 5100 5934 5112 5986
rect 5112 5934 5118 5986
rect 5142 5934 5164 5986
rect 5164 5934 5176 5986
rect 5176 5934 5198 5986
rect 5222 5934 5228 5986
rect 5228 5934 5240 5986
rect 5240 5934 5278 5986
rect 5302 5934 5304 5986
rect 5304 5934 5356 5986
rect 5356 5934 5358 5986
rect 4982 5932 5038 5934
rect 5062 5932 5118 5934
rect 5142 5932 5198 5934
rect 5222 5932 5278 5934
rect 5302 5932 5358 5934
rect 6913 5986 6969 5988
rect 6993 5986 7049 5988
rect 7073 5986 7129 5988
rect 7153 5986 7209 5988
rect 7233 5986 7289 5988
rect 6913 5934 6915 5986
rect 6915 5934 6967 5986
rect 6967 5934 6969 5986
rect 6993 5934 7031 5986
rect 7031 5934 7043 5986
rect 7043 5934 7049 5986
rect 7073 5934 7095 5986
rect 7095 5934 7107 5986
rect 7107 5934 7129 5986
rect 7153 5934 7159 5986
rect 7159 5934 7171 5986
rect 7171 5934 7209 5986
rect 7233 5934 7235 5986
rect 7235 5934 7287 5986
rect 7287 5934 7289 5986
rect 6913 5932 6969 5934
rect 6993 5932 7049 5934
rect 7073 5932 7129 5934
rect 7153 5932 7209 5934
rect 7233 5932 7289 5934
rect 4017 5442 4073 5444
rect 4097 5442 4153 5444
rect 4177 5442 4233 5444
rect 4257 5442 4313 5444
rect 4337 5442 4393 5444
rect 4017 5390 4019 5442
rect 4019 5390 4071 5442
rect 4071 5390 4073 5442
rect 4097 5390 4135 5442
rect 4135 5390 4147 5442
rect 4147 5390 4153 5442
rect 4177 5390 4199 5442
rect 4199 5390 4211 5442
rect 4211 5390 4233 5442
rect 4257 5390 4263 5442
rect 4263 5390 4275 5442
rect 4275 5390 4313 5442
rect 4337 5390 4339 5442
rect 4339 5390 4391 5442
rect 4391 5390 4393 5442
rect 4017 5388 4073 5390
rect 4097 5388 4153 5390
rect 4177 5388 4233 5390
rect 4257 5388 4313 5390
rect 4337 5388 4393 5390
rect 5948 5442 6004 5444
rect 6028 5442 6084 5444
rect 6108 5442 6164 5444
rect 6188 5442 6244 5444
rect 6268 5442 6324 5444
rect 5948 5390 5950 5442
rect 5950 5390 6002 5442
rect 6002 5390 6004 5442
rect 6028 5390 6066 5442
rect 6066 5390 6078 5442
rect 6078 5390 6084 5442
rect 6108 5390 6130 5442
rect 6130 5390 6142 5442
rect 6142 5390 6164 5442
rect 6188 5390 6194 5442
rect 6194 5390 6206 5442
rect 6206 5390 6244 5442
rect 6268 5390 6270 5442
rect 6270 5390 6322 5442
rect 6322 5390 6324 5442
rect 5948 5388 6004 5390
rect 6028 5388 6084 5390
rect 6108 5388 6164 5390
rect 6188 5388 6244 5390
rect 6268 5388 6324 5390
rect 4982 4898 5038 4900
rect 5062 4898 5118 4900
rect 5142 4898 5198 4900
rect 5222 4898 5278 4900
rect 5302 4898 5358 4900
rect 4982 4846 4984 4898
rect 4984 4846 5036 4898
rect 5036 4846 5038 4898
rect 5062 4846 5100 4898
rect 5100 4846 5112 4898
rect 5112 4846 5118 4898
rect 5142 4846 5164 4898
rect 5164 4846 5176 4898
rect 5176 4846 5198 4898
rect 5222 4846 5228 4898
rect 5228 4846 5240 4898
rect 5240 4846 5278 4898
rect 5302 4846 5304 4898
rect 5304 4846 5356 4898
rect 5356 4846 5358 4898
rect 4982 4844 5038 4846
rect 5062 4844 5118 4846
rect 5142 4844 5198 4846
rect 5222 4844 5278 4846
rect 5302 4844 5358 4846
rect 6913 4898 6969 4900
rect 6993 4898 7049 4900
rect 7073 4898 7129 4900
rect 7153 4898 7209 4900
rect 7233 4898 7289 4900
rect 6913 4846 6915 4898
rect 6915 4846 6967 4898
rect 6967 4846 6969 4898
rect 6993 4846 7031 4898
rect 7031 4846 7043 4898
rect 7043 4846 7049 4898
rect 7073 4846 7095 4898
rect 7095 4846 7107 4898
rect 7107 4846 7129 4898
rect 7153 4846 7159 4898
rect 7159 4846 7171 4898
rect 7171 4846 7209 4898
rect 7233 4846 7235 4898
rect 7235 4846 7287 4898
rect 7287 4846 7289 4898
rect 6913 4844 6969 4846
rect 6993 4844 7049 4846
rect 7073 4844 7129 4846
rect 7153 4844 7209 4846
rect 7233 4844 7289 4846
rect 7878 8706 7934 8708
rect 7958 8706 8014 8708
rect 8038 8706 8094 8708
rect 8118 8706 8174 8708
rect 8198 8706 8254 8708
rect 7878 8654 7880 8706
rect 7880 8654 7932 8706
rect 7932 8654 7934 8706
rect 7958 8654 7996 8706
rect 7996 8654 8008 8706
rect 8008 8654 8014 8706
rect 8038 8654 8060 8706
rect 8060 8654 8072 8706
rect 8072 8654 8094 8706
rect 8118 8654 8124 8706
rect 8124 8654 8136 8706
rect 8136 8654 8174 8706
rect 8198 8654 8200 8706
rect 8200 8654 8252 8706
rect 8252 8654 8254 8706
rect 7878 8652 7934 8654
rect 7958 8652 8014 8654
rect 8038 8652 8094 8654
rect 8118 8652 8174 8654
rect 8198 8652 8254 8654
rect 7878 7618 7934 7620
rect 7958 7618 8014 7620
rect 8038 7618 8094 7620
rect 8118 7618 8174 7620
rect 8198 7618 8254 7620
rect 7878 7566 7880 7618
rect 7880 7566 7932 7618
rect 7932 7566 7934 7618
rect 7958 7566 7996 7618
rect 7996 7566 8008 7618
rect 8008 7566 8014 7618
rect 8038 7566 8060 7618
rect 8060 7566 8072 7618
rect 8072 7566 8094 7618
rect 8118 7566 8124 7618
rect 8124 7566 8136 7618
rect 8136 7566 8174 7618
rect 8198 7566 8200 7618
rect 8200 7566 8252 7618
rect 8252 7566 8254 7618
rect 7878 7564 7934 7566
rect 7958 7564 8014 7566
rect 8038 7564 8094 7566
rect 8118 7564 8174 7566
rect 8198 7564 8254 7566
rect 7878 6530 7934 6532
rect 7958 6530 8014 6532
rect 8038 6530 8094 6532
rect 8118 6530 8174 6532
rect 8198 6530 8254 6532
rect 7878 6478 7880 6530
rect 7880 6478 7932 6530
rect 7932 6478 7934 6530
rect 7958 6478 7996 6530
rect 7996 6478 8008 6530
rect 8008 6478 8014 6530
rect 8038 6478 8060 6530
rect 8060 6478 8072 6530
rect 8072 6478 8094 6530
rect 8118 6478 8124 6530
rect 8124 6478 8136 6530
rect 8136 6478 8174 6530
rect 8198 6478 8200 6530
rect 8200 6478 8252 6530
rect 8252 6478 8254 6530
rect 7878 6476 7934 6478
rect 7958 6476 8014 6478
rect 8038 6476 8094 6478
rect 8118 6476 8174 6478
rect 8198 6476 8254 6478
rect 7878 5442 7934 5444
rect 7958 5442 8014 5444
rect 8038 5442 8094 5444
rect 8118 5442 8174 5444
rect 8198 5442 8254 5444
rect 7878 5390 7880 5442
rect 7880 5390 7932 5442
rect 7932 5390 7934 5442
rect 7958 5390 7996 5442
rect 7996 5390 8008 5442
rect 8008 5390 8014 5442
rect 8038 5390 8060 5442
rect 8060 5390 8072 5442
rect 8072 5390 8094 5442
rect 8118 5390 8124 5442
rect 8124 5390 8136 5442
rect 8136 5390 8174 5442
rect 8198 5390 8200 5442
rect 8200 5390 8252 5442
rect 8252 5390 8254 5442
rect 7878 5388 7934 5390
rect 7958 5388 8014 5390
rect 8038 5388 8094 5390
rect 8118 5388 8174 5390
rect 8198 5388 8254 5390
rect 4017 4354 4073 4356
rect 4097 4354 4153 4356
rect 4177 4354 4233 4356
rect 4257 4354 4313 4356
rect 4337 4354 4393 4356
rect 4017 4302 4019 4354
rect 4019 4302 4071 4354
rect 4071 4302 4073 4354
rect 4097 4302 4135 4354
rect 4135 4302 4147 4354
rect 4147 4302 4153 4354
rect 4177 4302 4199 4354
rect 4199 4302 4211 4354
rect 4211 4302 4233 4354
rect 4257 4302 4263 4354
rect 4263 4302 4275 4354
rect 4275 4302 4313 4354
rect 4337 4302 4339 4354
rect 4339 4302 4391 4354
rect 4391 4302 4393 4354
rect 4017 4300 4073 4302
rect 4097 4300 4153 4302
rect 4177 4300 4233 4302
rect 4257 4300 4313 4302
rect 4337 4300 4393 4302
rect 5948 4354 6004 4356
rect 6028 4354 6084 4356
rect 6108 4354 6164 4356
rect 6188 4354 6244 4356
rect 6268 4354 6324 4356
rect 5948 4302 5950 4354
rect 5950 4302 6002 4354
rect 6002 4302 6004 4354
rect 6028 4302 6066 4354
rect 6066 4302 6078 4354
rect 6078 4302 6084 4354
rect 6108 4302 6130 4354
rect 6130 4302 6142 4354
rect 6142 4302 6164 4354
rect 6188 4302 6194 4354
rect 6194 4302 6206 4354
rect 6206 4302 6244 4354
rect 6268 4302 6270 4354
rect 6270 4302 6322 4354
rect 6322 4302 6324 4354
rect 5948 4300 6004 4302
rect 6028 4300 6084 4302
rect 6108 4300 6164 4302
rect 6188 4300 6244 4302
rect 6268 4300 6324 4302
rect 7878 4354 7934 4356
rect 7958 4354 8014 4356
rect 8038 4354 8094 4356
rect 8118 4354 8174 4356
rect 8198 4354 8254 4356
rect 7878 4302 7880 4354
rect 7880 4302 7932 4354
rect 7932 4302 7934 4354
rect 7958 4302 7996 4354
rect 7996 4302 8008 4354
rect 8008 4302 8014 4354
rect 8038 4302 8060 4354
rect 8060 4302 8072 4354
rect 8072 4302 8094 4354
rect 8118 4302 8124 4354
rect 8124 4302 8136 4354
rect 8136 4302 8174 4354
rect 8198 4302 8200 4354
rect 8200 4302 8252 4354
rect 8252 4302 8254 4354
rect 7878 4300 7934 4302
rect 7958 4300 8014 4302
rect 8038 4300 8094 4302
rect 8118 4300 8174 4302
rect 8198 4300 8254 4302
rect 4982 3810 5038 3812
rect 5062 3810 5118 3812
rect 5142 3810 5198 3812
rect 5222 3810 5278 3812
rect 5302 3810 5358 3812
rect 4982 3758 4984 3810
rect 4984 3758 5036 3810
rect 5036 3758 5038 3810
rect 5062 3758 5100 3810
rect 5100 3758 5112 3810
rect 5112 3758 5118 3810
rect 5142 3758 5164 3810
rect 5164 3758 5176 3810
rect 5176 3758 5198 3810
rect 5222 3758 5228 3810
rect 5228 3758 5240 3810
rect 5240 3758 5278 3810
rect 5302 3758 5304 3810
rect 5304 3758 5356 3810
rect 5356 3758 5358 3810
rect 4982 3756 5038 3758
rect 5062 3756 5118 3758
rect 5142 3756 5198 3758
rect 5222 3756 5278 3758
rect 5302 3756 5358 3758
rect 6913 3810 6969 3812
rect 6993 3810 7049 3812
rect 7073 3810 7129 3812
rect 7153 3810 7209 3812
rect 7233 3810 7289 3812
rect 6913 3758 6915 3810
rect 6915 3758 6967 3810
rect 6967 3758 6969 3810
rect 6993 3758 7031 3810
rect 7031 3758 7043 3810
rect 7043 3758 7049 3810
rect 7073 3758 7095 3810
rect 7095 3758 7107 3810
rect 7107 3758 7129 3810
rect 7153 3758 7159 3810
rect 7159 3758 7171 3810
rect 7171 3758 7209 3810
rect 7233 3758 7235 3810
rect 7235 3758 7287 3810
rect 7287 3758 7289 3810
rect 6913 3756 6969 3758
rect 6993 3756 7049 3758
rect 7073 3756 7129 3758
rect 7153 3756 7209 3758
rect 7233 3756 7289 3758
rect 4017 3266 4073 3268
rect 4097 3266 4153 3268
rect 4177 3266 4233 3268
rect 4257 3266 4313 3268
rect 4337 3266 4393 3268
rect 4017 3214 4019 3266
rect 4019 3214 4071 3266
rect 4071 3214 4073 3266
rect 4097 3214 4135 3266
rect 4135 3214 4147 3266
rect 4147 3214 4153 3266
rect 4177 3214 4199 3266
rect 4199 3214 4211 3266
rect 4211 3214 4233 3266
rect 4257 3214 4263 3266
rect 4263 3214 4275 3266
rect 4275 3214 4313 3266
rect 4337 3214 4339 3266
rect 4339 3214 4391 3266
rect 4391 3214 4393 3266
rect 4017 3212 4073 3214
rect 4097 3212 4153 3214
rect 4177 3212 4233 3214
rect 4257 3212 4313 3214
rect 4337 3212 4393 3214
rect 5948 3266 6004 3268
rect 6028 3266 6084 3268
rect 6108 3266 6164 3268
rect 6188 3266 6244 3268
rect 6268 3266 6324 3268
rect 5948 3214 5950 3266
rect 5950 3214 6002 3266
rect 6002 3214 6004 3266
rect 6028 3214 6066 3266
rect 6066 3214 6078 3266
rect 6078 3214 6084 3266
rect 6108 3214 6130 3266
rect 6130 3214 6142 3266
rect 6142 3214 6164 3266
rect 6188 3214 6194 3266
rect 6194 3214 6206 3266
rect 6206 3214 6244 3266
rect 6268 3214 6270 3266
rect 6270 3214 6322 3266
rect 6322 3214 6324 3266
rect 5948 3212 6004 3214
rect 6028 3212 6084 3214
rect 6108 3212 6164 3214
rect 6188 3212 6244 3214
rect 6268 3212 6324 3214
rect 7878 3266 7934 3268
rect 7958 3266 8014 3268
rect 8038 3266 8094 3268
rect 8118 3266 8174 3268
rect 8198 3266 8254 3268
rect 7878 3214 7880 3266
rect 7880 3214 7932 3266
rect 7932 3214 7934 3266
rect 7958 3214 7996 3266
rect 7996 3214 8008 3266
rect 8008 3214 8014 3266
rect 8038 3214 8060 3266
rect 8060 3214 8072 3266
rect 8072 3214 8094 3266
rect 8118 3214 8124 3266
rect 8124 3214 8136 3266
rect 8136 3214 8174 3266
rect 8198 3214 8200 3266
rect 8200 3214 8252 3266
rect 8252 3214 8254 3266
rect 7878 3212 7934 3214
rect 7958 3212 8014 3214
rect 8038 3212 8094 3214
rect 8118 3212 8174 3214
rect 8198 3212 8254 3214
<< metal3 >>
rect 0 20072 12184 20080
rect 0 20008 8 20072
rect 72 20008 88 20072
rect 152 20008 168 20072
rect 232 20008 248 20072
rect 312 20008 328 20072
rect 392 20008 408 20072
rect 472 20008 488 20072
rect 552 20008 568 20072
rect 632 20008 648 20072
rect 712 20008 728 20072
rect 792 20008 4978 20072
rect 5042 20008 5058 20072
rect 5122 20008 5138 20072
rect 5202 20008 5218 20072
rect 5282 20008 5298 20072
rect 5362 20008 6909 20072
rect 6973 20008 6989 20072
rect 7053 20008 7069 20072
rect 7133 20008 7149 20072
rect 7213 20008 7229 20072
rect 7293 20008 11392 20072
rect 11456 20008 11472 20072
rect 11536 20008 11552 20072
rect 11616 20008 11632 20072
rect 11696 20008 11712 20072
rect 11776 20008 11792 20072
rect 11856 20008 11872 20072
rect 11936 20008 11952 20072
rect 12016 20008 12032 20072
rect 12096 20008 12112 20072
rect 12176 20008 12184 20072
rect 0 19992 12184 20008
rect 0 19928 8 19992
rect 72 19928 88 19992
rect 152 19928 168 19992
rect 232 19928 248 19992
rect 312 19928 328 19992
rect 392 19928 408 19992
rect 472 19928 488 19992
rect 552 19928 568 19992
rect 632 19928 648 19992
rect 712 19928 728 19992
rect 792 19928 4978 19992
rect 5042 19928 5058 19992
rect 5122 19928 5138 19992
rect 5202 19928 5218 19992
rect 5282 19928 5298 19992
rect 5362 19928 6909 19992
rect 6973 19928 6989 19992
rect 7053 19928 7069 19992
rect 7133 19928 7149 19992
rect 7213 19928 7229 19992
rect 7293 19928 11392 19992
rect 11456 19928 11472 19992
rect 11536 19928 11552 19992
rect 11616 19928 11632 19992
rect 11696 19928 11712 19992
rect 11776 19928 11792 19992
rect 11856 19928 11872 19992
rect 11936 19928 11952 19992
rect 12016 19928 12032 19992
rect 12096 19928 12112 19992
rect 12176 19928 12184 19992
rect 0 19912 12184 19928
rect 0 19848 8 19912
rect 72 19848 88 19912
rect 152 19848 168 19912
rect 232 19848 248 19912
rect 312 19848 328 19912
rect 392 19848 408 19912
rect 472 19848 488 19912
rect 552 19848 568 19912
rect 632 19848 648 19912
rect 712 19848 728 19912
rect 792 19848 4978 19912
rect 5042 19848 5058 19912
rect 5122 19848 5138 19912
rect 5202 19848 5218 19912
rect 5282 19848 5298 19912
rect 5362 19848 6909 19912
rect 6973 19848 6989 19912
rect 7053 19848 7069 19912
rect 7133 19848 7149 19912
rect 7213 19848 7229 19912
rect 7293 19848 11392 19912
rect 11456 19848 11472 19912
rect 11536 19848 11552 19912
rect 11616 19848 11632 19912
rect 11696 19848 11712 19912
rect 11776 19848 11792 19912
rect 11856 19848 11872 19912
rect 11936 19848 11952 19912
rect 12016 19848 12032 19912
rect 12096 19848 12112 19912
rect 12176 19848 12184 19912
rect 0 19832 12184 19848
rect 0 19768 8 19832
rect 72 19768 88 19832
rect 152 19768 168 19832
rect 232 19768 248 19832
rect 312 19768 328 19832
rect 392 19768 408 19832
rect 472 19768 488 19832
rect 552 19768 568 19832
rect 632 19768 648 19832
rect 712 19768 728 19832
rect 792 19768 4978 19832
rect 5042 19768 5058 19832
rect 5122 19768 5138 19832
rect 5202 19768 5218 19832
rect 5282 19768 5298 19832
rect 5362 19768 6909 19832
rect 6973 19768 6989 19832
rect 7053 19768 7069 19832
rect 7133 19768 7149 19832
rect 7213 19768 7229 19832
rect 7293 19768 11392 19832
rect 11456 19768 11472 19832
rect 11536 19768 11552 19832
rect 11616 19768 11632 19832
rect 11696 19768 11712 19832
rect 11776 19768 11792 19832
rect 11856 19768 11872 19832
rect 11936 19768 11952 19832
rect 12016 19768 12032 19832
rect 12096 19768 12112 19832
rect 12176 19768 12184 19832
rect 0 19752 12184 19768
rect 0 19688 8 19752
rect 72 19688 88 19752
rect 152 19688 168 19752
rect 232 19688 248 19752
rect 312 19688 328 19752
rect 392 19688 408 19752
rect 472 19688 488 19752
rect 552 19688 568 19752
rect 632 19688 648 19752
rect 712 19688 728 19752
rect 792 19688 4978 19752
rect 5042 19688 5058 19752
rect 5122 19688 5138 19752
rect 5202 19688 5218 19752
rect 5282 19688 5298 19752
rect 5362 19688 6909 19752
rect 6973 19688 6989 19752
rect 7053 19688 7069 19752
rect 7133 19688 7149 19752
rect 7213 19688 7229 19752
rect 7293 19688 11392 19752
rect 11456 19688 11472 19752
rect 11536 19688 11552 19752
rect 11616 19688 11632 19752
rect 11696 19688 11712 19752
rect 11776 19688 11792 19752
rect 11856 19688 11872 19752
rect 11936 19688 11952 19752
rect 12016 19688 12032 19752
rect 12096 19688 12112 19752
rect 12176 19688 12184 19752
rect 0 19672 12184 19688
rect 0 19608 8 19672
rect 72 19608 88 19672
rect 152 19608 168 19672
rect 232 19608 248 19672
rect 312 19608 328 19672
rect 392 19608 408 19672
rect 472 19608 488 19672
rect 552 19608 568 19672
rect 632 19608 648 19672
rect 712 19608 728 19672
rect 792 19608 4978 19672
rect 5042 19608 5058 19672
rect 5122 19608 5138 19672
rect 5202 19608 5218 19672
rect 5282 19608 5298 19672
rect 5362 19608 6909 19672
rect 6973 19608 6989 19672
rect 7053 19608 7069 19672
rect 7133 19608 7149 19672
rect 7213 19608 7229 19672
rect 7293 19608 11392 19672
rect 11456 19608 11472 19672
rect 11536 19608 11552 19672
rect 11616 19608 11632 19672
rect 11696 19608 11712 19672
rect 11776 19608 11792 19672
rect 11856 19608 11872 19672
rect 11936 19608 11952 19672
rect 12016 19608 12032 19672
rect 12096 19608 12112 19672
rect 12176 19608 12184 19672
rect 0 19592 12184 19608
rect 0 19528 8 19592
rect 72 19528 88 19592
rect 152 19528 168 19592
rect 232 19528 248 19592
rect 312 19528 328 19592
rect 392 19528 408 19592
rect 472 19528 488 19592
rect 552 19528 568 19592
rect 632 19528 648 19592
rect 712 19528 728 19592
rect 792 19528 4978 19592
rect 5042 19528 5058 19592
rect 5122 19528 5138 19592
rect 5202 19528 5218 19592
rect 5282 19528 5298 19592
rect 5362 19528 6909 19592
rect 6973 19528 6989 19592
rect 7053 19528 7069 19592
rect 7133 19528 7149 19592
rect 7213 19528 7229 19592
rect 7293 19528 11392 19592
rect 11456 19528 11472 19592
rect 11536 19528 11552 19592
rect 11616 19528 11632 19592
rect 11696 19528 11712 19592
rect 11776 19528 11792 19592
rect 11856 19528 11872 19592
rect 11936 19528 11952 19592
rect 12016 19528 12032 19592
rect 12096 19528 12112 19592
rect 12176 19528 12184 19592
rect 0 19512 12184 19528
rect 0 19448 8 19512
rect 72 19448 88 19512
rect 152 19448 168 19512
rect 232 19448 248 19512
rect 312 19448 328 19512
rect 392 19448 408 19512
rect 472 19448 488 19512
rect 552 19448 568 19512
rect 632 19448 648 19512
rect 712 19448 728 19512
rect 792 19448 4978 19512
rect 5042 19448 5058 19512
rect 5122 19448 5138 19512
rect 5202 19448 5218 19512
rect 5282 19448 5298 19512
rect 5362 19448 6909 19512
rect 6973 19448 6989 19512
rect 7053 19448 7069 19512
rect 7133 19448 7149 19512
rect 7213 19448 7229 19512
rect 7293 19448 11392 19512
rect 11456 19448 11472 19512
rect 11536 19448 11552 19512
rect 11616 19448 11632 19512
rect 11696 19448 11712 19512
rect 11776 19448 11792 19512
rect 11856 19448 11872 19512
rect 11936 19448 11952 19512
rect 12016 19448 12032 19512
rect 12096 19448 12112 19512
rect 12176 19448 12184 19512
rect 0 19432 12184 19448
rect 0 19368 8 19432
rect 72 19368 88 19432
rect 152 19368 168 19432
rect 232 19368 248 19432
rect 312 19368 328 19432
rect 392 19368 408 19432
rect 472 19368 488 19432
rect 552 19368 568 19432
rect 632 19368 648 19432
rect 712 19368 728 19432
rect 792 19368 4978 19432
rect 5042 19368 5058 19432
rect 5122 19368 5138 19432
rect 5202 19368 5218 19432
rect 5282 19368 5298 19432
rect 5362 19368 6909 19432
rect 6973 19368 6989 19432
rect 7053 19368 7069 19432
rect 7133 19368 7149 19432
rect 7213 19368 7229 19432
rect 7293 19368 11392 19432
rect 11456 19368 11472 19432
rect 11536 19368 11552 19432
rect 11616 19368 11632 19432
rect 11696 19368 11712 19432
rect 11776 19368 11792 19432
rect 11856 19368 11872 19432
rect 11936 19368 11952 19432
rect 12016 19368 12032 19432
rect 12096 19368 12112 19432
rect 12176 19368 12184 19432
rect 0 19352 12184 19368
rect 0 19288 8 19352
rect 72 19288 88 19352
rect 152 19288 168 19352
rect 232 19288 248 19352
rect 312 19288 328 19352
rect 392 19288 408 19352
rect 472 19288 488 19352
rect 552 19288 568 19352
rect 632 19288 648 19352
rect 712 19288 728 19352
rect 792 19288 4978 19352
rect 5042 19288 5058 19352
rect 5122 19288 5138 19352
rect 5202 19288 5218 19352
rect 5282 19288 5298 19352
rect 5362 19288 6909 19352
rect 6973 19288 6989 19352
rect 7053 19288 7069 19352
rect 7133 19288 7149 19352
rect 7213 19288 7229 19352
rect 7293 19288 11392 19352
rect 11456 19288 11472 19352
rect 11536 19288 11552 19352
rect 11616 19288 11632 19352
rect 11696 19288 11712 19352
rect 11776 19288 11792 19352
rect 11856 19288 11872 19352
rect 11936 19288 11952 19352
rect 12016 19288 12032 19352
rect 12096 19288 12112 19352
rect 12176 19288 12184 19352
rect 0 19280 12184 19288
rect 1140 18932 11044 18940
rect 1140 18868 1148 18932
rect 1212 18868 1228 18932
rect 1292 18868 1308 18932
rect 1372 18868 1388 18932
rect 1452 18868 1468 18932
rect 1532 18868 1548 18932
rect 1612 18868 1628 18932
rect 1692 18868 1708 18932
rect 1772 18868 1788 18932
rect 1852 18868 1868 18932
rect 1932 18868 4013 18932
rect 4077 18868 4093 18932
rect 4157 18868 4173 18932
rect 4237 18868 4253 18932
rect 4317 18868 4333 18932
rect 4397 18868 5944 18932
rect 6008 18868 6024 18932
rect 6088 18868 6104 18932
rect 6168 18868 6184 18932
rect 6248 18868 6264 18932
rect 6328 18868 7874 18932
rect 7938 18868 7954 18932
rect 8018 18868 8034 18932
rect 8098 18868 8114 18932
rect 8178 18868 8194 18932
rect 8258 18868 10252 18932
rect 10316 18868 10332 18932
rect 10396 18868 10412 18932
rect 10476 18868 10492 18932
rect 10556 18868 10572 18932
rect 10636 18868 10652 18932
rect 10716 18868 10732 18932
rect 10796 18868 10812 18932
rect 10876 18868 10892 18932
rect 10956 18868 10972 18932
rect 11036 18868 11044 18932
rect 1140 18852 11044 18868
rect 1140 18788 1148 18852
rect 1212 18788 1228 18852
rect 1292 18788 1308 18852
rect 1372 18788 1388 18852
rect 1452 18788 1468 18852
rect 1532 18788 1548 18852
rect 1612 18788 1628 18852
rect 1692 18788 1708 18852
rect 1772 18788 1788 18852
rect 1852 18788 1868 18852
rect 1932 18788 4013 18852
rect 4077 18788 4093 18852
rect 4157 18788 4173 18852
rect 4237 18788 4253 18852
rect 4317 18788 4333 18852
rect 4397 18788 5944 18852
rect 6008 18788 6024 18852
rect 6088 18788 6104 18852
rect 6168 18788 6184 18852
rect 6248 18788 6264 18852
rect 6328 18788 7874 18852
rect 7938 18788 7954 18852
rect 8018 18788 8034 18852
rect 8098 18788 8114 18852
rect 8178 18788 8194 18852
rect 8258 18788 10252 18852
rect 10316 18788 10332 18852
rect 10396 18788 10412 18852
rect 10476 18788 10492 18852
rect 10556 18788 10572 18852
rect 10636 18788 10652 18852
rect 10716 18788 10732 18852
rect 10796 18788 10812 18852
rect 10876 18788 10892 18852
rect 10956 18788 10972 18852
rect 11036 18788 11044 18852
rect 1140 18772 11044 18788
rect 1140 18708 1148 18772
rect 1212 18708 1228 18772
rect 1292 18708 1308 18772
rect 1372 18708 1388 18772
rect 1452 18708 1468 18772
rect 1532 18708 1548 18772
rect 1612 18708 1628 18772
rect 1692 18708 1708 18772
rect 1772 18708 1788 18772
rect 1852 18708 1868 18772
rect 1932 18708 4013 18772
rect 4077 18708 4093 18772
rect 4157 18708 4173 18772
rect 4237 18708 4253 18772
rect 4317 18708 4333 18772
rect 4397 18708 5944 18772
rect 6008 18708 6024 18772
rect 6088 18708 6104 18772
rect 6168 18708 6184 18772
rect 6248 18708 6264 18772
rect 6328 18708 7874 18772
rect 7938 18708 7954 18772
rect 8018 18708 8034 18772
rect 8098 18708 8114 18772
rect 8178 18708 8194 18772
rect 8258 18708 10252 18772
rect 10316 18708 10332 18772
rect 10396 18708 10412 18772
rect 10476 18708 10492 18772
rect 10556 18708 10572 18772
rect 10636 18708 10652 18772
rect 10716 18708 10732 18772
rect 10796 18708 10812 18772
rect 10876 18708 10892 18772
rect 10956 18708 10972 18772
rect 11036 18708 11044 18772
rect 1140 18692 11044 18708
rect 1140 18628 1148 18692
rect 1212 18628 1228 18692
rect 1292 18628 1308 18692
rect 1372 18628 1388 18692
rect 1452 18628 1468 18692
rect 1532 18628 1548 18692
rect 1612 18628 1628 18692
rect 1692 18628 1708 18692
rect 1772 18628 1788 18692
rect 1852 18628 1868 18692
rect 1932 18628 4013 18692
rect 4077 18628 4093 18692
rect 4157 18628 4173 18692
rect 4237 18628 4253 18692
rect 4317 18628 4333 18692
rect 4397 18628 5944 18692
rect 6008 18628 6024 18692
rect 6088 18628 6104 18692
rect 6168 18628 6184 18692
rect 6248 18628 6264 18692
rect 6328 18628 7874 18692
rect 7938 18628 7954 18692
rect 8018 18628 8034 18692
rect 8098 18628 8114 18692
rect 8178 18628 8194 18692
rect 8258 18628 10252 18692
rect 10316 18628 10332 18692
rect 10396 18628 10412 18692
rect 10476 18628 10492 18692
rect 10556 18628 10572 18692
rect 10636 18628 10652 18692
rect 10716 18628 10732 18692
rect 10796 18628 10812 18692
rect 10876 18628 10892 18692
rect 10956 18628 10972 18692
rect 11036 18628 11044 18692
rect 1140 18612 11044 18628
rect 1140 18548 1148 18612
rect 1212 18548 1228 18612
rect 1292 18548 1308 18612
rect 1372 18548 1388 18612
rect 1452 18548 1468 18612
rect 1532 18548 1548 18612
rect 1612 18548 1628 18612
rect 1692 18548 1708 18612
rect 1772 18548 1788 18612
rect 1852 18548 1868 18612
rect 1932 18548 4013 18612
rect 4077 18548 4093 18612
rect 4157 18548 4173 18612
rect 4237 18548 4253 18612
rect 4317 18548 4333 18612
rect 4397 18548 5944 18612
rect 6008 18548 6024 18612
rect 6088 18548 6104 18612
rect 6168 18548 6184 18612
rect 6248 18548 6264 18612
rect 6328 18548 7874 18612
rect 7938 18548 7954 18612
rect 8018 18548 8034 18612
rect 8098 18548 8114 18612
rect 8178 18548 8194 18612
rect 8258 18548 10252 18612
rect 10316 18548 10332 18612
rect 10396 18548 10412 18612
rect 10476 18548 10492 18612
rect 10556 18548 10572 18612
rect 10636 18548 10652 18612
rect 10716 18548 10732 18612
rect 10796 18548 10812 18612
rect 10876 18548 10892 18612
rect 10956 18548 10972 18612
rect 11036 18548 11044 18612
rect 1140 18532 11044 18548
rect 1140 18468 1148 18532
rect 1212 18468 1228 18532
rect 1292 18468 1308 18532
rect 1372 18468 1388 18532
rect 1452 18468 1468 18532
rect 1532 18468 1548 18532
rect 1612 18468 1628 18532
rect 1692 18468 1708 18532
rect 1772 18468 1788 18532
rect 1852 18468 1868 18532
rect 1932 18468 4013 18532
rect 4077 18468 4093 18532
rect 4157 18468 4173 18532
rect 4237 18468 4253 18532
rect 4317 18468 4333 18532
rect 4397 18468 5944 18532
rect 6008 18468 6024 18532
rect 6088 18468 6104 18532
rect 6168 18468 6184 18532
rect 6248 18468 6264 18532
rect 6328 18468 7874 18532
rect 7938 18468 7954 18532
rect 8018 18468 8034 18532
rect 8098 18468 8114 18532
rect 8178 18468 8194 18532
rect 8258 18468 10252 18532
rect 10316 18468 10332 18532
rect 10396 18468 10412 18532
rect 10476 18468 10492 18532
rect 10556 18468 10572 18532
rect 10636 18468 10652 18532
rect 10716 18468 10732 18532
rect 10796 18468 10812 18532
rect 10876 18468 10892 18532
rect 10956 18468 10972 18532
rect 11036 18468 11044 18532
rect 1140 18452 11044 18468
rect 1140 18388 1148 18452
rect 1212 18388 1228 18452
rect 1292 18388 1308 18452
rect 1372 18388 1388 18452
rect 1452 18388 1468 18452
rect 1532 18388 1548 18452
rect 1612 18388 1628 18452
rect 1692 18388 1708 18452
rect 1772 18388 1788 18452
rect 1852 18388 1868 18452
rect 1932 18388 4013 18452
rect 4077 18388 4093 18452
rect 4157 18388 4173 18452
rect 4237 18388 4253 18452
rect 4317 18388 4333 18452
rect 4397 18388 5944 18452
rect 6008 18388 6024 18452
rect 6088 18388 6104 18452
rect 6168 18388 6184 18452
rect 6248 18388 6264 18452
rect 6328 18388 7874 18452
rect 7938 18388 7954 18452
rect 8018 18388 8034 18452
rect 8098 18388 8114 18452
rect 8178 18388 8194 18452
rect 8258 18388 10252 18452
rect 10316 18388 10332 18452
rect 10396 18388 10412 18452
rect 10476 18388 10492 18452
rect 10556 18388 10572 18452
rect 10636 18388 10652 18452
rect 10716 18388 10732 18452
rect 10796 18388 10812 18452
rect 10876 18388 10892 18452
rect 10956 18388 10972 18452
rect 11036 18388 11044 18452
rect 1140 18372 11044 18388
rect 1140 18308 1148 18372
rect 1212 18308 1228 18372
rect 1292 18308 1308 18372
rect 1372 18308 1388 18372
rect 1452 18308 1468 18372
rect 1532 18308 1548 18372
rect 1612 18308 1628 18372
rect 1692 18308 1708 18372
rect 1772 18308 1788 18372
rect 1852 18308 1868 18372
rect 1932 18308 4013 18372
rect 4077 18308 4093 18372
rect 4157 18308 4173 18372
rect 4237 18308 4253 18372
rect 4317 18308 4333 18372
rect 4397 18308 5944 18372
rect 6008 18308 6024 18372
rect 6088 18308 6104 18372
rect 6168 18308 6184 18372
rect 6248 18308 6264 18372
rect 6328 18308 7874 18372
rect 7938 18308 7954 18372
rect 8018 18308 8034 18372
rect 8098 18308 8114 18372
rect 8178 18308 8194 18372
rect 8258 18308 10252 18372
rect 10316 18308 10332 18372
rect 10396 18308 10412 18372
rect 10476 18308 10492 18372
rect 10556 18308 10572 18372
rect 10636 18308 10652 18372
rect 10716 18308 10732 18372
rect 10796 18308 10812 18372
rect 10876 18308 10892 18372
rect 10956 18308 10972 18372
rect 11036 18308 11044 18372
rect 1140 18292 11044 18308
rect 1140 18228 1148 18292
rect 1212 18228 1228 18292
rect 1292 18228 1308 18292
rect 1372 18228 1388 18292
rect 1452 18228 1468 18292
rect 1532 18228 1548 18292
rect 1612 18228 1628 18292
rect 1692 18228 1708 18292
rect 1772 18228 1788 18292
rect 1852 18228 1868 18292
rect 1932 18228 4013 18292
rect 4077 18228 4093 18292
rect 4157 18228 4173 18292
rect 4237 18228 4253 18292
rect 4317 18228 4333 18292
rect 4397 18228 5944 18292
rect 6008 18228 6024 18292
rect 6088 18228 6104 18292
rect 6168 18228 6184 18292
rect 6248 18228 6264 18292
rect 6328 18228 7874 18292
rect 7938 18228 7954 18292
rect 8018 18228 8034 18292
rect 8098 18228 8114 18292
rect 8178 18228 8194 18292
rect 8258 18228 10252 18292
rect 10316 18228 10332 18292
rect 10396 18228 10412 18292
rect 10476 18228 10492 18292
rect 10556 18228 10572 18292
rect 10636 18228 10652 18292
rect 10716 18228 10732 18292
rect 10796 18228 10812 18292
rect 10876 18228 10892 18292
rect 10956 18228 10972 18292
rect 11036 18228 11044 18292
rect 1140 18212 11044 18228
rect 1140 18148 1148 18212
rect 1212 18148 1228 18212
rect 1292 18148 1308 18212
rect 1372 18148 1388 18212
rect 1452 18148 1468 18212
rect 1532 18148 1548 18212
rect 1612 18148 1628 18212
rect 1692 18148 1708 18212
rect 1772 18148 1788 18212
rect 1852 18148 1868 18212
rect 1932 18148 4013 18212
rect 4077 18148 4093 18212
rect 4157 18148 4173 18212
rect 4237 18148 4253 18212
rect 4317 18148 4333 18212
rect 4397 18148 5944 18212
rect 6008 18148 6024 18212
rect 6088 18148 6104 18212
rect 6168 18148 6184 18212
rect 6248 18148 6264 18212
rect 6328 18148 7874 18212
rect 7938 18148 7954 18212
rect 8018 18148 8034 18212
rect 8098 18148 8114 18212
rect 8178 18148 8194 18212
rect 8258 18148 10252 18212
rect 10316 18148 10332 18212
rect 10396 18148 10412 18212
rect 10476 18148 10492 18212
rect 10556 18148 10572 18212
rect 10636 18148 10652 18212
rect 10716 18148 10732 18212
rect 10796 18148 10812 18212
rect 10876 18148 10892 18212
rect 10956 18148 10972 18212
rect 11036 18148 11044 18212
rect 1140 18140 11044 18148
rect 4960 16872 5380 16873
rect 4960 16808 4978 16872
rect 5042 16808 5058 16872
rect 5122 16808 5138 16872
rect 5202 16808 5218 16872
rect 5282 16808 5298 16872
rect 5362 16808 5380 16872
rect 4960 16807 5380 16808
rect 6891 16872 7311 16873
rect 6891 16808 6909 16872
rect 6973 16808 6989 16872
rect 7053 16808 7069 16872
rect 7133 16808 7149 16872
rect 7213 16808 7229 16872
rect 7293 16808 7311 16872
rect 6891 16807 7311 16808
rect 3995 16328 4415 16329
rect 3995 16264 4013 16328
rect 4077 16264 4093 16328
rect 4157 16264 4173 16328
rect 4237 16264 4253 16328
rect 4317 16264 4333 16328
rect 4397 16264 4415 16328
rect 3995 16263 4415 16264
rect 5926 16328 6346 16329
rect 5926 16264 5944 16328
rect 6008 16264 6024 16328
rect 6088 16264 6104 16328
rect 6168 16264 6184 16328
rect 6248 16264 6264 16328
rect 6328 16264 6346 16328
rect 5926 16263 6346 16264
rect 7856 16328 8276 16329
rect 7856 16264 7874 16328
rect 7938 16264 7954 16328
rect 8018 16264 8034 16328
rect 8098 16264 8114 16328
rect 8178 16264 8194 16328
rect 8258 16264 8276 16328
rect 7856 16263 8276 16264
rect 4960 15784 5380 15785
rect 4960 15720 4978 15784
rect 5042 15720 5058 15784
rect 5122 15720 5138 15784
rect 5202 15720 5218 15784
rect 5282 15720 5298 15784
rect 5362 15720 5380 15784
rect 4960 15719 5380 15720
rect 6891 15784 7311 15785
rect 6891 15720 6909 15784
rect 6973 15720 6989 15784
rect 7053 15720 7069 15784
rect 7133 15720 7149 15784
rect 7213 15720 7229 15784
rect 7293 15720 7311 15784
rect 6891 15719 7311 15720
rect 3995 15240 4415 15241
rect 3995 15176 4013 15240
rect 4077 15176 4093 15240
rect 4157 15176 4173 15240
rect 4237 15176 4253 15240
rect 4317 15176 4333 15240
rect 4397 15176 4415 15240
rect 3995 15175 4415 15176
rect 5926 15240 6346 15241
rect 5926 15176 5944 15240
rect 6008 15176 6024 15240
rect 6088 15176 6104 15240
rect 6168 15176 6184 15240
rect 6248 15176 6264 15240
rect 6328 15176 6346 15240
rect 5926 15175 6346 15176
rect 7856 15240 8276 15241
rect 7856 15176 7874 15240
rect 7938 15176 7954 15240
rect 8018 15176 8034 15240
rect 8098 15176 8114 15240
rect 8178 15176 8194 15240
rect 8258 15176 8276 15240
rect 7856 15175 8276 15176
rect 4960 14696 5380 14697
rect 4960 14632 4978 14696
rect 5042 14632 5058 14696
rect 5122 14632 5138 14696
rect 5202 14632 5218 14696
rect 5282 14632 5298 14696
rect 5362 14632 5380 14696
rect 4960 14631 5380 14632
rect 6891 14696 7311 14697
rect 6891 14632 6909 14696
rect 6973 14632 6989 14696
rect 7053 14632 7069 14696
rect 7133 14632 7149 14696
rect 7213 14632 7229 14696
rect 7293 14632 7311 14696
rect 6891 14631 7311 14632
rect 3995 14152 4415 14153
rect 3995 14088 4013 14152
rect 4077 14088 4093 14152
rect 4157 14088 4173 14152
rect 4237 14088 4253 14152
rect 4317 14088 4333 14152
rect 4397 14088 4415 14152
rect 3995 14087 4415 14088
rect 5926 14152 6346 14153
rect 5926 14088 5944 14152
rect 6008 14088 6024 14152
rect 6088 14088 6104 14152
rect 6168 14088 6184 14152
rect 6248 14088 6264 14152
rect 6328 14088 6346 14152
rect 5926 14087 6346 14088
rect 7856 14152 8276 14153
rect 7856 14088 7874 14152
rect 7938 14088 7954 14152
rect 8018 14088 8034 14152
rect 8098 14088 8114 14152
rect 8178 14088 8194 14152
rect 8258 14088 8276 14152
rect 7856 14087 8276 14088
rect 4960 13608 5380 13609
rect 4960 13544 4978 13608
rect 5042 13544 5058 13608
rect 5122 13544 5138 13608
rect 5202 13544 5218 13608
rect 5282 13544 5298 13608
rect 5362 13544 5380 13608
rect 4960 13543 5380 13544
rect 6891 13608 7311 13609
rect 6891 13544 6909 13608
rect 6973 13544 6989 13608
rect 7053 13544 7069 13608
rect 7133 13544 7149 13608
rect 7213 13544 7229 13608
rect 7293 13544 7311 13608
rect 6891 13543 7311 13544
rect 3995 13064 4415 13065
rect 3995 13000 4013 13064
rect 4077 13000 4093 13064
rect 4157 13000 4173 13064
rect 4237 13000 4253 13064
rect 4317 13000 4333 13064
rect 4397 13000 4415 13064
rect 3995 12999 4415 13000
rect 5926 13064 6346 13065
rect 5926 13000 5944 13064
rect 6008 13000 6024 13064
rect 6088 13000 6104 13064
rect 6168 13000 6184 13064
rect 6248 13000 6264 13064
rect 6328 13000 6346 13064
rect 5926 12999 6346 13000
rect 7856 13064 8276 13065
rect 7856 13000 7874 13064
rect 7938 13000 7954 13064
rect 8018 13000 8034 13064
rect 8098 13000 8114 13064
rect 8178 13000 8194 13064
rect 8258 13000 8276 13064
rect 7856 12999 8276 13000
rect 4960 12520 5380 12521
rect 4960 12456 4978 12520
rect 5042 12456 5058 12520
rect 5122 12456 5138 12520
rect 5202 12456 5218 12520
rect 5282 12456 5298 12520
rect 5362 12456 5380 12520
rect 4960 12455 5380 12456
rect 6891 12520 7311 12521
rect 6891 12456 6909 12520
rect 6973 12456 6989 12520
rect 7053 12456 7069 12520
rect 7133 12456 7149 12520
rect 7213 12456 7229 12520
rect 7293 12456 7311 12520
rect 6891 12455 7311 12456
rect 3995 11976 4415 11977
rect 3995 11912 4013 11976
rect 4077 11912 4093 11976
rect 4157 11912 4173 11976
rect 4237 11912 4253 11976
rect 4317 11912 4333 11976
rect 4397 11912 4415 11976
rect 3995 11911 4415 11912
rect 5926 11976 6346 11977
rect 5926 11912 5944 11976
rect 6008 11912 6024 11976
rect 6088 11912 6104 11976
rect 6168 11912 6184 11976
rect 6248 11912 6264 11976
rect 6328 11912 6346 11976
rect 5926 11911 6346 11912
rect 7856 11976 8276 11977
rect 7856 11912 7874 11976
rect 7938 11912 7954 11976
rect 8018 11912 8034 11976
rect 8098 11912 8114 11976
rect 8178 11912 8194 11976
rect 8258 11912 8276 11976
rect 7856 11911 8276 11912
rect 4960 11432 5380 11433
rect 4960 11368 4978 11432
rect 5042 11368 5058 11432
rect 5122 11368 5138 11432
rect 5202 11368 5218 11432
rect 5282 11368 5298 11432
rect 5362 11368 5380 11432
rect 4960 11367 5380 11368
rect 6891 11432 7311 11433
rect 6891 11368 6909 11432
rect 6973 11368 6989 11432
rect 7053 11368 7069 11432
rect 7133 11368 7149 11432
rect 7213 11368 7229 11432
rect 7293 11368 7311 11432
rect 6891 11367 7311 11368
rect 3995 10888 4415 10889
rect 3995 10824 4013 10888
rect 4077 10824 4093 10888
rect 4157 10824 4173 10888
rect 4237 10824 4253 10888
rect 4317 10824 4333 10888
rect 4397 10824 4415 10888
rect 3995 10823 4415 10824
rect 5926 10888 6346 10889
rect 5926 10824 5944 10888
rect 6008 10824 6024 10888
rect 6088 10824 6104 10888
rect 6168 10824 6184 10888
rect 6248 10824 6264 10888
rect 6328 10824 6346 10888
rect 5926 10823 6346 10824
rect 7856 10888 8276 10889
rect 7856 10824 7874 10888
rect 7938 10824 7954 10888
rect 8018 10824 8034 10888
rect 8098 10824 8114 10888
rect 8178 10824 8194 10888
rect 8258 10824 8276 10888
rect 7856 10823 8276 10824
rect 7025 10546 7091 10549
rect 6614 10544 7091 10546
rect 6614 10488 7030 10544
rect 7086 10488 7091 10544
rect 6614 10486 7091 10488
rect 4960 10344 5380 10345
rect 4960 10280 4978 10344
rect 5042 10280 5058 10344
rect 5122 10280 5138 10344
rect 5202 10280 5218 10344
rect 5282 10280 5298 10344
rect 5362 10280 5380 10344
rect 4960 10279 5380 10280
rect 6614 10138 6674 10486
rect 7025 10483 7091 10486
rect 6891 10344 7311 10345
rect 6891 10280 6909 10344
rect 6973 10280 6989 10344
rect 7053 10280 7069 10344
rect 7133 10280 7149 10344
rect 7213 10280 7229 10344
rect 7293 10280 7311 10344
rect 6891 10279 7311 10280
rect 6841 10138 6907 10141
rect 6614 10136 6907 10138
rect 6614 10080 6846 10136
rect 6902 10080 6907 10136
rect 6614 10078 6907 10080
rect 6841 10075 6907 10078
rect 3995 9800 4415 9801
rect 3995 9736 4013 9800
rect 4077 9736 4093 9800
rect 4157 9736 4173 9800
rect 4237 9736 4253 9800
rect 4317 9736 4333 9800
rect 4397 9736 4415 9800
rect 3995 9735 4415 9736
rect 5926 9800 6346 9801
rect 5926 9736 5944 9800
rect 6008 9736 6024 9800
rect 6088 9736 6104 9800
rect 6168 9736 6184 9800
rect 6248 9736 6264 9800
rect 6328 9736 6346 9800
rect 5926 9735 6346 9736
rect 7856 9800 8276 9801
rect 7856 9736 7874 9800
rect 7938 9736 7954 9800
rect 8018 9736 8034 9800
rect 8098 9736 8114 9800
rect 8178 9736 8194 9800
rect 8258 9736 8276 9800
rect 7856 9735 8276 9736
rect 4960 9256 5380 9257
rect 4960 9192 4978 9256
rect 5042 9192 5058 9256
rect 5122 9192 5138 9256
rect 5202 9192 5218 9256
rect 5282 9192 5298 9256
rect 5362 9192 5380 9256
rect 4960 9191 5380 9192
rect 6891 9256 7311 9257
rect 6891 9192 6909 9256
rect 6973 9192 6989 9256
rect 7053 9192 7069 9256
rect 7133 9192 7149 9256
rect 7213 9192 7229 9256
rect 7293 9192 7311 9256
rect 6891 9191 7311 9192
rect 3995 8712 4415 8713
rect 3995 8648 4013 8712
rect 4077 8648 4093 8712
rect 4157 8648 4173 8712
rect 4237 8648 4253 8712
rect 4317 8648 4333 8712
rect 4397 8648 4415 8712
rect 3995 8647 4415 8648
rect 5926 8712 6346 8713
rect 5926 8648 5944 8712
rect 6008 8648 6024 8712
rect 6088 8648 6104 8712
rect 6168 8648 6184 8712
rect 6248 8648 6264 8712
rect 6328 8648 6346 8712
rect 5926 8647 6346 8648
rect 7856 8712 8276 8713
rect 7856 8648 7874 8712
rect 7938 8648 7954 8712
rect 8018 8648 8034 8712
rect 8098 8648 8114 8712
rect 8178 8648 8194 8712
rect 8258 8648 8276 8712
rect 7856 8647 8276 8648
rect 4960 8168 5380 8169
rect 4960 8104 4978 8168
rect 5042 8104 5058 8168
rect 5122 8104 5138 8168
rect 5202 8104 5218 8168
rect 5282 8104 5298 8168
rect 5362 8104 5380 8168
rect 4960 8103 5380 8104
rect 6891 8168 7311 8169
rect 6891 8104 6909 8168
rect 6973 8104 6989 8168
rect 7053 8104 7069 8168
rect 7133 8104 7149 8168
rect 7213 8104 7229 8168
rect 7293 8104 7311 8168
rect 6891 8103 7311 8104
rect 3995 7624 4415 7625
rect 3995 7560 4013 7624
rect 4077 7560 4093 7624
rect 4157 7560 4173 7624
rect 4237 7560 4253 7624
rect 4317 7560 4333 7624
rect 4397 7560 4415 7624
rect 3995 7559 4415 7560
rect 5926 7624 6346 7625
rect 5926 7560 5944 7624
rect 6008 7560 6024 7624
rect 6088 7560 6104 7624
rect 6168 7560 6184 7624
rect 6248 7560 6264 7624
rect 6328 7560 6346 7624
rect 5926 7559 6346 7560
rect 7856 7624 8276 7625
rect 7856 7560 7874 7624
rect 7938 7560 7954 7624
rect 8018 7560 8034 7624
rect 8098 7560 8114 7624
rect 8178 7560 8194 7624
rect 8258 7560 8276 7624
rect 7856 7559 8276 7560
rect 4960 7080 5380 7081
rect 4960 7016 4978 7080
rect 5042 7016 5058 7080
rect 5122 7016 5138 7080
rect 5202 7016 5218 7080
rect 5282 7016 5298 7080
rect 5362 7016 5380 7080
rect 4960 7015 5380 7016
rect 6891 7080 7311 7081
rect 6891 7016 6909 7080
rect 6973 7016 6989 7080
rect 7053 7016 7069 7080
rect 7133 7016 7149 7080
rect 7213 7016 7229 7080
rect 7293 7016 7311 7080
rect 6891 7015 7311 7016
rect 3995 6536 4415 6537
rect 3995 6472 4013 6536
rect 4077 6472 4093 6536
rect 4157 6472 4173 6536
rect 4237 6472 4253 6536
rect 4317 6472 4333 6536
rect 4397 6472 4415 6536
rect 3995 6471 4415 6472
rect 5926 6536 6346 6537
rect 5926 6472 5944 6536
rect 6008 6472 6024 6536
rect 6088 6472 6104 6536
rect 6168 6472 6184 6536
rect 6248 6472 6264 6536
rect 6328 6472 6346 6536
rect 5926 6471 6346 6472
rect 7856 6536 8276 6537
rect 7856 6472 7874 6536
rect 7938 6472 7954 6536
rect 8018 6472 8034 6536
rect 8098 6472 8114 6536
rect 8178 6472 8194 6536
rect 8258 6472 8276 6536
rect 7856 6471 8276 6472
rect 4960 5992 5380 5993
rect 4960 5928 4978 5992
rect 5042 5928 5058 5992
rect 5122 5928 5138 5992
rect 5202 5928 5218 5992
rect 5282 5928 5298 5992
rect 5362 5928 5380 5992
rect 4960 5927 5380 5928
rect 6891 5992 7311 5993
rect 6891 5928 6909 5992
rect 6973 5928 6989 5992
rect 7053 5928 7069 5992
rect 7133 5928 7149 5992
rect 7213 5928 7229 5992
rect 7293 5928 7311 5992
rect 6891 5927 7311 5928
rect 3995 5448 4415 5449
rect 3995 5384 4013 5448
rect 4077 5384 4093 5448
rect 4157 5384 4173 5448
rect 4237 5384 4253 5448
rect 4317 5384 4333 5448
rect 4397 5384 4415 5448
rect 3995 5383 4415 5384
rect 5926 5448 6346 5449
rect 5926 5384 5944 5448
rect 6008 5384 6024 5448
rect 6088 5384 6104 5448
rect 6168 5384 6184 5448
rect 6248 5384 6264 5448
rect 6328 5384 6346 5448
rect 5926 5383 6346 5384
rect 7856 5448 8276 5449
rect 7856 5384 7874 5448
rect 7938 5384 7954 5448
rect 8018 5384 8034 5448
rect 8098 5384 8114 5448
rect 8178 5384 8194 5448
rect 8258 5384 8276 5448
rect 7856 5383 8276 5384
rect 4960 4904 5380 4905
rect 4960 4840 4978 4904
rect 5042 4840 5058 4904
rect 5122 4840 5138 4904
rect 5202 4840 5218 4904
rect 5282 4840 5298 4904
rect 5362 4840 5380 4904
rect 4960 4839 5380 4840
rect 6891 4904 7311 4905
rect 6891 4840 6909 4904
rect 6973 4840 6989 4904
rect 7053 4840 7069 4904
rect 7133 4840 7149 4904
rect 7213 4840 7229 4904
rect 7293 4840 7311 4904
rect 6891 4839 7311 4840
rect 3995 4360 4415 4361
rect 3995 4296 4013 4360
rect 4077 4296 4093 4360
rect 4157 4296 4173 4360
rect 4237 4296 4253 4360
rect 4317 4296 4333 4360
rect 4397 4296 4415 4360
rect 3995 4295 4415 4296
rect 5926 4360 6346 4361
rect 5926 4296 5944 4360
rect 6008 4296 6024 4360
rect 6088 4296 6104 4360
rect 6168 4296 6184 4360
rect 6248 4296 6264 4360
rect 6328 4296 6346 4360
rect 5926 4295 6346 4296
rect 7856 4360 8276 4361
rect 7856 4296 7874 4360
rect 7938 4296 7954 4360
rect 8018 4296 8034 4360
rect 8098 4296 8114 4360
rect 8178 4296 8194 4360
rect 8258 4296 8276 4360
rect 7856 4295 8276 4296
rect 4960 3816 5380 3817
rect 4960 3752 4978 3816
rect 5042 3752 5058 3816
rect 5122 3752 5138 3816
rect 5202 3752 5218 3816
rect 5282 3752 5298 3816
rect 5362 3752 5380 3816
rect 4960 3751 5380 3752
rect 6891 3816 7311 3817
rect 6891 3752 6909 3816
rect 6973 3752 6989 3816
rect 7053 3752 7069 3816
rect 7133 3752 7149 3816
rect 7213 3752 7229 3816
rect 7293 3752 7311 3816
rect 6891 3751 7311 3752
rect 3995 3272 4415 3273
rect 3995 3208 4013 3272
rect 4077 3208 4093 3272
rect 4157 3208 4173 3272
rect 4237 3208 4253 3272
rect 4317 3208 4333 3272
rect 4397 3208 4415 3272
rect 3995 3207 4415 3208
rect 5926 3272 6346 3273
rect 5926 3208 5944 3272
rect 6008 3208 6024 3272
rect 6088 3208 6104 3272
rect 6168 3208 6184 3272
rect 6248 3208 6264 3272
rect 6328 3208 6346 3272
rect 5926 3207 6346 3208
rect 7856 3272 8276 3273
rect 7856 3208 7874 3272
rect 7938 3208 7954 3272
rect 8018 3208 8034 3272
rect 8098 3208 8114 3272
rect 8178 3208 8194 3272
rect 8258 3208 8276 3272
rect 7856 3207 8276 3208
rect 1140 1932 11044 1940
rect 1140 1868 1148 1932
rect 1212 1868 1228 1932
rect 1292 1868 1308 1932
rect 1372 1868 1388 1932
rect 1452 1868 1468 1932
rect 1532 1868 1548 1932
rect 1612 1868 1628 1932
rect 1692 1868 1708 1932
rect 1772 1868 1788 1932
rect 1852 1868 1868 1932
rect 1932 1868 4013 1932
rect 4077 1868 4093 1932
rect 4157 1868 4173 1932
rect 4237 1868 4253 1932
rect 4317 1868 4333 1932
rect 4397 1868 5944 1932
rect 6008 1868 6024 1932
rect 6088 1868 6104 1932
rect 6168 1868 6184 1932
rect 6248 1868 6264 1932
rect 6328 1868 7874 1932
rect 7938 1868 7954 1932
rect 8018 1868 8034 1932
rect 8098 1868 8114 1932
rect 8178 1868 8194 1932
rect 8258 1868 10252 1932
rect 10316 1868 10332 1932
rect 10396 1868 10412 1932
rect 10476 1868 10492 1932
rect 10556 1868 10572 1932
rect 10636 1868 10652 1932
rect 10716 1868 10732 1932
rect 10796 1868 10812 1932
rect 10876 1868 10892 1932
rect 10956 1868 10972 1932
rect 11036 1868 11044 1932
rect 1140 1852 11044 1868
rect 1140 1788 1148 1852
rect 1212 1788 1228 1852
rect 1292 1788 1308 1852
rect 1372 1788 1388 1852
rect 1452 1788 1468 1852
rect 1532 1788 1548 1852
rect 1612 1788 1628 1852
rect 1692 1788 1708 1852
rect 1772 1788 1788 1852
rect 1852 1788 1868 1852
rect 1932 1788 4013 1852
rect 4077 1788 4093 1852
rect 4157 1788 4173 1852
rect 4237 1788 4253 1852
rect 4317 1788 4333 1852
rect 4397 1788 5944 1852
rect 6008 1788 6024 1852
rect 6088 1788 6104 1852
rect 6168 1788 6184 1852
rect 6248 1788 6264 1852
rect 6328 1788 7874 1852
rect 7938 1788 7954 1852
rect 8018 1788 8034 1852
rect 8098 1788 8114 1852
rect 8178 1788 8194 1852
rect 8258 1788 10252 1852
rect 10316 1788 10332 1852
rect 10396 1788 10412 1852
rect 10476 1788 10492 1852
rect 10556 1788 10572 1852
rect 10636 1788 10652 1852
rect 10716 1788 10732 1852
rect 10796 1788 10812 1852
rect 10876 1788 10892 1852
rect 10956 1788 10972 1852
rect 11036 1788 11044 1852
rect 1140 1772 11044 1788
rect 1140 1708 1148 1772
rect 1212 1708 1228 1772
rect 1292 1708 1308 1772
rect 1372 1708 1388 1772
rect 1452 1708 1468 1772
rect 1532 1708 1548 1772
rect 1612 1708 1628 1772
rect 1692 1708 1708 1772
rect 1772 1708 1788 1772
rect 1852 1708 1868 1772
rect 1932 1708 4013 1772
rect 4077 1708 4093 1772
rect 4157 1708 4173 1772
rect 4237 1708 4253 1772
rect 4317 1708 4333 1772
rect 4397 1708 5944 1772
rect 6008 1708 6024 1772
rect 6088 1708 6104 1772
rect 6168 1708 6184 1772
rect 6248 1708 6264 1772
rect 6328 1708 7874 1772
rect 7938 1708 7954 1772
rect 8018 1708 8034 1772
rect 8098 1708 8114 1772
rect 8178 1708 8194 1772
rect 8258 1708 10252 1772
rect 10316 1708 10332 1772
rect 10396 1708 10412 1772
rect 10476 1708 10492 1772
rect 10556 1708 10572 1772
rect 10636 1708 10652 1772
rect 10716 1708 10732 1772
rect 10796 1708 10812 1772
rect 10876 1708 10892 1772
rect 10956 1708 10972 1772
rect 11036 1708 11044 1772
rect 1140 1692 11044 1708
rect 1140 1628 1148 1692
rect 1212 1628 1228 1692
rect 1292 1628 1308 1692
rect 1372 1628 1388 1692
rect 1452 1628 1468 1692
rect 1532 1628 1548 1692
rect 1612 1628 1628 1692
rect 1692 1628 1708 1692
rect 1772 1628 1788 1692
rect 1852 1628 1868 1692
rect 1932 1628 4013 1692
rect 4077 1628 4093 1692
rect 4157 1628 4173 1692
rect 4237 1628 4253 1692
rect 4317 1628 4333 1692
rect 4397 1628 5944 1692
rect 6008 1628 6024 1692
rect 6088 1628 6104 1692
rect 6168 1628 6184 1692
rect 6248 1628 6264 1692
rect 6328 1628 7874 1692
rect 7938 1628 7954 1692
rect 8018 1628 8034 1692
rect 8098 1628 8114 1692
rect 8178 1628 8194 1692
rect 8258 1628 10252 1692
rect 10316 1628 10332 1692
rect 10396 1628 10412 1692
rect 10476 1628 10492 1692
rect 10556 1628 10572 1692
rect 10636 1628 10652 1692
rect 10716 1628 10732 1692
rect 10796 1628 10812 1692
rect 10876 1628 10892 1692
rect 10956 1628 10972 1692
rect 11036 1628 11044 1692
rect 1140 1612 11044 1628
rect 1140 1548 1148 1612
rect 1212 1548 1228 1612
rect 1292 1548 1308 1612
rect 1372 1548 1388 1612
rect 1452 1548 1468 1612
rect 1532 1548 1548 1612
rect 1612 1548 1628 1612
rect 1692 1548 1708 1612
rect 1772 1548 1788 1612
rect 1852 1548 1868 1612
rect 1932 1548 4013 1612
rect 4077 1548 4093 1612
rect 4157 1548 4173 1612
rect 4237 1548 4253 1612
rect 4317 1548 4333 1612
rect 4397 1548 5944 1612
rect 6008 1548 6024 1612
rect 6088 1548 6104 1612
rect 6168 1548 6184 1612
rect 6248 1548 6264 1612
rect 6328 1548 7874 1612
rect 7938 1548 7954 1612
rect 8018 1548 8034 1612
rect 8098 1548 8114 1612
rect 8178 1548 8194 1612
rect 8258 1548 10252 1612
rect 10316 1548 10332 1612
rect 10396 1548 10412 1612
rect 10476 1548 10492 1612
rect 10556 1548 10572 1612
rect 10636 1548 10652 1612
rect 10716 1548 10732 1612
rect 10796 1548 10812 1612
rect 10876 1548 10892 1612
rect 10956 1548 10972 1612
rect 11036 1548 11044 1612
rect 1140 1532 11044 1548
rect 1140 1468 1148 1532
rect 1212 1468 1228 1532
rect 1292 1468 1308 1532
rect 1372 1468 1388 1532
rect 1452 1468 1468 1532
rect 1532 1468 1548 1532
rect 1612 1468 1628 1532
rect 1692 1468 1708 1532
rect 1772 1468 1788 1532
rect 1852 1468 1868 1532
rect 1932 1468 4013 1532
rect 4077 1468 4093 1532
rect 4157 1468 4173 1532
rect 4237 1468 4253 1532
rect 4317 1468 4333 1532
rect 4397 1468 5944 1532
rect 6008 1468 6024 1532
rect 6088 1468 6104 1532
rect 6168 1468 6184 1532
rect 6248 1468 6264 1532
rect 6328 1468 7874 1532
rect 7938 1468 7954 1532
rect 8018 1468 8034 1532
rect 8098 1468 8114 1532
rect 8178 1468 8194 1532
rect 8258 1468 10252 1532
rect 10316 1468 10332 1532
rect 10396 1468 10412 1532
rect 10476 1468 10492 1532
rect 10556 1468 10572 1532
rect 10636 1468 10652 1532
rect 10716 1468 10732 1532
rect 10796 1468 10812 1532
rect 10876 1468 10892 1532
rect 10956 1468 10972 1532
rect 11036 1468 11044 1532
rect 1140 1452 11044 1468
rect 1140 1388 1148 1452
rect 1212 1388 1228 1452
rect 1292 1388 1308 1452
rect 1372 1388 1388 1452
rect 1452 1388 1468 1452
rect 1532 1388 1548 1452
rect 1612 1388 1628 1452
rect 1692 1388 1708 1452
rect 1772 1388 1788 1452
rect 1852 1388 1868 1452
rect 1932 1388 4013 1452
rect 4077 1388 4093 1452
rect 4157 1388 4173 1452
rect 4237 1388 4253 1452
rect 4317 1388 4333 1452
rect 4397 1388 5944 1452
rect 6008 1388 6024 1452
rect 6088 1388 6104 1452
rect 6168 1388 6184 1452
rect 6248 1388 6264 1452
rect 6328 1388 7874 1452
rect 7938 1388 7954 1452
rect 8018 1388 8034 1452
rect 8098 1388 8114 1452
rect 8178 1388 8194 1452
rect 8258 1388 10252 1452
rect 10316 1388 10332 1452
rect 10396 1388 10412 1452
rect 10476 1388 10492 1452
rect 10556 1388 10572 1452
rect 10636 1388 10652 1452
rect 10716 1388 10732 1452
rect 10796 1388 10812 1452
rect 10876 1388 10892 1452
rect 10956 1388 10972 1452
rect 11036 1388 11044 1452
rect 1140 1372 11044 1388
rect 1140 1308 1148 1372
rect 1212 1308 1228 1372
rect 1292 1308 1308 1372
rect 1372 1308 1388 1372
rect 1452 1308 1468 1372
rect 1532 1308 1548 1372
rect 1612 1308 1628 1372
rect 1692 1308 1708 1372
rect 1772 1308 1788 1372
rect 1852 1308 1868 1372
rect 1932 1308 4013 1372
rect 4077 1308 4093 1372
rect 4157 1308 4173 1372
rect 4237 1308 4253 1372
rect 4317 1308 4333 1372
rect 4397 1308 5944 1372
rect 6008 1308 6024 1372
rect 6088 1308 6104 1372
rect 6168 1308 6184 1372
rect 6248 1308 6264 1372
rect 6328 1308 7874 1372
rect 7938 1308 7954 1372
rect 8018 1308 8034 1372
rect 8098 1308 8114 1372
rect 8178 1308 8194 1372
rect 8258 1308 10252 1372
rect 10316 1308 10332 1372
rect 10396 1308 10412 1372
rect 10476 1308 10492 1372
rect 10556 1308 10572 1372
rect 10636 1308 10652 1372
rect 10716 1308 10732 1372
rect 10796 1308 10812 1372
rect 10876 1308 10892 1372
rect 10956 1308 10972 1372
rect 11036 1308 11044 1372
rect 1140 1292 11044 1308
rect 1140 1228 1148 1292
rect 1212 1228 1228 1292
rect 1292 1228 1308 1292
rect 1372 1228 1388 1292
rect 1452 1228 1468 1292
rect 1532 1228 1548 1292
rect 1612 1228 1628 1292
rect 1692 1228 1708 1292
rect 1772 1228 1788 1292
rect 1852 1228 1868 1292
rect 1932 1228 4013 1292
rect 4077 1228 4093 1292
rect 4157 1228 4173 1292
rect 4237 1228 4253 1292
rect 4317 1228 4333 1292
rect 4397 1228 5944 1292
rect 6008 1228 6024 1292
rect 6088 1228 6104 1292
rect 6168 1228 6184 1292
rect 6248 1228 6264 1292
rect 6328 1228 7874 1292
rect 7938 1228 7954 1292
rect 8018 1228 8034 1292
rect 8098 1228 8114 1292
rect 8178 1228 8194 1292
rect 8258 1228 10252 1292
rect 10316 1228 10332 1292
rect 10396 1228 10412 1292
rect 10476 1228 10492 1292
rect 10556 1228 10572 1292
rect 10636 1228 10652 1292
rect 10716 1228 10732 1292
rect 10796 1228 10812 1292
rect 10876 1228 10892 1292
rect 10956 1228 10972 1292
rect 11036 1228 11044 1292
rect 1140 1212 11044 1228
rect 1140 1148 1148 1212
rect 1212 1148 1228 1212
rect 1292 1148 1308 1212
rect 1372 1148 1388 1212
rect 1452 1148 1468 1212
rect 1532 1148 1548 1212
rect 1612 1148 1628 1212
rect 1692 1148 1708 1212
rect 1772 1148 1788 1212
rect 1852 1148 1868 1212
rect 1932 1148 4013 1212
rect 4077 1148 4093 1212
rect 4157 1148 4173 1212
rect 4237 1148 4253 1212
rect 4317 1148 4333 1212
rect 4397 1148 5944 1212
rect 6008 1148 6024 1212
rect 6088 1148 6104 1212
rect 6168 1148 6184 1212
rect 6248 1148 6264 1212
rect 6328 1148 7874 1212
rect 7938 1148 7954 1212
rect 8018 1148 8034 1212
rect 8098 1148 8114 1212
rect 8178 1148 8194 1212
rect 8258 1148 10252 1212
rect 10316 1148 10332 1212
rect 10396 1148 10412 1212
rect 10476 1148 10492 1212
rect 10556 1148 10572 1212
rect 10636 1148 10652 1212
rect 10716 1148 10732 1212
rect 10796 1148 10812 1212
rect 10876 1148 10892 1212
rect 10956 1148 10972 1212
rect 11036 1148 11044 1212
rect 1140 1140 11044 1148
rect 0 792 12184 800
rect 0 728 8 792
rect 72 728 88 792
rect 152 728 168 792
rect 232 728 248 792
rect 312 728 328 792
rect 392 728 408 792
rect 472 728 488 792
rect 552 728 568 792
rect 632 728 648 792
rect 712 728 728 792
rect 792 728 4978 792
rect 5042 728 5058 792
rect 5122 728 5138 792
rect 5202 728 5218 792
rect 5282 728 5298 792
rect 5362 728 6909 792
rect 6973 728 6989 792
rect 7053 728 7069 792
rect 7133 728 7149 792
rect 7213 728 7229 792
rect 7293 728 11392 792
rect 11456 728 11472 792
rect 11536 728 11552 792
rect 11616 728 11632 792
rect 11696 728 11712 792
rect 11776 728 11792 792
rect 11856 728 11872 792
rect 11936 728 11952 792
rect 12016 728 12032 792
rect 12096 728 12112 792
rect 12176 728 12184 792
rect 0 712 12184 728
rect 0 648 8 712
rect 72 648 88 712
rect 152 648 168 712
rect 232 648 248 712
rect 312 648 328 712
rect 392 648 408 712
rect 472 648 488 712
rect 552 648 568 712
rect 632 648 648 712
rect 712 648 728 712
rect 792 648 4978 712
rect 5042 648 5058 712
rect 5122 648 5138 712
rect 5202 648 5218 712
rect 5282 648 5298 712
rect 5362 648 6909 712
rect 6973 648 6989 712
rect 7053 648 7069 712
rect 7133 648 7149 712
rect 7213 648 7229 712
rect 7293 648 11392 712
rect 11456 648 11472 712
rect 11536 648 11552 712
rect 11616 648 11632 712
rect 11696 648 11712 712
rect 11776 648 11792 712
rect 11856 648 11872 712
rect 11936 648 11952 712
rect 12016 648 12032 712
rect 12096 648 12112 712
rect 12176 648 12184 712
rect 0 632 12184 648
rect 0 568 8 632
rect 72 568 88 632
rect 152 568 168 632
rect 232 568 248 632
rect 312 568 328 632
rect 392 568 408 632
rect 472 568 488 632
rect 552 568 568 632
rect 632 568 648 632
rect 712 568 728 632
rect 792 568 4978 632
rect 5042 568 5058 632
rect 5122 568 5138 632
rect 5202 568 5218 632
rect 5282 568 5298 632
rect 5362 568 6909 632
rect 6973 568 6989 632
rect 7053 568 7069 632
rect 7133 568 7149 632
rect 7213 568 7229 632
rect 7293 568 11392 632
rect 11456 568 11472 632
rect 11536 568 11552 632
rect 11616 568 11632 632
rect 11696 568 11712 632
rect 11776 568 11792 632
rect 11856 568 11872 632
rect 11936 568 11952 632
rect 12016 568 12032 632
rect 12096 568 12112 632
rect 12176 568 12184 632
rect 0 552 12184 568
rect 0 488 8 552
rect 72 488 88 552
rect 152 488 168 552
rect 232 488 248 552
rect 312 488 328 552
rect 392 488 408 552
rect 472 488 488 552
rect 552 488 568 552
rect 632 488 648 552
rect 712 488 728 552
rect 792 488 4978 552
rect 5042 488 5058 552
rect 5122 488 5138 552
rect 5202 488 5218 552
rect 5282 488 5298 552
rect 5362 488 6909 552
rect 6973 488 6989 552
rect 7053 488 7069 552
rect 7133 488 7149 552
rect 7213 488 7229 552
rect 7293 488 11392 552
rect 11456 488 11472 552
rect 11536 488 11552 552
rect 11616 488 11632 552
rect 11696 488 11712 552
rect 11776 488 11792 552
rect 11856 488 11872 552
rect 11936 488 11952 552
rect 12016 488 12032 552
rect 12096 488 12112 552
rect 12176 488 12184 552
rect 0 472 12184 488
rect 0 408 8 472
rect 72 408 88 472
rect 152 408 168 472
rect 232 408 248 472
rect 312 408 328 472
rect 392 408 408 472
rect 472 408 488 472
rect 552 408 568 472
rect 632 408 648 472
rect 712 408 728 472
rect 792 408 4978 472
rect 5042 408 5058 472
rect 5122 408 5138 472
rect 5202 408 5218 472
rect 5282 408 5298 472
rect 5362 408 6909 472
rect 6973 408 6989 472
rect 7053 408 7069 472
rect 7133 408 7149 472
rect 7213 408 7229 472
rect 7293 408 11392 472
rect 11456 408 11472 472
rect 11536 408 11552 472
rect 11616 408 11632 472
rect 11696 408 11712 472
rect 11776 408 11792 472
rect 11856 408 11872 472
rect 11936 408 11952 472
rect 12016 408 12032 472
rect 12096 408 12112 472
rect 12176 408 12184 472
rect 0 392 12184 408
rect 0 328 8 392
rect 72 328 88 392
rect 152 328 168 392
rect 232 328 248 392
rect 312 328 328 392
rect 392 328 408 392
rect 472 328 488 392
rect 552 328 568 392
rect 632 328 648 392
rect 712 328 728 392
rect 792 328 4978 392
rect 5042 328 5058 392
rect 5122 328 5138 392
rect 5202 328 5218 392
rect 5282 328 5298 392
rect 5362 328 6909 392
rect 6973 328 6989 392
rect 7053 328 7069 392
rect 7133 328 7149 392
rect 7213 328 7229 392
rect 7293 328 11392 392
rect 11456 328 11472 392
rect 11536 328 11552 392
rect 11616 328 11632 392
rect 11696 328 11712 392
rect 11776 328 11792 392
rect 11856 328 11872 392
rect 11936 328 11952 392
rect 12016 328 12032 392
rect 12096 328 12112 392
rect 12176 328 12184 392
rect 0 312 12184 328
rect 0 248 8 312
rect 72 248 88 312
rect 152 248 168 312
rect 232 248 248 312
rect 312 248 328 312
rect 392 248 408 312
rect 472 248 488 312
rect 552 248 568 312
rect 632 248 648 312
rect 712 248 728 312
rect 792 248 4978 312
rect 5042 248 5058 312
rect 5122 248 5138 312
rect 5202 248 5218 312
rect 5282 248 5298 312
rect 5362 248 6909 312
rect 6973 248 6989 312
rect 7053 248 7069 312
rect 7133 248 7149 312
rect 7213 248 7229 312
rect 7293 248 11392 312
rect 11456 248 11472 312
rect 11536 248 11552 312
rect 11616 248 11632 312
rect 11696 248 11712 312
rect 11776 248 11792 312
rect 11856 248 11872 312
rect 11936 248 11952 312
rect 12016 248 12032 312
rect 12096 248 12112 312
rect 12176 248 12184 312
rect 0 232 12184 248
rect 0 168 8 232
rect 72 168 88 232
rect 152 168 168 232
rect 232 168 248 232
rect 312 168 328 232
rect 392 168 408 232
rect 472 168 488 232
rect 552 168 568 232
rect 632 168 648 232
rect 712 168 728 232
rect 792 168 4978 232
rect 5042 168 5058 232
rect 5122 168 5138 232
rect 5202 168 5218 232
rect 5282 168 5298 232
rect 5362 168 6909 232
rect 6973 168 6989 232
rect 7053 168 7069 232
rect 7133 168 7149 232
rect 7213 168 7229 232
rect 7293 168 11392 232
rect 11456 168 11472 232
rect 11536 168 11552 232
rect 11616 168 11632 232
rect 11696 168 11712 232
rect 11776 168 11792 232
rect 11856 168 11872 232
rect 11936 168 11952 232
rect 12016 168 12032 232
rect 12096 168 12112 232
rect 12176 168 12184 232
rect 0 152 12184 168
rect 0 88 8 152
rect 72 88 88 152
rect 152 88 168 152
rect 232 88 248 152
rect 312 88 328 152
rect 392 88 408 152
rect 472 88 488 152
rect 552 88 568 152
rect 632 88 648 152
rect 712 88 728 152
rect 792 88 4978 152
rect 5042 88 5058 152
rect 5122 88 5138 152
rect 5202 88 5218 152
rect 5282 88 5298 152
rect 5362 88 6909 152
rect 6973 88 6989 152
rect 7053 88 7069 152
rect 7133 88 7149 152
rect 7213 88 7229 152
rect 7293 88 11392 152
rect 11456 88 11472 152
rect 11536 88 11552 152
rect 11616 88 11632 152
rect 11696 88 11712 152
rect 11776 88 11792 152
rect 11856 88 11872 152
rect 11936 88 11952 152
rect 12016 88 12032 152
rect 12096 88 12112 152
rect 12176 88 12184 152
rect 0 72 12184 88
rect 0 8 8 72
rect 72 8 88 72
rect 152 8 168 72
rect 232 8 248 72
rect 312 8 328 72
rect 392 8 408 72
rect 472 8 488 72
rect 552 8 568 72
rect 632 8 648 72
rect 712 8 728 72
rect 792 8 4978 72
rect 5042 8 5058 72
rect 5122 8 5138 72
rect 5202 8 5218 72
rect 5282 8 5298 72
rect 5362 8 6909 72
rect 6973 8 6989 72
rect 7053 8 7069 72
rect 7133 8 7149 72
rect 7213 8 7229 72
rect 7293 8 11392 72
rect 11456 8 11472 72
rect 11536 8 11552 72
rect 11616 8 11632 72
rect 11696 8 11712 72
rect 11776 8 11792 72
rect 11856 8 11872 72
rect 11936 8 11952 72
rect 12016 8 12032 72
rect 12096 8 12112 72
rect 12176 8 12184 72
rect 0 0 12184 8
<< via3 >>
rect 8 20008 72 20072
rect 88 20008 152 20072
rect 168 20008 232 20072
rect 248 20008 312 20072
rect 328 20008 392 20072
rect 408 20008 472 20072
rect 488 20008 552 20072
rect 568 20008 632 20072
rect 648 20008 712 20072
rect 728 20008 792 20072
rect 4978 20008 5042 20072
rect 5058 20008 5122 20072
rect 5138 20008 5202 20072
rect 5218 20008 5282 20072
rect 5298 20008 5362 20072
rect 6909 20008 6973 20072
rect 6989 20008 7053 20072
rect 7069 20008 7133 20072
rect 7149 20008 7213 20072
rect 7229 20008 7293 20072
rect 11392 20008 11456 20072
rect 11472 20008 11536 20072
rect 11552 20008 11616 20072
rect 11632 20008 11696 20072
rect 11712 20008 11776 20072
rect 11792 20008 11856 20072
rect 11872 20008 11936 20072
rect 11952 20008 12016 20072
rect 12032 20008 12096 20072
rect 12112 20008 12176 20072
rect 8 19928 72 19992
rect 88 19928 152 19992
rect 168 19928 232 19992
rect 248 19928 312 19992
rect 328 19928 392 19992
rect 408 19928 472 19992
rect 488 19928 552 19992
rect 568 19928 632 19992
rect 648 19928 712 19992
rect 728 19928 792 19992
rect 4978 19928 5042 19992
rect 5058 19928 5122 19992
rect 5138 19928 5202 19992
rect 5218 19928 5282 19992
rect 5298 19928 5362 19992
rect 6909 19928 6973 19992
rect 6989 19928 7053 19992
rect 7069 19928 7133 19992
rect 7149 19928 7213 19992
rect 7229 19928 7293 19992
rect 11392 19928 11456 19992
rect 11472 19928 11536 19992
rect 11552 19928 11616 19992
rect 11632 19928 11696 19992
rect 11712 19928 11776 19992
rect 11792 19928 11856 19992
rect 11872 19928 11936 19992
rect 11952 19928 12016 19992
rect 12032 19928 12096 19992
rect 12112 19928 12176 19992
rect 8 19848 72 19912
rect 88 19848 152 19912
rect 168 19848 232 19912
rect 248 19848 312 19912
rect 328 19848 392 19912
rect 408 19848 472 19912
rect 488 19848 552 19912
rect 568 19848 632 19912
rect 648 19848 712 19912
rect 728 19848 792 19912
rect 4978 19848 5042 19912
rect 5058 19848 5122 19912
rect 5138 19848 5202 19912
rect 5218 19848 5282 19912
rect 5298 19848 5362 19912
rect 6909 19848 6973 19912
rect 6989 19848 7053 19912
rect 7069 19848 7133 19912
rect 7149 19848 7213 19912
rect 7229 19848 7293 19912
rect 11392 19848 11456 19912
rect 11472 19848 11536 19912
rect 11552 19848 11616 19912
rect 11632 19848 11696 19912
rect 11712 19848 11776 19912
rect 11792 19848 11856 19912
rect 11872 19848 11936 19912
rect 11952 19848 12016 19912
rect 12032 19848 12096 19912
rect 12112 19848 12176 19912
rect 8 19768 72 19832
rect 88 19768 152 19832
rect 168 19768 232 19832
rect 248 19768 312 19832
rect 328 19768 392 19832
rect 408 19768 472 19832
rect 488 19768 552 19832
rect 568 19768 632 19832
rect 648 19768 712 19832
rect 728 19768 792 19832
rect 4978 19768 5042 19832
rect 5058 19768 5122 19832
rect 5138 19768 5202 19832
rect 5218 19768 5282 19832
rect 5298 19768 5362 19832
rect 6909 19768 6973 19832
rect 6989 19768 7053 19832
rect 7069 19768 7133 19832
rect 7149 19768 7213 19832
rect 7229 19768 7293 19832
rect 11392 19768 11456 19832
rect 11472 19768 11536 19832
rect 11552 19768 11616 19832
rect 11632 19768 11696 19832
rect 11712 19768 11776 19832
rect 11792 19768 11856 19832
rect 11872 19768 11936 19832
rect 11952 19768 12016 19832
rect 12032 19768 12096 19832
rect 12112 19768 12176 19832
rect 8 19688 72 19752
rect 88 19688 152 19752
rect 168 19688 232 19752
rect 248 19688 312 19752
rect 328 19688 392 19752
rect 408 19688 472 19752
rect 488 19688 552 19752
rect 568 19688 632 19752
rect 648 19688 712 19752
rect 728 19688 792 19752
rect 4978 19688 5042 19752
rect 5058 19688 5122 19752
rect 5138 19688 5202 19752
rect 5218 19688 5282 19752
rect 5298 19688 5362 19752
rect 6909 19688 6973 19752
rect 6989 19688 7053 19752
rect 7069 19688 7133 19752
rect 7149 19688 7213 19752
rect 7229 19688 7293 19752
rect 11392 19688 11456 19752
rect 11472 19688 11536 19752
rect 11552 19688 11616 19752
rect 11632 19688 11696 19752
rect 11712 19688 11776 19752
rect 11792 19688 11856 19752
rect 11872 19688 11936 19752
rect 11952 19688 12016 19752
rect 12032 19688 12096 19752
rect 12112 19688 12176 19752
rect 8 19608 72 19672
rect 88 19608 152 19672
rect 168 19608 232 19672
rect 248 19608 312 19672
rect 328 19608 392 19672
rect 408 19608 472 19672
rect 488 19608 552 19672
rect 568 19608 632 19672
rect 648 19608 712 19672
rect 728 19608 792 19672
rect 4978 19608 5042 19672
rect 5058 19608 5122 19672
rect 5138 19608 5202 19672
rect 5218 19608 5282 19672
rect 5298 19608 5362 19672
rect 6909 19608 6973 19672
rect 6989 19608 7053 19672
rect 7069 19608 7133 19672
rect 7149 19608 7213 19672
rect 7229 19608 7293 19672
rect 11392 19608 11456 19672
rect 11472 19608 11536 19672
rect 11552 19608 11616 19672
rect 11632 19608 11696 19672
rect 11712 19608 11776 19672
rect 11792 19608 11856 19672
rect 11872 19608 11936 19672
rect 11952 19608 12016 19672
rect 12032 19608 12096 19672
rect 12112 19608 12176 19672
rect 8 19528 72 19592
rect 88 19528 152 19592
rect 168 19528 232 19592
rect 248 19528 312 19592
rect 328 19528 392 19592
rect 408 19528 472 19592
rect 488 19528 552 19592
rect 568 19528 632 19592
rect 648 19528 712 19592
rect 728 19528 792 19592
rect 4978 19528 5042 19592
rect 5058 19528 5122 19592
rect 5138 19528 5202 19592
rect 5218 19528 5282 19592
rect 5298 19528 5362 19592
rect 6909 19528 6973 19592
rect 6989 19528 7053 19592
rect 7069 19528 7133 19592
rect 7149 19528 7213 19592
rect 7229 19528 7293 19592
rect 11392 19528 11456 19592
rect 11472 19528 11536 19592
rect 11552 19528 11616 19592
rect 11632 19528 11696 19592
rect 11712 19528 11776 19592
rect 11792 19528 11856 19592
rect 11872 19528 11936 19592
rect 11952 19528 12016 19592
rect 12032 19528 12096 19592
rect 12112 19528 12176 19592
rect 8 19448 72 19512
rect 88 19448 152 19512
rect 168 19448 232 19512
rect 248 19448 312 19512
rect 328 19448 392 19512
rect 408 19448 472 19512
rect 488 19448 552 19512
rect 568 19448 632 19512
rect 648 19448 712 19512
rect 728 19448 792 19512
rect 4978 19448 5042 19512
rect 5058 19448 5122 19512
rect 5138 19448 5202 19512
rect 5218 19448 5282 19512
rect 5298 19448 5362 19512
rect 6909 19448 6973 19512
rect 6989 19448 7053 19512
rect 7069 19448 7133 19512
rect 7149 19448 7213 19512
rect 7229 19448 7293 19512
rect 11392 19448 11456 19512
rect 11472 19448 11536 19512
rect 11552 19448 11616 19512
rect 11632 19448 11696 19512
rect 11712 19448 11776 19512
rect 11792 19448 11856 19512
rect 11872 19448 11936 19512
rect 11952 19448 12016 19512
rect 12032 19448 12096 19512
rect 12112 19448 12176 19512
rect 8 19368 72 19432
rect 88 19368 152 19432
rect 168 19368 232 19432
rect 248 19368 312 19432
rect 328 19368 392 19432
rect 408 19368 472 19432
rect 488 19368 552 19432
rect 568 19368 632 19432
rect 648 19368 712 19432
rect 728 19368 792 19432
rect 4978 19368 5042 19432
rect 5058 19368 5122 19432
rect 5138 19368 5202 19432
rect 5218 19368 5282 19432
rect 5298 19368 5362 19432
rect 6909 19368 6973 19432
rect 6989 19368 7053 19432
rect 7069 19368 7133 19432
rect 7149 19368 7213 19432
rect 7229 19368 7293 19432
rect 11392 19368 11456 19432
rect 11472 19368 11536 19432
rect 11552 19368 11616 19432
rect 11632 19368 11696 19432
rect 11712 19368 11776 19432
rect 11792 19368 11856 19432
rect 11872 19368 11936 19432
rect 11952 19368 12016 19432
rect 12032 19368 12096 19432
rect 12112 19368 12176 19432
rect 8 19288 72 19352
rect 88 19288 152 19352
rect 168 19288 232 19352
rect 248 19288 312 19352
rect 328 19288 392 19352
rect 408 19288 472 19352
rect 488 19288 552 19352
rect 568 19288 632 19352
rect 648 19288 712 19352
rect 728 19288 792 19352
rect 4978 19288 5042 19352
rect 5058 19288 5122 19352
rect 5138 19288 5202 19352
rect 5218 19288 5282 19352
rect 5298 19288 5362 19352
rect 6909 19288 6973 19352
rect 6989 19288 7053 19352
rect 7069 19288 7133 19352
rect 7149 19288 7213 19352
rect 7229 19288 7293 19352
rect 11392 19288 11456 19352
rect 11472 19288 11536 19352
rect 11552 19288 11616 19352
rect 11632 19288 11696 19352
rect 11712 19288 11776 19352
rect 11792 19288 11856 19352
rect 11872 19288 11936 19352
rect 11952 19288 12016 19352
rect 12032 19288 12096 19352
rect 12112 19288 12176 19352
rect 1148 18868 1212 18932
rect 1228 18868 1292 18932
rect 1308 18868 1372 18932
rect 1388 18868 1452 18932
rect 1468 18868 1532 18932
rect 1548 18868 1612 18932
rect 1628 18868 1692 18932
rect 1708 18868 1772 18932
rect 1788 18868 1852 18932
rect 1868 18868 1932 18932
rect 4013 18868 4077 18932
rect 4093 18868 4157 18932
rect 4173 18868 4237 18932
rect 4253 18868 4317 18932
rect 4333 18868 4397 18932
rect 5944 18868 6008 18932
rect 6024 18868 6088 18932
rect 6104 18868 6168 18932
rect 6184 18868 6248 18932
rect 6264 18868 6328 18932
rect 7874 18868 7938 18932
rect 7954 18868 8018 18932
rect 8034 18868 8098 18932
rect 8114 18868 8178 18932
rect 8194 18868 8258 18932
rect 10252 18868 10316 18932
rect 10332 18868 10396 18932
rect 10412 18868 10476 18932
rect 10492 18868 10556 18932
rect 10572 18868 10636 18932
rect 10652 18868 10716 18932
rect 10732 18868 10796 18932
rect 10812 18868 10876 18932
rect 10892 18868 10956 18932
rect 10972 18868 11036 18932
rect 1148 18788 1212 18852
rect 1228 18788 1292 18852
rect 1308 18788 1372 18852
rect 1388 18788 1452 18852
rect 1468 18788 1532 18852
rect 1548 18788 1612 18852
rect 1628 18788 1692 18852
rect 1708 18788 1772 18852
rect 1788 18788 1852 18852
rect 1868 18788 1932 18852
rect 4013 18788 4077 18852
rect 4093 18788 4157 18852
rect 4173 18788 4237 18852
rect 4253 18788 4317 18852
rect 4333 18788 4397 18852
rect 5944 18788 6008 18852
rect 6024 18788 6088 18852
rect 6104 18788 6168 18852
rect 6184 18788 6248 18852
rect 6264 18788 6328 18852
rect 7874 18788 7938 18852
rect 7954 18788 8018 18852
rect 8034 18788 8098 18852
rect 8114 18788 8178 18852
rect 8194 18788 8258 18852
rect 10252 18788 10316 18852
rect 10332 18788 10396 18852
rect 10412 18788 10476 18852
rect 10492 18788 10556 18852
rect 10572 18788 10636 18852
rect 10652 18788 10716 18852
rect 10732 18788 10796 18852
rect 10812 18788 10876 18852
rect 10892 18788 10956 18852
rect 10972 18788 11036 18852
rect 1148 18708 1212 18772
rect 1228 18708 1292 18772
rect 1308 18708 1372 18772
rect 1388 18708 1452 18772
rect 1468 18708 1532 18772
rect 1548 18708 1612 18772
rect 1628 18708 1692 18772
rect 1708 18708 1772 18772
rect 1788 18708 1852 18772
rect 1868 18708 1932 18772
rect 4013 18708 4077 18772
rect 4093 18708 4157 18772
rect 4173 18708 4237 18772
rect 4253 18708 4317 18772
rect 4333 18708 4397 18772
rect 5944 18708 6008 18772
rect 6024 18708 6088 18772
rect 6104 18708 6168 18772
rect 6184 18708 6248 18772
rect 6264 18708 6328 18772
rect 7874 18708 7938 18772
rect 7954 18708 8018 18772
rect 8034 18708 8098 18772
rect 8114 18708 8178 18772
rect 8194 18708 8258 18772
rect 10252 18708 10316 18772
rect 10332 18708 10396 18772
rect 10412 18708 10476 18772
rect 10492 18708 10556 18772
rect 10572 18708 10636 18772
rect 10652 18708 10716 18772
rect 10732 18708 10796 18772
rect 10812 18708 10876 18772
rect 10892 18708 10956 18772
rect 10972 18708 11036 18772
rect 1148 18628 1212 18692
rect 1228 18628 1292 18692
rect 1308 18628 1372 18692
rect 1388 18628 1452 18692
rect 1468 18628 1532 18692
rect 1548 18628 1612 18692
rect 1628 18628 1692 18692
rect 1708 18628 1772 18692
rect 1788 18628 1852 18692
rect 1868 18628 1932 18692
rect 4013 18628 4077 18692
rect 4093 18628 4157 18692
rect 4173 18628 4237 18692
rect 4253 18628 4317 18692
rect 4333 18628 4397 18692
rect 5944 18628 6008 18692
rect 6024 18628 6088 18692
rect 6104 18628 6168 18692
rect 6184 18628 6248 18692
rect 6264 18628 6328 18692
rect 7874 18628 7938 18692
rect 7954 18628 8018 18692
rect 8034 18628 8098 18692
rect 8114 18628 8178 18692
rect 8194 18628 8258 18692
rect 10252 18628 10316 18692
rect 10332 18628 10396 18692
rect 10412 18628 10476 18692
rect 10492 18628 10556 18692
rect 10572 18628 10636 18692
rect 10652 18628 10716 18692
rect 10732 18628 10796 18692
rect 10812 18628 10876 18692
rect 10892 18628 10956 18692
rect 10972 18628 11036 18692
rect 1148 18548 1212 18612
rect 1228 18548 1292 18612
rect 1308 18548 1372 18612
rect 1388 18548 1452 18612
rect 1468 18548 1532 18612
rect 1548 18548 1612 18612
rect 1628 18548 1692 18612
rect 1708 18548 1772 18612
rect 1788 18548 1852 18612
rect 1868 18548 1932 18612
rect 4013 18548 4077 18612
rect 4093 18548 4157 18612
rect 4173 18548 4237 18612
rect 4253 18548 4317 18612
rect 4333 18548 4397 18612
rect 5944 18548 6008 18612
rect 6024 18548 6088 18612
rect 6104 18548 6168 18612
rect 6184 18548 6248 18612
rect 6264 18548 6328 18612
rect 7874 18548 7938 18612
rect 7954 18548 8018 18612
rect 8034 18548 8098 18612
rect 8114 18548 8178 18612
rect 8194 18548 8258 18612
rect 10252 18548 10316 18612
rect 10332 18548 10396 18612
rect 10412 18548 10476 18612
rect 10492 18548 10556 18612
rect 10572 18548 10636 18612
rect 10652 18548 10716 18612
rect 10732 18548 10796 18612
rect 10812 18548 10876 18612
rect 10892 18548 10956 18612
rect 10972 18548 11036 18612
rect 1148 18468 1212 18532
rect 1228 18468 1292 18532
rect 1308 18468 1372 18532
rect 1388 18468 1452 18532
rect 1468 18468 1532 18532
rect 1548 18468 1612 18532
rect 1628 18468 1692 18532
rect 1708 18468 1772 18532
rect 1788 18468 1852 18532
rect 1868 18468 1932 18532
rect 4013 18468 4077 18532
rect 4093 18468 4157 18532
rect 4173 18468 4237 18532
rect 4253 18468 4317 18532
rect 4333 18468 4397 18532
rect 5944 18468 6008 18532
rect 6024 18468 6088 18532
rect 6104 18468 6168 18532
rect 6184 18468 6248 18532
rect 6264 18468 6328 18532
rect 7874 18468 7938 18532
rect 7954 18468 8018 18532
rect 8034 18468 8098 18532
rect 8114 18468 8178 18532
rect 8194 18468 8258 18532
rect 10252 18468 10316 18532
rect 10332 18468 10396 18532
rect 10412 18468 10476 18532
rect 10492 18468 10556 18532
rect 10572 18468 10636 18532
rect 10652 18468 10716 18532
rect 10732 18468 10796 18532
rect 10812 18468 10876 18532
rect 10892 18468 10956 18532
rect 10972 18468 11036 18532
rect 1148 18388 1212 18452
rect 1228 18388 1292 18452
rect 1308 18388 1372 18452
rect 1388 18388 1452 18452
rect 1468 18388 1532 18452
rect 1548 18388 1612 18452
rect 1628 18388 1692 18452
rect 1708 18388 1772 18452
rect 1788 18388 1852 18452
rect 1868 18388 1932 18452
rect 4013 18388 4077 18452
rect 4093 18388 4157 18452
rect 4173 18388 4237 18452
rect 4253 18388 4317 18452
rect 4333 18388 4397 18452
rect 5944 18388 6008 18452
rect 6024 18388 6088 18452
rect 6104 18388 6168 18452
rect 6184 18388 6248 18452
rect 6264 18388 6328 18452
rect 7874 18388 7938 18452
rect 7954 18388 8018 18452
rect 8034 18388 8098 18452
rect 8114 18388 8178 18452
rect 8194 18388 8258 18452
rect 10252 18388 10316 18452
rect 10332 18388 10396 18452
rect 10412 18388 10476 18452
rect 10492 18388 10556 18452
rect 10572 18388 10636 18452
rect 10652 18388 10716 18452
rect 10732 18388 10796 18452
rect 10812 18388 10876 18452
rect 10892 18388 10956 18452
rect 10972 18388 11036 18452
rect 1148 18308 1212 18372
rect 1228 18308 1292 18372
rect 1308 18308 1372 18372
rect 1388 18308 1452 18372
rect 1468 18308 1532 18372
rect 1548 18308 1612 18372
rect 1628 18308 1692 18372
rect 1708 18308 1772 18372
rect 1788 18308 1852 18372
rect 1868 18308 1932 18372
rect 4013 18308 4077 18372
rect 4093 18308 4157 18372
rect 4173 18308 4237 18372
rect 4253 18308 4317 18372
rect 4333 18308 4397 18372
rect 5944 18308 6008 18372
rect 6024 18308 6088 18372
rect 6104 18308 6168 18372
rect 6184 18308 6248 18372
rect 6264 18308 6328 18372
rect 7874 18308 7938 18372
rect 7954 18308 8018 18372
rect 8034 18308 8098 18372
rect 8114 18308 8178 18372
rect 8194 18308 8258 18372
rect 10252 18308 10316 18372
rect 10332 18308 10396 18372
rect 10412 18308 10476 18372
rect 10492 18308 10556 18372
rect 10572 18308 10636 18372
rect 10652 18308 10716 18372
rect 10732 18308 10796 18372
rect 10812 18308 10876 18372
rect 10892 18308 10956 18372
rect 10972 18308 11036 18372
rect 1148 18228 1212 18292
rect 1228 18228 1292 18292
rect 1308 18228 1372 18292
rect 1388 18228 1452 18292
rect 1468 18228 1532 18292
rect 1548 18228 1612 18292
rect 1628 18228 1692 18292
rect 1708 18228 1772 18292
rect 1788 18228 1852 18292
rect 1868 18228 1932 18292
rect 4013 18228 4077 18292
rect 4093 18228 4157 18292
rect 4173 18228 4237 18292
rect 4253 18228 4317 18292
rect 4333 18228 4397 18292
rect 5944 18228 6008 18292
rect 6024 18228 6088 18292
rect 6104 18228 6168 18292
rect 6184 18228 6248 18292
rect 6264 18228 6328 18292
rect 7874 18228 7938 18292
rect 7954 18228 8018 18292
rect 8034 18228 8098 18292
rect 8114 18228 8178 18292
rect 8194 18228 8258 18292
rect 10252 18228 10316 18292
rect 10332 18228 10396 18292
rect 10412 18228 10476 18292
rect 10492 18228 10556 18292
rect 10572 18228 10636 18292
rect 10652 18228 10716 18292
rect 10732 18228 10796 18292
rect 10812 18228 10876 18292
rect 10892 18228 10956 18292
rect 10972 18228 11036 18292
rect 1148 18148 1212 18212
rect 1228 18148 1292 18212
rect 1308 18148 1372 18212
rect 1388 18148 1452 18212
rect 1468 18148 1532 18212
rect 1548 18148 1612 18212
rect 1628 18148 1692 18212
rect 1708 18148 1772 18212
rect 1788 18148 1852 18212
rect 1868 18148 1932 18212
rect 4013 18148 4077 18212
rect 4093 18148 4157 18212
rect 4173 18148 4237 18212
rect 4253 18148 4317 18212
rect 4333 18148 4397 18212
rect 5944 18148 6008 18212
rect 6024 18148 6088 18212
rect 6104 18148 6168 18212
rect 6184 18148 6248 18212
rect 6264 18148 6328 18212
rect 7874 18148 7938 18212
rect 7954 18148 8018 18212
rect 8034 18148 8098 18212
rect 8114 18148 8178 18212
rect 8194 18148 8258 18212
rect 10252 18148 10316 18212
rect 10332 18148 10396 18212
rect 10412 18148 10476 18212
rect 10492 18148 10556 18212
rect 10572 18148 10636 18212
rect 10652 18148 10716 18212
rect 10732 18148 10796 18212
rect 10812 18148 10876 18212
rect 10892 18148 10956 18212
rect 10972 18148 11036 18212
rect 4978 16868 5042 16872
rect 4978 16812 4982 16868
rect 4982 16812 5038 16868
rect 5038 16812 5042 16868
rect 4978 16808 5042 16812
rect 5058 16868 5122 16872
rect 5058 16812 5062 16868
rect 5062 16812 5118 16868
rect 5118 16812 5122 16868
rect 5058 16808 5122 16812
rect 5138 16868 5202 16872
rect 5138 16812 5142 16868
rect 5142 16812 5198 16868
rect 5198 16812 5202 16868
rect 5138 16808 5202 16812
rect 5218 16868 5282 16872
rect 5218 16812 5222 16868
rect 5222 16812 5278 16868
rect 5278 16812 5282 16868
rect 5218 16808 5282 16812
rect 5298 16868 5362 16872
rect 5298 16812 5302 16868
rect 5302 16812 5358 16868
rect 5358 16812 5362 16868
rect 5298 16808 5362 16812
rect 6909 16868 6973 16872
rect 6909 16812 6913 16868
rect 6913 16812 6969 16868
rect 6969 16812 6973 16868
rect 6909 16808 6973 16812
rect 6989 16868 7053 16872
rect 6989 16812 6993 16868
rect 6993 16812 7049 16868
rect 7049 16812 7053 16868
rect 6989 16808 7053 16812
rect 7069 16868 7133 16872
rect 7069 16812 7073 16868
rect 7073 16812 7129 16868
rect 7129 16812 7133 16868
rect 7069 16808 7133 16812
rect 7149 16868 7213 16872
rect 7149 16812 7153 16868
rect 7153 16812 7209 16868
rect 7209 16812 7213 16868
rect 7149 16808 7213 16812
rect 7229 16868 7293 16872
rect 7229 16812 7233 16868
rect 7233 16812 7289 16868
rect 7289 16812 7293 16868
rect 7229 16808 7293 16812
rect 4013 16324 4077 16328
rect 4013 16268 4017 16324
rect 4017 16268 4073 16324
rect 4073 16268 4077 16324
rect 4013 16264 4077 16268
rect 4093 16324 4157 16328
rect 4093 16268 4097 16324
rect 4097 16268 4153 16324
rect 4153 16268 4157 16324
rect 4093 16264 4157 16268
rect 4173 16324 4237 16328
rect 4173 16268 4177 16324
rect 4177 16268 4233 16324
rect 4233 16268 4237 16324
rect 4173 16264 4237 16268
rect 4253 16324 4317 16328
rect 4253 16268 4257 16324
rect 4257 16268 4313 16324
rect 4313 16268 4317 16324
rect 4253 16264 4317 16268
rect 4333 16324 4397 16328
rect 4333 16268 4337 16324
rect 4337 16268 4393 16324
rect 4393 16268 4397 16324
rect 4333 16264 4397 16268
rect 5944 16324 6008 16328
rect 5944 16268 5948 16324
rect 5948 16268 6004 16324
rect 6004 16268 6008 16324
rect 5944 16264 6008 16268
rect 6024 16324 6088 16328
rect 6024 16268 6028 16324
rect 6028 16268 6084 16324
rect 6084 16268 6088 16324
rect 6024 16264 6088 16268
rect 6104 16324 6168 16328
rect 6104 16268 6108 16324
rect 6108 16268 6164 16324
rect 6164 16268 6168 16324
rect 6104 16264 6168 16268
rect 6184 16324 6248 16328
rect 6184 16268 6188 16324
rect 6188 16268 6244 16324
rect 6244 16268 6248 16324
rect 6184 16264 6248 16268
rect 6264 16324 6328 16328
rect 6264 16268 6268 16324
rect 6268 16268 6324 16324
rect 6324 16268 6328 16324
rect 6264 16264 6328 16268
rect 7874 16324 7938 16328
rect 7874 16268 7878 16324
rect 7878 16268 7934 16324
rect 7934 16268 7938 16324
rect 7874 16264 7938 16268
rect 7954 16324 8018 16328
rect 7954 16268 7958 16324
rect 7958 16268 8014 16324
rect 8014 16268 8018 16324
rect 7954 16264 8018 16268
rect 8034 16324 8098 16328
rect 8034 16268 8038 16324
rect 8038 16268 8094 16324
rect 8094 16268 8098 16324
rect 8034 16264 8098 16268
rect 8114 16324 8178 16328
rect 8114 16268 8118 16324
rect 8118 16268 8174 16324
rect 8174 16268 8178 16324
rect 8114 16264 8178 16268
rect 8194 16324 8258 16328
rect 8194 16268 8198 16324
rect 8198 16268 8254 16324
rect 8254 16268 8258 16324
rect 8194 16264 8258 16268
rect 4978 15780 5042 15784
rect 4978 15724 4982 15780
rect 4982 15724 5038 15780
rect 5038 15724 5042 15780
rect 4978 15720 5042 15724
rect 5058 15780 5122 15784
rect 5058 15724 5062 15780
rect 5062 15724 5118 15780
rect 5118 15724 5122 15780
rect 5058 15720 5122 15724
rect 5138 15780 5202 15784
rect 5138 15724 5142 15780
rect 5142 15724 5198 15780
rect 5198 15724 5202 15780
rect 5138 15720 5202 15724
rect 5218 15780 5282 15784
rect 5218 15724 5222 15780
rect 5222 15724 5278 15780
rect 5278 15724 5282 15780
rect 5218 15720 5282 15724
rect 5298 15780 5362 15784
rect 5298 15724 5302 15780
rect 5302 15724 5358 15780
rect 5358 15724 5362 15780
rect 5298 15720 5362 15724
rect 6909 15780 6973 15784
rect 6909 15724 6913 15780
rect 6913 15724 6969 15780
rect 6969 15724 6973 15780
rect 6909 15720 6973 15724
rect 6989 15780 7053 15784
rect 6989 15724 6993 15780
rect 6993 15724 7049 15780
rect 7049 15724 7053 15780
rect 6989 15720 7053 15724
rect 7069 15780 7133 15784
rect 7069 15724 7073 15780
rect 7073 15724 7129 15780
rect 7129 15724 7133 15780
rect 7069 15720 7133 15724
rect 7149 15780 7213 15784
rect 7149 15724 7153 15780
rect 7153 15724 7209 15780
rect 7209 15724 7213 15780
rect 7149 15720 7213 15724
rect 7229 15780 7293 15784
rect 7229 15724 7233 15780
rect 7233 15724 7289 15780
rect 7289 15724 7293 15780
rect 7229 15720 7293 15724
rect 4013 15236 4077 15240
rect 4013 15180 4017 15236
rect 4017 15180 4073 15236
rect 4073 15180 4077 15236
rect 4013 15176 4077 15180
rect 4093 15236 4157 15240
rect 4093 15180 4097 15236
rect 4097 15180 4153 15236
rect 4153 15180 4157 15236
rect 4093 15176 4157 15180
rect 4173 15236 4237 15240
rect 4173 15180 4177 15236
rect 4177 15180 4233 15236
rect 4233 15180 4237 15236
rect 4173 15176 4237 15180
rect 4253 15236 4317 15240
rect 4253 15180 4257 15236
rect 4257 15180 4313 15236
rect 4313 15180 4317 15236
rect 4253 15176 4317 15180
rect 4333 15236 4397 15240
rect 4333 15180 4337 15236
rect 4337 15180 4393 15236
rect 4393 15180 4397 15236
rect 4333 15176 4397 15180
rect 5944 15236 6008 15240
rect 5944 15180 5948 15236
rect 5948 15180 6004 15236
rect 6004 15180 6008 15236
rect 5944 15176 6008 15180
rect 6024 15236 6088 15240
rect 6024 15180 6028 15236
rect 6028 15180 6084 15236
rect 6084 15180 6088 15236
rect 6024 15176 6088 15180
rect 6104 15236 6168 15240
rect 6104 15180 6108 15236
rect 6108 15180 6164 15236
rect 6164 15180 6168 15236
rect 6104 15176 6168 15180
rect 6184 15236 6248 15240
rect 6184 15180 6188 15236
rect 6188 15180 6244 15236
rect 6244 15180 6248 15236
rect 6184 15176 6248 15180
rect 6264 15236 6328 15240
rect 6264 15180 6268 15236
rect 6268 15180 6324 15236
rect 6324 15180 6328 15236
rect 6264 15176 6328 15180
rect 7874 15236 7938 15240
rect 7874 15180 7878 15236
rect 7878 15180 7934 15236
rect 7934 15180 7938 15236
rect 7874 15176 7938 15180
rect 7954 15236 8018 15240
rect 7954 15180 7958 15236
rect 7958 15180 8014 15236
rect 8014 15180 8018 15236
rect 7954 15176 8018 15180
rect 8034 15236 8098 15240
rect 8034 15180 8038 15236
rect 8038 15180 8094 15236
rect 8094 15180 8098 15236
rect 8034 15176 8098 15180
rect 8114 15236 8178 15240
rect 8114 15180 8118 15236
rect 8118 15180 8174 15236
rect 8174 15180 8178 15236
rect 8114 15176 8178 15180
rect 8194 15236 8258 15240
rect 8194 15180 8198 15236
rect 8198 15180 8254 15236
rect 8254 15180 8258 15236
rect 8194 15176 8258 15180
rect 4978 14692 5042 14696
rect 4978 14636 4982 14692
rect 4982 14636 5038 14692
rect 5038 14636 5042 14692
rect 4978 14632 5042 14636
rect 5058 14692 5122 14696
rect 5058 14636 5062 14692
rect 5062 14636 5118 14692
rect 5118 14636 5122 14692
rect 5058 14632 5122 14636
rect 5138 14692 5202 14696
rect 5138 14636 5142 14692
rect 5142 14636 5198 14692
rect 5198 14636 5202 14692
rect 5138 14632 5202 14636
rect 5218 14692 5282 14696
rect 5218 14636 5222 14692
rect 5222 14636 5278 14692
rect 5278 14636 5282 14692
rect 5218 14632 5282 14636
rect 5298 14692 5362 14696
rect 5298 14636 5302 14692
rect 5302 14636 5358 14692
rect 5358 14636 5362 14692
rect 5298 14632 5362 14636
rect 6909 14692 6973 14696
rect 6909 14636 6913 14692
rect 6913 14636 6969 14692
rect 6969 14636 6973 14692
rect 6909 14632 6973 14636
rect 6989 14692 7053 14696
rect 6989 14636 6993 14692
rect 6993 14636 7049 14692
rect 7049 14636 7053 14692
rect 6989 14632 7053 14636
rect 7069 14692 7133 14696
rect 7069 14636 7073 14692
rect 7073 14636 7129 14692
rect 7129 14636 7133 14692
rect 7069 14632 7133 14636
rect 7149 14692 7213 14696
rect 7149 14636 7153 14692
rect 7153 14636 7209 14692
rect 7209 14636 7213 14692
rect 7149 14632 7213 14636
rect 7229 14692 7293 14696
rect 7229 14636 7233 14692
rect 7233 14636 7289 14692
rect 7289 14636 7293 14692
rect 7229 14632 7293 14636
rect 4013 14148 4077 14152
rect 4013 14092 4017 14148
rect 4017 14092 4073 14148
rect 4073 14092 4077 14148
rect 4013 14088 4077 14092
rect 4093 14148 4157 14152
rect 4093 14092 4097 14148
rect 4097 14092 4153 14148
rect 4153 14092 4157 14148
rect 4093 14088 4157 14092
rect 4173 14148 4237 14152
rect 4173 14092 4177 14148
rect 4177 14092 4233 14148
rect 4233 14092 4237 14148
rect 4173 14088 4237 14092
rect 4253 14148 4317 14152
rect 4253 14092 4257 14148
rect 4257 14092 4313 14148
rect 4313 14092 4317 14148
rect 4253 14088 4317 14092
rect 4333 14148 4397 14152
rect 4333 14092 4337 14148
rect 4337 14092 4393 14148
rect 4393 14092 4397 14148
rect 4333 14088 4397 14092
rect 5944 14148 6008 14152
rect 5944 14092 5948 14148
rect 5948 14092 6004 14148
rect 6004 14092 6008 14148
rect 5944 14088 6008 14092
rect 6024 14148 6088 14152
rect 6024 14092 6028 14148
rect 6028 14092 6084 14148
rect 6084 14092 6088 14148
rect 6024 14088 6088 14092
rect 6104 14148 6168 14152
rect 6104 14092 6108 14148
rect 6108 14092 6164 14148
rect 6164 14092 6168 14148
rect 6104 14088 6168 14092
rect 6184 14148 6248 14152
rect 6184 14092 6188 14148
rect 6188 14092 6244 14148
rect 6244 14092 6248 14148
rect 6184 14088 6248 14092
rect 6264 14148 6328 14152
rect 6264 14092 6268 14148
rect 6268 14092 6324 14148
rect 6324 14092 6328 14148
rect 6264 14088 6328 14092
rect 7874 14148 7938 14152
rect 7874 14092 7878 14148
rect 7878 14092 7934 14148
rect 7934 14092 7938 14148
rect 7874 14088 7938 14092
rect 7954 14148 8018 14152
rect 7954 14092 7958 14148
rect 7958 14092 8014 14148
rect 8014 14092 8018 14148
rect 7954 14088 8018 14092
rect 8034 14148 8098 14152
rect 8034 14092 8038 14148
rect 8038 14092 8094 14148
rect 8094 14092 8098 14148
rect 8034 14088 8098 14092
rect 8114 14148 8178 14152
rect 8114 14092 8118 14148
rect 8118 14092 8174 14148
rect 8174 14092 8178 14148
rect 8114 14088 8178 14092
rect 8194 14148 8258 14152
rect 8194 14092 8198 14148
rect 8198 14092 8254 14148
rect 8254 14092 8258 14148
rect 8194 14088 8258 14092
rect 4978 13604 5042 13608
rect 4978 13548 4982 13604
rect 4982 13548 5038 13604
rect 5038 13548 5042 13604
rect 4978 13544 5042 13548
rect 5058 13604 5122 13608
rect 5058 13548 5062 13604
rect 5062 13548 5118 13604
rect 5118 13548 5122 13604
rect 5058 13544 5122 13548
rect 5138 13604 5202 13608
rect 5138 13548 5142 13604
rect 5142 13548 5198 13604
rect 5198 13548 5202 13604
rect 5138 13544 5202 13548
rect 5218 13604 5282 13608
rect 5218 13548 5222 13604
rect 5222 13548 5278 13604
rect 5278 13548 5282 13604
rect 5218 13544 5282 13548
rect 5298 13604 5362 13608
rect 5298 13548 5302 13604
rect 5302 13548 5358 13604
rect 5358 13548 5362 13604
rect 5298 13544 5362 13548
rect 6909 13604 6973 13608
rect 6909 13548 6913 13604
rect 6913 13548 6969 13604
rect 6969 13548 6973 13604
rect 6909 13544 6973 13548
rect 6989 13604 7053 13608
rect 6989 13548 6993 13604
rect 6993 13548 7049 13604
rect 7049 13548 7053 13604
rect 6989 13544 7053 13548
rect 7069 13604 7133 13608
rect 7069 13548 7073 13604
rect 7073 13548 7129 13604
rect 7129 13548 7133 13604
rect 7069 13544 7133 13548
rect 7149 13604 7213 13608
rect 7149 13548 7153 13604
rect 7153 13548 7209 13604
rect 7209 13548 7213 13604
rect 7149 13544 7213 13548
rect 7229 13604 7293 13608
rect 7229 13548 7233 13604
rect 7233 13548 7289 13604
rect 7289 13548 7293 13604
rect 7229 13544 7293 13548
rect 4013 13060 4077 13064
rect 4013 13004 4017 13060
rect 4017 13004 4073 13060
rect 4073 13004 4077 13060
rect 4013 13000 4077 13004
rect 4093 13060 4157 13064
rect 4093 13004 4097 13060
rect 4097 13004 4153 13060
rect 4153 13004 4157 13060
rect 4093 13000 4157 13004
rect 4173 13060 4237 13064
rect 4173 13004 4177 13060
rect 4177 13004 4233 13060
rect 4233 13004 4237 13060
rect 4173 13000 4237 13004
rect 4253 13060 4317 13064
rect 4253 13004 4257 13060
rect 4257 13004 4313 13060
rect 4313 13004 4317 13060
rect 4253 13000 4317 13004
rect 4333 13060 4397 13064
rect 4333 13004 4337 13060
rect 4337 13004 4393 13060
rect 4393 13004 4397 13060
rect 4333 13000 4397 13004
rect 5944 13060 6008 13064
rect 5944 13004 5948 13060
rect 5948 13004 6004 13060
rect 6004 13004 6008 13060
rect 5944 13000 6008 13004
rect 6024 13060 6088 13064
rect 6024 13004 6028 13060
rect 6028 13004 6084 13060
rect 6084 13004 6088 13060
rect 6024 13000 6088 13004
rect 6104 13060 6168 13064
rect 6104 13004 6108 13060
rect 6108 13004 6164 13060
rect 6164 13004 6168 13060
rect 6104 13000 6168 13004
rect 6184 13060 6248 13064
rect 6184 13004 6188 13060
rect 6188 13004 6244 13060
rect 6244 13004 6248 13060
rect 6184 13000 6248 13004
rect 6264 13060 6328 13064
rect 6264 13004 6268 13060
rect 6268 13004 6324 13060
rect 6324 13004 6328 13060
rect 6264 13000 6328 13004
rect 7874 13060 7938 13064
rect 7874 13004 7878 13060
rect 7878 13004 7934 13060
rect 7934 13004 7938 13060
rect 7874 13000 7938 13004
rect 7954 13060 8018 13064
rect 7954 13004 7958 13060
rect 7958 13004 8014 13060
rect 8014 13004 8018 13060
rect 7954 13000 8018 13004
rect 8034 13060 8098 13064
rect 8034 13004 8038 13060
rect 8038 13004 8094 13060
rect 8094 13004 8098 13060
rect 8034 13000 8098 13004
rect 8114 13060 8178 13064
rect 8114 13004 8118 13060
rect 8118 13004 8174 13060
rect 8174 13004 8178 13060
rect 8114 13000 8178 13004
rect 8194 13060 8258 13064
rect 8194 13004 8198 13060
rect 8198 13004 8254 13060
rect 8254 13004 8258 13060
rect 8194 13000 8258 13004
rect 4978 12516 5042 12520
rect 4978 12460 4982 12516
rect 4982 12460 5038 12516
rect 5038 12460 5042 12516
rect 4978 12456 5042 12460
rect 5058 12516 5122 12520
rect 5058 12460 5062 12516
rect 5062 12460 5118 12516
rect 5118 12460 5122 12516
rect 5058 12456 5122 12460
rect 5138 12516 5202 12520
rect 5138 12460 5142 12516
rect 5142 12460 5198 12516
rect 5198 12460 5202 12516
rect 5138 12456 5202 12460
rect 5218 12516 5282 12520
rect 5218 12460 5222 12516
rect 5222 12460 5278 12516
rect 5278 12460 5282 12516
rect 5218 12456 5282 12460
rect 5298 12516 5362 12520
rect 5298 12460 5302 12516
rect 5302 12460 5358 12516
rect 5358 12460 5362 12516
rect 5298 12456 5362 12460
rect 6909 12516 6973 12520
rect 6909 12460 6913 12516
rect 6913 12460 6969 12516
rect 6969 12460 6973 12516
rect 6909 12456 6973 12460
rect 6989 12516 7053 12520
rect 6989 12460 6993 12516
rect 6993 12460 7049 12516
rect 7049 12460 7053 12516
rect 6989 12456 7053 12460
rect 7069 12516 7133 12520
rect 7069 12460 7073 12516
rect 7073 12460 7129 12516
rect 7129 12460 7133 12516
rect 7069 12456 7133 12460
rect 7149 12516 7213 12520
rect 7149 12460 7153 12516
rect 7153 12460 7209 12516
rect 7209 12460 7213 12516
rect 7149 12456 7213 12460
rect 7229 12516 7293 12520
rect 7229 12460 7233 12516
rect 7233 12460 7289 12516
rect 7289 12460 7293 12516
rect 7229 12456 7293 12460
rect 4013 11972 4077 11976
rect 4013 11916 4017 11972
rect 4017 11916 4073 11972
rect 4073 11916 4077 11972
rect 4013 11912 4077 11916
rect 4093 11972 4157 11976
rect 4093 11916 4097 11972
rect 4097 11916 4153 11972
rect 4153 11916 4157 11972
rect 4093 11912 4157 11916
rect 4173 11972 4237 11976
rect 4173 11916 4177 11972
rect 4177 11916 4233 11972
rect 4233 11916 4237 11972
rect 4173 11912 4237 11916
rect 4253 11972 4317 11976
rect 4253 11916 4257 11972
rect 4257 11916 4313 11972
rect 4313 11916 4317 11972
rect 4253 11912 4317 11916
rect 4333 11972 4397 11976
rect 4333 11916 4337 11972
rect 4337 11916 4393 11972
rect 4393 11916 4397 11972
rect 4333 11912 4397 11916
rect 5944 11972 6008 11976
rect 5944 11916 5948 11972
rect 5948 11916 6004 11972
rect 6004 11916 6008 11972
rect 5944 11912 6008 11916
rect 6024 11972 6088 11976
rect 6024 11916 6028 11972
rect 6028 11916 6084 11972
rect 6084 11916 6088 11972
rect 6024 11912 6088 11916
rect 6104 11972 6168 11976
rect 6104 11916 6108 11972
rect 6108 11916 6164 11972
rect 6164 11916 6168 11972
rect 6104 11912 6168 11916
rect 6184 11972 6248 11976
rect 6184 11916 6188 11972
rect 6188 11916 6244 11972
rect 6244 11916 6248 11972
rect 6184 11912 6248 11916
rect 6264 11972 6328 11976
rect 6264 11916 6268 11972
rect 6268 11916 6324 11972
rect 6324 11916 6328 11972
rect 6264 11912 6328 11916
rect 7874 11972 7938 11976
rect 7874 11916 7878 11972
rect 7878 11916 7934 11972
rect 7934 11916 7938 11972
rect 7874 11912 7938 11916
rect 7954 11972 8018 11976
rect 7954 11916 7958 11972
rect 7958 11916 8014 11972
rect 8014 11916 8018 11972
rect 7954 11912 8018 11916
rect 8034 11972 8098 11976
rect 8034 11916 8038 11972
rect 8038 11916 8094 11972
rect 8094 11916 8098 11972
rect 8034 11912 8098 11916
rect 8114 11972 8178 11976
rect 8114 11916 8118 11972
rect 8118 11916 8174 11972
rect 8174 11916 8178 11972
rect 8114 11912 8178 11916
rect 8194 11972 8258 11976
rect 8194 11916 8198 11972
rect 8198 11916 8254 11972
rect 8254 11916 8258 11972
rect 8194 11912 8258 11916
rect 4978 11428 5042 11432
rect 4978 11372 4982 11428
rect 4982 11372 5038 11428
rect 5038 11372 5042 11428
rect 4978 11368 5042 11372
rect 5058 11428 5122 11432
rect 5058 11372 5062 11428
rect 5062 11372 5118 11428
rect 5118 11372 5122 11428
rect 5058 11368 5122 11372
rect 5138 11428 5202 11432
rect 5138 11372 5142 11428
rect 5142 11372 5198 11428
rect 5198 11372 5202 11428
rect 5138 11368 5202 11372
rect 5218 11428 5282 11432
rect 5218 11372 5222 11428
rect 5222 11372 5278 11428
rect 5278 11372 5282 11428
rect 5218 11368 5282 11372
rect 5298 11428 5362 11432
rect 5298 11372 5302 11428
rect 5302 11372 5358 11428
rect 5358 11372 5362 11428
rect 5298 11368 5362 11372
rect 6909 11428 6973 11432
rect 6909 11372 6913 11428
rect 6913 11372 6969 11428
rect 6969 11372 6973 11428
rect 6909 11368 6973 11372
rect 6989 11428 7053 11432
rect 6989 11372 6993 11428
rect 6993 11372 7049 11428
rect 7049 11372 7053 11428
rect 6989 11368 7053 11372
rect 7069 11428 7133 11432
rect 7069 11372 7073 11428
rect 7073 11372 7129 11428
rect 7129 11372 7133 11428
rect 7069 11368 7133 11372
rect 7149 11428 7213 11432
rect 7149 11372 7153 11428
rect 7153 11372 7209 11428
rect 7209 11372 7213 11428
rect 7149 11368 7213 11372
rect 7229 11428 7293 11432
rect 7229 11372 7233 11428
rect 7233 11372 7289 11428
rect 7289 11372 7293 11428
rect 7229 11368 7293 11372
rect 4013 10884 4077 10888
rect 4013 10828 4017 10884
rect 4017 10828 4073 10884
rect 4073 10828 4077 10884
rect 4013 10824 4077 10828
rect 4093 10884 4157 10888
rect 4093 10828 4097 10884
rect 4097 10828 4153 10884
rect 4153 10828 4157 10884
rect 4093 10824 4157 10828
rect 4173 10884 4237 10888
rect 4173 10828 4177 10884
rect 4177 10828 4233 10884
rect 4233 10828 4237 10884
rect 4173 10824 4237 10828
rect 4253 10884 4317 10888
rect 4253 10828 4257 10884
rect 4257 10828 4313 10884
rect 4313 10828 4317 10884
rect 4253 10824 4317 10828
rect 4333 10884 4397 10888
rect 4333 10828 4337 10884
rect 4337 10828 4393 10884
rect 4393 10828 4397 10884
rect 4333 10824 4397 10828
rect 5944 10884 6008 10888
rect 5944 10828 5948 10884
rect 5948 10828 6004 10884
rect 6004 10828 6008 10884
rect 5944 10824 6008 10828
rect 6024 10884 6088 10888
rect 6024 10828 6028 10884
rect 6028 10828 6084 10884
rect 6084 10828 6088 10884
rect 6024 10824 6088 10828
rect 6104 10884 6168 10888
rect 6104 10828 6108 10884
rect 6108 10828 6164 10884
rect 6164 10828 6168 10884
rect 6104 10824 6168 10828
rect 6184 10884 6248 10888
rect 6184 10828 6188 10884
rect 6188 10828 6244 10884
rect 6244 10828 6248 10884
rect 6184 10824 6248 10828
rect 6264 10884 6328 10888
rect 6264 10828 6268 10884
rect 6268 10828 6324 10884
rect 6324 10828 6328 10884
rect 6264 10824 6328 10828
rect 7874 10884 7938 10888
rect 7874 10828 7878 10884
rect 7878 10828 7934 10884
rect 7934 10828 7938 10884
rect 7874 10824 7938 10828
rect 7954 10884 8018 10888
rect 7954 10828 7958 10884
rect 7958 10828 8014 10884
rect 8014 10828 8018 10884
rect 7954 10824 8018 10828
rect 8034 10884 8098 10888
rect 8034 10828 8038 10884
rect 8038 10828 8094 10884
rect 8094 10828 8098 10884
rect 8034 10824 8098 10828
rect 8114 10884 8178 10888
rect 8114 10828 8118 10884
rect 8118 10828 8174 10884
rect 8174 10828 8178 10884
rect 8114 10824 8178 10828
rect 8194 10884 8258 10888
rect 8194 10828 8198 10884
rect 8198 10828 8254 10884
rect 8254 10828 8258 10884
rect 8194 10824 8258 10828
rect 4978 10340 5042 10344
rect 4978 10284 4982 10340
rect 4982 10284 5038 10340
rect 5038 10284 5042 10340
rect 4978 10280 5042 10284
rect 5058 10340 5122 10344
rect 5058 10284 5062 10340
rect 5062 10284 5118 10340
rect 5118 10284 5122 10340
rect 5058 10280 5122 10284
rect 5138 10340 5202 10344
rect 5138 10284 5142 10340
rect 5142 10284 5198 10340
rect 5198 10284 5202 10340
rect 5138 10280 5202 10284
rect 5218 10340 5282 10344
rect 5218 10284 5222 10340
rect 5222 10284 5278 10340
rect 5278 10284 5282 10340
rect 5218 10280 5282 10284
rect 5298 10340 5362 10344
rect 5298 10284 5302 10340
rect 5302 10284 5358 10340
rect 5358 10284 5362 10340
rect 5298 10280 5362 10284
rect 6909 10340 6973 10344
rect 6909 10284 6913 10340
rect 6913 10284 6969 10340
rect 6969 10284 6973 10340
rect 6909 10280 6973 10284
rect 6989 10340 7053 10344
rect 6989 10284 6993 10340
rect 6993 10284 7049 10340
rect 7049 10284 7053 10340
rect 6989 10280 7053 10284
rect 7069 10340 7133 10344
rect 7069 10284 7073 10340
rect 7073 10284 7129 10340
rect 7129 10284 7133 10340
rect 7069 10280 7133 10284
rect 7149 10340 7213 10344
rect 7149 10284 7153 10340
rect 7153 10284 7209 10340
rect 7209 10284 7213 10340
rect 7149 10280 7213 10284
rect 7229 10340 7293 10344
rect 7229 10284 7233 10340
rect 7233 10284 7289 10340
rect 7289 10284 7293 10340
rect 7229 10280 7293 10284
rect 4013 9796 4077 9800
rect 4013 9740 4017 9796
rect 4017 9740 4073 9796
rect 4073 9740 4077 9796
rect 4013 9736 4077 9740
rect 4093 9796 4157 9800
rect 4093 9740 4097 9796
rect 4097 9740 4153 9796
rect 4153 9740 4157 9796
rect 4093 9736 4157 9740
rect 4173 9796 4237 9800
rect 4173 9740 4177 9796
rect 4177 9740 4233 9796
rect 4233 9740 4237 9796
rect 4173 9736 4237 9740
rect 4253 9796 4317 9800
rect 4253 9740 4257 9796
rect 4257 9740 4313 9796
rect 4313 9740 4317 9796
rect 4253 9736 4317 9740
rect 4333 9796 4397 9800
rect 4333 9740 4337 9796
rect 4337 9740 4393 9796
rect 4393 9740 4397 9796
rect 4333 9736 4397 9740
rect 5944 9796 6008 9800
rect 5944 9740 5948 9796
rect 5948 9740 6004 9796
rect 6004 9740 6008 9796
rect 5944 9736 6008 9740
rect 6024 9796 6088 9800
rect 6024 9740 6028 9796
rect 6028 9740 6084 9796
rect 6084 9740 6088 9796
rect 6024 9736 6088 9740
rect 6104 9796 6168 9800
rect 6104 9740 6108 9796
rect 6108 9740 6164 9796
rect 6164 9740 6168 9796
rect 6104 9736 6168 9740
rect 6184 9796 6248 9800
rect 6184 9740 6188 9796
rect 6188 9740 6244 9796
rect 6244 9740 6248 9796
rect 6184 9736 6248 9740
rect 6264 9796 6328 9800
rect 6264 9740 6268 9796
rect 6268 9740 6324 9796
rect 6324 9740 6328 9796
rect 6264 9736 6328 9740
rect 7874 9796 7938 9800
rect 7874 9740 7878 9796
rect 7878 9740 7934 9796
rect 7934 9740 7938 9796
rect 7874 9736 7938 9740
rect 7954 9796 8018 9800
rect 7954 9740 7958 9796
rect 7958 9740 8014 9796
rect 8014 9740 8018 9796
rect 7954 9736 8018 9740
rect 8034 9796 8098 9800
rect 8034 9740 8038 9796
rect 8038 9740 8094 9796
rect 8094 9740 8098 9796
rect 8034 9736 8098 9740
rect 8114 9796 8178 9800
rect 8114 9740 8118 9796
rect 8118 9740 8174 9796
rect 8174 9740 8178 9796
rect 8114 9736 8178 9740
rect 8194 9796 8258 9800
rect 8194 9740 8198 9796
rect 8198 9740 8254 9796
rect 8254 9740 8258 9796
rect 8194 9736 8258 9740
rect 4978 9252 5042 9256
rect 4978 9196 4982 9252
rect 4982 9196 5038 9252
rect 5038 9196 5042 9252
rect 4978 9192 5042 9196
rect 5058 9252 5122 9256
rect 5058 9196 5062 9252
rect 5062 9196 5118 9252
rect 5118 9196 5122 9252
rect 5058 9192 5122 9196
rect 5138 9252 5202 9256
rect 5138 9196 5142 9252
rect 5142 9196 5198 9252
rect 5198 9196 5202 9252
rect 5138 9192 5202 9196
rect 5218 9252 5282 9256
rect 5218 9196 5222 9252
rect 5222 9196 5278 9252
rect 5278 9196 5282 9252
rect 5218 9192 5282 9196
rect 5298 9252 5362 9256
rect 5298 9196 5302 9252
rect 5302 9196 5358 9252
rect 5358 9196 5362 9252
rect 5298 9192 5362 9196
rect 6909 9252 6973 9256
rect 6909 9196 6913 9252
rect 6913 9196 6969 9252
rect 6969 9196 6973 9252
rect 6909 9192 6973 9196
rect 6989 9252 7053 9256
rect 6989 9196 6993 9252
rect 6993 9196 7049 9252
rect 7049 9196 7053 9252
rect 6989 9192 7053 9196
rect 7069 9252 7133 9256
rect 7069 9196 7073 9252
rect 7073 9196 7129 9252
rect 7129 9196 7133 9252
rect 7069 9192 7133 9196
rect 7149 9252 7213 9256
rect 7149 9196 7153 9252
rect 7153 9196 7209 9252
rect 7209 9196 7213 9252
rect 7149 9192 7213 9196
rect 7229 9252 7293 9256
rect 7229 9196 7233 9252
rect 7233 9196 7289 9252
rect 7289 9196 7293 9252
rect 7229 9192 7293 9196
rect 4013 8708 4077 8712
rect 4013 8652 4017 8708
rect 4017 8652 4073 8708
rect 4073 8652 4077 8708
rect 4013 8648 4077 8652
rect 4093 8708 4157 8712
rect 4093 8652 4097 8708
rect 4097 8652 4153 8708
rect 4153 8652 4157 8708
rect 4093 8648 4157 8652
rect 4173 8708 4237 8712
rect 4173 8652 4177 8708
rect 4177 8652 4233 8708
rect 4233 8652 4237 8708
rect 4173 8648 4237 8652
rect 4253 8708 4317 8712
rect 4253 8652 4257 8708
rect 4257 8652 4313 8708
rect 4313 8652 4317 8708
rect 4253 8648 4317 8652
rect 4333 8708 4397 8712
rect 4333 8652 4337 8708
rect 4337 8652 4393 8708
rect 4393 8652 4397 8708
rect 4333 8648 4397 8652
rect 5944 8708 6008 8712
rect 5944 8652 5948 8708
rect 5948 8652 6004 8708
rect 6004 8652 6008 8708
rect 5944 8648 6008 8652
rect 6024 8708 6088 8712
rect 6024 8652 6028 8708
rect 6028 8652 6084 8708
rect 6084 8652 6088 8708
rect 6024 8648 6088 8652
rect 6104 8708 6168 8712
rect 6104 8652 6108 8708
rect 6108 8652 6164 8708
rect 6164 8652 6168 8708
rect 6104 8648 6168 8652
rect 6184 8708 6248 8712
rect 6184 8652 6188 8708
rect 6188 8652 6244 8708
rect 6244 8652 6248 8708
rect 6184 8648 6248 8652
rect 6264 8708 6328 8712
rect 6264 8652 6268 8708
rect 6268 8652 6324 8708
rect 6324 8652 6328 8708
rect 6264 8648 6328 8652
rect 7874 8708 7938 8712
rect 7874 8652 7878 8708
rect 7878 8652 7934 8708
rect 7934 8652 7938 8708
rect 7874 8648 7938 8652
rect 7954 8708 8018 8712
rect 7954 8652 7958 8708
rect 7958 8652 8014 8708
rect 8014 8652 8018 8708
rect 7954 8648 8018 8652
rect 8034 8708 8098 8712
rect 8034 8652 8038 8708
rect 8038 8652 8094 8708
rect 8094 8652 8098 8708
rect 8034 8648 8098 8652
rect 8114 8708 8178 8712
rect 8114 8652 8118 8708
rect 8118 8652 8174 8708
rect 8174 8652 8178 8708
rect 8114 8648 8178 8652
rect 8194 8708 8258 8712
rect 8194 8652 8198 8708
rect 8198 8652 8254 8708
rect 8254 8652 8258 8708
rect 8194 8648 8258 8652
rect 4978 8164 5042 8168
rect 4978 8108 4982 8164
rect 4982 8108 5038 8164
rect 5038 8108 5042 8164
rect 4978 8104 5042 8108
rect 5058 8164 5122 8168
rect 5058 8108 5062 8164
rect 5062 8108 5118 8164
rect 5118 8108 5122 8164
rect 5058 8104 5122 8108
rect 5138 8164 5202 8168
rect 5138 8108 5142 8164
rect 5142 8108 5198 8164
rect 5198 8108 5202 8164
rect 5138 8104 5202 8108
rect 5218 8164 5282 8168
rect 5218 8108 5222 8164
rect 5222 8108 5278 8164
rect 5278 8108 5282 8164
rect 5218 8104 5282 8108
rect 5298 8164 5362 8168
rect 5298 8108 5302 8164
rect 5302 8108 5358 8164
rect 5358 8108 5362 8164
rect 5298 8104 5362 8108
rect 6909 8164 6973 8168
rect 6909 8108 6913 8164
rect 6913 8108 6969 8164
rect 6969 8108 6973 8164
rect 6909 8104 6973 8108
rect 6989 8164 7053 8168
rect 6989 8108 6993 8164
rect 6993 8108 7049 8164
rect 7049 8108 7053 8164
rect 6989 8104 7053 8108
rect 7069 8164 7133 8168
rect 7069 8108 7073 8164
rect 7073 8108 7129 8164
rect 7129 8108 7133 8164
rect 7069 8104 7133 8108
rect 7149 8164 7213 8168
rect 7149 8108 7153 8164
rect 7153 8108 7209 8164
rect 7209 8108 7213 8164
rect 7149 8104 7213 8108
rect 7229 8164 7293 8168
rect 7229 8108 7233 8164
rect 7233 8108 7289 8164
rect 7289 8108 7293 8164
rect 7229 8104 7293 8108
rect 4013 7620 4077 7624
rect 4013 7564 4017 7620
rect 4017 7564 4073 7620
rect 4073 7564 4077 7620
rect 4013 7560 4077 7564
rect 4093 7620 4157 7624
rect 4093 7564 4097 7620
rect 4097 7564 4153 7620
rect 4153 7564 4157 7620
rect 4093 7560 4157 7564
rect 4173 7620 4237 7624
rect 4173 7564 4177 7620
rect 4177 7564 4233 7620
rect 4233 7564 4237 7620
rect 4173 7560 4237 7564
rect 4253 7620 4317 7624
rect 4253 7564 4257 7620
rect 4257 7564 4313 7620
rect 4313 7564 4317 7620
rect 4253 7560 4317 7564
rect 4333 7620 4397 7624
rect 4333 7564 4337 7620
rect 4337 7564 4393 7620
rect 4393 7564 4397 7620
rect 4333 7560 4397 7564
rect 5944 7620 6008 7624
rect 5944 7564 5948 7620
rect 5948 7564 6004 7620
rect 6004 7564 6008 7620
rect 5944 7560 6008 7564
rect 6024 7620 6088 7624
rect 6024 7564 6028 7620
rect 6028 7564 6084 7620
rect 6084 7564 6088 7620
rect 6024 7560 6088 7564
rect 6104 7620 6168 7624
rect 6104 7564 6108 7620
rect 6108 7564 6164 7620
rect 6164 7564 6168 7620
rect 6104 7560 6168 7564
rect 6184 7620 6248 7624
rect 6184 7564 6188 7620
rect 6188 7564 6244 7620
rect 6244 7564 6248 7620
rect 6184 7560 6248 7564
rect 6264 7620 6328 7624
rect 6264 7564 6268 7620
rect 6268 7564 6324 7620
rect 6324 7564 6328 7620
rect 6264 7560 6328 7564
rect 7874 7620 7938 7624
rect 7874 7564 7878 7620
rect 7878 7564 7934 7620
rect 7934 7564 7938 7620
rect 7874 7560 7938 7564
rect 7954 7620 8018 7624
rect 7954 7564 7958 7620
rect 7958 7564 8014 7620
rect 8014 7564 8018 7620
rect 7954 7560 8018 7564
rect 8034 7620 8098 7624
rect 8034 7564 8038 7620
rect 8038 7564 8094 7620
rect 8094 7564 8098 7620
rect 8034 7560 8098 7564
rect 8114 7620 8178 7624
rect 8114 7564 8118 7620
rect 8118 7564 8174 7620
rect 8174 7564 8178 7620
rect 8114 7560 8178 7564
rect 8194 7620 8258 7624
rect 8194 7564 8198 7620
rect 8198 7564 8254 7620
rect 8254 7564 8258 7620
rect 8194 7560 8258 7564
rect 4978 7076 5042 7080
rect 4978 7020 4982 7076
rect 4982 7020 5038 7076
rect 5038 7020 5042 7076
rect 4978 7016 5042 7020
rect 5058 7076 5122 7080
rect 5058 7020 5062 7076
rect 5062 7020 5118 7076
rect 5118 7020 5122 7076
rect 5058 7016 5122 7020
rect 5138 7076 5202 7080
rect 5138 7020 5142 7076
rect 5142 7020 5198 7076
rect 5198 7020 5202 7076
rect 5138 7016 5202 7020
rect 5218 7076 5282 7080
rect 5218 7020 5222 7076
rect 5222 7020 5278 7076
rect 5278 7020 5282 7076
rect 5218 7016 5282 7020
rect 5298 7076 5362 7080
rect 5298 7020 5302 7076
rect 5302 7020 5358 7076
rect 5358 7020 5362 7076
rect 5298 7016 5362 7020
rect 6909 7076 6973 7080
rect 6909 7020 6913 7076
rect 6913 7020 6969 7076
rect 6969 7020 6973 7076
rect 6909 7016 6973 7020
rect 6989 7076 7053 7080
rect 6989 7020 6993 7076
rect 6993 7020 7049 7076
rect 7049 7020 7053 7076
rect 6989 7016 7053 7020
rect 7069 7076 7133 7080
rect 7069 7020 7073 7076
rect 7073 7020 7129 7076
rect 7129 7020 7133 7076
rect 7069 7016 7133 7020
rect 7149 7076 7213 7080
rect 7149 7020 7153 7076
rect 7153 7020 7209 7076
rect 7209 7020 7213 7076
rect 7149 7016 7213 7020
rect 7229 7076 7293 7080
rect 7229 7020 7233 7076
rect 7233 7020 7289 7076
rect 7289 7020 7293 7076
rect 7229 7016 7293 7020
rect 4013 6532 4077 6536
rect 4013 6476 4017 6532
rect 4017 6476 4073 6532
rect 4073 6476 4077 6532
rect 4013 6472 4077 6476
rect 4093 6532 4157 6536
rect 4093 6476 4097 6532
rect 4097 6476 4153 6532
rect 4153 6476 4157 6532
rect 4093 6472 4157 6476
rect 4173 6532 4237 6536
rect 4173 6476 4177 6532
rect 4177 6476 4233 6532
rect 4233 6476 4237 6532
rect 4173 6472 4237 6476
rect 4253 6532 4317 6536
rect 4253 6476 4257 6532
rect 4257 6476 4313 6532
rect 4313 6476 4317 6532
rect 4253 6472 4317 6476
rect 4333 6532 4397 6536
rect 4333 6476 4337 6532
rect 4337 6476 4393 6532
rect 4393 6476 4397 6532
rect 4333 6472 4397 6476
rect 5944 6532 6008 6536
rect 5944 6476 5948 6532
rect 5948 6476 6004 6532
rect 6004 6476 6008 6532
rect 5944 6472 6008 6476
rect 6024 6532 6088 6536
rect 6024 6476 6028 6532
rect 6028 6476 6084 6532
rect 6084 6476 6088 6532
rect 6024 6472 6088 6476
rect 6104 6532 6168 6536
rect 6104 6476 6108 6532
rect 6108 6476 6164 6532
rect 6164 6476 6168 6532
rect 6104 6472 6168 6476
rect 6184 6532 6248 6536
rect 6184 6476 6188 6532
rect 6188 6476 6244 6532
rect 6244 6476 6248 6532
rect 6184 6472 6248 6476
rect 6264 6532 6328 6536
rect 6264 6476 6268 6532
rect 6268 6476 6324 6532
rect 6324 6476 6328 6532
rect 6264 6472 6328 6476
rect 7874 6532 7938 6536
rect 7874 6476 7878 6532
rect 7878 6476 7934 6532
rect 7934 6476 7938 6532
rect 7874 6472 7938 6476
rect 7954 6532 8018 6536
rect 7954 6476 7958 6532
rect 7958 6476 8014 6532
rect 8014 6476 8018 6532
rect 7954 6472 8018 6476
rect 8034 6532 8098 6536
rect 8034 6476 8038 6532
rect 8038 6476 8094 6532
rect 8094 6476 8098 6532
rect 8034 6472 8098 6476
rect 8114 6532 8178 6536
rect 8114 6476 8118 6532
rect 8118 6476 8174 6532
rect 8174 6476 8178 6532
rect 8114 6472 8178 6476
rect 8194 6532 8258 6536
rect 8194 6476 8198 6532
rect 8198 6476 8254 6532
rect 8254 6476 8258 6532
rect 8194 6472 8258 6476
rect 4978 5988 5042 5992
rect 4978 5932 4982 5988
rect 4982 5932 5038 5988
rect 5038 5932 5042 5988
rect 4978 5928 5042 5932
rect 5058 5988 5122 5992
rect 5058 5932 5062 5988
rect 5062 5932 5118 5988
rect 5118 5932 5122 5988
rect 5058 5928 5122 5932
rect 5138 5988 5202 5992
rect 5138 5932 5142 5988
rect 5142 5932 5198 5988
rect 5198 5932 5202 5988
rect 5138 5928 5202 5932
rect 5218 5988 5282 5992
rect 5218 5932 5222 5988
rect 5222 5932 5278 5988
rect 5278 5932 5282 5988
rect 5218 5928 5282 5932
rect 5298 5988 5362 5992
rect 5298 5932 5302 5988
rect 5302 5932 5358 5988
rect 5358 5932 5362 5988
rect 5298 5928 5362 5932
rect 6909 5988 6973 5992
rect 6909 5932 6913 5988
rect 6913 5932 6969 5988
rect 6969 5932 6973 5988
rect 6909 5928 6973 5932
rect 6989 5988 7053 5992
rect 6989 5932 6993 5988
rect 6993 5932 7049 5988
rect 7049 5932 7053 5988
rect 6989 5928 7053 5932
rect 7069 5988 7133 5992
rect 7069 5932 7073 5988
rect 7073 5932 7129 5988
rect 7129 5932 7133 5988
rect 7069 5928 7133 5932
rect 7149 5988 7213 5992
rect 7149 5932 7153 5988
rect 7153 5932 7209 5988
rect 7209 5932 7213 5988
rect 7149 5928 7213 5932
rect 7229 5988 7293 5992
rect 7229 5932 7233 5988
rect 7233 5932 7289 5988
rect 7289 5932 7293 5988
rect 7229 5928 7293 5932
rect 4013 5444 4077 5448
rect 4013 5388 4017 5444
rect 4017 5388 4073 5444
rect 4073 5388 4077 5444
rect 4013 5384 4077 5388
rect 4093 5444 4157 5448
rect 4093 5388 4097 5444
rect 4097 5388 4153 5444
rect 4153 5388 4157 5444
rect 4093 5384 4157 5388
rect 4173 5444 4237 5448
rect 4173 5388 4177 5444
rect 4177 5388 4233 5444
rect 4233 5388 4237 5444
rect 4173 5384 4237 5388
rect 4253 5444 4317 5448
rect 4253 5388 4257 5444
rect 4257 5388 4313 5444
rect 4313 5388 4317 5444
rect 4253 5384 4317 5388
rect 4333 5444 4397 5448
rect 4333 5388 4337 5444
rect 4337 5388 4393 5444
rect 4393 5388 4397 5444
rect 4333 5384 4397 5388
rect 5944 5444 6008 5448
rect 5944 5388 5948 5444
rect 5948 5388 6004 5444
rect 6004 5388 6008 5444
rect 5944 5384 6008 5388
rect 6024 5444 6088 5448
rect 6024 5388 6028 5444
rect 6028 5388 6084 5444
rect 6084 5388 6088 5444
rect 6024 5384 6088 5388
rect 6104 5444 6168 5448
rect 6104 5388 6108 5444
rect 6108 5388 6164 5444
rect 6164 5388 6168 5444
rect 6104 5384 6168 5388
rect 6184 5444 6248 5448
rect 6184 5388 6188 5444
rect 6188 5388 6244 5444
rect 6244 5388 6248 5444
rect 6184 5384 6248 5388
rect 6264 5444 6328 5448
rect 6264 5388 6268 5444
rect 6268 5388 6324 5444
rect 6324 5388 6328 5444
rect 6264 5384 6328 5388
rect 7874 5444 7938 5448
rect 7874 5388 7878 5444
rect 7878 5388 7934 5444
rect 7934 5388 7938 5444
rect 7874 5384 7938 5388
rect 7954 5444 8018 5448
rect 7954 5388 7958 5444
rect 7958 5388 8014 5444
rect 8014 5388 8018 5444
rect 7954 5384 8018 5388
rect 8034 5444 8098 5448
rect 8034 5388 8038 5444
rect 8038 5388 8094 5444
rect 8094 5388 8098 5444
rect 8034 5384 8098 5388
rect 8114 5444 8178 5448
rect 8114 5388 8118 5444
rect 8118 5388 8174 5444
rect 8174 5388 8178 5444
rect 8114 5384 8178 5388
rect 8194 5444 8258 5448
rect 8194 5388 8198 5444
rect 8198 5388 8254 5444
rect 8254 5388 8258 5444
rect 8194 5384 8258 5388
rect 4978 4900 5042 4904
rect 4978 4844 4982 4900
rect 4982 4844 5038 4900
rect 5038 4844 5042 4900
rect 4978 4840 5042 4844
rect 5058 4900 5122 4904
rect 5058 4844 5062 4900
rect 5062 4844 5118 4900
rect 5118 4844 5122 4900
rect 5058 4840 5122 4844
rect 5138 4900 5202 4904
rect 5138 4844 5142 4900
rect 5142 4844 5198 4900
rect 5198 4844 5202 4900
rect 5138 4840 5202 4844
rect 5218 4900 5282 4904
rect 5218 4844 5222 4900
rect 5222 4844 5278 4900
rect 5278 4844 5282 4900
rect 5218 4840 5282 4844
rect 5298 4900 5362 4904
rect 5298 4844 5302 4900
rect 5302 4844 5358 4900
rect 5358 4844 5362 4900
rect 5298 4840 5362 4844
rect 6909 4900 6973 4904
rect 6909 4844 6913 4900
rect 6913 4844 6969 4900
rect 6969 4844 6973 4900
rect 6909 4840 6973 4844
rect 6989 4900 7053 4904
rect 6989 4844 6993 4900
rect 6993 4844 7049 4900
rect 7049 4844 7053 4900
rect 6989 4840 7053 4844
rect 7069 4900 7133 4904
rect 7069 4844 7073 4900
rect 7073 4844 7129 4900
rect 7129 4844 7133 4900
rect 7069 4840 7133 4844
rect 7149 4900 7213 4904
rect 7149 4844 7153 4900
rect 7153 4844 7209 4900
rect 7209 4844 7213 4900
rect 7149 4840 7213 4844
rect 7229 4900 7293 4904
rect 7229 4844 7233 4900
rect 7233 4844 7289 4900
rect 7289 4844 7293 4900
rect 7229 4840 7293 4844
rect 4013 4356 4077 4360
rect 4013 4300 4017 4356
rect 4017 4300 4073 4356
rect 4073 4300 4077 4356
rect 4013 4296 4077 4300
rect 4093 4356 4157 4360
rect 4093 4300 4097 4356
rect 4097 4300 4153 4356
rect 4153 4300 4157 4356
rect 4093 4296 4157 4300
rect 4173 4356 4237 4360
rect 4173 4300 4177 4356
rect 4177 4300 4233 4356
rect 4233 4300 4237 4356
rect 4173 4296 4237 4300
rect 4253 4356 4317 4360
rect 4253 4300 4257 4356
rect 4257 4300 4313 4356
rect 4313 4300 4317 4356
rect 4253 4296 4317 4300
rect 4333 4356 4397 4360
rect 4333 4300 4337 4356
rect 4337 4300 4393 4356
rect 4393 4300 4397 4356
rect 4333 4296 4397 4300
rect 5944 4356 6008 4360
rect 5944 4300 5948 4356
rect 5948 4300 6004 4356
rect 6004 4300 6008 4356
rect 5944 4296 6008 4300
rect 6024 4356 6088 4360
rect 6024 4300 6028 4356
rect 6028 4300 6084 4356
rect 6084 4300 6088 4356
rect 6024 4296 6088 4300
rect 6104 4356 6168 4360
rect 6104 4300 6108 4356
rect 6108 4300 6164 4356
rect 6164 4300 6168 4356
rect 6104 4296 6168 4300
rect 6184 4356 6248 4360
rect 6184 4300 6188 4356
rect 6188 4300 6244 4356
rect 6244 4300 6248 4356
rect 6184 4296 6248 4300
rect 6264 4356 6328 4360
rect 6264 4300 6268 4356
rect 6268 4300 6324 4356
rect 6324 4300 6328 4356
rect 6264 4296 6328 4300
rect 7874 4356 7938 4360
rect 7874 4300 7878 4356
rect 7878 4300 7934 4356
rect 7934 4300 7938 4356
rect 7874 4296 7938 4300
rect 7954 4356 8018 4360
rect 7954 4300 7958 4356
rect 7958 4300 8014 4356
rect 8014 4300 8018 4356
rect 7954 4296 8018 4300
rect 8034 4356 8098 4360
rect 8034 4300 8038 4356
rect 8038 4300 8094 4356
rect 8094 4300 8098 4356
rect 8034 4296 8098 4300
rect 8114 4356 8178 4360
rect 8114 4300 8118 4356
rect 8118 4300 8174 4356
rect 8174 4300 8178 4356
rect 8114 4296 8178 4300
rect 8194 4356 8258 4360
rect 8194 4300 8198 4356
rect 8198 4300 8254 4356
rect 8254 4300 8258 4356
rect 8194 4296 8258 4300
rect 4978 3812 5042 3816
rect 4978 3756 4982 3812
rect 4982 3756 5038 3812
rect 5038 3756 5042 3812
rect 4978 3752 5042 3756
rect 5058 3812 5122 3816
rect 5058 3756 5062 3812
rect 5062 3756 5118 3812
rect 5118 3756 5122 3812
rect 5058 3752 5122 3756
rect 5138 3812 5202 3816
rect 5138 3756 5142 3812
rect 5142 3756 5198 3812
rect 5198 3756 5202 3812
rect 5138 3752 5202 3756
rect 5218 3812 5282 3816
rect 5218 3756 5222 3812
rect 5222 3756 5278 3812
rect 5278 3756 5282 3812
rect 5218 3752 5282 3756
rect 5298 3812 5362 3816
rect 5298 3756 5302 3812
rect 5302 3756 5358 3812
rect 5358 3756 5362 3812
rect 5298 3752 5362 3756
rect 6909 3812 6973 3816
rect 6909 3756 6913 3812
rect 6913 3756 6969 3812
rect 6969 3756 6973 3812
rect 6909 3752 6973 3756
rect 6989 3812 7053 3816
rect 6989 3756 6993 3812
rect 6993 3756 7049 3812
rect 7049 3756 7053 3812
rect 6989 3752 7053 3756
rect 7069 3812 7133 3816
rect 7069 3756 7073 3812
rect 7073 3756 7129 3812
rect 7129 3756 7133 3812
rect 7069 3752 7133 3756
rect 7149 3812 7213 3816
rect 7149 3756 7153 3812
rect 7153 3756 7209 3812
rect 7209 3756 7213 3812
rect 7149 3752 7213 3756
rect 7229 3812 7293 3816
rect 7229 3756 7233 3812
rect 7233 3756 7289 3812
rect 7289 3756 7293 3812
rect 7229 3752 7293 3756
rect 4013 3268 4077 3272
rect 4013 3212 4017 3268
rect 4017 3212 4073 3268
rect 4073 3212 4077 3268
rect 4013 3208 4077 3212
rect 4093 3268 4157 3272
rect 4093 3212 4097 3268
rect 4097 3212 4153 3268
rect 4153 3212 4157 3268
rect 4093 3208 4157 3212
rect 4173 3268 4237 3272
rect 4173 3212 4177 3268
rect 4177 3212 4233 3268
rect 4233 3212 4237 3268
rect 4173 3208 4237 3212
rect 4253 3268 4317 3272
rect 4253 3212 4257 3268
rect 4257 3212 4313 3268
rect 4313 3212 4317 3268
rect 4253 3208 4317 3212
rect 4333 3268 4397 3272
rect 4333 3212 4337 3268
rect 4337 3212 4393 3268
rect 4393 3212 4397 3268
rect 4333 3208 4397 3212
rect 5944 3268 6008 3272
rect 5944 3212 5948 3268
rect 5948 3212 6004 3268
rect 6004 3212 6008 3268
rect 5944 3208 6008 3212
rect 6024 3268 6088 3272
rect 6024 3212 6028 3268
rect 6028 3212 6084 3268
rect 6084 3212 6088 3268
rect 6024 3208 6088 3212
rect 6104 3268 6168 3272
rect 6104 3212 6108 3268
rect 6108 3212 6164 3268
rect 6164 3212 6168 3268
rect 6104 3208 6168 3212
rect 6184 3268 6248 3272
rect 6184 3212 6188 3268
rect 6188 3212 6244 3268
rect 6244 3212 6248 3268
rect 6184 3208 6248 3212
rect 6264 3268 6328 3272
rect 6264 3212 6268 3268
rect 6268 3212 6324 3268
rect 6324 3212 6328 3268
rect 6264 3208 6328 3212
rect 7874 3268 7938 3272
rect 7874 3212 7878 3268
rect 7878 3212 7934 3268
rect 7934 3212 7938 3268
rect 7874 3208 7938 3212
rect 7954 3268 8018 3272
rect 7954 3212 7958 3268
rect 7958 3212 8014 3268
rect 8014 3212 8018 3268
rect 7954 3208 8018 3212
rect 8034 3268 8098 3272
rect 8034 3212 8038 3268
rect 8038 3212 8094 3268
rect 8094 3212 8098 3268
rect 8034 3208 8098 3212
rect 8114 3268 8178 3272
rect 8114 3212 8118 3268
rect 8118 3212 8174 3268
rect 8174 3212 8178 3268
rect 8114 3208 8178 3212
rect 8194 3268 8258 3272
rect 8194 3212 8198 3268
rect 8198 3212 8254 3268
rect 8254 3212 8258 3268
rect 8194 3208 8258 3212
rect 1148 1868 1212 1932
rect 1228 1868 1292 1932
rect 1308 1868 1372 1932
rect 1388 1868 1452 1932
rect 1468 1868 1532 1932
rect 1548 1868 1612 1932
rect 1628 1868 1692 1932
rect 1708 1868 1772 1932
rect 1788 1868 1852 1932
rect 1868 1868 1932 1932
rect 4013 1868 4077 1932
rect 4093 1868 4157 1932
rect 4173 1868 4237 1932
rect 4253 1868 4317 1932
rect 4333 1868 4397 1932
rect 5944 1868 6008 1932
rect 6024 1868 6088 1932
rect 6104 1868 6168 1932
rect 6184 1868 6248 1932
rect 6264 1868 6328 1932
rect 7874 1868 7938 1932
rect 7954 1868 8018 1932
rect 8034 1868 8098 1932
rect 8114 1868 8178 1932
rect 8194 1868 8258 1932
rect 10252 1868 10316 1932
rect 10332 1868 10396 1932
rect 10412 1868 10476 1932
rect 10492 1868 10556 1932
rect 10572 1868 10636 1932
rect 10652 1868 10716 1932
rect 10732 1868 10796 1932
rect 10812 1868 10876 1932
rect 10892 1868 10956 1932
rect 10972 1868 11036 1932
rect 1148 1788 1212 1852
rect 1228 1788 1292 1852
rect 1308 1788 1372 1852
rect 1388 1788 1452 1852
rect 1468 1788 1532 1852
rect 1548 1788 1612 1852
rect 1628 1788 1692 1852
rect 1708 1788 1772 1852
rect 1788 1788 1852 1852
rect 1868 1788 1932 1852
rect 4013 1788 4077 1852
rect 4093 1788 4157 1852
rect 4173 1788 4237 1852
rect 4253 1788 4317 1852
rect 4333 1788 4397 1852
rect 5944 1788 6008 1852
rect 6024 1788 6088 1852
rect 6104 1788 6168 1852
rect 6184 1788 6248 1852
rect 6264 1788 6328 1852
rect 7874 1788 7938 1852
rect 7954 1788 8018 1852
rect 8034 1788 8098 1852
rect 8114 1788 8178 1852
rect 8194 1788 8258 1852
rect 10252 1788 10316 1852
rect 10332 1788 10396 1852
rect 10412 1788 10476 1852
rect 10492 1788 10556 1852
rect 10572 1788 10636 1852
rect 10652 1788 10716 1852
rect 10732 1788 10796 1852
rect 10812 1788 10876 1852
rect 10892 1788 10956 1852
rect 10972 1788 11036 1852
rect 1148 1708 1212 1772
rect 1228 1708 1292 1772
rect 1308 1708 1372 1772
rect 1388 1708 1452 1772
rect 1468 1708 1532 1772
rect 1548 1708 1612 1772
rect 1628 1708 1692 1772
rect 1708 1708 1772 1772
rect 1788 1708 1852 1772
rect 1868 1708 1932 1772
rect 4013 1708 4077 1772
rect 4093 1708 4157 1772
rect 4173 1708 4237 1772
rect 4253 1708 4317 1772
rect 4333 1708 4397 1772
rect 5944 1708 6008 1772
rect 6024 1708 6088 1772
rect 6104 1708 6168 1772
rect 6184 1708 6248 1772
rect 6264 1708 6328 1772
rect 7874 1708 7938 1772
rect 7954 1708 8018 1772
rect 8034 1708 8098 1772
rect 8114 1708 8178 1772
rect 8194 1708 8258 1772
rect 10252 1708 10316 1772
rect 10332 1708 10396 1772
rect 10412 1708 10476 1772
rect 10492 1708 10556 1772
rect 10572 1708 10636 1772
rect 10652 1708 10716 1772
rect 10732 1708 10796 1772
rect 10812 1708 10876 1772
rect 10892 1708 10956 1772
rect 10972 1708 11036 1772
rect 1148 1628 1212 1692
rect 1228 1628 1292 1692
rect 1308 1628 1372 1692
rect 1388 1628 1452 1692
rect 1468 1628 1532 1692
rect 1548 1628 1612 1692
rect 1628 1628 1692 1692
rect 1708 1628 1772 1692
rect 1788 1628 1852 1692
rect 1868 1628 1932 1692
rect 4013 1628 4077 1692
rect 4093 1628 4157 1692
rect 4173 1628 4237 1692
rect 4253 1628 4317 1692
rect 4333 1628 4397 1692
rect 5944 1628 6008 1692
rect 6024 1628 6088 1692
rect 6104 1628 6168 1692
rect 6184 1628 6248 1692
rect 6264 1628 6328 1692
rect 7874 1628 7938 1692
rect 7954 1628 8018 1692
rect 8034 1628 8098 1692
rect 8114 1628 8178 1692
rect 8194 1628 8258 1692
rect 10252 1628 10316 1692
rect 10332 1628 10396 1692
rect 10412 1628 10476 1692
rect 10492 1628 10556 1692
rect 10572 1628 10636 1692
rect 10652 1628 10716 1692
rect 10732 1628 10796 1692
rect 10812 1628 10876 1692
rect 10892 1628 10956 1692
rect 10972 1628 11036 1692
rect 1148 1548 1212 1612
rect 1228 1548 1292 1612
rect 1308 1548 1372 1612
rect 1388 1548 1452 1612
rect 1468 1548 1532 1612
rect 1548 1548 1612 1612
rect 1628 1548 1692 1612
rect 1708 1548 1772 1612
rect 1788 1548 1852 1612
rect 1868 1548 1932 1612
rect 4013 1548 4077 1612
rect 4093 1548 4157 1612
rect 4173 1548 4237 1612
rect 4253 1548 4317 1612
rect 4333 1548 4397 1612
rect 5944 1548 6008 1612
rect 6024 1548 6088 1612
rect 6104 1548 6168 1612
rect 6184 1548 6248 1612
rect 6264 1548 6328 1612
rect 7874 1548 7938 1612
rect 7954 1548 8018 1612
rect 8034 1548 8098 1612
rect 8114 1548 8178 1612
rect 8194 1548 8258 1612
rect 10252 1548 10316 1612
rect 10332 1548 10396 1612
rect 10412 1548 10476 1612
rect 10492 1548 10556 1612
rect 10572 1548 10636 1612
rect 10652 1548 10716 1612
rect 10732 1548 10796 1612
rect 10812 1548 10876 1612
rect 10892 1548 10956 1612
rect 10972 1548 11036 1612
rect 1148 1468 1212 1532
rect 1228 1468 1292 1532
rect 1308 1468 1372 1532
rect 1388 1468 1452 1532
rect 1468 1468 1532 1532
rect 1548 1468 1612 1532
rect 1628 1468 1692 1532
rect 1708 1468 1772 1532
rect 1788 1468 1852 1532
rect 1868 1468 1932 1532
rect 4013 1468 4077 1532
rect 4093 1468 4157 1532
rect 4173 1468 4237 1532
rect 4253 1468 4317 1532
rect 4333 1468 4397 1532
rect 5944 1468 6008 1532
rect 6024 1468 6088 1532
rect 6104 1468 6168 1532
rect 6184 1468 6248 1532
rect 6264 1468 6328 1532
rect 7874 1468 7938 1532
rect 7954 1468 8018 1532
rect 8034 1468 8098 1532
rect 8114 1468 8178 1532
rect 8194 1468 8258 1532
rect 10252 1468 10316 1532
rect 10332 1468 10396 1532
rect 10412 1468 10476 1532
rect 10492 1468 10556 1532
rect 10572 1468 10636 1532
rect 10652 1468 10716 1532
rect 10732 1468 10796 1532
rect 10812 1468 10876 1532
rect 10892 1468 10956 1532
rect 10972 1468 11036 1532
rect 1148 1388 1212 1452
rect 1228 1388 1292 1452
rect 1308 1388 1372 1452
rect 1388 1388 1452 1452
rect 1468 1388 1532 1452
rect 1548 1388 1612 1452
rect 1628 1388 1692 1452
rect 1708 1388 1772 1452
rect 1788 1388 1852 1452
rect 1868 1388 1932 1452
rect 4013 1388 4077 1452
rect 4093 1388 4157 1452
rect 4173 1388 4237 1452
rect 4253 1388 4317 1452
rect 4333 1388 4397 1452
rect 5944 1388 6008 1452
rect 6024 1388 6088 1452
rect 6104 1388 6168 1452
rect 6184 1388 6248 1452
rect 6264 1388 6328 1452
rect 7874 1388 7938 1452
rect 7954 1388 8018 1452
rect 8034 1388 8098 1452
rect 8114 1388 8178 1452
rect 8194 1388 8258 1452
rect 10252 1388 10316 1452
rect 10332 1388 10396 1452
rect 10412 1388 10476 1452
rect 10492 1388 10556 1452
rect 10572 1388 10636 1452
rect 10652 1388 10716 1452
rect 10732 1388 10796 1452
rect 10812 1388 10876 1452
rect 10892 1388 10956 1452
rect 10972 1388 11036 1452
rect 1148 1308 1212 1372
rect 1228 1308 1292 1372
rect 1308 1308 1372 1372
rect 1388 1308 1452 1372
rect 1468 1308 1532 1372
rect 1548 1308 1612 1372
rect 1628 1308 1692 1372
rect 1708 1308 1772 1372
rect 1788 1308 1852 1372
rect 1868 1308 1932 1372
rect 4013 1308 4077 1372
rect 4093 1308 4157 1372
rect 4173 1308 4237 1372
rect 4253 1308 4317 1372
rect 4333 1308 4397 1372
rect 5944 1308 6008 1372
rect 6024 1308 6088 1372
rect 6104 1308 6168 1372
rect 6184 1308 6248 1372
rect 6264 1308 6328 1372
rect 7874 1308 7938 1372
rect 7954 1308 8018 1372
rect 8034 1308 8098 1372
rect 8114 1308 8178 1372
rect 8194 1308 8258 1372
rect 10252 1308 10316 1372
rect 10332 1308 10396 1372
rect 10412 1308 10476 1372
rect 10492 1308 10556 1372
rect 10572 1308 10636 1372
rect 10652 1308 10716 1372
rect 10732 1308 10796 1372
rect 10812 1308 10876 1372
rect 10892 1308 10956 1372
rect 10972 1308 11036 1372
rect 1148 1228 1212 1292
rect 1228 1228 1292 1292
rect 1308 1228 1372 1292
rect 1388 1228 1452 1292
rect 1468 1228 1532 1292
rect 1548 1228 1612 1292
rect 1628 1228 1692 1292
rect 1708 1228 1772 1292
rect 1788 1228 1852 1292
rect 1868 1228 1932 1292
rect 4013 1228 4077 1292
rect 4093 1228 4157 1292
rect 4173 1228 4237 1292
rect 4253 1228 4317 1292
rect 4333 1228 4397 1292
rect 5944 1228 6008 1292
rect 6024 1228 6088 1292
rect 6104 1228 6168 1292
rect 6184 1228 6248 1292
rect 6264 1228 6328 1292
rect 7874 1228 7938 1292
rect 7954 1228 8018 1292
rect 8034 1228 8098 1292
rect 8114 1228 8178 1292
rect 8194 1228 8258 1292
rect 10252 1228 10316 1292
rect 10332 1228 10396 1292
rect 10412 1228 10476 1292
rect 10492 1228 10556 1292
rect 10572 1228 10636 1292
rect 10652 1228 10716 1292
rect 10732 1228 10796 1292
rect 10812 1228 10876 1292
rect 10892 1228 10956 1292
rect 10972 1228 11036 1292
rect 1148 1148 1212 1212
rect 1228 1148 1292 1212
rect 1308 1148 1372 1212
rect 1388 1148 1452 1212
rect 1468 1148 1532 1212
rect 1548 1148 1612 1212
rect 1628 1148 1692 1212
rect 1708 1148 1772 1212
rect 1788 1148 1852 1212
rect 1868 1148 1932 1212
rect 4013 1148 4077 1212
rect 4093 1148 4157 1212
rect 4173 1148 4237 1212
rect 4253 1148 4317 1212
rect 4333 1148 4397 1212
rect 5944 1148 6008 1212
rect 6024 1148 6088 1212
rect 6104 1148 6168 1212
rect 6184 1148 6248 1212
rect 6264 1148 6328 1212
rect 7874 1148 7938 1212
rect 7954 1148 8018 1212
rect 8034 1148 8098 1212
rect 8114 1148 8178 1212
rect 8194 1148 8258 1212
rect 10252 1148 10316 1212
rect 10332 1148 10396 1212
rect 10412 1148 10476 1212
rect 10492 1148 10556 1212
rect 10572 1148 10636 1212
rect 10652 1148 10716 1212
rect 10732 1148 10796 1212
rect 10812 1148 10876 1212
rect 10892 1148 10956 1212
rect 10972 1148 11036 1212
rect 8 728 72 792
rect 88 728 152 792
rect 168 728 232 792
rect 248 728 312 792
rect 328 728 392 792
rect 408 728 472 792
rect 488 728 552 792
rect 568 728 632 792
rect 648 728 712 792
rect 728 728 792 792
rect 4978 728 5042 792
rect 5058 728 5122 792
rect 5138 728 5202 792
rect 5218 728 5282 792
rect 5298 728 5362 792
rect 6909 728 6973 792
rect 6989 728 7053 792
rect 7069 728 7133 792
rect 7149 728 7213 792
rect 7229 728 7293 792
rect 11392 728 11456 792
rect 11472 728 11536 792
rect 11552 728 11616 792
rect 11632 728 11696 792
rect 11712 728 11776 792
rect 11792 728 11856 792
rect 11872 728 11936 792
rect 11952 728 12016 792
rect 12032 728 12096 792
rect 12112 728 12176 792
rect 8 648 72 712
rect 88 648 152 712
rect 168 648 232 712
rect 248 648 312 712
rect 328 648 392 712
rect 408 648 472 712
rect 488 648 552 712
rect 568 648 632 712
rect 648 648 712 712
rect 728 648 792 712
rect 4978 648 5042 712
rect 5058 648 5122 712
rect 5138 648 5202 712
rect 5218 648 5282 712
rect 5298 648 5362 712
rect 6909 648 6973 712
rect 6989 648 7053 712
rect 7069 648 7133 712
rect 7149 648 7213 712
rect 7229 648 7293 712
rect 11392 648 11456 712
rect 11472 648 11536 712
rect 11552 648 11616 712
rect 11632 648 11696 712
rect 11712 648 11776 712
rect 11792 648 11856 712
rect 11872 648 11936 712
rect 11952 648 12016 712
rect 12032 648 12096 712
rect 12112 648 12176 712
rect 8 568 72 632
rect 88 568 152 632
rect 168 568 232 632
rect 248 568 312 632
rect 328 568 392 632
rect 408 568 472 632
rect 488 568 552 632
rect 568 568 632 632
rect 648 568 712 632
rect 728 568 792 632
rect 4978 568 5042 632
rect 5058 568 5122 632
rect 5138 568 5202 632
rect 5218 568 5282 632
rect 5298 568 5362 632
rect 6909 568 6973 632
rect 6989 568 7053 632
rect 7069 568 7133 632
rect 7149 568 7213 632
rect 7229 568 7293 632
rect 11392 568 11456 632
rect 11472 568 11536 632
rect 11552 568 11616 632
rect 11632 568 11696 632
rect 11712 568 11776 632
rect 11792 568 11856 632
rect 11872 568 11936 632
rect 11952 568 12016 632
rect 12032 568 12096 632
rect 12112 568 12176 632
rect 8 488 72 552
rect 88 488 152 552
rect 168 488 232 552
rect 248 488 312 552
rect 328 488 392 552
rect 408 488 472 552
rect 488 488 552 552
rect 568 488 632 552
rect 648 488 712 552
rect 728 488 792 552
rect 4978 488 5042 552
rect 5058 488 5122 552
rect 5138 488 5202 552
rect 5218 488 5282 552
rect 5298 488 5362 552
rect 6909 488 6973 552
rect 6989 488 7053 552
rect 7069 488 7133 552
rect 7149 488 7213 552
rect 7229 488 7293 552
rect 11392 488 11456 552
rect 11472 488 11536 552
rect 11552 488 11616 552
rect 11632 488 11696 552
rect 11712 488 11776 552
rect 11792 488 11856 552
rect 11872 488 11936 552
rect 11952 488 12016 552
rect 12032 488 12096 552
rect 12112 488 12176 552
rect 8 408 72 472
rect 88 408 152 472
rect 168 408 232 472
rect 248 408 312 472
rect 328 408 392 472
rect 408 408 472 472
rect 488 408 552 472
rect 568 408 632 472
rect 648 408 712 472
rect 728 408 792 472
rect 4978 408 5042 472
rect 5058 408 5122 472
rect 5138 408 5202 472
rect 5218 408 5282 472
rect 5298 408 5362 472
rect 6909 408 6973 472
rect 6989 408 7053 472
rect 7069 408 7133 472
rect 7149 408 7213 472
rect 7229 408 7293 472
rect 11392 408 11456 472
rect 11472 408 11536 472
rect 11552 408 11616 472
rect 11632 408 11696 472
rect 11712 408 11776 472
rect 11792 408 11856 472
rect 11872 408 11936 472
rect 11952 408 12016 472
rect 12032 408 12096 472
rect 12112 408 12176 472
rect 8 328 72 392
rect 88 328 152 392
rect 168 328 232 392
rect 248 328 312 392
rect 328 328 392 392
rect 408 328 472 392
rect 488 328 552 392
rect 568 328 632 392
rect 648 328 712 392
rect 728 328 792 392
rect 4978 328 5042 392
rect 5058 328 5122 392
rect 5138 328 5202 392
rect 5218 328 5282 392
rect 5298 328 5362 392
rect 6909 328 6973 392
rect 6989 328 7053 392
rect 7069 328 7133 392
rect 7149 328 7213 392
rect 7229 328 7293 392
rect 11392 328 11456 392
rect 11472 328 11536 392
rect 11552 328 11616 392
rect 11632 328 11696 392
rect 11712 328 11776 392
rect 11792 328 11856 392
rect 11872 328 11936 392
rect 11952 328 12016 392
rect 12032 328 12096 392
rect 12112 328 12176 392
rect 8 248 72 312
rect 88 248 152 312
rect 168 248 232 312
rect 248 248 312 312
rect 328 248 392 312
rect 408 248 472 312
rect 488 248 552 312
rect 568 248 632 312
rect 648 248 712 312
rect 728 248 792 312
rect 4978 248 5042 312
rect 5058 248 5122 312
rect 5138 248 5202 312
rect 5218 248 5282 312
rect 5298 248 5362 312
rect 6909 248 6973 312
rect 6989 248 7053 312
rect 7069 248 7133 312
rect 7149 248 7213 312
rect 7229 248 7293 312
rect 11392 248 11456 312
rect 11472 248 11536 312
rect 11552 248 11616 312
rect 11632 248 11696 312
rect 11712 248 11776 312
rect 11792 248 11856 312
rect 11872 248 11936 312
rect 11952 248 12016 312
rect 12032 248 12096 312
rect 12112 248 12176 312
rect 8 168 72 232
rect 88 168 152 232
rect 168 168 232 232
rect 248 168 312 232
rect 328 168 392 232
rect 408 168 472 232
rect 488 168 552 232
rect 568 168 632 232
rect 648 168 712 232
rect 728 168 792 232
rect 4978 168 5042 232
rect 5058 168 5122 232
rect 5138 168 5202 232
rect 5218 168 5282 232
rect 5298 168 5362 232
rect 6909 168 6973 232
rect 6989 168 7053 232
rect 7069 168 7133 232
rect 7149 168 7213 232
rect 7229 168 7293 232
rect 11392 168 11456 232
rect 11472 168 11536 232
rect 11552 168 11616 232
rect 11632 168 11696 232
rect 11712 168 11776 232
rect 11792 168 11856 232
rect 11872 168 11936 232
rect 11952 168 12016 232
rect 12032 168 12096 232
rect 12112 168 12176 232
rect 8 88 72 152
rect 88 88 152 152
rect 168 88 232 152
rect 248 88 312 152
rect 328 88 392 152
rect 408 88 472 152
rect 488 88 552 152
rect 568 88 632 152
rect 648 88 712 152
rect 728 88 792 152
rect 4978 88 5042 152
rect 5058 88 5122 152
rect 5138 88 5202 152
rect 5218 88 5282 152
rect 5298 88 5362 152
rect 6909 88 6973 152
rect 6989 88 7053 152
rect 7069 88 7133 152
rect 7149 88 7213 152
rect 7229 88 7293 152
rect 11392 88 11456 152
rect 11472 88 11536 152
rect 11552 88 11616 152
rect 11632 88 11696 152
rect 11712 88 11776 152
rect 11792 88 11856 152
rect 11872 88 11936 152
rect 11952 88 12016 152
rect 12032 88 12096 152
rect 12112 88 12176 152
rect 8 8 72 72
rect 88 8 152 72
rect 168 8 232 72
rect 248 8 312 72
rect 328 8 392 72
rect 408 8 472 72
rect 488 8 552 72
rect 568 8 632 72
rect 648 8 712 72
rect 728 8 792 72
rect 4978 8 5042 72
rect 5058 8 5122 72
rect 5138 8 5202 72
rect 5218 8 5282 72
rect 5298 8 5362 72
rect 6909 8 6973 72
rect 6989 8 7053 72
rect 7069 8 7133 72
rect 7149 8 7213 72
rect 7229 8 7293 72
rect 11392 8 11456 72
rect 11472 8 11536 72
rect 11552 8 11616 72
rect 11632 8 11696 72
rect 11712 8 11776 72
rect 11792 8 11856 72
rect 11872 8 11936 72
rect 11952 8 12016 72
rect 12032 8 12096 72
rect 12112 8 12176 72
<< metal4 >>
rect 0 20072 800 20080
rect 0 20008 8 20072
rect 72 20008 88 20072
rect 152 20008 168 20072
rect 232 20008 248 20072
rect 312 20008 328 20072
rect 392 20008 408 20072
rect 472 20008 488 20072
rect 552 20008 568 20072
rect 632 20008 648 20072
rect 712 20008 728 20072
rect 792 20008 800 20072
rect 0 19992 800 20008
rect 0 19928 8 19992
rect 72 19928 88 19992
rect 152 19928 168 19992
rect 232 19928 248 19992
rect 312 19928 328 19992
rect 392 19928 408 19992
rect 472 19928 488 19992
rect 552 19928 568 19992
rect 632 19928 648 19992
rect 712 19928 728 19992
rect 792 19928 800 19992
rect 0 19912 800 19928
rect 0 19848 8 19912
rect 72 19848 88 19912
rect 152 19848 168 19912
rect 232 19848 248 19912
rect 312 19848 328 19912
rect 392 19848 408 19912
rect 472 19848 488 19912
rect 552 19848 568 19912
rect 632 19848 648 19912
rect 712 19848 728 19912
rect 792 19848 800 19912
rect 0 19832 800 19848
rect 0 19768 8 19832
rect 72 19768 88 19832
rect 152 19768 168 19832
rect 232 19768 248 19832
rect 312 19768 328 19832
rect 392 19768 408 19832
rect 472 19768 488 19832
rect 552 19768 568 19832
rect 632 19768 648 19832
rect 712 19768 728 19832
rect 792 19768 800 19832
rect 0 19752 800 19768
rect 0 19688 8 19752
rect 72 19688 88 19752
rect 152 19688 168 19752
rect 232 19688 248 19752
rect 312 19688 328 19752
rect 392 19688 408 19752
rect 472 19688 488 19752
rect 552 19688 568 19752
rect 632 19688 648 19752
rect 712 19688 728 19752
rect 792 19688 800 19752
rect 0 19672 800 19688
rect 0 19608 8 19672
rect 72 19608 88 19672
rect 152 19608 168 19672
rect 232 19608 248 19672
rect 312 19608 328 19672
rect 392 19608 408 19672
rect 472 19608 488 19672
rect 552 19608 568 19672
rect 632 19608 648 19672
rect 712 19608 728 19672
rect 792 19608 800 19672
rect 0 19592 800 19608
rect 0 19528 8 19592
rect 72 19528 88 19592
rect 152 19528 168 19592
rect 232 19528 248 19592
rect 312 19528 328 19592
rect 392 19528 408 19592
rect 472 19528 488 19592
rect 552 19528 568 19592
rect 632 19528 648 19592
rect 712 19528 728 19592
rect 792 19528 800 19592
rect 0 19512 800 19528
rect 0 19448 8 19512
rect 72 19448 88 19512
rect 152 19448 168 19512
rect 232 19448 248 19512
rect 312 19448 328 19512
rect 392 19448 408 19512
rect 472 19448 488 19512
rect 552 19448 568 19512
rect 632 19448 648 19512
rect 712 19448 728 19512
rect 792 19448 800 19512
rect 0 19432 800 19448
rect 0 19368 8 19432
rect 72 19368 88 19432
rect 152 19368 168 19432
rect 232 19368 248 19432
rect 312 19368 328 19432
rect 392 19368 408 19432
rect 472 19368 488 19432
rect 552 19368 568 19432
rect 632 19368 648 19432
rect 712 19368 728 19432
rect 792 19368 800 19432
rect 0 19352 800 19368
rect 0 19288 8 19352
rect 72 19288 88 19352
rect 152 19288 168 19352
rect 232 19288 248 19352
rect 312 19288 328 19352
rect 392 19288 408 19352
rect 472 19288 488 19352
rect 552 19288 568 19352
rect 632 19288 648 19352
rect 712 19288 728 19352
rect 792 19288 800 19352
rect 0 792 800 19288
rect 1140 18932 1940 18940
rect 1140 18868 1148 18932
rect 1212 18868 1228 18932
rect 1292 18868 1308 18932
rect 1372 18868 1388 18932
rect 1452 18868 1468 18932
rect 1532 18868 1548 18932
rect 1612 18868 1628 18932
rect 1692 18868 1708 18932
rect 1772 18868 1788 18932
rect 1852 18868 1868 18932
rect 1932 18868 1940 18932
rect 1140 18852 1940 18868
rect 1140 18788 1148 18852
rect 1212 18788 1228 18852
rect 1292 18788 1308 18852
rect 1372 18788 1388 18852
rect 1452 18788 1468 18852
rect 1532 18788 1548 18852
rect 1612 18788 1628 18852
rect 1692 18788 1708 18852
rect 1772 18788 1788 18852
rect 1852 18788 1868 18852
rect 1932 18788 1940 18852
rect 1140 18772 1940 18788
rect 1140 18708 1148 18772
rect 1212 18708 1228 18772
rect 1292 18708 1308 18772
rect 1372 18708 1388 18772
rect 1452 18708 1468 18772
rect 1532 18708 1548 18772
rect 1612 18708 1628 18772
rect 1692 18708 1708 18772
rect 1772 18708 1788 18772
rect 1852 18708 1868 18772
rect 1932 18708 1940 18772
rect 1140 18692 1940 18708
rect 1140 18628 1148 18692
rect 1212 18628 1228 18692
rect 1292 18628 1308 18692
rect 1372 18628 1388 18692
rect 1452 18628 1468 18692
rect 1532 18628 1548 18692
rect 1612 18628 1628 18692
rect 1692 18628 1708 18692
rect 1772 18628 1788 18692
rect 1852 18628 1868 18692
rect 1932 18628 1940 18692
rect 1140 18612 1940 18628
rect 1140 18548 1148 18612
rect 1212 18548 1228 18612
rect 1292 18548 1308 18612
rect 1372 18548 1388 18612
rect 1452 18548 1468 18612
rect 1532 18548 1548 18612
rect 1612 18548 1628 18612
rect 1692 18548 1708 18612
rect 1772 18548 1788 18612
rect 1852 18548 1868 18612
rect 1932 18548 1940 18612
rect 1140 18532 1940 18548
rect 1140 18468 1148 18532
rect 1212 18468 1228 18532
rect 1292 18468 1308 18532
rect 1372 18468 1388 18532
rect 1452 18468 1468 18532
rect 1532 18468 1548 18532
rect 1612 18468 1628 18532
rect 1692 18468 1708 18532
rect 1772 18468 1788 18532
rect 1852 18468 1868 18532
rect 1932 18468 1940 18532
rect 1140 18452 1940 18468
rect 1140 18388 1148 18452
rect 1212 18388 1228 18452
rect 1292 18388 1308 18452
rect 1372 18388 1388 18452
rect 1452 18388 1468 18452
rect 1532 18388 1548 18452
rect 1612 18388 1628 18452
rect 1692 18388 1708 18452
rect 1772 18388 1788 18452
rect 1852 18388 1868 18452
rect 1932 18388 1940 18452
rect 1140 18372 1940 18388
rect 1140 18308 1148 18372
rect 1212 18308 1228 18372
rect 1292 18308 1308 18372
rect 1372 18308 1388 18372
rect 1452 18308 1468 18372
rect 1532 18308 1548 18372
rect 1612 18308 1628 18372
rect 1692 18308 1708 18372
rect 1772 18308 1788 18372
rect 1852 18308 1868 18372
rect 1932 18308 1940 18372
rect 1140 18292 1940 18308
rect 1140 18228 1148 18292
rect 1212 18228 1228 18292
rect 1292 18228 1308 18292
rect 1372 18228 1388 18292
rect 1452 18228 1468 18292
rect 1532 18228 1548 18292
rect 1612 18228 1628 18292
rect 1692 18228 1708 18292
rect 1772 18228 1788 18292
rect 1852 18228 1868 18292
rect 1932 18228 1940 18292
rect 1140 18212 1940 18228
rect 1140 18148 1148 18212
rect 1212 18148 1228 18212
rect 1292 18148 1308 18212
rect 1372 18148 1388 18212
rect 1452 18148 1468 18212
rect 1532 18148 1548 18212
rect 1612 18148 1628 18212
rect 1692 18148 1708 18212
rect 1772 18148 1788 18212
rect 1852 18148 1868 18212
rect 1932 18148 1940 18212
rect 1140 1932 1940 18148
rect 1140 1868 1148 1932
rect 1212 1868 1228 1932
rect 1292 1868 1308 1932
rect 1372 1868 1388 1932
rect 1452 1868 1468 1932
rect 1532 1868 1548 1932
rect 1612 1868 1628 1932
rect 1692 1868 1708 1932
rect 1772 1868 1788 1932
rect 1852 1868 1868 1932
rect 1932 1868 1940 1932
rect 1140 1852 1940 1868
rect 1140 1788 1148 1852
rect 1212 1788 1228 1852
rect 1292 1788 1308 1852
rect 1372 1788 1388 1852
rect 1452 1788 1468 1852
rect 1532 1788 1548 1852
rect 1612 1788 1628 1852
rect 1692 1788 1708 1852
rect 1772 1788 1788 1852
rect 1852 1788 1868 1852
rect 1932 1788 1940 1852
rect 1140 1772 1940 1788
rect 1140 1708 1148 1772
rect 1212 1708 1228 1772
rect 1292 1708 1308 1772
rect 1372 1708 1388 1772
rect 1452 1708 1468 1772
rect 1532 1708 1548 1772
rect 1612 1708 1628 1772
rect 1692 1708 1708 1772
rect 1772 1708 1788 1772
rect 1852 1708 1868 1772
rect 1932 1708 1940 1772
rect 1140 1692 1940 1708
rect 1140 1628 1148 1692
rect 1212 1628 1228 1692
rect 1292 1628 1308 1692
rect 1372 1628 1388 1692
rect 1452 1628 1468 1692
rect 1532 1628 1548 1692
rect 1612 1628 1628 1692
rect 1692 1628 1708 1692
rect 1772 1628 1788 1692
rect 1852 1628 1868 1692
rect 1932 1628 1940 1692
rect 1140 1612 1940 1628
rect 1140 1548 1148 1612
rect 1212 1548 1228 1612
rect 1292 1548 1308 1612
rect 1372 1548 1388 1612
rect 1452 1548 1468 1612
rect 1532 1548 1548 1612
rect 1612 1548 1628 1612
rect 1692 1548 1708 1612
rect 1772 1548 1788 1612
rect 1852 1548 1868 1612
rect 1932 1548 1940 1612
rect 1140 1532 1940 1548
rect 1140 1468 1148 1532
rect 1212 1468 1228 1532
rect 1292 1468 1308 1532
rect 1372 1468 1388 1532
rect 1452 1468 1468 1532
rect 1532 1468 1548 1532
rect 1612 1468 1628 1532
rect 1692 1468 1708 1532
rect 1772 1468 1788 1532
rect 1852 1468 1868 1532
rect 1932 1468 1940 1532
rect 1140 1452 1940 1468
rect 1140 1388 1148 1452
rect 1212 1388 1228 1452
rect 1292 1388 1308 1452
rect 1372 1388 1388 1452
rect 1452 1388 1468 1452
rect 1532 1388 1548 1452
rect 1612 1388 1628 1452
rect 1692 1388 1708 1452
rect 1772 1388 1788 1452
rect 1852 1388 1868 1452
rect 1932 1388 1940 1452
rect 1140 1372 1940 1388
rect 1140 1308 1148 1372
rect 1212 1308 1228 1372
rect 1292 1308 1308 1372
rect 1372 1308 1388 1372
rect 1452 1308 1468 1372
rect 1532 1308 1548 1372
rect 1612 1308 1628 1372
rect 1692 1308 1708 1372
rect 1772 1308 1788 1372
rect 1852 1308 1868 1372
rect 1932 1308 1940 1372
rect 1140 1292 1940 1308
rect 1140 1228 1148 1292
rect 1212 1228 1228 1292
rect 1292 1228 1308 1292
rect 1372 1228 1388 1292
rect 1452 1228 1468 1292
rect 1532 1228 1548 1292
rect 1612 1228 1628 1292
rect 1692 1228 1708 1292
rect 1772 1228 1788 1292
rect 1852 1228 1868 1292
rect 1932 1228 1940 1292
rect 1140 1212 1940 1228
rect 1140 1148 1148 1212
rect 1212 1148 1228 1212
rect 1292 1148 1308 1212
rect 1372 1148 1388 1212
rect 1452 1148 1468 1212
rect 1532 1148 1548 1212
rect 1612 1148 1628 1212
rect 1692 1148 1708 1212
rect 1772 1148 1788 1212
rect 1852 1148 1868 1212
rect 1932 1148 1940 1212
rect 1140 1140 1940 1148
rect 3995 18932 4415 20080
rect 3995 18868 4013 18932
rect 4077 18868 4093 18932
rect 4157 18868 4173 18932
rect 4237 18868 4253 18932
rect 4317 18868 4333 18932
rect 4397 18868 4415 18932
rect 3995 18852 4415 18868
rect 3995 18788 4013 18852
rect 4077 18788 4093 18852
rect 4157 18788 4173 18852
rect 4237 18788 4253 18852
rect 4317 18788 4333 18852
rect 4397 18788 4415 18852
rect 3995 18772 4415 18788
rect 3995 18708 4013 18772
rect 4077 18708 4093 18772
rect 4157 18708 4173 18772
rect 4237 18708 4253 18772
rect 4317 18708 4333 18772
rect 4397 18708 4415 18772
rect 3995 18692 4415 18708
rect 3995 18628 4013 18692
rect 4077 18628 4093 18692
rect 4157 18628 4173 18692
rect 4237 18628 4253 18692
rect 4317 18628 4333 18692
rect 4397 18628 4415 18692
rect 3995 18612 4415 18628
rect 3995 18548 4013 18612
rect 4077 18548 4093 18612
rect 4157 18548 4173 18612
rect 4237 18548 4253 18612
rect 4317 18548 4333 18612
rect 4397 18548 4415 18612
rect 3995 18532 4415 18548
rect 3995 18468 4013 18532
rect 4077 18468 4093 18532
rect 4157 18468 4173 18532
rect 4237 18468 4253 18532
rect 4317 18468 4333 18532
rect 4397 18468 4415 18532
rect 3995 18452 4415 18468
rect 3995 18388 4013 18452
rect 4077 18388 4093 18452
rect 4157 18388 4173 18452
rect 4237 18388 4253 18452
rect 4317 18388 4333 18452
rect 4397 18388 4415 18452
rect 3995 18372 4415 18388
rect 3995 18308 4013 18372
rect 4077 18308 4093 18372
rect 4157 18308 4173 18372
rect 4237 18308 4253 18372
rect 4317 18308 4333 18372
rect 4397 18308 4415 18372
rect 3995 18292 4415 18308
rect 3995 18228 4013 18292
rect 4077 18228 4093 18292
rect 4157 18228 4173 18292
rect 4237 18228 4253 18292
rect 4317 18228 4333 18292
rect 4397 18228 4415 18292
rect 3995 18212 4415 18228
rect 3995 18148 4013 18212
rect 4077 18148 4093 18212
rect 4157 18148 4173 18212
rect 4237 18148 4253 18212
rect 4317 18148 4333 18212
rect 4397 18148 4415 18212
rect 3995 16328 4415 18148
rect 3995 16264 4013 16328
rect 4077 16264 4093 16328
rect 4157 16264 4173 16328
rect 4237 16264 4253 16328
rect 4317 16264 4333 16328
rect 4397 16264 4415 16328
rect 3995 15240 4415 16264
rect 3995 15176 4013 15240
rect 4077 15176 4093 15240
rect 4157 15176 4173 15240
rect 4237 15176 4253 15240
rect 4317 15176 4333 15240
rect 4397 15176 4415 15240
rect 3995 14152 4415 15176
rect 3995 14088 4013 14152
rect 4077 14088 4093 14152
rect 4157 14088 4173 14152
rect 4237 14088 4253 14152
rect 4317 14088 4333 14152
rect 4397 14088 4415 14152
rect 3995 13064 4415 14088
rect 3995 13000 4013 13064
rect 4077 13000 4093 13064
rect 4157 13000 4173 13064
rect 4237 13000 4253 13064
rect 4317 13000 4333 13064
rect 4397 13000 4415 13064
rect 3995 11976 4415 13000
rect 3995 11912 4013 11976
rect 4077 11912 4093 11976
rect 4157 11912 4173 11976
rect 4237 11912 4253 11976
rect 4317 11912 4333 11976
rect 4397 11912 4415 11976
rect 3995 10888 4415 11912
rect 3995 10824 4013 10888
rect 4077 10824 4093 10888
rect 4157 10824 4173 10888
rect 4237 10824 4253 10888
rect 4317 10824 4333 10888
rect 4397 10824 4415 10888
rect 3995 9800 4415 10824
rect 3995 9736 4013 9800
rect 4077 9736 4093 9800
rect 4157 9736 4173 9800
rect 4237 9736 4253 9800
rect 4317 9736 4333 9800
rect 4397 9736 4415 9800
rect 3995 8712 4415 9736
rect 3995 8648 4013 8712
rect 4077 8648 4093 8712
rect 4157 8648 4173 8712
rect 4237 8648 4253 8712
rect 4317 8648 4333 8712
rect 4397 8648 4415 8712
rect 3995 7624 4415 8648
rect 3995 7560 4013 7624
rect 4077 7560 4093 7624
rect 4157 7560 4173 7624
rect 4237 7560 4253 7624
rect 4317 7560 4333 7624
rect 4397 7560 4415 7624
rect 3995 6536 4415 7560
rect 3995 6472 4013 6536
rect 4077 6472 4093 6536
rect 4157 6472 4173 6536
rect 4237 6472 4253 6536
rect 4317 6472 4333 6536
rect 4397 6472 4415 6536
rect 3995 5448 4415 6472
rect 3995 5384 4013 5448
rect 4077 5384 4093 5448
rect 4157 5384 4173 5448
rect 4237 5384 4253 5448
rect 4317 5384 4333 5448
rect 4397 5384 4415 5448
rect 3995 4360 4415 5384
rect 3995 4296 4013 4360
rect 4077 4296 4093 4360
rect 4157 4296 4173 4360
rect 4237 4296 4253 4360
rect 4317 4296 4333 4360
rect 4397 4296 4415 4360
rect 3995 3272 4415 4296
rect 3995 3208 4013 3272
rect 4077 3208 4093 3272
rect 4157 3208 4173 3272
rect 4237 3208 4253 3272
rect 4317 3208 4333 3272
rect 4397 3208 4415 3272
rect 3995 1932 4415 3208
rect 3995 1868 4013 1932
rect 4077 1868 4093 1932
rect 4157 1868 4173 1932
rect 4237 1868 4253 1932
rect 4317 1868 4333 1932
rect 4397 1868 4415 1932
rect 3995 1852 4415 1868
rect 3995 1788 4013 1852
rect 4077 1788 4093 1852
rect 4157 1788 4173 1852
rect 4237 1788 4253 1852
rect 4317 1788 4333 1852
rect 4397 1788 4415 1852
rect 3995 1772 4415 1788
rect 3995 1708 4013 1772
rect 4077 1708 4093 1772
rect 4157 1708 4173 1772
rect 4237 1708 4253 1772
rect 4317 1708 4333 1772
rect 4397 1708 4415 1772
rect 3995 1692 4415 1708
rect 3995 1628 4013 1692
rect 4077 1628 4093 1692
rect 4157 1628 4173 1692
rect 4237 1628 4253 1692
rect 4317 1628 4333 1692
rect 4397 1628 4415 1692
rect 3995 1612 4415 1628
rect 3995 1548 4013 1612
rect 4077 1548 4093 1612
rect 4157 1548 4173 1612
rect 4237 1548 4253 1612
rect 4317 1548 4333 1612
rect 4397 1548 4415 1612
rect 3995 1532 4415 1548
rect 3995 1468 4013 1532
rect 4077 1468 4093 1532
rect 4157 1468 4173 1532
rect 4237 1468 4253 1532
rect 4317 1468 4333 1532
rect 4397 1468 4415 1532
rect 3995 1452 4415 1468
rect 3995 1388 4013 1452
rect 4077 1388 4093 1452
rect 4157 1388 4173 1452
rect 4237 1388 4253 1452
rect 4317 1388 4333 1452
rect 4397 1388 4415 1452
rect 3995 1372 4415 1388
rect 3995 1308 4013 1372
rect 4077 1308 4093 1372
rect 4157 1308 4173 1372
rect 4237 1308 4253 1372
rect 4317 1308 4333 1372
rect 4397 1308 4415 1372
rect 3995 1292 4415 1308
rect 3995 1228 4013 1292
rect 4077 1228 4093 1292
rect 4157 1228 4173 1292
rect 4237 1228 4253 1292
rect 4317 1228 4333 1292
rect 4397 1228 4415 1292
rect 3995 1212 4415 1228
rect 3995 1148 4013 1212
rect 4077 1148 4093 1212
rect 4157 1148 4173 1212
rect 4237 1148 4253 1212
rect 4317 1148 4333 1212
rect 4397 1148 4415 1212
rect 0 728 8 792
rect 72 728 88 792
rect 152 728 168 792
rect 232 728 248 792
rect 312 728 328 792
rect 392 728 408 792
rect 472 728 488 792
rect 552 728 568 792
rect 632 728 648 792
rect 712 728 728 792
rect 792 728 800 792
rect 0 712 800 728
rect 0 648 8 712
rect 72 648 88 712
rect 152 648 168 712
rect 232 648 248 712
rect 312 648 328 712
rect 392 648 408 712
rect 472 648 488 712
rect 552 648 568 712
rect 632 648 648 712
rect 712 648 728 712
rect 792 648 800 712
rect 0 632 800 648
rect 0 568 8 632
rect 72 568 88 632
rect 152 568 168 632
rect 232 568 248 632
rect 312 568 328 632
rect 392 568 408 632
rect 472 568 488 632
rect 552 568 568 632
rect 632 568 648 632
rect 712 568 728 632
rect 792 568 800 632
rect 0 552 800 568
rect 0 488 8 552
rect 72 488 88 552
rect 152 488 168 552
rect 232 488 248 552
rect 312 488 328 552
rect 392 488 408 552
rect 472 488 488 552
rect 552 488 568 552
rect 632 488 648 552
rect 712 488 728 552
rect 792 488 800 552
rect 0 472 800 488
rect 0 408 8 472
rect 72 408 88 472
rect 152 408 168 472
rect 232 408 248 472
rect 312 408 328 472
rect 392 408 408 472
rect 472 408 488 472
rect 552 408 568 472
rect 632 408 648 472
rect 712 408 728 472
rect 792 408 800 472
rect 0 392 800 408
rect 0 328 8 392
rect 72 328 88 392
rect 152 328 168 392
rect 232 328 248 392
rect 312 328 328 392
rect 392 328 408 392
rect 472 328 488 392
rect 552 328 568 392
rect 632 328 648 392
rect 712 328 728 392
rect 792 328 800 392
rect 0 312 800 328
rect 0 248 8 312
rect 72 248 88 312
rect 152 248 168 312
rect 232 248 248 312
rect 312 248 328 312
rect 392 248 408 312
rect 472 248 488 312
rect 552 248 568 312
rect 632 248 648 312
rect 712 248 728 312
rect 792 248 800 312
rect 0 232 800 248
rect 0 168 8 232
rect 72 168 88 232
rect 152 168 168 232
rect 232 168 248 232
rect 312 168 328 232
rect 392 168 408 232
rect 472 168 488 232
rect 552 168 568 232
rect 632 168 648 232
rect 712 168 728 232
rect 792 168 800 232
rect 0 152 800 168
rect 0 88 8 152
rect 72 88 88 152
rect 152 88 168 152
rect 232 88 248 152
rect 312 88 328 152
rect 392 88 408 152
rect 472 88 488 152
rect 552 88 568 152
rect 632 88 648 152
rect 712 88 728 152
rect 792 88 800 152
rect 0 72 800 88
rect 0 8 8 72
rect 72 8 88 72
rect 152 8 168 72
rect 232 8 248 72
rect 312 8 328 72
rect 392 8 408 72
rect 472 8 488 72
rect 552 8 568 72
rect 632 8 648 72
rect 712 8 728 72
rect 792 8 800 72
rect 0 0 800 8
rect 3995 0 4415 1148
rect 4960 20072 5381 20080
rect 4960 20008 4978 20072
rect 5042 20008 5058 20072
rect 5122 20008 5138 20072
rect 5202 20008 5218 20072
rect 5282 20008 5298 20072
rect 5362 20008 5381 20072
rect 4960 19992 5381 20008
rect 4960 19928 4978 19992
rect 5042 19928 5058 19992
rect 5122 19928 5138 19992
rect 5202 19928 5218 19992
rect 5282 19928 5298 19992
rect 5362 19928 5381 19992
rect 4960 19912 5381 19928
rect 4960 19848 4978 19912
rect 5042 19848 5058 19912
rect 5122 19848 5138 19912
rect 5202 19848 5218 19912
rect 5282 19848 5298 19912
rect 5362 19848 5381 19912
rect 4960 19832 5381 19848
rect 4960 19768 4978 19832
rect 5042 19768 5058 19832
rect 5122 19768 5138 19832
rect 5202 19768 5218 19832
rect 5282 19768 5298 19832
rect 5362 19768 5381 19832
rect 4960 19752 5381 19768
rect 4960 19688 4978 19752
rect 5042 19688 5058 19752
rect 5122 19688 5138 19752
rect 5202 19688 5218 19752
rect 5282 19688 5298 19752
rect 5362 19688 5381 19752
rect 4960 19672 5381 19688
rect 4960 19608 4978 19672
rect 5042 19608 5058 19672
rect 5122 19608 5138 19672
rect 5202 19608 5218 19672
rect 5282 19608 5298 19672
rect 5362 19608 5381 19672
rect 4960 19592 5381 19608
rect 4960 19528 4978 19592
rect 5042 19528 5058 19592
rect 5122 19528 5138 19592
rect 5202 19528 5218 19592
rect 5282 19528 5298 19592
rect 5362 19528 5381 19592
rect 4960 19512 5381 19528
rect 4960 19448 4978 19512
rect 5042 19448 5058 19512
rect 5122 19448 5138 19512
rect 5202 19448 5218 19512
rect 5282 19448 5298 19512
rect 5362 19448 5381 19512
rect 4960 19432 5381 19448
rect 4960 19368 4978 19432
rect 5042 19368 5058 19432
rect 5122 19368 5138 19432
rect 5202 19368 5218 19432
rect 5282 19368 5298 19432
rect 5362 19368 5381 19432
rect 4960 19352 5381 19368
rect 4960 19288 4978 19352
rect 5042 19288 5058 19352
rect 5122 19288 5138 19352
rect 5202 19288 5218 19352
rect 5282 19288 5298 19352
rect 5362 19288 5381 19352
rect 4960 16872 5381 19288
rect 4960 16808 4978 16872
rect 5042 16808 5058 16872
rect 5122 16808 5138 16872
rect 5202 16808 5218 16872
rect 5282 16808 5298 16872
rect 5362 16808 5381 16872
rect 4960 15784 5381 16808
rect 4960 15720 4978 15784
rect 5042 15720 5058 15784
rect 5122 15720 5138 15784
rect 5202 15720 5218 15784
rect 5282 15720 5298 15784
rect 5362 15720 5381 15784
rect 4960 14696 5381 15720
rect 4960 14632 4978 14696
rect 5042 14632 5058 14696
rect 5122 14632 5138 14696
rect 5202 14632 5218 14696
rect 5282 14632 5298 14696
rect 5362 14632 5381 14696
rect 4960 13608 5381 14632
rect 4960 13544 4978 13608
rect 5042 13544 5058 13608
rect 5122 13544 5138 13608
rect 5202 13544 5218 13608
rect 5282 13544 5298 13608
rect 5362 13544 5381 13608
rect 4960 12520 5381 13544
rect 4960 12456 4978 12520
rect 5042 12456 5058 12520
rect 5122 12456 5138 12520
rect 5202 12456 5218 12520
rect 5282 12456 5298 12520
rect 5362 12456 5381 12520
rect 4960 11432 5381 12456
rect 4960 11368 4978 11432
rect 5042 11368 5058 11432
rect 5122 11368 5138 11432
rect 5202 11368 5218 11432
rect 5282 11368 5298 11432
rect 5362 11368 5381 11432
rect 4960 10344 5381 11368
rect 4960 10280 4978 10344
rect 5042 10280 5058 10344
rect 5122 10280 5138 10344
rect 5202 10280 5218 10344
rect 5282 10280 5298 10344
rect 5362 10280 5381 10344
rect 4960 9256 5381 10280
rect 4960 9192 4978 9256
rect 5042 9192 5058 9256
rect 5122 9192 5138 9256
rect 5202 9192 5218 9256
rect 5282 9192 5298 9256
rect 5362 9192 5381 9256
rect 4960 8168 5381 9192
rect 4960 8104 4978 8168
rect 5042 8104 5058 8168
rect 5122 8104 5138 8168
rect 5202 8104 5218 8168
rect 5282 8104 5298 8168
rect 5362 8104 5381 8168
rect 4960 7080 5381 8104
rect 4960 7016 4978 7080
rect 5042 7016 5058 7080
rect 5122 7016 5138 7080
rect 5202 7016 5218 7080
rect 5282 7016 5298 7080
rect 5362 7016 5381 7080
rect 4960 5992 5381 7016
rect 4960 5928 4978 5992
rect 5042 5928 5058 5992
rect 5122 5928 5138 5992
rect 5202 5928 5218 5992
rect 5282 5928 5298 5992
rect 5362 5928 5381 5992
rect 4960 4904 5381 5928
rect 4960 4840 4978 4904
rect 5042 4840 5058 4904
rect 5122 4840 5138 4904
rect 5202 4840 5218 4904
rect 5282 4840 5298 4904
rect 5362 4840 5381 4904
rect 4960 3816 5381 4840
rect 4960 3752 4978 3816
rect 5042 3752 5058 3816
rect 5122 3752 5138 3816
rect 5202 3752 5218 3816
rect 5282 3752 5298 3816
rect 5362 3752 5381 3816
rect 4960 792 5381 3752
rect 4960 728 4978 792
rect 5042 728 5058 792
rect 5122 728 5138 792
rect 5202 728 5218 792
rect 5282 728 5298 792
rect 5362 728 5381 792
rect 4960 712 5381 728
rect 4960 648 4978 712
rect 5042 648 5058 712
rect 5122 648 5138 712
rect 5202 648 5218 712
rect 5282 648 5298 712
rect 5362 648 5381 712
rect 4960 632 5381 648
rect 4960 568 4978 632
rect 5042 568 5058 632
rect 5122 568 5138 632
rect 5202 568 5218 632
rect 5282 568 5298 632
rect 5362 568 5381 632
rect 4960 552 5381 568
rect 4960 488 4978 552
rect 5042 488 5058 552
rect 5122 488 5138 552
rect 5202 488 5218 552
rect 5282 488 5298 552
rect 5362 488 5381 552
rect 4960 472 5381 488
rect 4960 408 4978 472
rect 5042 408 5058 472
rect 5122 408 5138 472
rect 5202 408 5218 472
rect 5282 408 5298 472
rect 5362 408 5381 472
rect 4960 392 5381 408
rect 4960 328 4978 392
rect 5042 328 5058 392
rect 5122 328 5138 392
rect 5202 328 5218 392
rect 5282 328 5298 392
rect 5362 328 5381 392
rect 4960 312 5381 328
rect 4960 248 4978 312
rect 5042 248 5058 312
rect 5122 248 5138 312
rect 5202 248 5218 312
rect 5282 248 5298 312
rect 5362 248 5381 312
rect 4960 232 5381 248
rect 4960 168 4978 232
rect 5042 168 5058 232
rect 5122 168 5138 232
rect 5202 168 5218 232
rect 5282 168 5298 232
rect 5362 168 5381 232
rect 4960 152 5381 168
rect 4960 88 4978 152
rect 5042 88 5058 152
rect 5122 88 5138 152
rect 5202 88 5218 152
rect 5282 88 5298 152
rect 5362 88 5381 152
rect 4960 72 5381 88
rect 4960 8 4978 72
rect 5042 8 5058 72
rect 5122 8 5138 72
rect 5202 8 5218 72
rect 5282 8 5298 72
rect 5362 8 5381 72
rect 4960 0 5381 8
rect 5926 18932 6346 20080
rect 5926 18868 5944 18932
rect 6008 18868 6024 18932
rect 6088 18868 6104 18932
rect 6168 18868 6184 18932
rect 6248 18868 6264 18932
rect 6328 18868 6346 18932
rect 5926 18852 6346 18868
rect 5926 18788 5944 18852
rect 6008 18788 6024 18852
rect 6088 18788 6104 18852
rect 6168 18788 6184 18852
rect 6248 18788 6264 18852
rect 6328 18788 6346 18852
rect 5926 18772 6346 18788
rect 5926 18708 5944 18772
rect 6008 18708 6024 18772
rect 6088 18708 6104 18772
rect 6168 18708 6184 18772
rect 6248 18708 6264 18772
rect 6328 18708 6346 18772
rect 5926 18692 6346 18708
rect 5926 18628 5944 18692
rect 6008 18628 6024 18692
rect 6088 18628 6104 18692
rect 6168 18628 6184 18692
rect 6248 18628 6264 18692
rect 6328 18628 6346 18692
rect 5926 18612 6346 18628
rect 5926 18548 5944 18612
rect 6008 18548 6024 18612
rect 6088 18548 6104 18612
rect 6168 18548 6184 18612
rect 6248 18548 6264 18612
rect 6328 18548 6346 18612
rect 5926 18532 6346 18548
rect 5926 18468 5944 18532
rect 6008 18468 6024 18532
rect 6088 18468 6104 18532
rect 6168 18468 6184 18532
rect 6248 18468 6264 18532
rect 6328 18468 6346 18532
rect 5926 18452 6346 18468
rect 5926 18388 5944 18452
rect 6008 18388 6024 18452
rect 6088 18388 6104 18452
rect 6168 18388 6184 18452
rect 6248 18388 6264 18452
rect 6328 18388 6346 18452
rect 5926 18372 6346 18388
rect 5926 18308 5944 18372
rect 6008 18308 6024 18372
rect 6088 18308 6104 18372
rect 6168 18308 6184 18372
rect 6248 18308 6264 18372
rect 6328 18308 6346 18372
rect 5926 18292 6346 18308
rect 5926 18228 5944 18292
rect 6008 18228 6024 18292
rect 6088 18228 6104 18292
rect 6168 18228 6184 18292
rect 6248 18228 6264 18292
rect 6328 18228 6346 18292
rect 5926 18212 6346 18228
rect 5926 18148 5944 18212
rect 6008 18148 6024 18212
rect 6088 18148 6104 18212
rect 6168 18148 6184 18212
rect 6248 18148 6264 18212
rect 6328 18148 6346 18212
rect 5926 16328 6346 18148
rect 5926 16264 5944 16328
rect 6008 16264 6024 16328
rect 6088 16264 6104 16328
rect 6168 16264 6184 16328
rect 6248 16264 6264 16328
rect 6328 16264 6346 16328
rect 5926 15240 6346 16264
rect 5926 15176 5944 15240
rect 6008 15176 6024 15240
rect 6088 15176 6104 15240
rect 6168 15176 6184 15240
rect 6248 15176 6264 15240
rect 6328 15176 6346 15240
rect 5926 14152 6346 15176
rect 5926 14088 5944 14152
rect 6008 14088 6024 14152
rect 6088 14088 6104 14152
rect 6168 14088 6184 14152
rect 6248 14088 6264 14152
rect 6328 14088 6346 14152
rect 5926 13064 6346 14088
rect 5926 13000 5944 13064
rect 6008 13000 6024 13064
rect 6088 13000 6104 13064
rect 6168 13000 6184 13064
rect 6248 13000 6264 13064
rect 6328 13000 6346 13064
rect 5926 11976 6346 13000
rect 5926 11912 5944 11976
rect 6008 11912 6024 11976
rect 6088 11912 6104 11976
rect 6168 11912 6184 11976
rect 6248 11912 6264 11976
rect 6328 11912 6346 11976
rect 5926 10888 6346 11912
rect 5926 10824 5944 10888
rect 6008 10824 6024 10888
rect 6088 10824 6104 10888
rect 6168 10824 6184 10888
rect 6248 10824 6264 10888
rect 6328 10824 6346 10888
rect 5926 9800 6346 10824
rect 5926 9736 5944 9800
rect 6008 9736 6024 9800
rect 6088 9736 6104 9800
rect 6168 9736 6184 9800
rect 6248 9736 6264 9800
rect 6328 9736 6346 9800
rect 5926 8712 6346 9736
rect 5926 8648 5944 8712
rect 6008 8648 6024 8712
rect 6088 8648 6104 8712
rect 6168 8648 6184 8712
rect 6248 8648 6264 8712
rect 6328 8648 6346 8712
rect 5926 7624 6346 8648
rect 5926 7560 5944 7624
rect 6008 7560 6024 7624
rect 6088 7560 6104 7624
rect 6168 7560 6184 7624
rect 6248 7560 6264 7624
rect 6328 7560 6346 7624
rect 5926 6536 6346 7560
rect 5926 6472 5944 6536
rect 6008 6472 6024 6536
rect 6088 6472 6104 6536
rect 6168 6472 6184 6536
rect 6248 6472 6264 6536
rect 6328 6472 6346 6536
rect 5926 5448 6346 6472
rect 5926 5384 5944 5448
rect 6008 5384 6024 5448
rect 6088 5384 6104 5448
rect 6168 5384 6184 5448
rect 6248 5384 6264 5448
rect 6328 5384 6346 5448
rect 5926 4360 6346 5384
rect 5926 4296 5944 4360
rect 6008 4296 6024 4360
rect 6088 4296 6104 4360
rect 6168 4296 6184 4360
rect 6248 4296 6264 4360
rect 6328 4296 6346 4360
rect 5926 3272 6346 4296
rect 5926 3208 5944 3272
rect 6008 3208 6024 3272
rect 6088 3208 6104 3272
rect 6168 3208 6184 3272
rect 6248 3208 6264 3272
rect 6328 3208 6346 3272
rect 5926 1932 6346 3208
rect 5926 1868 5944 1932
rect 6008 1868 6024 1932
rect 6088 1868 6104 1932
rect 6168 1868 6184 1932
rect 6248 1868 6264 1932
rect 6328 1868 6346 1932
rect 5926 1852 6346 1868
rect 5926 1788 5944 1852
rect 6008 1788 6024 1852
rect 6088 1788 6104 1852
rect 6168 1788 6184 1852
rect 6248 1788 6264 1852
rect 6328 1788 6346 1852
rect 5926 1772 6346 1788
rect 5926 1708 5944 1772
rect 6008 1708 6024 1772
rect 6088 1708 6104 1772
rect 6168 1708 6184 1772
rect 6248 1708 6264 1772
rect 6328 1708 6346 1772
rect 5926 1692 6346 1708
rect 5926 1628 5944 1692
rect 6008 1628 6024 1692
rect 6088 1628 6104 1692
rect 6168 1628 6184 1692
rect 6248 1628 6264 1692
rect 6328 1628 6346 1692
rect 5926 1612 6346 1628
rect 5926 1548 5944 1612
rect 6008 1548 6024 1612
rect 6088 1548 6104 1612
rect 6168 1548 6184 1612
rect 6248 1548 6264 1612
rect 6328 1548 6346 1612
rect 5926 1532 6346 1548
rect 5926 1468 5944 1532
rect 6008 1468 6024 1532
rect 6088 1468 6104 1532
rect 6168 1468 6184 1532
rect 6248 1468 6264 1532
rect 6328 1468 6346 1532
rect 5926 1452 6346 1468
rect 5926 1388 5944 1452
rect 6008 1388 6024 1452
rect 6088 1388 6104 1452
rect 6168 1388 6184 1452
rect 6248 1388 6264 1452
rect 6328 1388 6346 1452
rect 5926 1372 6346 1388
rect 5926 1308 5944 1372
rect 6008 1308 6024 1372
rect 6088 1308 6104 1372
rect 6168 1308 6184 1372
rect 6248 1308 6264 1372
rect 6328 1308 6346 1372
rect 5926 1292 6346 1308
rect 5926 1228 5944 1292
rect 6008 1228 6024 1292
rect 6088 1228 6104 1292
rect 6168 1228 6184 1292
rect 6248 1228 6264 1292
rect 6328 1228 6346 1292
rect 5926 1212 6346 1228
rect 5926 1148 5944 1212
rect 6008 1148 6024 1212
rect 6088 1148 6104 1212
rect 6168 1148 6184 1212
rect 6248 1148 6264 1212
rect 6328 1148 6346 1212
rect 5926 0 6346 1148
rect 6891 20072 7311 20080
rect 6891 20008 6909 20072
rect 6973 20008 6989 20072
rect 7053 20008 7069 20072
rect 7133 20008 7149 20072
rect 7213 20008 7229 20072
rect 7293 20008 7311 20072
rect 6891 19992 7311 20008
rect 6891 19928 6909 19992
rect 6973 19928 6989 19992
rect 7053 19928 7069 19992
rect 7133 19928 7149 19992
rect 7213 19928 7229 19992
rect 7293 19928 7311 19992
rect 6891 19912 7311 19928
rect 6891 19848 6909 19912
rect 6973 19848 6989 19912
rect 7053 19848 7069 19912
rect 7133 19848 7149 19912
rect 7213 19848 7229 19912
rect 7293 19848 7311 19912
rect 6891 19832 7311 19848
rect 6891 19768 6909 19832
rect 6973 19768 6989 19832
rect 7053 19768 7069 19832
rect 7133 19768 7149 19832
rect 7213 19768 7229 19832
rect 7293 19768 7311 19832
rect 6891 19752 7311 19768
rect 6891 19688 6909 19752
rect 6973 19688 6989 19752
rect 7053 19688 7069 19752
rect 7133 19688 7149 19752
rect 7213 19688 7229 19752
rect 7293 19688 7311 19752
rect 6891 19672 7311 19688
rect 6891 19608 6909 19672
rect 6973 19608 6989 19672
rect 7053 19608 7069 19672
rect 7133 19608 7149 19672
rect 7213 19608 7229 19672
rect 7293 19608 7311 19672
rect 6891 19592 7311 19608
rect 6891 19528 6909 19592
rect 6973 19528 6989 19592
rect 7053 19528 7069 19592
rect 7133 19528 7149 19592
rect 7213 19528 7229 19592
rect 7293 19528 7311 19592
rect 6891 19512 7311 19528
rect 6891 19448 6909 19512
rect 6973 19448 6989 19512
rect 7053 19448 7069 19512
rect 7133 19448 7149 19512
rect 7213 19448 7229 19512
rect 7293 19448 7311 19512
rect 6891 19432 7311 19448
rect 6891 19368 6909 19432
rect 6973 19368 6989 19432
rect 7053 19368 7069 19432
rect 7133 19368 7149 19432
rect 7213 19368 7229 19432
rect 7293 19368 7311 19432
rect 6891 19352 7311 19368
rect 6891 19288 6909 19352
rect 6973 19288 6989 19352
rect 7053 19288 7069 19352
rect 7133 19288 7149 19352
rect 7213 19288 7229 19352
rect 7293 19288 7311 19352
rect 6891 16872 7311 19288
rect 6891 16808 6909 16872
rect 6973 16808 6989 16872
rect 7053 16808 7069 16872
rect 7133 16808 7149 16872
rect 7213 16808 7229 16872
rect 7293 16808 7311 16872
rect 6891 15784 7311 16808
rect 6891 15720 6909 15784
rect 6973 15720 6989 15784
rect 7053 15720 7069 15784
rect 7133 15720 7149 15784
rect 7213 15720 7229 15784
rect 7293 15720 7311 15784
rect 6891 14696 7311 15720
rect 6891 14632 6909 14696
rect 6973 14632 6989 14696
rect 7053 14632 7069 14696
rect 7133 14632 7149 14696
rect 7213 14632 7229 14696
rect 7293 14632 7311 14696
rect 6891 13608 7311 14632
rect 6891 13544 6909 13608
rect 6973 13544 6989 13608
rect 7053 13544 7069 13608
rect 7133 13544 7149 13608
rect 7213 13544 7229 13608
rect 7293 13544 7311 13608
rect 6891 12520 7311 13544
rect 6891 12456 6909 12520
rect 6973 12456 6989 12520
rect 7053 12456 7069 12520
rect 7133 12456 7149 12520
rect 7213 12456 7229 12520
rect 7293 12456 7311 12520
rect 6891 11432 7311 12456
rect 6891 11368 6909 11432
rect 6973 11368 6989 11432
rect 7053 11368 7069 11432
rect 7133 11368 7149 11432
rect 7213 11368 7229 11432
rect 7293 11368 7311 11432
rect 6891 10344 7311 11368
rect 6891 10280 6909 10344
rect 6973 10280 6989 10344
rect 7053 10280 7069 10344
rect 7133 10280 7149 10344
rect 7213 10280 7229 10344
rect 7293 10280 7311 10344
rect 6891 9256 7311 10280
rect 6891 9192 6909 9256
rect 6973 9192 6989 9256
rect 7053 9192 7069 9256
rect 7133 9192 7149 9256
rect 7213 9192 7229 9256
rect 7293 9192 7311 9256
rect 6891 8168 7311 9192
rect 6891 8104 6909 8168
rect 6973 8104 6989 8168
rect 7053 8104 7069 8168
rect 7133 8104 7149 8168
rect 7213 8104 7229 8168
rect 7293 8104 7311 8168
rect 6891 7080 7311 8104
rect 6891 7016 6909 7080
rect 6973 7016 6989 7080
rect 7053 7016 7069 7080
rect 7133 7016 7149 7080
rect 7213 7016 7229 7080
rect 7293 7016 7311 7080
rect 6891 5992 7311 7016
rect 6891 5928 6909 5992
rect 6973 5928 6989 5992
rect 7053 5928 7069 5992
rect 7133 5928 7149 5992
rect 7213 5928 7229 5992
rect 7293 5928 7311 5992
rect 6891 4904 7311 5928
rect 6891 4840 6909 4904
rect 6973 4840 6989 4904
rect 7053 4840 7069 4904
rect 7133 4840 7149 4904
rect 7213 4840 7229 4904
rect 7293 4840 7311 4904
rect 6891 3816 7311 4840
rect 6891 3752 6909 3816
rect 6973 3752 6989 3816
rect 7053 3752 7069 3816
rect 7133 3752 7149 3816
rect 7213 3752 7229 3816
rect 7293 3752 7311 3816
rect 6891 792 7311 3752
rect 6891 728 6909 792
rect 6973 728 6989 792
rect 7053 728 7069 792
rect 7133 728 7149 792
rect 7213 728 7229 792
rect 7293 728 7311 792
rect 6891 712 7311 728
rect 6891 648 6909 712
rect 6973 648 6989 712
rect 7053 648 7069 712
rect 7133 648 7149 712
rect 7213 648 7229 712
rect 7293 648 7311 712
rect 6891 632 7311 648
rect 6891 568 6909 632
rect 6973 568 6989 632
rect 7053 568 7069 632
rect 7133 568 7149 632
rect 7213 568 7229 632
rect 7293 568 7311 632
rect 6891 552 7311 568
rect 6891 488 6909 552
rect 6973 488 6989 552
rect 7053 488 7069 552
rect 7133 488 7149 552
rect 7213 488 7229 552
rect 7293 488 7311 552
rect 6891 472 7311 488
rect 6891 408 6909 472
rect 6973 408 6989 472
rect 7053 408 7069 472
rect 7133 408 7149 472
rect 7213 408 7229 472
rect 7293 408 7311 472
rect 6891 392 7311 408
rect 6891 328 6909 392
rect 6973 328 6989 392
rect 7053 328 7069 392
rect 7133 328 7149 392
rect 7213 328 7229 392
rect 7293 328 7311 392
rect 6891 312 7311 328
rect 6891 248 6909 312
rect 6973 248 6989 312
rect 7053 248 7069 312
rect 7133 248 7149 312
rect 7213 248 7229 312
rect 7293 248 7311 312
rect 6891 232 7311 248
rect 6891 168 6909 232
rect 6973 168 6989 232
rect 7053 168 7069 232
rect 7133 168 7149 232
rect 7213 168 7229 232
rect 7293 168 7311 232
rect 6891 152 7311 168
rect 6891 88 6909 152
rect 6973 88 6989 152
rect 7053 88 7069 152
rect 7133 88 7149 152
rect 7213 88 7229 152
rect 7293 88 7311 152
rect 6891 72 7311 88
rect 6891 8 6909 72
rect 6973 8 6989 72
rect 7053 8 7069 72
rect 7133 8 7149 72
rect 7213 8 7229 72
rect 7293 8 7311 72
rect 6891 0 7311 8
rect 7856 18932 8277 20080
rect 11384 20072 12184 20080
rect 11384 20008 11392 20072
rect 11456 20008 11472 20072
rect 11536 20008 11552 20072
rect 11616 20008 11632 20072
rect 11696 20008 11712 20072
rect 11776 20008 11792 20072
rect 11856 20008 11872 20072
rect 11936 20008 11952 20072
rect 12016 20008 12032 20072
rect 12096 20008 12112 20072
rect 12176 20008 12184 20072
rect 11384 19992 12184 20008
rect 11384 19928 11392 19992
rect 11456 19928 11472 19992
rect 11536 19928 11552 19992
rect 11616 19928 11632 19992
rect 11696 19928 11712 19992
rect 11776 19928 11792 19992
rect 11856 19928 11872 19992
rect 11936 19928 11952 19992
rect 12016 19928 12032 19992
rect 12096 19928 12112 19992
rect 12176 19928 12184 19992
rect 11384 19912 12184 19928
rect 11384 19848 11392 19912
rect 11456 19848 11472 19912
rect 11536 19848 11552 19912
rect 11616 19848 11632 19912
rect 11696 19848 11712 19912
rect 11776 19848 11792 19912
rect 11856 19848 11872 19912
rect 11936 19848 11952 19912
rect 12016 19848 12032 19912
rect 12096 19848 12112 19912
rect 12176 19848 12184 19912
rect 11384 19832 12184 19848
rect 11384 19768 11392 19832
rect 11456 19768 11472 19832
rect 11536 19768 11552 19832
rect 11616 19768 11632 19832
rect 11696 19768 11712 19832
rect 11776 19768 11792 19832
rect 11856 19768 11872 19832
rect 11936 19768 11952 19832
rect 12016 19768 12032 19832
rect 12096 19768 12112 19832
rect 12176 19768 12184 19832
rect 11384 19752 12184 19768
rect 11384 19688 11392 19752
rect 11456 19688 11472 19752
rect 11536 19688 11552 19752
rect 11616 19688 11632 19752
rect 11696 19688 11712 19752
rect 11776 19688 11792 19752
rect 11856 19688 11872 19752
rect 11936 19688 11952 19752
rect 12016 19688 12032 19752
rect 12096 19688 12112 19752
rect 12176 19688 12184 19752
rect 11384 19672 12184 19688
rect 11384 19608 11392 19672
rect 11456 19608 11472 19672
rect 11536 19608 11552 19672
rect 11616 19608 11632 19672
rect 11696 19608 11712 19672
rect 11776 19608 11792 19672
rect 11856 19608 11872 19672
rect 11936 19608 11952 19672
rect 12016 19608 12032 19672
rect 12096 19608 12112 19672
rect 12176 19608 12184 19672
rect 11384 19592 12184 19608
rect 11384 19528 11392 19592
rect 11456 19528 11472 19592
rect 11536 19528 11552 19592
rect 11616 19528 11632 19592
rect 11696 19528 11712 19592
rect 11776 19528 11792 19592
rect 11856 19528 11872 19592
rect 11936 19528 11952 19592
rect 12016 19528 12032 19592
rect 12096 19528 12112 19592
rect 12176 19528 12184 19592
rect 11384 19512 12184 19528
rect 11384 19448 11392 19512
rect 11456 19448 11472 19512
rect 11536 19448 11552 19512
rect 11616 19448 11632 19512
rect 11696 19448 11712 19512
rect 11776 19448 11792 19512
rect 11856 19448 11872 19512
rect 11936 19448 11952 19512
rect 12016 19448 12032 19512
rect 12096 19448 12112 19512
rect 12176 19448 12184 19512
rect 11384 19432 12184 19448
rect 11384 19368 11392 19432
rect 11456 19368 11472 19432
rect 11536 19368 11552 19432
rect 11616 19368 11632 19432
rect 11696 19368 11712 19432
rect 11776 19368 11792 19432
rect 11856 19368 11872 19432
rect 11936 19368 11952 19432
rect 12016 19368 12032 19432
rect 12096 19368 12112 19432
rect 12176 19368 12184 19432
rect 11384 19352 12184 19368
rect 11384 19288 11392 19352
rect 11456 19288 11472 19352
rect 11536 19288 11552 19352
rect 11616 19288 11632 19352
rect 11696 19288 11712 19352
rect 11776 19288 11792 19352
rect 11856 19288 11872 19352
rect 11936 19288 11952 19352
rect 12016 19288 12032 19352
rect 12096 19288 12112 19352
rect 12176 19288 12184 19352
rect 7856 18868 7874 18932
rect 7938 18868 7954 18932
rect 8018 18868 8034 18932
rect 8098 18868 8114 18932
rect 8178 18868 8194 18932
rect 8258 18868 8277 18932
rect 7856 18852 8277 18868
rect 7856 18788 7874 18852
rect 7938 18788 7954 18852
rect 8018 18788 8034 18852
rect 8098 18788 8114 18852
rect 8178 18788 8194 18852
rect 8258 18788 8277 18852
rect 7856 18772 8277 18788
rect 7856 18708 7874 18772
rect 7938 18708 7954 18772
rect 8018 18708 8034 18772
rect 8098 18708 8114 18772
rect 8178 18708 8194 18772
rect 8258 18708 8277 18772
rect 7856 18692 8277 18708
rect 7856 18628 7874 18692
rect 7938 18628 7954 18692
rect 8018 18628 8034 18692
rect 8098 18628 8114 18692
rect 8178 18628 8194 18692
rect 8258 18628 8277 18692
rect 7856 18612 8277 18628
rect 7856 18548 7874 18612
rect 7938 18548 7954 18612
rect 8018 18548 8034 18612
rect 8098 18548 8114 18612
rect 8178 18548 8194 18612
rect 8258 18548 8277 18612
rect 7856 18532 8277 18548
rect 7856 18468 7874 18532
rect 7938 18468 7954 18532
rect 8018 18468 8034 18532
rect 8098 18468 8114 18532
rect 8178 18468 8194 18532
rect 8258 18468 8277 18532
rect 7856 18452 8277 18468
rect 7856 18388 7874 18452
rect 7938 18388 7954 18452
rect 8018 18388 8034 18452
rect 8098 18388 8114 18452
rect 8178 18388 8194 18452
rect 8258 18388 8277 18452
rect 7856 18372 8277 18388
rect 7856 18308 7874 18372
rect 7938 18308 7954 18372
rect 8018 18308 8034 18372
rect 8098 18308 8114 18372
rect 8178 18308 8194 18372
rect 8258 18308 8277 18372
rect 7856 18292 8277 18308
rect 7856 18228 7874 18292
rect 7938 18228 7954 18292
rect 8018 18228 8034 18292
rect 8098 18228 8114 18292
rect 8178 18228 8194 18292
rect 8258 18228 8277 18292
rect 7856 18212 8277 18228
rect 7856 18148 7874 18212
rect 7938 18148 7954 18212
rect 8018 18148 8034 18212
rect 8098 18148 8114 18212
rect 8178 18148 8194 18212
rect 8258 18148 8277 18212
rect 7856 16328 8277 18148
rect 7856 16264 7874 16328
rect 7938 16264 7954 16328
rect 8018 16264 8034 16328
rect 8098 16264 8114 16328
rect 8178 16264 8194 16328
rect 8258 16264 8277 16328
rect 7856 15240 8277 16264
rect 7856 15176 7874 15240
rect 7938 15176 7954 15240
rect 8018 15176 8034 15240
rect 8098 15176 8114 15240
rect 8178 15176 8194 15240
rect 8258 15176 8277 15240
rect 7856 14152 8277 15176
rect 7856 14088 7874 14152
rect 7938 14088 7954 14152
rect 8018 14088 8034 14152
rect 8098 14088 8114 14152
rect 8178 14088 8194 14152
rect 8258 14088 8277 14152
rect 7856 13064 8277 14088
rect 7856 13000 7874 13064
rect 7938 13000 7954 13064
rect 8018 13000 8034 13064
rect 8098 13000 8114 13064
rect 8178 13000 8194 13064
rect 8258 13000 8277 13064
rect 7856 11976 8277 13000
rect 7856 11912 7874 11976
rect 7938 11912 7954 11976
rect 8018 11912 8034 11976
rect 8098 11912 8114 11976
rect 8178 11912 8194 11976
rect 8258 11912 8277 11976
rect 7856 10888 8277 11912
rect 7856 10824 7874 10888
rect 7938 10824 7954 10888
rect 8018 10824 8034 10888
rect 8098 10824 8114 10888
rect 8178 10824 8194 10888
rect 8258 10824 8277 10888
rect 7856 9800 8277 10824
rect 7856 9736 7874 9800
rect 7938 9736 7954 9800
rect 8018 9736 8034 9800
rect 8098 9736 8114 9800
rect 8178 9736 8194 9800
rect 8258 9736 8277 9800
rect 7856 8712 8277 9736
rect 7856 8648 7874 8712
rect 7938 8648 7954 8712
rect 8018 8648 8034 8712
rect 8098 8648 8114 8712
rect 8178 8648 8194 8712
rect 8258 8648 8277 8712
rect 7856 7624 8277 8648
rect 7856 7560 7874 7624
rect 7938 7560 7954 7624
rect 8018 7560 8034 7624
rect 8098 7560 8114 7624
rect 8178 7560 8194 7624
rect 8258 7560 8277 7624
rect 7856 6536 8277 7560
rect 7856 6472 7874 6536
rect 7938 6472 7954 6536
rect 8018 6472 8034 6536
rect 8098 6472 8114 6536
rect 8178 6472 8194 6536
rect 8258 6472 8277 6536
rect 7856 5448 8277 6472
rect 7856 5384 7874 5448
rect 7938 5384 7954 5448
rect 8018 5384 8034 5448
rect 8098 5384 8114 5448
rect 8178 5384 8194 5448
rect 8258 5384 8277 5448
rect 7856 4360 8277 5384
rect 7856 4296 7874 4360
rect 7938 4296 7954 4360
rect 8018 4296 8034 4360
rect 8098 4296 8114 4360
rect 8178 4296 8194 4360
rect 8258 4296 8277 4360
rect 7856 3272 8277 4296
rect 7856 3208 7874 3272
rect 7938 3208 7954 3272
rect 8018 3208 8034 3272
rect 8098 3208 8114 3272
rect 8178 3208 8194 3272
rect 8258 3208 8277 3272
rect 7856 1932 8277 3208
rect 7856 1868 7874 1932
rect 7938 1868 7954 1932
rect 8018 1868 8034 1932
rect 8098 1868 8114 1932
rect 8178 1868 8194 1932
rect 8258 1868 8277 1932
rect 7856 1852 8277 1868
rect 7856 1788 7874 1852
rect 7938 1788 7954 1852
rect 8018 1788 8034 1852
rect 8098 1788 8114 1852
rect 8178 1788 8194 1852
rect 8258 1788 8277 1852
rect 7856 1772 8277 1788
rect 7856 1708 7874 1772
rect 7938 1708 7954 1772
rect 8018 1708 8034 1772
rect 8098 1708 8114 1772
rect 8178 1708 8194 1772
rect 8258 1708 8277 1772
rect 7856 1692 8277 1708
rect 7856 1628 7874 1692
rect 7938 1628 7954 1692
rect 8018 1628 8034 1692
rect 8098 1628 8114 1692
rect 8178 1628 8194 1692
rect 8258 1628 8277 1692
rect 7856 1612 8277 1628
rect 7856 1548 7874 1612
rect 7938 1548 7954 1612
rect 8018 1548 8034 1612
rect 8098 1548 8114 1612
rect 8178 1548 8194 1612
rect 8258 1548 8277 1612
rect 7856 1532 8277 1548
rect 7856 1468 7874 1532
rect 7938 1468 7954 1532
rect 8018 1468 8034 1532
rect 8098 1468 8114 1532
rect 8178 1468 8194 1532
rect 8258 1468 8277 1532
rect 7856 1452 8277 1468
rect 7856 1388 7874 1452
rect 7938 1388 7954 1452
rect 8018 1388 8034 1452
rect 8098 1388 8114 1452
rect 8178 1388 8194 1452
rect 8258 1388 8277 1452
rect 7856 1372 8277 1388
rect 7856 1308 7874 1372
rect 7938 1308 7954 1372
rect 8018 1308 8034 1372
rect 8098 1308 8114 1372
rect 8178 1308 8194 1372
rect 8258 1308 8277 1372
rect 7856 1292 8277 1308
rect 7856 1228 7874 1292
rect 7938 1228 7954 1292
rect 8018 1228 8034 1292
rect 8098 1228 8114 1292
rect 8178 1228 8194 1292
rect 8258 1228 8277 1292
rect 7856 1212 8277 1228
rect 7856 1148 7874 1212
rect 7938 1148 7954 1212
rect 8018 1148 8034 1212
rect 8098 1148 8114 1212
rect 8178 1148 8194 1212
rect 8258 1148 8277 1212
rect 7856 0 8277 1148
rect 10244 18932 11044 18940
rect 10244 18868 10252 18932
rect 10316 18868 10332 18932
rect 10396 18868 10412 18932
rect 10476 18868 10492 18932
rect 10556 18868 10572 18932
rect 10636 18868 10652 18932
rect 10716 18868 10732 18932
rect 10796 18868 10812 18932
rect 10876 18868 10892 18932
rect 10956 18868 10972 18932
rect 11036 18868 11044 18932
rect 10244 18852 11044 18868
rect 10244 18788 10252 18852
rect 10316 18788 10332 18852
rect 10396 18788 10412 18852
rect 10476 18788 10492 18852
rect 10556 18788 10572 18852
rect 10636 18788 10652 18852
rect 10716 18788 10732 18852
rect 10796 18788 10812 18852
rect 10876 18788 10892 18852
rect 10956 18788 10972 18852
rect 11036 18788 11044 18852
rect 10244 18772 11044 18788
rect 10244 18708 10252 18772
rect 10316 18708 10332 18772
rect 10396 18708 10412 18772
rect 10476 18708 10492 18772
rect 10556 18708 10572 18772
rect 10636 18708 10652 18772
rect 10716 18708 10732 18772
rect 10796 18708 10812 18772
rect 10876 18708 10892 18772
rect 10956 18708 10972 18772
rect 11036 18708 11044 18772
rect 10244 18692 11044 18708
rect 10244 18628 10252 18692
rect 10316 18628 10332 18692
rect 10396 18628 10412 18692
rect 10476 18628 10492 18692
rect 10556 18628 10572 18692
rect 10636 18628 10652 18692
rect 10716 18628 10732 18692
rect 10796 18628 10812 18692
rect 10876 18628 10892 18692
rect 10956 18628 10972 18692
rect 11036 18628 11044 18692
rect 10244 18612 11044 18628
rect 10244 18548 10252 18612
rect 10316 18548 10332 18612
rect 10396 18548 10412 18612
rect 10476 18548 10492 18612
rect 10556 18548 10572 18612
rect 10636 18548 10652 18612
rect 10716 18548 10732 18612
rect 10796 18548 10812 18612
rect 10876 18548 10892 18612
rect 10956 18548 10972 18612
rect 11036 18548 11044 18612
rect 10244 18532 11044 18548
rect 10244 18468 10252 18532
rect 10316 18468 10332 18532
rect 10396 18468 10412 18532
rect 10476 18468 10492 18532
rect 10556 18468 10572 18532
rect 10636 18468 10652 18532
rect 10716 18468 10732 18532
rect 10796 18468 10812 18532
rect 10876 18468 10892 18532
rect 10956 18468 10972 18532
rect 11036 18468 11044 18532
rect 10244 18452 11044 18468
rect 10244 18388 10252 18452
rect 10316 18388 10332 18452
rect 10396 18388 10412 18452
rect 10476 18388 10492 18452
rect 10556 18388 10572 18452
rect 10636 18388 10652 18452
rect 10716 18388 10732 18452
rect 10796 18388 10812 18452
rect 10876 18388 10892 18452
rect 10956 18388 10972 18452
rect 11036 18388 11044 18452
rect 10244 18372 11044 18388
rect 10244 18308 10252 18372
rect 10316 18308 10332 18372
rect 10396 18308 10412 18372
rect 10476 18308 10492 18372
rect 10556 18308 10572 18372
rect 10636 18308 10652 18372
rect 10716 18308 10732 18372
rect 10796 18308 10812 18372
rect 10876 18308 10892 18372
rect 10956 18308 10972 18372
rect 11036 18308 11044 18372
rect 10244 18292 11044 18308
rect 10244 18228 10252 18292
rect 10316 18228 10332 18292
rect 10396 18228 10412 18292
rect 10476 18228 10492 18292
rect 10556 18228 10572 18292
rect 10636 18228 10652 18292
rect 10716 18228 10732 18292
rect 10796 18228 10812 18292
rect 10876 18228 10892 18292
rect 10956 18228 10972 18292
rect 11036 18228 11044 18292
rect 10244 18212 11044 18228
rect 10244 18148 10252 18212
rect 10316 18148 10332 18212
rect 10396 18148 10412 18212
rect 10476 18148 10492 18212
rect 10556 18148 10572 18212
rect 10636 18148 10652 18212
rect 10716 18148 10732 18212
rect 10796 18148 10812 18212
rect 10876 18148 10892 18212
rect 10956 18148 10972 18212
rect 11036 18148 11044 18212
rect 10244 1932 11044 18148
rect 10244 1868 10252 1932
rect 10316 1868 10332 1932
rect 10396 1868 10412 1932
rect 10476 1868 10492 1932
rect 10556 1868 10572 1932
rect 10636 1868 10652 1932
rect 10716 1868 10732 1932
rect 10796 1868 10812 1932
rect 10876 1868 10892 1932
rect 10956 1868 10972 1932
rect 11036 1868 11044 1932
rect 10244 1852 11044 1868
rect 10244 1788 10252 1852
rect 10316 1788 10332 1852
rect 10396 1788 10412 1852
rect 10476 1788 10492 1852
rect 10556 1788 10572 1852
rect 10636 1788 10652 1852
rect 10716 1788 10732 1852
rect 10796 1788 10812 1852
rect 10876 1788 10892 1852
rect 10956 1788 10972 1852
rect 11036 1788 11044 1852
rect 10244 1772 11044 1788
rect 10244 1708 10252 1772
rect 10316 1708 10332 1772
rect 10396 1708 10412 1772
rect 10476 1708 10492 1772
rect 10556 1708 10572 1772
rect 10636 1708 10652 1772
rect 10716 1708 10732 1772
rect 10796 1708 10812 1772
rect 10876 1708 10892 1772
rect 10956 1708 10972 1772
rect 11036 1708 11044 1772
rect 10244 1692 11044 1708
rect 10244 1628 10252 1692
rect 10316 1628 10332 1692
rect 10396 1628 10412 1692
rect 10476 1628 10492 1692
rect 10556 1628 10572 1692
rect 10636 1628 10652 1692
rect 10716 1628 10732 1692
rect 10796 1628 10812 1692
rect 10876 1628 10892 1692
rect 10956 1628 10972 1692
rect 11036 1628 11044 1692
rect 10244 1612 11044 1628
rect 10244 1548 10252 1612
rect 10316 1548 10332 1612
rect 10396 1548 10412 1612
rect 10476 1548 10492 1612
rect 10556 1548 10572 1612
rect 10636 1548 10652 1612
rect 10716 1548 10732 1612
rect 10796 1548 10812 1612
rect 10876 1548 10892 1612
rect 10956 1548 10972 1612
rect 11036 1548 11044 1612
rect 10244 1532 11044 1548
rect 10244 1468 10252 1532
rect 10316 1468 10332 1532
rect 10396 1468 10412 1532
rect 10476 1468 10492 1532
rect 10556 1468 10572 1532
rect 10636 1468 10652 1532
rect 10716 1468 10732 1532
rect 10796 1468 10812 1532
rect 10876 1468 10892 1532
rect 10956 1468 10972 1532
rect 11036 1468 11044 1532
rect 10244 1452 11044 1468
rect 10244 1388 10252 1452
rect 10316 1388 10332 1452
rect 10396 1388 10412 1452
rect 10476 1388 10492 1452
rect 10556 1388 10572 1452
rect 10636 1388 10652 1452
rect 10716 1388 10732 1452
rect 10796 1388 10812 1452
rect 10876 1388 10892 1452
rect 10956 1388 10972 1452
rect 11036 1388 11044 1452
rect 10244 1372 11044 1388
rect 10244 1308 10252 1372
rect 10316 1308 10332 1372
rect 10396 1308 10412 1372
rect 10476 1308 10492 1372
rect 10556 1308 10572 1372
rect 10636 1308 10652 1372
rect 10716 1308 10732 1372
rect 10796 1308 10812 1372
rect 10876 1308 10892 1372
rect 10956 1308 10972 1372
rect 11036 1308 11044 1372
rect 10244 1292 11044 1308
rect 10244 1228 10252 1292
rect 10316 1228 10332 1292
rect 10396 1228 10412 1292
rect 10476 1228 10492 1292
rect 10556 1228 10572 1292
rect 10636 1228 10652 1292
rect 10716 1228 10732 1292
rect 10796 1228 10812 1292
rect 10876 1228 10892 1292
rect 10956 1228 10972 1292
rect 11036 1228 11044 1292
rect 10244 1212 11044 1228
rect 10244 1148 10252 1212
rect 10316 1148 10332 1212
rect 10396 1148 10412 1212
rect 10476 1148 10492 1212
rect 10556 1148 10572 1212
rect 10636 1148 10652 1212
rect 10716 1148 10732 1212
rect 10796 1148 10812 1212
rect 10876 1148 10892 1212
rect 10956 1148 10972 1212
rect 11036 1148 11044 1212
rect 10244 1140 11044 1148
rect 11384 792 12184 19288
rect 11384 728 11392 792
rect 11456 728 11472 792
rect 11536 728 11552 792
rect 11616 728 11632 792
rect 11696 728 11712 792
rect 11776 728 11792 792
rect 11856 728 11872 792
rect 11936 728 11952 792
rect 12016 728 12032 792
rect 12096 728 12112 792
rect 12176 728 12184 792
rect 11384 712 12184 728
rect 11384 648 11392 712
rect 11456 648 11472 712
rect 11536 648 11552 712
rect 11616 648 11632 712
rect 11696 648 11712 712
rect 11776 648 11792 712
rect 11856 648 11872 712
rect 11936 648 11952 712
rect 12016 648 12032 712
rect 12096 648 12112 712
rect 12176 648 12184 712
rect 11384 632 12184 648
rect 11384 568 11392 632
rect 11456 568 11472 632
rect 11536 568 11552 632
rect 11616 568 11632 632
rect 11696 568 11712 632
rect 11776 568 11792 632
rect 11856 568 11872 632
rect 11936 568 11952 632
rect 12016 568 12032 632
rect 12096 568 12112 632
rect 12176 568 12184 632
rect 11384 552 12184 568
rect 11384 488 11392 552
rect 11456 488 11472 552
rect 11536 488 11552 552
rect 11616 488 11632 552
rect 11696 488 11712 552
rect 11776 488 11792 552
rect 11856 488 11872 552
rect 11936 488 11952 552
rect 12016 488 12032 552
rect 12096 488 12112 552
rect 12176 488 12184 552
rect 11384 472 12184 488
rect 11384 408 11392 472
rect 11456 408 11472 472
rect 11536 408 11552 472
rect 11616 408 11632 472
rect 11696 408 11712 472
rect 11776 408 11792 472
rect 11856 408 11872 472
rect 11936 408 11952 472
rect 12016 408 12032 472
rect 12096 408 12112 472
rect 12176 408 12184 472
rect 11384 392 12184 408
rect 11384 328 11392 392
rect 11456 328 11472 392
rect 11536 328 11552 392
rect 11616 328 11632 392
rect 11696 328 11712 392
rect 11776 328 11792 392
rect 11856 328 11872 392
rect 11936 328 11952 392
rect 12016 328 12032 392
rect 12096 328 12112 392
rect 12176 328 12184 392
rect 11384 312 12184 328
rect 11384 248 11392 312
rect 11456 248 11472 312
rect 11536 248 11552 312
rect 11616 248 11632 312
rect 11696 248 11712 312
rect 11776 248 11792 312
rect 11856 248 11872 312
rect 11936 248 11952 312
rect 12016 248 12032 312
rect 12096 248 12112 312
rect 12176 248 12184 312
rect 11384 232 12184 248
rect 11384 168 11392 232
rect 11456 168 11472 232
rect 11536 168 11552 232
rect 11616 168 11632 232
rect 11696 168 11712 232
rect 11776 168 11792 232
rect 11856 168 11872 232
rect 11936 168 11952 232
rect 12016 168 12032 232
rect 12096 168 12112 232
rect 12176 168 12184 232
rect 11384 152 12184 168
rect 11384 88 11392 152
rect 11456 88 11472 152
rect 11536 88 11552 152
rect 11616 88 11632 152
rect 11696 88 11712 152
rect 11776 88 11792 152
rect 11856 88 11872 152
rect 11936 88 11952 152
rect 12016 88 12032 152
rect 12096 88 12112 152
rect 12176 88 12184 152
rect 11384 72 12184 88
rect 11384 8 11392 72
rect 11456 8 11472 72
rect 11536 8 11552 72
rect 11616 8 11632 72
rect 11696 8 11712 72
rect 11776 8 11792 72
rect 11856 8 11872 72
rect 11936 8 11952 72
rect 12016 8 12032 72
rect 12096 8 12112 72
rect 12176 8 12184 72
rect 11384 0 12184 8
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3516 0 1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1624635492
transform 1 0 3516 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3240 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 3240 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1624635492
transform 1 0 4620 0 1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1624635492
transform 1 0 4620 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1624635492
transform 1 0 5724 0 1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1624635492
transform 1 0 6000 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5724 0 -1 3784
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5908 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7932 0 1 3784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1624635492
transform 1 0 6828 0 1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1624635492
transform 1 0 7104 0 -1 3784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8576 0 1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8208 0 -1 3784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1624635492
transform 1 0 8484 0 1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1624635492
transform 1 0 8576 0 -1 3784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 8944 0 1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 8944 0 -1 3784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 3516 0 -1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 3240 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1624635492
transform 1 0 4620 0 -1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 6000 0 -1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1624635492
transform 1 0 5724 0 -1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1624635492
transform 1 0 5908 0 -1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1624635492
transform 1 0 7656 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_42
timestamp 1624635492
transform 1 0 7104 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7656 0 -1 4872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1624635492
transform 1 0 8300 0 -1 4872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8300 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 8944 0 -1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 3516 0 1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 3240 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1624635492
transform 1 0 4620 0 1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1624635492
transform 1 0 5724 0 1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1624635492
transform 1 0 7932 0 1 4872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1624635492
transform 1 0 6828 0 1 4872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1624635492
transform 1 0 8576 0 1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1624635492
transform 1 0 8484 0 1 4872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 8944 0 1 4872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 3516 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 3240 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 4620 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 6000 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 5724 0 -1 5960
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1624635492
transform 1 0 5908 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 7104 0 -1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1624635492
transform 1 0 8576 0 -1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1624635492
transform 1 0 8208 0 -1 5960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 8944 0 -1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624635492
transform 1 0 3516 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 3240 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624635492
transform 1 0 4620 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1624635492
transform 1 0 5724 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1624635492
transform 1 0 7932 0 1 5960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1624635492
transform 1 0 6828 0 1 5960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1624635492
transform 1 0 8576 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1624635492
transform 1 0 8484 0 1 5960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 8944 0 1 5960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 3516 0 1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624635492
transform 1 0 3516 0 -1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 3240 0 1 7048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 3240 0 -1 7048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 4620 0 1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624635492
transform 1 0 4620 0 -1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624635492
transform 1 0 5724 0 1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 6000 0 -1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 5724 0 -1 7048
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 5908 0 -1 7048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1624635492
transform 1 0 7932 0 1 7048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1624635492
transform 1 0 6828 0 1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624635492
transform 1 0 7104 0 -1 7048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1624635492
transform 1 0 8576 0 1 7048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_58
timestamp 1624635492
transform 1 0 8576 0 -1 7048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_54
timestamp 1624635492
transform 1 0 8208 0 -1 7048
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 8484 0 1 7048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 8944 0 1 7048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 8944 0 -1 7048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 3516 0 -1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 3240 0 -1 8136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 4620 0 -1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624635492
transform 1 0 6000 0 -1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 5724 0 -1 8136
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 5908 0 -1 8136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624635492
transform 1 0 7104 0 -1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_58
timestamp 1624635492
transform 1 0 8576 0 -1 8136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1624635492
transform 1 0 8208 0 -1 8136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 8944 0 -1 8136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 3516 0 1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 3240 0 1 8136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 4620 0 1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624635492
transform 1 0 5724 0 1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1624635492
transform 1 0 7932 0 1 8136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1624635492
transform 1 0 6828 0 1 8136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_58
timestamp 1624635492
transform 1 0 8576 0 1 8136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 8484 0 1 8136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 8944 0 1 8136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 3516 0 -1 9224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 3240 0 -1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 4620 0 -1 9224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_35
timestamp 1624635492
transform 1 0 6460 0 -1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_30
timestamp 1624635492
transform 1 0 6000 0 -1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 5724 0 -1 9224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x15_A
timestamp 1624635492
transform 1 0 6276 0 -1 9224
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 5908 0 -1 9224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1624635492
transform 1 0 7656 0 -1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_42
timestamp 1624635492
transform 1 0 7104 0 -1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 7656 0 -1 9224
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6828 0 -1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1624635492
transform 1 0 8300 0 -1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform -1 0 8300 0 -1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 8944 0 -1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624635492
transform 1 0 3516 0 1 9224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 3240 0 1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624635492
transform 1 0 4620 0 1 9224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1624635492
transform 1 0 6460 0 1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_27
timestamp 1624635492
transform 1 0 5724 0 1 9224
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x6_B1
timestamp 1624635492
transform 1 0 6276 0 1 9224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_46
timestamp 1624635492
transform 1 0 7472 0 1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6828 0 1 9224
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1624635492
transform 1 0 7840 0 1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_58
timestamp 1624635492
transform 1 0 8576 0 1 9224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_53
timestamp 1624635492
transform 1 0 8116 0 1 9224
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 8484 0 1 9224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 8944 0 1 9224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_12
timestamp 1624635492
transform 1 0 4344 0 -1 10312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1624635492
transform 1 0 3792 0 -1 10312
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 4344 0 -1 10312
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3792 0 -1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 3240 0 -1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1624635492
transform 1 0 5448 0 -1 10312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1624635492
transform 1 0 6736 0 -1 10312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_34
timestamp 1624635492
transform 1 0 6368 0 -1 10312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_30
timestamp 1624635492
transform 1 0 6000 0 -1 10312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1624635492
transform 1 0 5816 0 -1 10312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 5908 0 -1 10312
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1624635492
transform 1 0 6460 0 -1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7748 0 -1 10312
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7104 0 -1 10312
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1624635492
transform 1 0 8484 0 -1 10312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 8944 0 -1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624635492
transform 1 0 3516 0 -1 11400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 3516 0 1 10312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 3240 0 -1 11400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 3240 0 1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624635492
transform 1 0 4620 0 -1 11400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 4620 0 1 10312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_35
timestamp 1624635492
transform 1 0 6460 0 -1 11400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_30
timestamp 1624635492
transform 1 0 6000 0 -1 11400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 5724 0 -1 11400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624635492
transform 1 0 5724 0 1 10312
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x9_B1
timestamp 1624635492
transform 1 0 6276 0 -1 11400
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 5908 0 -1 11400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1624635492
transform 1 0 7472 0 -1 11400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_49
timestamp 1624635492
transform 1 0 7748 0 1 10312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_39
timestamp 1624635492
transform 1 0 6828 0 1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  x9
timestamp 1624635492
transform 1 0 6828 0 -1 11400
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  x8
timestamp 1624635492
transform 1 0 7104 0 1 10312
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  x10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7840 0 -1 11400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1624635492
transform 1 0 8576 0 -1 11400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1624635492
transform 1 0 8208 0 -1 11400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_58
timestamp 1624635492
transform 1 0 8576 0 1 10312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 8484 0 1 10312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 8944 0 -1 11400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 8944 0 1 10312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 3516 0 1 11400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 3240 0 1 11400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624635492
transform 1 0 4620 0 1 11400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624635492
transform 1 0 5724 0 1 11400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_49
timestamp 1624635492
transform 1 0 7748 0 1 11400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1624635492
transform 1 0 6828 0 1 11400
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  x11
timestamp 1624635492
transform 1 0 7380 0 1 11400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_58
timestamp 1624635492
transform 1 0 8576 0 1 11400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 8484 0 1 11400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 8944 0 1 11400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624635492
transform 1 0 3516 0 -1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 3240 0 -1 12488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624635492
transform 1 0 4620 0 -1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 6000 0 -1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 5724 0 -1 12488
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 5908 0 -1 12488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 7104 0 -1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1624635492
transform 1 0 8576 0 -1 12488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1624635492
transform 1 0 8208 0 -1 12488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 8944 0 -1 12488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1624635492
transform 1 0 3516 0 1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 3240 0 1 12488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1624635492
transform 1 0 4620 0 1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1624635492
transform 1 0 5724 0 1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1624635492
transform 1 0 7932 0 1 12488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1624635492
transform 1 0 6828 0 1 12488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_58
timestamp 1624635492
transform 1 0 8576 0 1 12488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 8484 0 1 12488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 8944 0 1 12488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 3516 0 -1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 3240 0 -1 13576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624635492
transform 1 0 4620 0 -1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1624635492
transform 1 0 6000 0 -1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624635492
transform 1 0 5724 0 -1 13576
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 5908 0 -1 13576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1624635492
transform 1 0 7104 0 -1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1624635492
transform 1 0 8576 0 -1 13576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1624635492
transform 1 0 8208 0 -1 13576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 8944 0 -1 13576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624635492
transform 1 0 3516 0 -1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624635492
transform 1 0 3516 0 1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 3240 0 -1 14664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 3240 0 1 13576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1624635492
transform 1 0 4620 0 -1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1624635492
transform 1 0 4620 0 1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1624635492
transform 1 0 6000 0 -1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1624635492
transform 1 0 5724 0 -1 14664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1624635492
transform 1 0 5724 0 1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 5908 0 -1 14664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1624635492
transform 1 0 7104 0 -1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1624635492
transform 1 0 7932 0 1 13576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1624635492
transform 1 0 6828 0 1 13576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_58
timestamp 1624635492
transform 1 0 8576 0 -1 14664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_54
timestamp 1624635492
transform 1 0 8208 0 -1 14664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_58
timestamp 1624635492
transform 1 0 8576 0 1 13576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 8484 0 1 13576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 8944 0 -1 14664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 8944 0 1 13576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 3516 0 1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 3240 0 1 14664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624635492
transform 1 0 4620 0 1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1624635492
transform 1 0 5724 0 1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1624635492
transform 1 0 7932 0 1 14664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1624635492
transform 1 0 6828 0 1 14664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_58
timestamp 1624635492
transform 1 0 8576 0 1 14664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 8484 0 1 14664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 8944 0 1 14664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624635492
transform 1 0 3516 0 -1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 3240 0 -1 15752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1624635492
transform 1 0 4620 0 -1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1624635492
transform 1 0 6000 0 -1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 5724 0 -1 15752
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 5908 0 -1 15752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1624635492
transform 1 0 7104 0 -1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_58
timestamp 1624635492
transform 1 0 8576 0 -1 15752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_54
timestamp 1624635492
transform 1 0 8208 0 -1 15752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 8944 0 -1 15752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_12
timestamp 1624635492
transform 1 0 4344 0 1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_6
timestamp 1624635492
transform 1 0 3792 0 1 15752
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 4344 0 1 15752
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 3516 0 1 15752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 3240 0 1 15752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_24
timestamp 1624635492
transform 1 0 5448 0 1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1624635492
transform 1 0 6552 0 1 15752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_48
timestamp 1624635492
transform 1 0 7656 0 1 15752
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1624635492
transform 1 0 7840 0 1 15752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_58
timestamp 1624635492
transform 1 0 8576 0 1 15752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1624635492
transform 1 0 8116 0 1 15752
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 8484 0 1 15752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 8944 0 1 15752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1624635492
transform 1 0 3516 0 -1 16840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 3240 0 -1 16840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1624635492
transform 1 0 4620 0 -1 16840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1624635492
transform 1 0 6000 0 -1 16840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624635492
transform 1 0 5724 0 -1 16840
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 5908 0 -1 16840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1624635492
transform 1 0 7104 0 -1 16840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1624635492
transform 1 0 8208 0 -1 16840
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 8576 0 -1 16840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 8944 0 -1 16840
box -38 -48 314 592
<< labels >>
rlabel metal2 s 9336 9922 10136 10146 6 INN
port 0 nsew signal input
rlabel metal2 s 9336 3942 10136 4166 6 INP
port 1 nsew signal input
rlabel metal2 s 9336 15902 10136 16126 6 Q
port 2 nsew signal tristate
rlabel metal2 s 2136 15902 2936 16126 6 VDD
port 3 nsew signal input
rlabel metal2 s 2136 9922 2936 10146 6 VSS
port 4 nsew signal input
rlabel metal2 s 2136 3942 2936 4166 6 clk
port 5 nsew signal input
rlabel metal3 s 1140 18140 11044 18940 6 vccd2
port 6 nsew power bidirectional
rlabel metal3 s 1140 1140 11044 1940 6 vccd2
port 7 nsew power bidirectional
rlabel metal4 s 7857 0 8277 20080 6 vccd2
port 8 nsew power bidirectional
rlabel metal4 s 5926 0 6346 20080 6 vccd2
port 9 nsew power bidirectional
rlabel metal4 s 3995 0 4415 20080 6 vccd2
port 10 nsew power bidirectional
rlabel metal4 s 10244 1140 11044 18940 6 vccd2
port 11 nsew power bidirectional
rlabel metal4 s 1140 1140 1940 18940 4 vccd2
port 12 nsew power bidirectional
rlabel metal3 s 0 19280 12184 20080 6 vssd2
port 13 nsew ground bidirectional
rlabel metal3 s 0 0 12184 800 8 vssd2
port 14 nsew ground bidirectional
rlabel metal4 s 11384 0 12184 20080 6 vssd2
port 15 nsew ground bidirectional
rlabel metal4 s 6891 0 7311 20080 6 vssd2
port 16 nsew ground bidirectional
rlabel metal4 s 4961 0 5381 20080 6 vssd2
port 17 nsew ground bidirectional
rlabel metal4 s 0 0 800 20080 4 vssd2
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12184 20080
<< end >>
