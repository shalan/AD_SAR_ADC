magic
tech sky130A
magscale 1 2
timestamp 1626642740
<< obsli1 >>
rect 3240 3223 8944 16857
<< obsm1 >>
rect 3162 3192 9206 16888
<< metal2 >>
rect 2136 15902 2936 16126
rect 9336 15902 10136 16126
rect 2136 9922 2936 10146
rect 9336 9922 10136 10146
rect 2136 3942 2936 4166
rect 9336 3942 10136 4166
<< obsm2 >>
rect 2936 16182 9336 16888
rect 2992 15846 9280 16182
rect 2936 10202 9336 15846
rect 2992 9866 9280 10202
rect 2936 4222 9336 9866
rect 2992 3886 9280 4222
rect 2936 3192 9336 3886
<< metal3 >>
rect 0 19280 12184 20080
rect 1140 18140 11044 18940
rect 1140 1140 11044 1940
rect 0 0 12184 800
<< obsm3 >>
rect 3995 3207 8276 16873
<< metal4 >>
rect 0 0 800 20080
rect 1140 1140 1940 18940
rect 3995 0 4415 20080
rect 4961 0 5381 20080
rect 5926 0 6346 20080
rect 6891 0 7311 20080
rect 7857 0 8277 20080
rect 10244 1140 11044 18940
rect 11384 0 12184 20080
<< obsm4 >>
rect 5461 0 5846 20080
rect 6426 0 6811 20080
rect 7391 0 7777 20080
<< labels >>
rlabel metal2 s 9336 9922 10136 10146 6 INN
port 1 nsew signal input
rlabel metal2 s 9336 3942 10136 4166 6 INP
port 2 nsew signal input
rlabel metal2 s 9336 15902 10136 16126 6 Q
port 3 nsew signal output
rlabel metal2 s 2136 15902 2936 16126 6 VDD
port 4 nsew signal input
rlabel metal2 s 2136 9922 2936 10146 6 VSS
port 5 nsew signal input
rlabel metal2 s 2136 3942 2936 4166 6 clk
port 6 nsew signal input
rlabel metal3 s 1140 18140 11044 18940 6 vccd2
port 7 nsew power bidirectional
rlabel metal3 s 1140 1140 11044 1940 6 vccd2
port 8 nsew power bidirectional
rlabel metal4 s 7857 0 8277 20080 6 vccd2
port 9 nsew power bidirectional
rlabel metal4 s 5926 0 6346 20080 6 vccd2
port 10 nsew power bidirectional
rlabel metal4 s 3995 0 4415 20080 6 vccd2
port 11 nsew power bidirectional
rlabel metal4 s 10244 1140 11044 18940 6 vccd2
port 12 nsew power bidirectional
rlabel metal4 s 1140 1140 1940 18940 6 vccd2
port 13 nsew power bidirectional
rlabel metal3 s 0 19280 12184 20080 6 vssd2
port 14 nsew ground bidirectional
rlabel metal3 s 0 0 12184 800 6 vssd2
port 15 nsew ground bidirectional
rlabel metal4 s 11384 0 12184 20080 6 vssd2
port 16 nsew ground bidirectional
rlabel metal4 s 6891 0 7311 20080 6 vssd2
port 17 nsew ground bidirectional
rlabel metal4 s 4961 0 5381 20080 6 vssd2
port 18 nsew ground bidirectional
rlabel metal4 s 0 0 800 20080 6 vssd2
port 19 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 12184 20080
string LEFview TRUE
string GDS_FILE /project/openlane/ACMP/runs/ACMP/results/magic/ACMP.gds
string GDS_END 269770
string GDS_START 52858
<< end >>

