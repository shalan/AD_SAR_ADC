magic
tech sky130A
magscale 1 2
timestamp 1626123697
<< locali >>
rect 3525 410363 3559 410737
rect 236101 336107 236135 337909
rect 239045 330259 239079 337841
rect 239413 335767 239447 336617
rect 244105 335835 244139 337841
rect 248981 336243 249015 336549
rect 249073 336379 249107 336617
rect 254409 336243 254443 337841
rect 275569 336515 275603 337841
rect 249717 330803 249751 330973
rect 249809 330735 249843 330905
rect 254593 329035 254627 336413
rect 258733 335835 258767 336073
rect 258825 335903 258859 336073
rect 257353 334883 257387 335053
rect 277961 332163 277995 337841
rect 278145 336175 278179 336277
rect 278237 336243 278271 337773
rect 278053 335563 278087 336073
rect 280813 330395 280847 337773
rect 284769 336175 284803 336277
rect 282469 335359 282503 335733
rect 287621 335631 287655 336413
rect 287713 335971 287747 336617
rect 285873 334407 285907 335529
rect 290841 331959 290875 337773
rect 292497 335495 292531 336549
rect 296637 335835 296671 336209
rect 300317 334747 300351 335801
rect 298845 330463 298879 330905
rect 300685 330259 300719 337841
rect 307033 335903 307067 339745
rect 302065 335631 302099 335869
rect 302341 335699 302375 335801
rect 302065 335597 302157 335631
rect 302433 335427 302467 335665
rect 302617 335631 302651 335869
rect 302375 335393 302467 335427
rect 292129 326247 292163 326485
rect 295165 12019 295199 12257
rect 295257 11951 295291 12325
rect 249257 5151 249291 5525
rect 304641 4471 304675 4641
rect 229661 3451 229695 4165
rect 233801 3451 233835 3689
rect 233893 3587 233927 3689
rect 233709 3383 233743 3417
rect 233985 3383 234019 3553
rect 260573 3519 260607 3825
rect 263057 3587 263091 3757
rect 233709 3349 234019 3383
rect 102241 3179 102275 3281
rect 102183 3145 102275 3179
rect 110429 3043 110463 3145
rect 119997 2907 120031 3009
rect 415443 2941 415627 2975
rect 415593 2907 415627 2941
rect 122205 2839 122239 2873
rect 122205 2805 122423 2839
rect 127023 2805 127173 2839
rect 122389 2771 122423 2805
<< viali >>
rect 3525 410737 3559 410771
rect 3525 410329 3559 410363
rect 307033 339745 307067 339779
rect 236101 337909 236135 337943
rect 236101 336073 236135 336107
rect 239045 337841 239079 337875
rect 244105 337841 244139 337875
rect 239413 336617 239447 336651
rect 254409 337841 254443 337875
rect 249073 336617 249107 336651
rect 248981 336549 249015 336583
rect 249073 336345 249107 336379
rect 248981 336209 249015 336243
rect 275569 337841 275603 337875
rect 275569 336481 275603 336515
rect 277961 337841 277995 337875
rect 254409 336209 254443 336243
rect 254593 336413 254627 336447
rect 244105 335801 244139 335835
rect 239413 335733 239447 335767
rect 249717 330973 249751 331007
rect 249717 330769 249751 330803
rect 249809 330905 249843 330939
rect 249809 330701 249843 330735
rect 239045 330225 239079 330259
rect 258733 336073 258767 336107
rect 258825 336073 258859 336107
rect 258825 335869 258859 335903
rect 258733 335801 258767 335835
rect 257353 335053 257387 335087
rect 257353 334849 257387 334883
rect 300685 337841 300719 337875
rect 278237 337773 278271 337807
rect 278145 336277 278179 336311
rect 278237 336209 278271 336243
rect 280813 337773 280847 337807
rect 278145 336141 278179 336175
rect 278053 336073 278087 336107
rect 278053 335529 278087 335563
rect 277961 332129 277995 332163
rect 290841 337773 290875 337807
rect 287713 336617 287747 336651
rect 287621 336413 287655 336447
rect 284769 336277 284803 336311
rect 284769 336141 284803 336175
rect 282469 335733 282503 335767
rect 287713 335937 287747 335971
rect 287621 335597 287655 335631
rect 282469 335325 282503 335359
rect 285873 335529 285907 335563
rect 285873 334373 285907 334407
rect 292497 336549 292531 336583
rect 296637 336209 296671 336243
rect 296637 335801 296671 335835
rect 300317 335801 300351 335835
rect 292497 335461 292531 335495
rect 300317 334713 300351 334747
rect 290841 331925 290875 331959
rect 298845 330905 298879 330939
rect 298845 330429 298879 330463
rect 280813 330361 280847 330395
rect 302065 335869 302099 335903
rect 302617 335869 302651 335903
rect 307033 335869 307067 335903
rect 302341 335801 302375 335835
rect 302341 335665 302375 335699
rect 302433 335665 302467 335699
rect 302157 335597 302191 335631
rect 302617 335597 302651 335631
rect 302341 335393 302375 335427
rect 300685 330225 300719 330259
rect 254593 329001 254627 329035
rect 292129 326485 292163 326519
rect 292129 326213 292163 326247
rect 295257 12325 295291 12359
rect 295165 12257 295199 12291
rect 295165 11985 295199 12019
rect 295257 11917 295291 11951
rect 249257 5525 249291 5559
rect 249257 5117 249291 5151
rect 304641 4641 304675 4675
rect 304641 4437 304675 4471
rect 229661 4165 229695 4199
rect 260573 3825 260607 3859
rect 233801 3689 233835 3723
rect 233893 3689 233927 3723
rect 233893 3553 233927 3587
rect 233985 3553 234019 3587
rect 229661 3417 229695 3451
rect 233709 3417 233743 3451
rect 233801 3417 233835 3451
rect 263057 3757 263091 3791
rect 263057 3553 263091 3587
rect 260573 3485 260607 3519
rect 102241 3281 102275 3315
rect 102149 3145 102183 3179
rect 110429 3145 110463 3179
rect 110429 3009 110463 3043
rect 119997 3009 120031 3043
rect 415409 2941 415443 2975
rect 119997 2873 120031 2907
rect 122205 2873 122239 2907
rect 415593 2873 415627 2907
rect 126989 2805 127023 2839
rect 127173 2805 127207 2839
rect 122389 2737 122423 2771
<< metal1 >>
rect 285582 700952 285588 701004
rect 285640 700992 285646 701004
rect 413646 700992 413652 701004
rect 285640 700964 413652 700992
rect 285640 700952 285646 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 286962 700884 286968 700936
rect 287020 700924 287026 700936
rect 429838 700924 429844 700936
rect 287020 700896 429844 700924
rect 287020 700884 287026 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 288342 700816 288348 700868
rect 288400 700856 288406 700868
rect 446122 700856 446128 700868
rect 288400 700828 446128 700856
rect 288400 700816 288406 700828
rect 446122 700816 446128 700828
rect 446180 700816 446186 700868
rect 291102 700748 291108 700800
rect 291160 700788 291166 700800
rect 462314 700788 462320 700800
rect 291160 700760 462320 700788
rect 291160 700748 291166 700760
rect 462314 700748 462320 700760
rect 462372 700748 462378 700800
rect 292482 700680 292488 700732
rect 292540 700720 292546 700732
rect 478506 700720 478512 700732
rect 292540 700692 478512 700720
rect 292540 700680 292546 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 295242 700612 295248 700664
rect 295300 700652 295306 700664
rect 494790 700652 494796 700664
rect 295300 700624 494796 700652
rect 295300 700612 295306 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 296622 700544 296628 700596
rect 296680 700584 296686 700596
rect 510982 700584 510988 700596
rect 296680 700556 510988 700584
rect 296680 700544 296686 700556
rect 510982 700544 510988 700556
rect 511040 700544 511046 700596
rect 299382 700476 299388 700528
rect 299440 700516 299446 700528
rect 527174 700516 527180 700528
rect 299440 700488 527180 700516
rect 299440 700476 299446 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 300762 700408 300768 700460
rect 300820 700448 300826 700460
rect 543458 700448 543464 700460
rect 300820 700420 543464 700448
rect 300820 700408 300826 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 235902 700380 235908 700392
rect 235224 700352 235908 700380
rect 235224 700340 235230 700352
rect 235902 700340 235908 700352
rect 235960 700340 235966 700392
rect 269022 700340 269028 700392
rect 269080 700380 269086 700392
rect 283834 700380 283840 700392
rect 269080 700352 283840 700380
rect 269080 700340 269086 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 302142 700340 302148 700392
rect 302200 700380 302206 700392
rect 559650 700380 559656 700392
rect 302200 700352 559656 700380
rect 302200 700340 302206 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 271782 700272 271788 700324
rect 271840 700312 271846 700324
rect 300118 700312 300124 700324
rect 271840 700284 300124 700312
rect 271840 700272 271846 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 304902 700272 304908 700324
rect 304960 700312 304966 700324
rect 575842 700312 575848 700324
rect 304960 700284 575848 700312
rect 304960 700272 304966 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 282822 700204 282828 700256
rect 282880 700244 282886 700256
rect 397454 700244 397460 700256
rect 282880 700216 397460 700244
rect 282880 700204 282886 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 56778 700136 56784 700188
rect 56836 700176 56842 700188
rect 57882 700176 57888 700188
rect 56836 700148 57888 700176
rect 56836 700136 56842 700148
rect 57882 700136 57888 700148
rect 57940 700136 57946 700188
rect 186498 700136 186504 700188
rect 186556 700176 186562 700188
rect 187602 700176 187608 700188
rect 186556 700148 187608 700176
rect 186556 700136 186562 700148
rect 187602 700136 187608 700148
rect 187660 700136 187666 700188
rect 281442 700136 281448 700188
rect 281500 700176 281506 700188
rect 381170 700176 381176 700188
rect 281500 700148 381176 700176
rect 281500 700136 281506 700148
rect 381170 700136 381176 700148
rect 381228 700136 381234 700188
rect 251450 700068 251456 700120
rect 251508 700108 251514 700120
rect 252462 700108 252468 700120
rect 251508 700080 252468 700108
rect 251508 700068 251514 700080
rect 252462 700068 252468 700080
rect 252520 700068 252526 700120
rect 278682 700068 278688 700120
rect 278740 700108 278746 700120
rect 364978 700108 364984 700120
rect 278740 700080 364984 700108
rect 278740 700068 278746 700080
rect 364978 700068 364984 700080
rect 365036 700068 365042 700120
rect 277302 700000 277308 700052
rect 277360 700040 277366 700052
rect 348786 700040 348792 700052
rect 277360 700012 348792 700040
rect 277360 700000 277366 700012
rect 348786 700000 348792 700012
rect 348844 700000 348850 700052
rect 275922 699932 275928 699984
rect 275980 699972 275986 699984
rect 332502 699972 332508 699984
rect 275980 699944 332508 699972
rect 275980 699932 275986 699944
rect 332502 699932 332508 699944
rect 332560 699932 332566 699984
rect 273162 699864 273168 699916
rect 273220 699904 273226 699916
rect 316310 699904 316316 699916
rect 273220 699876 316316 699904
rect 273220 699864 273226 699876
rect 316310 699864 316316 699876
rect 316368 699864 316374 699916
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 122742 699700 122748 699712
rect 121696 699672 122748 699700
rect 121696 699660 121702 699672
rect 122742 699660 122748 699672
rect 122800 699660 122806 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 266354 699660 266360 699712
rect 266412 699700 266418 699712
rect 267642 699700 267648 699712
rect 266412 699672 267648 699700
rect 266412 699660 266418 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 3418 696940 3424 696992
rect 3476 696980 3482 696992
rect 184198 696980 184204 696992
rect 3476 696952 184204 696980
rect 3476 696940 3482 696952
rect 184198 696940 184204 696952
rect 184256 696940 184262 696992
rect 307018 696940 307024 696992
rect 307076 696980 307082 696992
rect 580166 696980 580172 696992
rect 307076 696952 580172 696980
rect 307076 696940 307082 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 307110 683136 307116 683188
rect 307168 683176 307174 683188
rect 580166 683176 580172 683188
rect 307168 683148 580172 683176
rect 307168 683136 307174 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 307202 670692 307208 670744
rect 307260 670732 307266 670744
rect 580166 670732 580172 670744
rect 307260 670704 580172 670732
rect 307260 670692 307266 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3326 644444 3332 644496
rect 3384 644484 3390 644496
rect 195238 644484 195244 644496
rect 3384 644456 195244 644484
rect 3384 644444 3390 644456
rect 195238 644444 195244 644456
rect 195296 644444 195302 644496
rect 307294 643084 307300 643136
rect 307352 643124 307358 643136
rect 580166 643124 580172 643136
rect 307352 643096 580172 643124
rect 307352 643084 307358 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 309778 630640 309784 630692
rect 309836 630680 309842 630692
rect 579982 630680 579988 630692
rect 309836 630652 579988 630680
rect 309836 630640 309842 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 2774 619080 2780 619132
rect 2832 619120 2838 619132
rect 4798 619120 4804 619132
rect 2832 619092 4804 619120
rect 2832 619080 2838 619092
rect 4798 619080 4804 619092
rect 4856 619080 4862 619132
rect 2958 592016 2964 592068
rect 3016 592056 3022 592068
rect 197998 592056 198004 592068
rect 3016 592028 198004 592056
rect 3016 592016 3022 592028
rect 197998 592016 198004 592028
rect 198056 592016 198062 592068
rect 307386 590656 307392 590708
rect 307444 590696 307450 590708
rect 580166 590696 580172 590708
rect 307444 590668 580172 590696
rect 307444 590656 307450 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 307478 576852 307484 576904
rect 307536 576892 307542 576904
rect 579982 576892 579988 576904
rect 307536 576864 579988 576892
rect 307536 576852 307542 576864
rect 579982 576852 579988 576864
rect 580040 576852 580046 576904
rect 2866 539588 2872 539640
rect 2924 539628 2930 539640
rect 220078 539628 220084 539640
rect 2924 539600 220084 539628
rect 2924 539588 2930 539600
rect 220078 539588 220084 539600
rect 220136 539588 220142 539640
rect 307570 536800 307576 536852
rect 307628 536840 307634 536852
rect 580166 536840 580172 536852
rect 307628 536812 580172 536840
rect 307628 536800 307634 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 307662 524424 307668 524476
rect 307720 524464 307726 524476
rect 580166 524464 580172 524476
rect 307720 524436 580172 524464
rect 307720 524424 307726 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 10318 514808 10324 514820
rect 3384 514780 10324 514808
rect 3384 514768 3390 514780
rect 10318 514768 10324 514780
rect 10376 514768 10382 514820
rect 306926 484372 306932 484424
rect 306984 484412 306990 484424
rect 580166 484412 580172 484424
rect 306984 484384 580172 484412
rect 306984 484372 306990 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 306834 470568 306840 470620
rect 306892 470608 306898 470620
rect 579982 470608 579988 470620
rect 306892 470580 579988 470608
rect 306892 470568 306898 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 306742 430584 306748 430636
rect 306800 430624 306806 430636
rect 580074 430624 580080 430636
rect 306800 430596 580080 430624
rect 306800 430584 306806 430596
rect 580074 430584 580080 430596
rect 580132 430584 580138 430636
rect 312538 418140 312544 418192
rect 312596 418180 312602 418192
rect 580074 418180 580080 418192
rect 312596 418152 580080 418180
rect 312596 418140 312602 418152
rect 580074 418140 580080 418152
rect 580132 418140 580138 418192
rect 171042 411204 171048 411256
rect 171100 411244 171106 411256
rect 255314 411244 255320 411256
rect 171100 411216 255320 411244
rect 171100 411204 171106 411216
rect 255314 411204 255320 411216
rect 255372 411204 255378 411256
rect 154482 411136 154488 411188
rect 154540 411176 154546 411188
rect 253106 411176 253112 411188
rect 154540 411148 253112 411176
rect 154540 411136 154546 411148
rect 253106 411136 253112 411148
rect 253164 411136 253170 411188
rect 137922 411068 137928 411120
rect 137980 411108 137986 411120
rect 251174 411108 251180 411120
rect 137980 411080 251180 411108
rect 137980 411068 137986 411080
rect 251174 411068 251180 411080
rect 251232 411068 251238 411120
rect 122742 411000 122748 411052
rect 122800 411040 122806 411052
rect 249150 411040 249156 411052
rect 122800 411012 249156 411040
rect 122800 411000 122806 411012
rect 249150 411000 249156 411012
rect 249208 411000 249214 411052
rect 106182 410932 106188 410984
rect 106240 410972 106246 410984
rect 247218 410972 247224 410984
rect 106240 410944 247224 410972
rect 106240 410932 106246 410944
rect 247218 410932 247224 410944
rect 247276 410932 247282 410984
rect 89622 410864 89628 410916
rect 89680 410904 89686 410916
rect 245286 410904 245292 410916
rect 89680 410876 245292 410904
rect 89680 410864 89686 410876
rect 245286 410864 245292 410876
rect 245344 410864 245350 410916
rect 73062 410796 73068 410848
rect 73120 410836 73126 410848
rect 243354 410836 243360 410848
rect 73120 410808 243360 410836
rect 73120 410796 73126 410808
rect 243354 410796 243360 410808
rect 243412 410796 243418 410848
rect 3510 410768 3516 410780
rect 3471 410740 3516 410768
rect 3510 410728 3516 410740
rect 3568 410728 3574 410780
rect 57882 410728 57888 410780
rect 57940 410768 57946 410780
rect 241514 410768 241520 410780
rect 57940 410740 241520 410768
rect 57940 410728 57946 410740
rect 241514 410728 241520 410740
rect 241572 410728 241578 410780
rect 41322 410660 41328 410712
rect 41380 410700 41386 410712
rect 239490 410700 239496 410712
rect 41380 410672 239496 410700
rect 41380 410660 41386 410672
rect 239490 410660 239496 410672
rect 239548 410660 239554 410712
rect 24762 410592 24768 410644
rect 24820 410632 24826 410644
rect 237558 410632 237564 410644
rect 24820 410604 237564 410632
rect 24820 410592 24826 410604
rect 237558 410592 237564 410604
rect 237616 410592 237622 410644
rect 252462 410592 252468 410644
rect 252520 410632 252526 410644
rect 264974 410632 264980 410644
rect 252520 410604 264980 410632
rect 252520 410592 252526 410604
rect 264974 410592 264980 410604
rect 265032 410592 265038 410644
rect 8202 410524 8208 410576
rect 8260 410564 8266 410576
rect 235626 410564 235632 410576
rect 8260 410536 235632 410564
rect 8260 410524 8266 410536
rect 235626 410524 235632 410536
rect 235684 410524 235690 410576
rect 235902 410524 235908 410576
rect 235960 410564 235966 410576
rect 262766 410564 262772 410576
rect 235960 410536 262772 410564
rect 235960 410524 235966 410536
rect 262766 410524 262772 410536
rect 262824 410524 262830 410576
rect 3418 410456 3424 410508
rect 3476 410496 3482 410508
rect 7558 410496 7564 410508
rect 3476 410468 7564 410496
rect 3476 410456 3482 410468
rect 7558 410456 7564 410468
rect 7616 410456 7622 410508
rect 187602 410456 187608 410508
rect 187660 410496 187666 410508
rect 256970 410496 256976 410508
rect 187660 410468 256976 410496
rect 187660 410456 187666 410468
rect 256970 410456 256976 410468
rect 257028 410456 257034 410508
rect 202782 410388 202788 410440
rect 202840 410428 202846 410440
rect 258902 410428 258908 410440
rect 202840 410400 258908 410428
rect 202840 410388 202846 410400
rect 258902 410388 258908 410400
rect 258960 410388 258966 410440
rect 3418 410320 3424 410372
rect 3476 410360 3482 410372
rect 3513 410363 3571 410369
rect 3513 410360 3525 410363
rect 3476 410332 3525 410360
rect 3476 410320 3482 410332
rect 3513 410329 3525 410332
rect 3559 410329 3571 410363
rect 3513 410323 3571 410329
rect 219342 410320 219348 410372
rect 219400 410360 219406 410372
rect 260834 410360 260840 410372
rect 219400 410332 260840 410360
rect 219400 410320 219406 410332
rect 260834 410320 260840 410332
rect 260892 410320 260898 410372
rect 271230 409912 271236 409964
rect 271288 409952 271294 409964
rect 271782 409952 271788 409964
rect 271288 409924 271788 409952
rect 271288 409912 271294 409924
rect 271782 409912 271788 409924
rect 271840 409912 271846 409964
rect 275094 409912 275100 409964
rect 275152 409952 275158 409964
rect 275922 409952 275928 409964
rect 275152 409924 275928 409952
rect 275152 409912 275158 409924
rect 275922 409912 275928 409924
rect 275980 409912 275986 409964
rect 280982 409912 280988 409964
rect 281040 409952 281046 409964
rect 281442 409952 281448 409964
rect 281040 409924 281448 409952
rect 281040 409912 281046 409924
rect 281442 409912 281448 409924
rect 281500 409912 281506 409964
rect 284846 409912 284852 409964
rect 284904 409952 284910 409964
rect 285582 409952 285588 409964
rect 284904 409924 285588 409952
rect 284904 409912 284910 409924
rect 285582 409912 285588 409924
rect 285640 409912 285646 409964
rect 290642 409912 290648 409964
rect 290700 409952 290706 409964
rect 291102 409952 291108 409964
rect 290700 409924 291108 409952
rect 290700 409912 290706 409924
rect 291102 409912 291108 409924
rect 291160 409912 291166 409964
rect 294598 409912 294604 409964
rect 294656 409952 294662 409964
rect 295242 409952 295248 409964
rect 294656 409924 295248 409952
rect 294656 409912 294662 409924
rect 295242 409912 295248 409924
rect 295300 409912 295306 409964
rect 298462 409912 298468 409964
rect 298520 409952 298526 409964
rect 299382 409952 299388 409964
rect 298520 409924 299388 409952
rect 298520 409912 298526 409924
rect 299382 409912 299388 409924
rect 299440 409912 299446 409964
rect 304258 409912 304264 409964
rect 304316 409952 304322 409964
rect 304902 409952 304908 409964
rect 304316 409924 304908 409952
rect 304316 409912 304322 409924
rect 304902 409912 304908 409924
rect 304960 409912 304966 409964
rect 184198 408416 184204 408468
rect 184256 408456 184262 408468
rect 232038 408456 232044 408468
rect 184256 408428 232044 408456
rect 184256 408416 184262 408428
rect 232038 408416 232044 408428
rect 232096 408416 232102 408468
rect 3510 405628 3516 405680
rect 3568 405668 3574 405680
rect 232038 405668 232044 405680
rect 3568 405640 232044 405668
rect 3568 405628 3574 405640
rect 232038 405628 232044 405640
rect 232096 405628 232102 405680
rect 307018 404336 307024 404388
rect 307076 404376 307082 404388
rect 580074 404376 580080 404388
rect 307076 404348 580080 404376
rect 307076 404336 307082 404348
rect 580074 404336 580080 404348
rect 580132 404336 580138 404388
rect 3418 404268 3424 404320
rect 3476 404308 3482 404320
rect 232038 404308 232044 404320
rect 3476 404280 232044 404308
rect 3476 404268 3482 404280
rect 232038 404268 232044 404280
rect 232096 404268 232102 404320
rect 307202 404268 307208 404320
rect 307260 404308 307266 404320
rect 580258 404308 580264 404320
rect 307260 404280 580264 404308
rect 307260 404268 307266 404280
rect 580258 404268 580264 404280
rect 580316 404268 580322 404320
rect 580074 404200 580080 404252
rect 580132 404240 580138 404252
rect 580442 404240 580448 404252
rect 580132 404212 580448 404240
rect 580132 404200 580138 404212
rect 580442 404200 580448 404212
rect 580500 404200 580506 404252
rect 195238 402908 195244 402960
rect 195296 402948 195302 402960
rect 232038 402948 232044 402960
rect 195296 402920 232044 402948
rect 195296 402908 195302 402920
rect 232038 402908 232044 402920
rect 232096 402908 232102 402960
rect 3602 401548 3608 401600
rect 3660 401588 3666 401600
rect 232038 401588 232044 401600
rect 3660 401560 232044 401588
rect 3660 401548 3666 401560
rect 232038 401548 232044 401560
rect 232096 401548 232102 401600
rect 307294 401276 307300 401328
rect 307352 401316 307358 401328
rect 309778 401316 309784 401328
rect 307352 401288 309784 401316
rect 307352 401276 307358 401288
rect 309778 401276 309784 401288
rect 309836 401276 309842 401328
rect 4798 400120 4804 400172
rect 4856 400160 4862 400172
rect 232038 400160 232044 400172
rect 4856 400132 232044 400160
rect 4856 400120 4862 400132
rect 232038 400120 232044 400132
rect 232096 400120 232102 400172
rect 307202 400120 307208 400172
rect 307260 400160 307266 400172
rect 580350 400160 580356 400172
rect 307260 400132 580356 400160
rect 307260 400120 307266 400132
rect 580350 400120 580356 400132
rect 580408 400120 580414 400172
rect 307294 398896 307300 398948
rect 307352 398936 307358 398948
rect 307478 398936 307484 398948
rect 307352 398908 307484 398936
rect 307352 398896 307358 398908
rect 307478 398896 307484 398908
rect 307536 398896 307542 398948
rect 3694 398760 3700 398812
rect 3752 398800 3758 398812
rect 232038 398800 232044 398812
rect 3752 398772 232044 398800
rect 3752 398760 3758 398772
rect 232038 398760 232044 398772
rect 232096 398760 232102 398812
rect 307478 398760 307484 398812
rect 307536 398800 307542 398812
rect 580074 398800 580080 398812
rect 307536 398772 580080 398800
rect 307536 398760 307542 398772
rect 580074 398760 580080 398772
rect 580132 398760 580138 398812
rect 197998 397400 198004 397452
rect 198056 397440 198062 397452
rect 232038 397440 232044 397452
rect 198056 397412 232044 397440
rect 198056 397400 198062 397412
rect 232038 397400 232044 397412
rect 232096 397400 232102 397452
rect 3786 395972 3792 396024
rect 3844 396012 3850 396024
rect 232038 396012 232044 396024
rect 3844 395984 232044 396012
rect 3844 395972 3850 395984
rect 232038 395972 232044 395984
rect 232096 395972 232102 396024
rect 3878 394612 3884 394664
rect 3936 394652 3942 394664
rect 231946 394652 231952 394664
rect 3936 394624 231952 394652
rect 3936 394612 3942 394624
rect 231946 394612 231952 394624
rect 232004 394612 232010 394664
rect 307478 394612 307484 394664
rect 307536 394652 307542 394664
rect 580534 394652 580540 394664
rect 307536 394624 580540 394652
rect 307536 394612 307542 394624
rect 580534 394612 580540 394624
rect 580592 394612 580598 394664
rect 3970 393252 3976 393304
rect 4028 393292 4034 393304
rect 232038 393292 232044 393304
rect 4028 393264 232044 393292
rect 4028 393252 4034 393264
rect 232038 393252 232044 393264
rect 232096 393252 232102 393304
rect 307478 393252 307484 393304
rect 307536 393292 307542 393304
rect 580626 393292 580632 393304
rect 307536 393264 580632 393292
rect 307536 393252 307542 393264
rect 580626 393252 580632 393264
rect 580684 393252 580690 393304
rect 220078 391892 220084 391944
rect 220136 391932 220142 391944
rect 232038 391932 232044 391944
rect 220136 391904 232044 391932
rect 220136 391892 220142 391904
rect 232038 391892 232044 391904
rect 232096 391892 232102 391944
rect 307110 390532 307116 390584
rect 307168 390572 307174 390584
rect 580074 390572 580080 390584
rect 307168 390544 580080 390572
rect 307168 390532 307174 390544
rect 580074 390532 580080 390544
rect 580132 390532 580138 390584
rect 4062 390464 4068 390516
rect 4120 390504 4126 390516
rect 232038 390504 232044 390516
rect 4120 390476 232044 390504
rect 4120 390464 4126 390476
rect 232038 390464 232044 390476
rect 232096 390464 232102 390516
rect 3326 389104 3332 389156
rect 3384 389144 3390 389156
rect 231946 389144 231952 389156
rect 3384 389116 231952 389144
rect 3384 389104 3390 389116
rect 231946 389104 231952 389116
rect 232004 389104 232010 389156
rect 307662 389104 307668 389156
rect 307720 389144 307726 389156
rect 580718 389144 580724 389156
rect 307720 389116 580724 389144
rect 307720 389104 307726 389116
rect 580718 389104 580724 389116
rect 580776 389104 580782 389156
rect 10318 389036 10324 389088
rect 10376 389076 10382 389088
rect 232038 389076 232044 389088
rect 10376 389048 232044 389076
rect 10376 389036 10382 389048
rect 232038 389036 232044 389048
rect 232096 389036 232102 389088
rect 3234 387744 3240 387796
rect 3292 387784 3298 387796
rect 232038 387784 232044 387796
rect 3292 387756 232044 387784
rect 3292 387744 3298 387756
rect 232038 387744 232044 387756
rect 232096 387744 232102 387796
rect 307662 387744 307668 387796
rect 307720 387784 307726 387796
rect 580810 387784 580816 387796
rect 307720 387756 580816 387784
rect 307720 387744 307726 387756
rect 580810 387744 580816 387756
rect 580868 387744 580874 387796
rect 3142 386316 3148 386368
rect 3200 386356 3206 386368
rect 232038 386356 232044 386368
rect 3200 386328 232044 386356
rect 3200 386316 3206 386328
rect 232038 386316 232044 386328
rect 232096 386316 232102 386368
rect 3050 384956 3056 385008
rect 3108 384996 3114 385008
rect 232038 384996 232044 385008
rect 3108 384968 232044 384996
rect 3108 384956 3114 384968
rect 232038 384956 232044 384968
rect 232096 384956 232102 385008
rect 2958 383596 2964 383648
rect 3016 383636 3022 383648
rect 231854 383636 231860 383648
rect 3016 383608 231860 383636
rect 3016 383596 3022 383608
rect 231854 383596 231860 383608
rect 231912 383596 231918 383648
rect 307662 383596 307668 383648
rect 307720 383636 307726 383648
rect 580902 383636 580908 383648
rect 307720 383608 580908 383636
rect 307720 383596 307726 383608
rect 580902 383596 580908 383608
rect 580960 383596 580966 383648
rect 2866 382168 2872 382220
rect 2924 382208 2930 382220
rect 232038 382208 232044 382220
rect 2924 382180 232044 382208
rect 2924 382168 2930 382180
rect 232038 382168 232044 382180
rect 232096 382168 232102 382220
rect 307662 382168 307668 382220
rect 307720 382208 307726 382220
rect 580166 382208 580172 382220
rect 307720 382180 580172 382208
rect 307720 382168 307726 382180
rect 580166 382168 580172 382180
rect 580224 382168 580230 382220
rect 2774 380808 2780 380860
rect 2832 380848 2838 380860
rect 232038 380848 232044 380860
rect 2832 380820 232044 380848
rect 2832 380808 2838 380820
rect 232038 380808 232044 380820
rect 232096 380808 232102 380860
rect 306834 380808 306840 380860
rect 306892 380848 306898 380860
rect 312538 380848 312544 380860
rect 306892 380820 312544 380848
rect 306892 380808 306898 380820
rect 312538 380808 312544 380820
rect 312596 380808 312602 380860
rect 7558 379448 7564 379500
rect 7616 379488 7622 379500
rect 232038 379488 232044 379500
rect 7616 379460 232044 379488
rect 7616 379448 7622 379460
rect 232038 379448 232044 379460
rect 232096 379448 232102 379500
rect 307662 378156 307668 378208
rect 307720 378196 307726 378208
rect 580166 378196 580172 378208
rect 307720 378168 580172 378196
rect 307720 378156 307726 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3418 378088 3424 378140
rect 3476 378128 3482 378140
rect 232038 378128 232044 378140
rect 3476 378100 232044 378128
rect 3476 378088 3482 378100
rect 232038 378088 232044 378100
rect 232096 378088 232102 378140
rect 3510 376660 3516 376712
rect 3568 376700 3574 376712
rect 232038 376700 232044 376712
rect 3568 376672 232044 376700
rect 3568 376660 3574 376672
rect 232038 376660 232044 376672
rect 232096 376660 232102 376712
rect 3510 374008 3516 374060
rect 3568 374048 3574 374060
rect 232038 374048 232044 374060
rect 3568 374020 232044 374048
rect 3568 374008 3574 374020
rect 232038 374008 232044 374020
rect 232096 374008 232102 374060
rect 3602 372580 3608 372632
rect 3660 372620 3666 372632
rect 232038 372620 232044 372632
rect 3660 372592 232044 372620
rect 3660 372580 3666 372592
rect 232038 372580 232044 372592
rect 232096 372580 232102 372632
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 232038 371260 232044 371272
rect 3476 371232 232044 371260
rect 3476 371220 3482 371232
rect 232038 371220 232044 371232
rect 232096 371220 232102 371272
rect 307662 371220 307668 371272
rect 307720 371260 307726 371272
rect 320818 371260 320824 371272
rect 307720 371232 320824 371260
rect 307720 371220 307726 371232
rect 320818 371220 320824 371232
rect 320876 371220 320882 371272
rect 3142 367072 3148 367124
rect 3200 367112 3206 367124
rect 232038 367112 232044 367124
rect 3200 367084 232044 367112
rect 3200 367072 3206 367084
rect 232038 367072 232044 367084
rect 232096 367072 232102 367124
rect 7558 365712 7564 365764
rect 7616 365752 7622 365764
rect 232038 365752 232044 365764
rect 7616 365724 232044 365752
rect 7616 365712 7622 365724
rect 232038 365712 232044 365724
rect 232096 365712 232102 365764
rect 307662 365712 307668 365764
rect 307720 365752 307726 365764
rect 461578 365752 461584 365764
rect 307720 365724 461584 365752
rect 307720 365712 307726 365724
rect 461578 365712 461584 365724
rect 461636 365712 461642 365764
rect 307110 365644 307116 365696
rect 307168 365684 307174 365696
rect 580166 365684 580172 365696
rect 307168 365656 580172 365684
rect 307168 365644 307174 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 307662 364352 307668 364404
rect 307720 364392 307726 364404
rect 316678 364392 316684 364404
rect 307720 364364 316684 364392
rect 307720 364352 307726 364364
rect 316678 364352 316684 364364
rect 316736 364352 316742 364404
rect 22830 362924 22836 362976
rect 22888 362964 22894 362976
rect 232038 362964 232044 362976
rect 22888 362936 232044 362964
rect 22888 362924 22894 362936
rect 232038 362924 232044 362936
rect 232096 362924 232102 362976
rect 307294 362924 307300 362976
rect 307352 362964 307358 362976
rect 331858 362964 331864 362976
rect 307352 362936 331864 362964
rect 307352 362924 307358 362936
rect 331858 362924 331864 362936
rect 331916 362924 331922 362976
rect 3234 361564 3240 361616
rect 3292 361604 3298 361616
rect 232038 361604 232044 361616
rect 3292 361576 232044 361604
rect 3292 361564 3298 361576
rect 232038 361564 232044 361576
rect 232096 361564 232102 361616
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 232038 357456 232044 357468
rect 3384 357428 232044 357456
rect 3384 357416 3390 357428
rect 232038 357416 232044 357428
rect 232096 357416 232102 357468
rect 307662 356328 307668 356380
rect 307720 356368 307726 356380
rect 309778 356368 309784 356380
rect 307720 356340 309784 356368
rect 307720 356328 307726 356340
rect 309778 356328 309784 356340
rect 309836 356328 309842 356380
rect 14550 356056 14556 356108
rect 14608 356096 14614 356108
rect 232038 356096 232044 356108
rect 14608 356068 232044 356096
rect 14608 356056 14614 356068
rect 232038 356056 232044 356068
rect 232096 356056 232102 356108
rect 307662 354696 307668 354748
rect 307720 354736 307726 354748
rect 324958 354736 324964 354748
rect 307720 354708 324964 354736
rect 307720 354696 307726 354708
rect 324958 354696 324964 354708
rect 325016 354696 325022 354748
rect 4062 353268 4068 353320
rect 4120 353308 4126 353320
rect 232038 353308 232044 353320
rect 4120 353280 232044 353308
rect 4120 353268 4126 353280
rect 232038 353268 232044 353280
rect 232096 353268 232102 353320
rect 307110 353200 307116 353252
rect 307168 353240 307174 353252
rect 580166 353240 580172 353252
rect 307168 353212 580172 353240
rect 307168 353200 307174 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 25498 351908 25504 351960
rect 25556 351948 25562 351960
rect 232038 351948 232044 351960
rect 25556 351920 232044 351948
rect 25556 351908 25562 351920
rect 232038 351908 232044 351920
rect 232096 351908 232102 351960
rect 3970 350548 3976 350600
rect 4028 350588 4034 350600
rect 232038 350588 232044 350600
rect 4028 350560 232044 350588
rect 4028 350548 4034 350560
rect 232038 350548 232044 350560
rect 232096 350548 232102 350600
rect 3878 347760 3884 347812
rect 3936 347800 3942 347812
rect 232038 347800 232044 347812
rect 3936 347772 232044 347800
rect 3936 347760 3942 347772
rect 232038 347760 232044 347772
rect 232096 347760 232102 347812
rect 307662 347760 307668 347812
rect 307720 347800 307726 347812
rect 323578 347800 323584 347812
rect 307720 347772 323584 347800
rect 307720 347760 307726 347772
rect 323578 347760 323584 347772
rect 323636 347760 323642 347812
rect 3786 346400 3792 346452
rect 3844 346440 3850 346452
rect 232038 346440 232044 346452
rect 3844 346412 232044 346440
rect 3844 346400 3850 346412
rect 232038 346400 232044 346412
rect 232096 346400 232102 346452
rect 15838 345040 15844 345092
rect 15896 345080 15902 345092
rect 232038 345080 232044 345092
rect 15896 345052 232044 345080
rect 15896 345040 15902 345052
rect 232038 345040 232044 345052
rect 232096 345040 232102 345092
rect 32398 343680 32404 343732
rect 32456 343720 32462 343732
rect 232038 343720 232044 343732
rect 32456 343692 232044 343720
rect 32456 343680 32462 343692
rect 232038 343680 232044 343692
rect 232096 343680 232102 343732
rect 3694 343612 3700 343664
rect 3752 343652 3758 343664
rect 231854 343652 231860 343664
rect 3752 343624 231860 343652
rect 3752 343612 3758 343624
rect 231854 343612 231860 343624
rect 231912 343612 231918 343664
rect 3602 342252 3608 342304
rect 3660 342292 3666 342304
rect 232038 342292 232044 342304
rect 3660 342264 232044 342292
rect 3660 342252 3666 342264
rect 232038 342252 232044 342264
rect 232096 342252 232102 342304
rect 306282 342252 306288 342304
rect 306340 342292 306346 342304
rect 460198 342292 460204 342304
rect 306340 342264 460204 342292
rect 306340 342252 306346 342264
rect 460198 342252 460204 342264
rect 460256 342252 460262 342304
rect 3510 340892 3516 340944
rect 3568 340932 3574 340944
rect 232038 340932 232044 340944
rect 3568 340904 232044 340932
rect 3568 340892 3574 340904
rect 232038 340892 232044 340904
rect 232096 340892 232102 340944
rect 320818 340144 320824 340196
rect 320876 340184 320882 340196
rect 580166 340184 580172 340196
rect 320876 340156 580172 340184
rect 320876 340144 320882 340156
rect 580166 340144 580172 340156
rect 580224 340144 580230 340196
rect 307021 339779 307079 339785
rect 307021 339745 307033 339779
rect 307067 339776 307079 339779
rect 307202 339776 307208 339788
rect 307067 339748 307208 339776
rect 307067 339745 307079 339748
rect 307021 339739 307079 339745
rect 307202 339736 307208 339748
rect 307260 339736 307266 339788
rect 3418 339464 3424 339516
rect 3476 339504 3482 339516
rect 232038 339504 232044 339516
rect 3476 339476 232044 339504
rect 3476 339464 3482 339476
rect 232038 339464 232044 339476
rect 232096 339464 232102 339516
rect 307202 339464 307208 339516
rect 307260 339504 307266 339516
rect 318058 339504 318064 339516
rect 307260 339476 318064 339504
rect 307260 339464 307266 339476
rect 318058 339464 318064 339476
rect 318116 339464 318122 339516
rect 17218 338104 17224 338156
rect 17276 338144 17282 338156
rect 232038 338144 232044 338156
rect 17276 338116 232044 338144
rect 17276 338104 17282 338116
rect 232038 338104 232044 338116
rect 232096 338104 232102 338156
rect 307202 338104 307208 338156
rect 307260 338144 307266 338156
rect 406378 338144 406384 338156
rect 307260 338116 406384 338144
rect 307260 338104 307266 338116
rect 406378 338104 406384 338116
rect 406436 338104 406442 338156
rect 234798 337900 234804 337952
rect 234856 337940 234862 337952
rect 235120 337940 235126 337952
rect 234856 337912 235126 337940
rect 234856 337900 234862 337912
rect 235120 337900 235126 337912
rect 235178 337900 235184 337952
rect 236086 337940 236092 337952
rect 236047 337912 236092 337940
rect 236086 337900 236092 337912
rect 236144 337900 236150 337952
rect 262444 337900 262450 337952
rect 262502 337900 262508 337952
rect 303844 337900 303850 337952
rect 303902 337940 303908 337952
rect 305822 337940 305828 337952
rect 303902 337912 305828 337940
rect 303902 337900 303908 337912
rect 305822 337900 305828 337912
rect 305880 337900 305886 337952
rect 235258 337872 235264 337884
rect 234908 337844 235264 337872
rect 234908 337748 234936 337844
rect 235258 337832 235264 337844
rect 235316 337832 235322 337884
rect 239076 337881 239082 337884
rect 239033 337875 239082 337881
rect 239033 337841 239045 337875
rect 239079 337841 239082 337875
rect 239033 337835 239082 337841
rect 239076 337832 239082 337835
rect 239134 337832 239140 337884
rect 241652 337832 241658 337884
rect 241710 337832 241716 337884
rect 244093 337875 244151 337881
rect 244093 337841 244105 337875
rect 244139 337872 244151 337875
rect 244596 337872 244602 337884
rect 244139 337844 244602 337872
rect 244139 337841 244151 337844
rect 244093 337835 244151 337841
rect 244596 337832 244602 337844
rect 244654 337832 244660 337884
rect 246344 337832 246350 337884
rect 246402 337832 246408 337884
rect 247448 337832 247454 337884
rect 247506 337832 247512 337884
rect 254397 337875 254455 337881
rect 254397 337841 254409 337875
rect 254443 337872 254455 337875
rect 257200 337872 257206 337884
rect 254443 337844 257206 337872
rect 254443 337841 254455 337844
rect 254397 337835 254455 337841
rect 257200 337832 257206 337844
rect 257258 337832 257264 337884
rect 262462 337872 262490 337900
rect 262416 337844 262490 337872
rect 236086 337764 236092 337816
rect 236144 337804 236150 337816
rect 236960 337804 236966 337816
rect 236144 337776 236966 337804
rect 236144 337764 236150 337776
rect 236960 337764 236966 337776
rect 237018 337764 237024 337816
rect 240134 337764 240140 337816
rect 240192 337804 240198 337816
rect 240916 337804 240922 337816
rect 240192 337776 240922 337804
rect 240192 337764 240198 337776
rect 240916 337764 240922 337776
rect 240974 337764 240980 337816
rect 241670 337804 241698 337832
rect 242158 337804 242164 337816
rect 241670 337776 242164 337804
rect 242158 337764 242164 337776
rect 242216 337764 242222 337816
rect 243262 337764 243268 337816
rect 243320 337804 243326 337816
rect 243584 337804 243590 337816
rect 243320 337776 243590 337804
rect 243320 337764 243326 337776
rect 243584 337764 243590 337776
rect 243642 337764 243648 337816
rect 246114 337764 246120 337816
rect 246172 337804 246178 337816
rect 246362 337804 246390 337832
rect 246172 337776 246390 337804
rect 246172 337764 246178 337776
rect 247126 337764 247132 337816
rect 247184 337804 247190 337816
rect 247466 337804 247494 337832
rect 247184 337776 247494 337804
rect 247184 337764 247190 337776
rect 251588 337764 251594 337816
rect 251646 337804 251652 337816
rect 251910 337804 251916 337816
rect 251646 337776 251916 337804
rect 251646 337764 251652 337776
rect 251910 337764 251916 337776
rect 251968 337764 251974 337816
rect 253980 337764 253986 337816
rect 254038 337804 254044 337816
rect 254486 337804 254492 337816
rect 254038 337776 254492 337804
rect 254038 337764 254044 337776
rect 254486 337764 254492 337776
rect 254544 337764 254550 337816
rect 255636 337764 255642 337816
rect 255694 337804 255700 337816
rect 256142 337804 256148 337816
rect 255694 337776 256148 337804
rect 255694 337764 255700 337776
rect 256142 337764 256148 337776
rect 256200 337764 256206 337816
rect 258166 337764 258172 337816
rect 258224 337804 258230 337816
rect 259316 337804 259322 337816
rect 258224 337776 259322 337804
rect 258224 337764 258230 337776
rect 259316 337764 259322 337776
rect 259374 337764 259380 337816
rect 261386 337764 261392 337816
rect 261444 337804 261450 337816
rect 262168 337804 262174 337816
rect 261444 337776 262174 337804
rect 261444 337764 261450 337776
rect 262168 337764 262174 337776
rect 262226 337764 262232 337816
rect 234890 337696 234896 337748
rect 234948 337696 234954 337748
rect 262306 337628 262312 337680
rect 262364 337668 262370 337680
rect 262416 337668 262444 337844
rect 275508 337832 275514 337884
rect 275566 337881 275572 337884
rect 275566 337875 275615 337881
rect 275566 337841 275569 337875
rect 275603 337841 275615 337875
rect 275566 337835 275615 337841
rect 275566 337832 275572 337835
rect 276060 337832 276066 337884
rect 276118 337872 276124 337884
rect 277949 337875 278007 337881
rect 277949 337872 277961 337875
rect 276118 337844 277961 337872
rect 276118 337832 276124 337844
rect 277949 337841 277961 337844
rect 277995 337841 278007 337875
rect 277949 337835 278007 337841
rect 280292 337832 280298 337884
rect 280350 337832 280356 337884
rect 300440 337832 300446 337884
rect 300498 337832 300504 337884
rect 300716 337881 300722 337884
rect 300673 337875 300722 337881
rect 300673 337841 300685 337875
rect 300719 337841 300722 337875
rect 300673 337835 300722 337841
rect 300716 337832 300722 337835
rect 300774 337832 300780 337884
rect 301728 337832 301734 337884
rect 301786 337872 301792 337884
rect 305914 337872 305920 337884
rect 301786 337844 305920 337872
rect 301786 337832 301792 337844
rect 305914 337832 305920 337844
rect 305972 337832 305978 337884
rect 262490 337764 262496 337816
rect 262548 337804 262554 337816
rect 263456 337804 263462 337816
rect 262548 337776 263462 337804
rect 262548 337764 262554 337776
rect 263456 337764 263462 337776
rect 263514 337764 263520 337816
rect 267964 337764 267970 337816
rect 268022 337804 268028 337816
rect 268930 337804 268936 337816
rect 268022 337776 268936 337804
rect 268022 337764 268028 337776
rect 268930 337764 268936 337776
rect 268988 337764 268994 337816
rect 271644 337764 271650 337816
rect 271702 337804 271708 337816
rect 278225 337807 278283 337813
rect 278225 337804 278237 337807
rect 271702 337776 278237 337804
rect 271702 337764 271708 337776
rect 278225 337773 278237 337776
rect 278271 337773 278283 337807
rect 278225 337767 278283 337773
rect 278912 337764 278918 337816
rect 278970 337804 278976 337816
rect 279970 337804 279976 337816
rect 278970 337776 279976 337804
rect 278970 337764 278976 337776
rect 279970 337764 279976 337776
rect 280028 337764 280034 337816
rect 280310 337736 280338 337832
rect 280801 337807 280859 337813
rect 280801 337773 280813 337807
rect 280847 337804 280859 337807
rect 281304 337804 281310 337816
rect 280847 337776 281310 337804
rect 280847 337773 280859 337776
rect 280801 337767 280859 337773
rect 281304 337764 281310 337776
rect 281362 337764 281368 337816
rect 281580 337764 281586 337816
rect 281638 337804 281644 337816
rect 282546 337804 282552 337816
rect 281638 337776 282552 337804
rect 281638 337764 281644 337776
rect 282546 337764 282552 337776
rect 282604 337764 282610 337816
rect 285674 337764 285680 337816
rect 285732 337804 285738 337816
rect 286548 337804 286554 337816
rect 285732 337776 286554 337804
rect 285732 337764 285738 337776
rect 286548 337764 286554 337776
rect 286606 337764 286612 337816
rect 287330 337764 287336 337816
rect 287388 337804 287394 337816
rect 288112 337804 288118 337816
rect 287388 337776 288118 337804
rect 287388 337764 287394 337776
rect 288112 337764 288118 337776
rect 288170 337764 288176 337816
rect 289354 337764 289360 337816
rect 289412 337804 289418 337816
rect 289676 337804 289682 337816
rect 289412 337776 289682 337804
rect 289412 337764 289418 337776
rect 289676 337764 289682 337776
rect 289734 337764 289740 337816
rect 290780 337764 290786 337816
rect 290838 337813 290844 337816
rect 290838 337807 290887 337813
rect 290838 337773 290841 337807
rect 290875 337773 290887 337807
rect 290838 337767 290887 337773
rect 290838 337764 290844 337767
rect 292804 337764 292810 337816
rect 292862 337804 292868 337816
rect 293586 337804 293592 337816
rect 292862 337776 293592 337804
rect 292862 337764 292868 337776
rect 293586 337764 293592 337776
rect 293644 337764 293650 337816
rect 296162 337764 296168 337816
rect 296220 337804 296226 337816
rect 296484 337804 296490 337816
rect 296220 337776 296490 337804
rect 296220 337764 296226 337776
rect 296484 337764 296490 337776
rect 296542 337764 296548 337816
rect 280982 337736 280988 337748
rect 280310 337708 280988 337736
rect 280982 337696 280988 337708
rect 281040 337696 281046 337748
rect 262364 337640 262444 337668
rect 262364 337628 262370 337640
rect 300026 337628 300032 337680
rect 300084 337668 300090 337680
rect 300458 337668 300486 337832
rect 302280 337764 302286 337816
rect 302338 337804 302344 337816
rect 303338 337804 303344 337816
rect 302338 337776 303344 337804
rect 302338 337764 302344 337776
rect 303338 337764 303344 337776
rect 303396 337764 303402 337816
rect 304396 337764 304402 337816
rect 304454 337804 304460 337816
rect 304994 337804 305000 337816
rect 304454 337776 305000 337804
rect 304454 337764 304460 337776
rect 304994 337764 305000 337776
rect 305052 337764 305058 337816
rect 300084 337640 300486 337668
rect 300084 337628 300090 337640
rect 277854 337152 277860 337204
rect 277912 337192 277918 337204
rect 278406 337192 278412 337204
rect 277912 337164 278412 337192
rect 277912 337152 277918 337164
rect 278406 337152 278412 337164
rect 278464 337152 278470 337204
rect 254670 336716 254676 336728
rect 234586 336688 254676 336716
rect 231118 336608 231124 336660
rect 231176 336648 231182 336660
rect 234586 336648 234614 336688
rect 254670 336676 254676 336688
rect 254728 336676 254734 336728
rect 262950 336676 262956 336728
rect 263008 336716 263014 336728
rect 265710 336716 265716 336728
rect 263008 336688 265716 336716
rect 263008 336676 263014 336688
rect 265710 336676 265716 336688
rect 265768 336676 265774 336728
rect 293402 336676 293408 336728
rect 293460 336716 293466 336728
rect 312538 336716 312544 336728
rect 293460 336688 312544 336716
rect 293460 336676 293466 336688
rect 312538 336676 312544 336688
rect 312596 336676 312602 336728
rect 231176 336620 234614 336648
rect 239401 336651 239459 336657
rect 231176 336608 231182 336620
rect 239401 336617 239413 336651
rect 239447 336648 239459 336651
rect 249061 336651 249119 336657
rect 249061 336648 249073 336651
rect 239447 336620 249073 336648
rect 239447 336617 239459 336620
rect 239401 336611 239459 336617
rect 249061 336617 249073 336620
rect 249107 336617 249119 336651
rect 249061 336611 249119 336617
rect 272518 336608 272524 336660
rect 272576 336648 272582 336660
rect 272576 336620 273254 336648
rect 272576 336608 272582 336620
rect 226978 336540 226984 336592
rect 227036 336580 227042 336592
rect 248969 336583 249027 336589
rect 248969 336580 248981 336583
rect 227036 336552 248981 336580
rect 227036 336540 227042 336552
rect 248969 336549 248981 336552
rect 249015 336549 249027 336583
rect 273226 336580 273254 336620
rect 274634 336608 274640 336660
rect 274692 336648 274698 336660
rect 287701 336651 287759 336657
rect 287701 336648 287713 336651
rect 274692 336620 287713 336648
rect 274692 336608 274698 336620
rect 287701 336617 287713 336620
rect 287747 336617 287759 336651
rect 287701 336611 287759 336617
rect 292485 336583 292543 336589
rect 292485 336580 292497 336583
rect 273226 336552 292497 336580
rect 248969 336543 249027 336549
rect 292485 336549 292497 336552
rect 292531 336549 292543 336583
rect 292485 336543 292543 336549
rect 224218 336472 224224 336524
rect 224276 336512 224282 336524
rect 261478 336512 261484 336524
rect 224276 336484 261484 336512
rect 224276 336472 224282 336484
rect 261478 336472 261484 336484
rect 261536 336472 261542 336524
rect 275557 336515 275615 336521
rect 275557 336481 275569 336515
rect 275603 336512 275615 336515
rect 288434 336512 288440 336524
rect 275603 336484 288440 336512
rect 275603 336481 275615 336484
rect 275557 336475 275615 336481
rect 288434 336472 288440 336484
rect 288492 336472 288498 336524
rect 294690 336472 294696 336524
rect 294748 336512 294754 336524
rect 320818 336512 320824 336524
rect 294748 336484 320824 336512
rect 294748 336472 294754 336484
rect 320818 336472 320824 336484
rect 320876 336472 320882 336524
rect 125502 336404 125508 336456
rect 125560 336444 125566 336456
rect 249794 336444 249800 336456
rect 125560 336416 249800 336444
rect 125560 336404 125566 336416
rect 249794 336404 249800 336416
rect 249852 336404 249858 336456
rect 254581 336447 254639 336453
rect 254581 336413 254593 336447
rect 254627 336444 254639 336447
rect 263778 336444 263784 336456
rect 254627 336416 263784 336444
rect 254627 336413 254639 336416
rect 254581 336407 254639 336413
rect 263778 336404 263784 336416
rect 263836 336404 263842 336456
rect 271138 336404 271144 336456
rect 271196 336444 271202 336456
rect 287609 336447 287667 336453
rect 287609 336444 287621 336447
rect 271196 336416 287621 336444
rect 271196 336404 271202 336416
rect 287609 336413 287621 336416
rect 287655 336413 287667 336447
rect 287609 336407 287667 336413
rect 295518 336404 295524 336456
rect 295576 336444 295582 336456
rect 322198 336444 322204 336456
rect 295576 336416 322204 336444
rect 295576 336404 295582 336416
rect 322198 336404 322204 336416
rect 322256 336404 322262 336456
rect 114462 336336 114468 336388
rect 114520 336376 114526 336388
rect 248598 336376 248604 336388
rect 114520 336348 248604 336376
rect 114520 336336 114526 336348
rect 248598 336336 248604 336348
rect 248656 336336 248662 336388
rect 249061 336379 249119 336385
rect 249061 336345 249073 336379
rect 249107 336376 249119 336379
rect 255498 336376 255504 336388
rect 249107 336348 255504 336376
rect 249107 336345 249119 336348
rect 249061 336339 249119 336345
rect 255498 336336 255504 336348
rect 255556 336336 255562 336388
rect 297266 336376 297272 336388
rect 278056 336348 297272 336376
rect 35158 336268 35164 336320
rect 35216 336308 35222 336320
rect 238386 336308 238392 336320
rect 35216 336280 238392 336308
rect 35216 336268 35222 336280
rect 238386 336268 238392 336280
rect 238444 336268 238450 336320
rect 253198 336268 253204 336320
rect 253256 336308 253262 336320
rect 253256 336280 256326 336308
rect 253256 336268 253262 336280
rect 28258 336200 28264 336252
rect 28316 336240 28322 336252
rect 236270 336240 236276 336252
rect 28316 336212 236276 336240
rect 28316 336200 28322 336212
rect 236270 336200 236276 336212
rect 236328 336200 236334 336252
rect 248969 336243 249027 336249
rect 248969 336209 248981 336243
rect 249015 336240 249027 336243
rect 254397 336243 254455 336249
rect 254397 336240 254409 336243
rect 249015 336212 254409 336240
rect 249015 336209 249027 336212
rect 248969 336203 249027 336209
rect 254397 336209 254409 336212
rect 254443 336209 254455 336243
rect 256298 336240 256326 336280
rect 261478 336268 261484 336320
rect 261536 336308 261542 336320
rect 263962 336308 263968 336320
rect 261536 336280 263968 336308
rect 261536 336268 261542 336280
rect 263962 336268 263968 336280
rect 264020 336268 264026 336320
rect 270678 336268 270684 336320
rect 270736 336308 270742 336320
rect 278056 336308 278084 336348
rect 297266 336336 297272 336348
rect 297324 336336 297330 336388
rect 307018 336336 307024 336388
rect 307076 336376 307082 336388
rect 307202 336376 307208 336388
rect 307076 336348 307208 336376
rect 307076 336336 307082 336348
rect 307202 336336 307208 336348
rect 307260 336336 307266 336388
rect 270736 336280 278084 336308
rect 278133 336311 278191 336317
rect 270736 336268 270742 336280
rect 278133 336277 278145 336311
rect 278179 336308 278191 336311
rect 284757 336311 284815 336317
rect 284757 336308 284769 336311
rect 278179 336280 284769 336308
rect 278179 336277 278191 336280
rect 278133 336271 278191 336277
rect 284757 336277 284769 336280
rect 284803 336277 284815 336311
rect 284757 336271 284815 336277
rect 290366 336268 290372 336320
rect 290424 336308 290430 336320
rect 327718 336308 327724 336320
rect 290424 336280 297404 336308
rect 290424 336268 290430 336280
rect 264146 336240 264152 336252
rect 256298 336212 264152 336240
rect 254397 336203 254455 336209
rect 264146 336200 264152 336212
rect 264204 336200 264210 336252
rect 278225 336243 278283 336249
rect 278225 336209 278237 336243
rect 278271 336240 278283 336243
rect 296625 336243 296683 336249
rect 296625 336240 296637 336243
rect 278271 336212 296637 336240
rect 278271 336209 278283 336212
rect 278225 336203 278283 336209
rect 296625 336209 296637 336212
rect 296671 336209 296683 336243
rect 296625 336203 296683 336209
rect 21358 336132 21364 336184
rect 21416 336172 21422 336184
rect 237190 336172 237196 336184
rect 21416 336144 237196 336172
rect 21416 336132 21422 336144
rect 237190 336132 237196 336144
rect 237248 336132 237254 336184
rect 249610 336132 249616 336184
rect 249668 336172 249674 336184
rect 264698 336172 264704 336184
rect 249668 336144 264704 336172
rect 249668 336132 249674 336144
rect 264698 336132 264704 336144
rect 264756 336132 264762 336184
rect 270218 336132 270224 336184
rect 270276 336172 270282 336184
rect 278133 336175 278191 336181
rect 278133 336172 278145 336175
rect 270276 336144 278145 336172
rect 270276 336132 270282 336144
rect 278133 336141 278145 336144
rect 278179 336141 278191 336175
rect 278133 336135 278191 336141
rect 284757 336175 284815 336181
rect 284757 336141 284769 336175
rect 284803 336172 284815 336175
rect 292942 336172 292948 336184
rect 284803 336144 292948 336172
rect 284803 336141 284815 336144
rect 284757 336135 284815 336141
rect 292942 336132 292948 336144
rect 293000 336132 293006 336184
rect 297376 336172 297404 336280
rect 311866 336280 327724 336308
rect 297634 336200 297640 336252
rect 297692 336240 297698 336252
rect 311866 336240 311894 336280
rect 327718 336268 327724 336280
rect 327776 336268 327782 336320
rect 297692 336212 311894 336240
rect 297692 336200 297698 336212
rect 335998 336172 336004 336184
rect 297376 336144 336004 336172
rect 335998 336132 336004 336144
rect 336056 336132 336062 336184
rect 18598 336064 18604 336116
rect 18656 336104 18662 336116
rect 236089 336107 236147 336113
rect 236089 336104 236101 336107
rect 18656 336076 236101 336104
rect 18656 336064 18662 336076
rect 236089 336073 236101 336076
rect 236135 336073 236147 336107
rect 236089 336067 236147 336073
rect 252462 336064 252468 336116
rect 252520 336104 252526 336116
rect 258721 336107 258779 336113
rect 258721 336104 258733 336107
rect 252520 336076 258733 336104
rect 252520 336064 252526 336076
rect 258721 336073 258733 336076
rect 258767 336073 258779 336107
rect 258721 336067 258779 336073
rect 258813 336107 258871 336113
rect 258813 336073 258825 336107
rect 258859 336104 258871 336107
rect 265250 336104 265256 336116
rect 258859 336076 265256 336104
rect 258859 336073 258871 336076
rect 258813 336067 258871 336073
rect 265250 336064 265256 336076
rect 265308 336064 265314 336116
rect 269390 336064 269396 336116
rect 269448 336104 269454 336116
rect 278041 336107 278099 336113
rect 278041 336104 278053 336107
rect 269448 336076 278053 336104
rect 269448 336064 269454 336076
rect 278041 336073 278053 336076
rect 278087 336073 278099 336107
rect 278041 336067 278099 336073
rect 284018 336064 284024 336116
rect 284076 336104 284082 336116
rect 400858 336104 400864 336116
rect 284076 336076 400864 336104
rect 284076 336064 284082 336076
rect 400858 336064 400864 336076
rect 400916 336064 400922 336116
rect 10318 335996 10324 336048
rect 10376 336036 10382 336048
rect 235534 336036 235540 336048
rect 10376 336008 235540 336036
rect 10376 335996 10382 336008
rect 235534 335996 235540 336008
rect 235592 335996 235598 336048
rect 245470 335996 245476 336048
rect 245528 336036 245534 336048
rect 264238 336036 264244 336048
rect 245528 336008 258672 336036
rect 245528 335996 245534 336008
rect 233970 335928 233976 335980
rect 234028 335968 234034 335980
rect 257614 335968 257620 335980
rect 234028 335940 257620 335968
rect 234028 335928 234034 335940
rect 257614 335928 257620 335940
rect 257672 335928 257678 335980
rect 258644 335968 258672 336008
rect 258828 336008 264244 336036
rect 258828 335968 258856 336008
rect 264238 335996 264244 336008
rect 264296 335996 264302 336048
rect 269942 335996 269948 336048
rect 270000 336036 270006 336048
rect 287054 336036 287060 336048
rect 270000 336008 287060 336036
rect 270000 335996 270006 336008
rect 287054 335996 287060 336008
rect 287112 335996 287118 336048
rect 292574 335996 292580 336048
rect 292632 336036 292638 336048
rect 479518 336036 479524 336048
rect 292632 336008 479524 336036
rect 292632 335996 292638 336008
rect 479518 335996 479524 336008
rect 479576 335996 479582 336048
rect 265158 335968 265164 335980
rect 258644 335940 258856 335968
rect 263566 335940 265164 335968
rect 233878 335860 233884 335912
rect 233936 335900 233942 335912
rect 254210 335900 254216 335912
rect 233936 335872 254216 335900
rect 233936 335860 233942 335872
rect 254210 335860 254216 335872
rect 254268 335860 254274 335912
rect 255866 335860 255872 335912
rect 255924 335900 255930 335912
rect 258813 335903 258871 335909
rect 258813 335900 258825 335903
rect 255924 335872 258825 335900
rect 255924 335860 255930 335872
rect 258813 335869 258825 335872
rect 258859 335869 258871 335903
rect 258813 335863 258871 335869
rect 234062 335792 234068 335844
rect 234120 335832 234126 335844
rect 244093 335835 244151 335841
rect 244093 335832 244105 335835
rect 234120 335804 244105 335832
rect 234120 335792 234126 335804
rect 244093 335801 244105 335804
rect 244139 335801 244151 335835
rect 244093 335795 244151 335801
rect 258721 335835 258779 335841
rect 258721 335801 258733 335835
rect 258767 335832 258779 335835
rect 263566 335832 263594 335940
rect 265158 335928 265164 335940
rect 265216 335928 265222 335980
rect 287701 335971 287759 335977
rect 287701 335937 287713 335971
rect 287747 335968 287759 335971
rect 294138 335968 294144 335980
rect 287747 335940 294144 335968
rect 287747 335937 287759 335940
rect 287701 335931 287759 335937
rect 294138 335928 294144 335940
rect 294196 335928 294202 335980
rect 294230 335928 294236 335980
rect 294288 335968 294294 335980
rect 313918 335968 313924 335980
rect 294288 335940 313924 335968
rect 294288 335928 294294 335940
rect 313918 335928 313924 335940
rect 313976 335928 313982 335980
rect 268470 335860 268476 335912
rect 268528 335900 268534 335912
rect 273898 335900 273904 335912
rect 268528 335872 273904 335900
rect 268528 335860 268534 335872
rect 273898 335860 273904 335872
rect 273956 335860 273962 335912
rect 293034 335860 293040 335912
rect 293092 335900 293098 335912
rect 302053 335903 302111 335909
rect 302053 335900 302065 335903
rect 293092 335872 302065 335900
rect 293092 335860 293098 335872
rect 302053 335869 302065 335872
rect 302099 335869 302111 335903
rect 302053 335863 302111 335869
rect 302605 335903 302663 335909
rect 302605 335869 302617 335903
rect 302651 335900 302663 335903
rect 305730 335900 305736 335912
rect 302651 335872 305736 335900
rect 302651 335869 302663 335872
rect 302605 335863 302663 335869
rect 305730 335860 305736 335872
rect 305788 335860 305794 335912
rect 307018 335900 307024 335912
rect 306979 335872 307024 335900
rect 307018 335860 307024 335872
rect 307076 335860 307082 335912
rect 258767 335804 263594 335832
rect 258767 335801 258779 335804
rect 258721 335795 258779 335801
rect 268562 335792 268568 335844
rect 268620 335832 268626 335844
rect 276658 335832 276664 335844
rect 268620 335804 276664 335832
rect 268620 335792 268626 335804
rect 276658 335792 276664 335804
rect 276716 335792 276722 335844
rect 282362 335792 282368 335844
rect 282420 335832 282426 335844
rect 282822 335832 282828 335844
rect 282420 335804 282828 335832
rect 282420 335792 282426 335804
rect 282822 335792 282828 335804
rect 282880 335792 282886 335844
rect 284478 335792 284484 335844
rect 284536 335832 284542 335844
rect 294414 335832 294420 335844
rect 284536 335804 294420 335832
rect 284536 335792 284542 335804
rect 294414 335792 294420 335804
rect 294472 335792 294478 335844
rect 296625 335835 296683 335841
rect 296625 335801 296637 335835
rect 296671 335832 296683 335835
rect 300305 335835 300363 335841
rect 300305 335832 300317 335835
rect 296671 335804 300317 335832
rect 296671 335801 296683 335804
rect 296625 335795 296683 335801
rect 300305 335801 300317 335804
rect 300351 335801 300363 335835
rect 300305 335795 300363 335801
rect 301590 335792 301596 335844
rect 301648 335832 301654 335844
rect 302142 335832 302148 335844
rect 301648 335804 302148 335832
rect 301648 335792 301654 335804
rect 302142 335792 302148 335804
rect 302200 335792 302206 335844
rect 302329 335835 302387 335841
rect 302329 335801 302341 335835
rect 302375 335832 302387 335835
rect 305086 335832 305092 335844
rect 302375 335804 305092 335832
rect 302375 335801 302387 335804
rect 302329 335795 302387 335801
rect 305086 335792 305092 335804
rect 305144 335792 305150 335844
rect 229738 335724 229744 335776
rect 229796 335764 229802 335776
rect 239401 335767 239459 335773
rect 239401 335764 239413 335767
rect 229796 335736 239413 335764
rect 229796 335724 229802 335736
rect 239401 335733 239413 335736
rect 239447 335733 239459 335767
rect 239401 335727 239459 335733
rect 267458 335724 267464 335776
rect 267516 335764 267522 335776
rect 270494 335764 270500 335776
rect 267516 335736 270500 335764
rect 267516 335724 267522 335736
rect 270494 335724 270500 335736
rect 270552 335724 270558 335776
rect 278774 335724 278780 335776
rect 278832 335764 278838 335776
rect 282457 335767 282515 335773
rect 282457 335764 282469 335767
rect 278832 335736 282469 335764
rect 278832 335724 278838 335736
rect 282457 335733 282469 335736
rect 282503 335733 282515 335767
rect 282457 335727 282515 335733
rect 283006 335724 283012 335776
rect 283064 335764 283070 335776
rect 283650 335764 283656 335776
rect 283064 335736 283656 335764
rect 283064 335724 283070 335736
rect 283650 335724 283656 335736
rect 283708 335724 283714 335776
rect 293770 335724 293776 335776
rect 293828 335764 293834 335776
rect 306282 335764 306288 335776
rect 293828 335736 306288 335764
rect 293828 335724 293834 335736
rect 306282 335724 306288 335736
rect 306340 335724 306346 335776
rect 283374 335656 283380 335708
rect 283432 335696 283438 335708
rect 283558 335696 283564 335708
rect 283432 335668 283564 335696
rect 283432 335656 283438 335668
rect 283558 335656 283564 335668
rect 283616 335656 283622 335708
rect 290090 335656 290096 335708
rect 290148 335696 290154 335708
rect 292758 335696 292764 335708
rect 290148 335668 292764 335696
rect 290148 335656 290154 335668
rect 292758 335656 292764 335668
rect 292816 335656 292822 335708
rect 296806 335656 296812 335708
rect 296864 335696 296870 335708
rect 302329 335699 302387 335705
rect 302329 335696 302341 335699
rect 296864 335668 302341 335696
rect 296864 335656 296870 335668
rect 302329 335665 302341 335668
rect 302375 335665 302387 335699
rect 302329 335659 302387 335665
rect 302421 335699 302479 335705
rect 302421 335665 302433 335699
rect 302467 335696 302479 335699
rect 305178 335696 305184 335708
rect 302467 335668 305184 335696
rect 302467 335665 302479 335668
rect 302421 335659 302479 335665
rect 305178 335656 305184 335668
rect 305236 335656 305242 335708
rect 273530 335588 273536 335640
rect 273588 335628 273594 335640
rect 273806 335628 273812 335640
rect 273588 335600 273812 335628
rect 273588 335588 273594 335600
rect 273806 335588 273812 335600
rect 273864 335588 273870 335640
rect 280614 335588 280620 335640
rect 280672 335628 280678 335640
rect 281258 335628 281264 335640
rect 280672 335600 281264 335628
rect 280672 335588 280678 335600
rect 281258 335588 281264 335600
rect 281316 335588 281322 335640
rect 281718 335588 281724 335640
rect 281776 335628 281782 335640
rect 284662 335628 284668 335640
rect 281776 335600 284668 335628
rect 281776 335588 281782 335600
rect 284662 335588 284668 335600
rect 284720 335588 284726 335640
rect 287609 335631 287667 335637
rect 287609 335597 287621 335631
rect 287655 335628 287667 335631
rect 293402 335628 293408 335640
rect 287655 335600 293408 335628
rect 287655 335597 287667 335600
rect 287609 335591 287667 335597
rect 293402 335588 293408 335600
rect 293460 335588 293466 335640
rect 302145 335631 302203 335637
rect 302145 335597 302157 335631
rect 302191 335628 302203 335631
rect 302605 335631 302663 335637
rect 302605 335628 302617 335631
rect 302191 335600 302617 335628
rect 302191 335597 302203 335600
rect 302145 335591 302203 335597
rect 302605 335597 302617 335600
rect 302651 335597 302663 335631
rect 302605 335591 302663 335597
rect 302694 335588 302700 335640
rect 302752 335628 302758 335640
rect 303522 335628 303528 335640
rect 302752 335600 303528 335628
rect 302752 335588 302758 335600
rect 303522 335588 303528 335600
rect 303580 335588 303586 335640
rect 267550 335520 267556 335572
rect 267608 335560 267614 335572
rect 268378 335560 268384 335572
rect 267608 335532 268384 335560
rect 267608 335520 267614 335532
rect 268378 335520 268384 335532
rect 268436 335520 268442 335572
rect 278041 335563 278099 335569
rect 278041 335529 278053 335563
rect 278087 335560 278099 335563
rect 285861 335563 285919 335569
rect 285861 335560 285873 335563
rect 278087 335532 285873 335560
rect 278087 335529 278099 335532
rect 278041 335523 278099 335529
rect 285861 335529 285873 335532
rect 285907 335529 285919 335563
rect 285861 335523 285919 335529
rect 294782 335520 294788 335572
rect 294840 335560 294846 335572
rect 295242 335560 295248 335572
rect 294840 335532 295248 335560
rect 294840 335520 294846 335532
rect 295242 335520 295248 335532
rect 295300 335520 295306 335572
rect 297174 335520 297180 335572
rect 297232 335560 297238 335572
rect 297232 335532 300532 335560
rect 297232 335520 297238 335532
rect 272610 335452 272616 335504
rect 272668 335492 272674 335504
rect 273070 335492 273076 335504
rect 272668 335464 273076 335492
rect 272668 335452 272674 335464
rect 273070 335452 273076 335464
rect 273128 335452 273134 335504
rect 273806 335452 273812 335504
rect 273864 335492 273870 335504
rect 274358 335492 274364 335504
rect 273864 335464 274364 335492
rect 273864 335452 273870 335464
rect 274358 335452 274364 335464
rect 274416 335452 274422 335504
rect 283926 335492 283932 335504
rect 283024 335464 283932 335492
rect 236730 335384 236736 335436
rect 236788 335424 236794 335436
rect 243446 335424 243452 335436
rect 236788 335396 243452 335424
rect 236788 335384 236794 335396
rect 243446 335384 243452 335396
rect 243504 335384 243510 335436
rect 257338 335384 257344 335436
rect 257396 335424 257402 335436
rect 263318 335424 263324 335436
rect 257396 335396 263324 335424
rect 257396 335384 257402 335396
rect 263318 335384 263324 335396
rect 263376 335384 263382 335436
rect 266998 335384 267004 335436
rect 267056 335424 267062 335436
rect 267550 335424 267556 335436
rect 267056 335396 267556 335424
rect 267056 335384 267062 335396
rect 267550 335384 267556 335396
rect 267608 335384 267614 335436
rect 268286 335384 268292 335436
rect 268344 335424 268350 335436
rect 268746 335424 268752 335436
rect 268344 335396 268752 335424
rect 268344 335384 268350 335396
rect 268746 335384 268752 335396
rect 268804 335384 268810 335436
rect 272242 335384 272248 335436
rect 272300 335424 272306 335436
rect 272978 335424 272984 335436
rect 272300 335396 272984 335424
rect 272300 335384 272306 335396
rect 272978 335384 272984 335396
rect 273036 335384 273042 335436
rect 274910 335384 274916 335436
rect 274968 335424 274974 335436
rect 275738 335424 275744 335436
rect 274968 335396 275744 335424
rect 274968 335384 274974 335396
rect 275738 335384 275744 335396
rect 275796 335384 275802 335436
rect 276474 335384 276480 335436
rect 276532 335424 276538 335436
rect 277302 335424 277308 335436
rect 276532 335396 277308 335424
rect 276532 335384 276538 335396
rect 277302 335384 277308 335396
rect 277360 335384 277366 335436
rect 277486 335384 277492 335436
rect 277544 335424 277550 335436
rect 278222 335424 278228 335436
rect 277544 335396 278228 335424
rect 277544 335384 277550 335396
rect 278222 335384 278228 335396
rect 278280 335384 278286 335436
rect 255314 335316 255320 335368
rect 255372 335356 255378 335368
rect 256786 335356 256792 335368
rect 255372 335328 256792 335356
rect 255372 335316 255378 335328
rect 256786 335316 256792 335328
rect 256844 335316 256850 335368
rect 261018 335356 261024 335368
rect 257494 335328 261024 335356
rect 226242 335044 226248 335096
rect 226300 335084 226306 335096
rect 257341 335087 257399 335093
rect 257341 335084 257353 335087
rect 226300 335056 257353 335084
rect 226300 335044 226306 335056
rect 257341 335053 257353 335056
rect 257387 335053 257399 335087
rect 257341 335047 257399 335053
rect 219342 334976 219348 335028
rect 219400 335016 219406 335028
rect 257494 335016 257522 335328
rect 261018 335316 261024 335328
rect 261076 335316 261082 335368
rect 261570 335316 261576 335368
rect 261628 335356 261634 335368
rect 263042 335356 263048 335368
rect 261628 335328 263048 335356
rect 261628 335316 261634 335328
rect 263042 335316 263048 335328
rect 263100 335316 263106 335368
rect 267826 335316 267832 335368
rect 267884 335356 267890 335368
rect 268562 335356 268568 335368
rect 267884 335328 268568 335356
rect 267884 335316 267890 335328
rect 268562 335316 268568 335328
rect 268620 335316 268626 335368
rect 269942 335316 269948 335368
rect 270000 335356 270006 335368
rect 270402 335356 270408 335368
rect 270000 335328 270408 335356
rect 270000 335316 270006 335328
rect 270402 335316 270408 335328
rect 270460 335316 270466 335368
rect 271506 335316 271512 335368
rect 271564 335356 271570 335368
rect 271782 335356 271788 335368
rect 271564 335328 271788 335356
rect 271564 335316 271570 335328
rect 271782 335316 271788 335328
rect 271840 335316 271846 335368
rect 275462 335316 275468 335368
rect 275520 335356 275526 335368
rect 275922 335356 275928 335368
rect 275520 335328 275928 335356
rect 275520 335316 275526 335328
rect 275922 335316 275928 335328
rect 275980 335316 275986 335368
rect 276198 335316 276204 335368
rect 276256 335356 276262 335368
rect 276934 335356 276940 335368
rect 276256 335328 276940 335356
rect 276256 335316 276262 335328
rect 276934 335316 276940 335328
rect 276992 335316 276998 335368
rect 280706 335316 280712 335368
rect 280764 335356 280770 335368
rect 280890 335356 280896 335368
rect 280764 335328 280896 335356
rect 280764 335316 280770 335328
rect 280890 335316 280896 335328
rect 280948 335316 280954 335368
rect 281994 335316 282000 335368
rect 282052 335356 282058 335368
rect 282270 335356 282276 335368
rect 282052 335328 282276 335356
rect 282052 335316 282058 335328
rect 282270 335316 282276 335328
rect 282328 335316 282334 335368
rect 282457 335359 282515 335365
rect 282457 335325 282469 335359
rect 282503 335356 282515 335359
rect 283024 335356 283052 335464
rect 283926 335452 283932 335464
rect 283984 335452 283990 335504
rect 284478 335452 284484 335504
rect 284536 335492 284542 335504
rect 284846 335492 284852 335504
rect 284536 335464 284852 335492
rect 284536 335452 284542 335464
rect 284846 335452 284852 335464
rect 284904 335452 284910 335504
rect 287790 335452 287796 335504
rect 287848 335492 287854 335504
rect 288342 335492 288348 335504
rect 287848 335464 288348 335492
rect 287848 335452 287854 335464
rect 288342 335452 288348 335464
rect 288400 335452 288406 335504
rect 291930 335452 291936 335504
rect 291988 335492 291994 335504
rect 292298 335492 292304 335504
rect 291988 335464 292304 335492
rect 291988 335452 291994 335464
rect 292298 335452 292304 335464
rect 292356 335452 292362 335504
rect 292485 335495 292543 335501
rect 292485 335461 292497 335495
rect 292531 335492 292543 335495
rect 292531 335464 295288 335492
rect 292531 335461 292543 335464
rect 292485 335455 292543 335461
rect 283282 335384 283288 335436
rect 283340 335424 283346 335436
rect 284202 335424 284208 335436
rect 283340 335396 284208 335424
rect 283340 335384 283346 335396
rect 284202 335384 284208 335396
rect 284260 335384 284266 335436
rect 286502 335384 286508 335436
rect 286560 335424 286566 335436
rect 286962 335424 286968 335436
rect 286560 335396 286968 335424
rect 286560 335384 286566 335396
rect 286962 335384 286968 335396
rect 287020 335384 287026 335436
rect 289814 335384 289820 335436
rect 289872 335424 289878 335436
rect 290826 335424 290832 335436
rect 289872 335396 290832 335424
rect 289872 335384 289878 335396
rect 290826 335384 290832 335396
rect 290884 335384 290890 335436
rect 291654 335384 291660 335436
rect 291712 335424 291718 335436
rect 292022 335424 292028 335436
rect 291712 335396 292028 335424
rect 291712 335384 291718 335396
rect 292022 335384 292028 335396
rect 292080 335384 292086 335436
rect 282503 335328 283052 335356
rect 282503 335325 282515 335328
rect 282457 335319 282515 335325
rect 284570 335316 284576 335368
rect 284628 335356 284634 335368
rect 284628 335328 284892 335356
rect 284628 335316 284634 335328
rect 284864 335220 284892 335328
rect 284938 335316 284944 335368
rect 284996 335356 285002 335368
rect 285122 335356 285128 335368
rect 284996 335328 285128 335356
rect 284996 335316 285002 335328
rect 285122 335316 285128 335328
rect 285180 335316 285186 335368
rect 285214 335316 285220 335368
rect 285272 335356 285278 335368
rect 285398 335356 285404 335368
rect 285272 335328 285404 335356
rect 285272 335316 285278 335328
rect 285398 335316 285404 335328
rect 285456 335316 285462 335368
rect 286134 335316 286140 335368
rect 286192 335356 286198 335368
rect 286192 335328 286364 335356
rect 286192 335316 286198 335328
rect 285122 335220 285128 335232
rect 284864 335192 285128 335220
rect 285122 335180 285128 335192
rect 285180 335180 285186 335232
rect 286336 335220 286364 335328
rect 286410 335316 286416 335368
rect 286468 335356 286474 335368
rect 286778 335356 286784 335368
rect 286468 335328 286784 335356
rect 286468 335316 286474 335328
rect 286778 335316 286784 335328
rect 286836 335316 286842 335368
rect 287238 335316 287244 335368
rect 287296 335356 287302 335368
rect 287296 335328 287468 335356
rect 287296 335316 287302 335328
rect 287440 335288 287468 335328
rect 287514 335316 287520 335368
rect 287572 335356 287578 335368
rect 287698 335356 287704 335368
rect 287572 335328 287704 335356
rect 287572 335316 287578 335328
rect 287698 335316 287704 335328
rect 287756 335316 287762 335368
rect 287974 335316 287980 335368
rect 288032 335356 288038 335368
rect 288342 335356 288348 335368
rect 288032 335328 288348 335356
rect 288032 335316 288038 335328
rect 288342 335316 288348 335328
rect 288400 335316 288406 335368
rect 289078 335316 289084 335368
rect 289136 335356 289142 335368
rect 289262 335356 289268 335368
rect 289136 335328 289268 335356
rect 289136 335316 289142 335328
rect 289262 335316 289268 335328
rect 289320 335316 289326 335368
rect 290642 335316 290648 335368
rect 290700 335356 290706 335368
rect 291010 335356 291016 335368
rect 290700 335328 291016 335356
rect 290700 335316 290706 335328
rect 291010 335316 291016 335328
rect 291068 335316 291074 335368
rect 291378 335316 291384 335368
rect 291436 335356 291442 335368
rect 291838 335356 291844 335368
rect 291436 335328 291844 335356
rect 291436 335316 291442 335328
rect 291838 335316 291844 335328
rect 291896 335316 291902 335368
rect 291930 335316 291936 335368
rect 291988 335356 291994 335368
rect 292206 335356 292212 335368
rect 291988 335328 292212 335356
rect 291988 335316 291994 335328
rect 292206 335316 292212 335328
rect 292264 335316 292270 335368
rect 294046 335316 294052 335368
rect 294104 335356 294110 335368
rect 294690 335356 294696 335368
rect 294104 335328 294696 335356
rect 294104 335316 294110 335328
rect 294690 335316 294696 335328
rect 294748 335316 294754 335368
rect 288158 335288 288164 335300
rect 287440 335260 288164 335288
rect 288158 335248 288164 335260
rect 288216 335248 288222 335300
rect 295260 335288 295288 335464
rect 295886 335452 295892 335504
rect 295944 335492 295950 335504
rect 296438 335492 296444 335504
rect 295944 335464 296444 335492
rect 295944 335452 295950 335464
rect 296438 335452 296444 335464
rect 296496 335452 296502 335504
rect 298462 335452 298468 335504
rect 298520 335492 298526 335504
rect 299474 335492 299480 335504
rect 298520 335464 299480 335492
rect 298520 335452 298526 335464
rect 299474 335452 299480 335464
rect 299532 335452 299538 335504
rect 299566 335452 299572 335504
rect 299624 335492 299630 335504
rect 300302 335492 300308 335504
rect 299624 335464 300308 335492
rect 299624 335452 299630 335464
rect 300302 335452 300308 335464
rect 300360 335452 300366 335504
rect 295978 335384 295984 335436
rect 296036 335424 296042 335436
rect 296346 335424 296352 335436
rect 296036 335396 296352 335424
rect 296036 335384 296042 335396
rect 296346 335384 296352 335396
rect 296404 335384 296410 335436
rect 298738 335384 298744 335436
rect 298796 335424 298802 335436
rect 299014 335424 299020 335436
rect 298796 335396 299020 335424
rect 298796 335384 298802 335396
rect 299014 335384 299020 335396
rect 299072 335384 299078 335436
rect 300504 335424 300532 335532
rect 301406 335520 301412 335572
rect 301464 335560 301470 335572
rect 302050 335560 302056 335572
rect 301464 335532 302056 335560
rect 301464 335520 301470 335532
rect 302050 335520 302056 335532
rect 302108 335520 302114 335572
rect 301130 335452 301136 335504
rect 301188 335492 301194 335504
rect 301774 335492 301780 335504
rect 301188 335464 301780 335492
rect 301188 335452 301194 335464
rect 301774 335452 301780 335464
rect 301832 335452 301838 335504
rect 302970 335452 302976 335504
rect 303028 335492 303034 335504
rect 303522 335492 303528 335504
rect 303028 335464 303528 335492
rect 303028 335452 303034 335464
rect 303522 335452 303528 335464
rect 303580 335452 303586 335504
rect 302329 335427 302387 335433
rect 302329 335424 302341 335427
rect 300504 335396 302341 335424
rect 302329 335393 302341 335396
rect 302375 335393 302387 335427
rect 302329 335387 302387 335393
rect 302418 335384 302424 335436
rect 302476 335424 302482 335436
rect 303062 335424 303068 335436
rect 302476 335396 303068 335424
rect 302476 335384 302482 335396
rect 303062 335384 303068 335396
rect 303120 335384 303126 335436
rect 304534 335384 304540 335436
rect 304592 335424 304598 335436
rect 304902 335424 304908 335436
rect 304592 335396 304908 335424
rect 304592 335384 304598 335396
rect 304902 335384 304908 335396
rect 304960 335384 304966 335436
rect 295334 335316 295340 335368
rect 295392 335356 295398 335368
rect 295886 335356 295892 335368
rect 295392 335328 295892 335356
rect 295392 335316 295398 335328
rect 295886 335316 295892 335328
rect 295944 335316 295950 335368
rect 297450 335316 297456 335368
rect 297508 335356 297514 335368
rect 297910 335356 297916 335368
rect 297508 335328 297916 335356
rect 297508 335316 297514 335328
rect 297910 335316 297916 335328
rect 297968 335316 297974 335368
rect 299198 335316 299204 335368
rect 299256 335356 299262 335368
rect 299382 335356 299388 335368
rect 299256 335328 299388 335356
rect 299256 335316 299262 335328
rect 299382 335316 299388 335328
rect 299440 335316 299446 335368
rect 300854 335316 300860 335368
rect 300912 335356 300918 335368
rect 301406 335356 301412 335368
rect 300912 335328 301412 335356
rect 300912 335316 300918 335328
rect 301406 335316 301412 335328
rect 301464 335316 301470 335368
rect 301866 335316 301872 335368
rect 301924 335356 301930 335368
rect 302142 335356 302148 335368
rect 301924 335328 302148 335356
rect 301924 335316 301930 335328
rect 302142 335316 302148 335328
rect 302200 335316 302206 335368
rect 302970 335316 302976 335368
rect 303028 335356 303034 335368
rect 303246 335356 303252 335368
rect 303028 335328 303252 335356
rect 303028 335316 303034 335328
rect 303246 335316 303252 335328
rect 303304 335316 303310 335368
rect 304166 335316 304172 335368
rect 304224 335356 304230 335368
rect 304350 335356 304356 335368
rect 304224 335328 304356 335356
rect 304224 335316 304230 335328
rect 304350 335316 304356 335328
rect 304408 335316 304414 335368
rect 295260 335260 302234 335288
rect 286410 335220 286416 335232
rect 286336 335192 286416 335220
rect 286410 335180 286416 335192
rect 286468 335180 286474 335232
rect 289998 335180 290004 335232
rect 290056 335220 290062 335232
rect 294598 335220 294604 335232
rect 290056 335192 294604 335220
rect 290056 335180 290062 335192
rect 294598 335180 294604 335192
rect 294656 335180 294662 335232
rect 302206 335152 302234 335260
rect 313274 335152 313280 335164
rect 302206 335124 313280 335152
rect 313274 335112 313280 335124
rect 313332 335112 313338 335164
rect 271966 335044 271972 335096
rect 272024 335084 272030 335096
rect 307754 335084 307760 335096
rect 272024 335056 307760 335084
rect 272024 335044 272030 335056
rect 307754 335044 307760 335056
rect 307812 335044 307818 335096
rect 219400 334988 257522 335016
rect 219400 334976 219406 334988
rect 272150 334976 272156 335028
rect 272208 335016 272214 335028
rect 309134 335016 309140 335028
rect 272208 334988 309140 335016
rect 272208 334976 272214 334988
rect 309134 334976 309140 334988
rect 309192 334976 309198 335028
rect 210970 334908 210976 334960
rect 211028 334948 211034 334960
rect 260006 334948 260012 334960
rect 211028 334920 260012 334948
rect 211028 334908 211034 334920
rect 260006 334908 260012 334920
rect 260064 334908 260070 334960
rect 275094 334908 275100 334960
rect 275152 334948 275158 334960
rect 333974 334948 333980 334960
rect 275152 334920 333980 334948
rect 275152 334908 275158 334920
rect 333974 334908 333980 334920
rect 334032 334908 334038 334960
rect 176562 334840 176568 334892
rect 176620 334880 176626 334892
rect 255958 334880 255964 334892
rect 176620 334852 255964 334880
rect 176620 334840 176626 334852
rect 255958 334840 255964 334852
rect 256016 334840 256022 334892
rect 257341 334883 257399 334889
rect 257341 334849 257353 334883
rect 257387 334880 257399 334883
rect 261846 334880 261852 334892
rect 257387 334852 261852 334880
rect 257387 334849 257399 334852
rect 257341 334843 257399 334849
rect 261846 334840 261852 334852
rect 261904 334840 261910 334892
rect 275278 334840 275284 334892
rect 275336 334880 275342 334892
rect 335354 334880 335360 334892
rect 275336 334852 335360 334880
rect 275336 334840 275342 334852
rect 335354 334840 335360 334852
rect 335412 334840 335418 334892
rect 158622 334772 158628 334824
rect 158680 334812 158686 334824
rect 253842 334812 253848 334824
rect 158680 334784 253848 334812
rect 158680 334772 158686 334784
rect 253842 334772 253848 334784
rect 253900 334772 253906 334824
rect 279142 334772 279148 334824
rect 279200 334812 279206 334824
rect 368474 334812 368480 334824
rect 279200 334784 368480 334812
rect 279200 334772 279206 334784
rect 368474 334772 368480 334784
rect 368532 334772 368538 334824
rect 126882 334704 126888 334756
rect 126940 334744 126946 334756
rect 249978 334744 249984 334756
rect 126940 334716 249984 334744
rect 126940 334704 126946 334716
rect 249978 334704 249984 334716
rect 250036 334704 250042 334756
rect 293126 334704 293132 334756
rect 293184 334744 293190 334756
rect 293770 334744 293776 334756
rect 293184 334716 293776 334744
rect 293184 334704 293190 334716
rect 293770 334704 293776 334716
rect 293828 334704 293834 334756
rect 300305 334747 300363 334753
rect 300305 334713 300317 334747
rect 300351 334744 300363 334747
rect 305638 334744 305644 334756
rect 300351 334716 305644 334744
rect 300351 334713 300363 334716
rect 300305 334707 300363 334713
rect 305638 334704 305644 334716
rect 305696 334704 305702 334756
rect 306282 334704 306288 334756
rect 306340 334744 306346 334756
rect 489914 334744 489920 334756
rect 306340 334716 489920 334744
rect 306340 334704 306346 334716
rect 489914 334704 489920 334716
rect 489972 334704 489978 334756
rect 97902 334636 97908 334688
rect 97960 334676 97966 334688
rect 246574 334676 246580 334688
rect 97960 334648 246580 334676
rect 97960 334636 97966 334648
rect 246574 334636 246580 334648
rect 246632 334636 246638 334688
rect 298186 334636 298192 334688
rect 298244 334676 298250 334688
rect 525058 334676 525064 334688
rect 298244 334648 525064 334676
rect 298244 334636 298250 334648
rect 525058 334636 525064 334648
rect 525116 334636 525122 334688
rect 39298 334568 39304 334620
rect 39356 334608 39362 334620
rect 39356 334580 234614 334608
rect 39356 334568 39362 334580
rect 234586 334540 234614 334580
rect 236454 334568 236460 334620
rect 236512 334608 236518 334620
rect 236638 334608 236644 334620
rect 236512 334580 236644 334608
rect 236512 334568 236518 334580
rect 236638 334568 236644 334580
rect 236696 334568 236702 334620
rect 242894 334568 242900 334620
rect 242952 334608 242958 334620
rect 243998 334608 244004 334620
rect 242952 334580 244004 334608
rect 242952 334568 242958 334580
rect 243998 334568 244004 334580
rect 244056 334568 244062 334620
rect 248690 334568 248696 334620
rect 248748 334608 248754 334620
rect 249518 334608 249524 334620
rect 248748 334580 249524 334608
rect 248748 334568 248754 334580
rect 249518 334568 249524 334580
rect 249576 334568 249582 334620
rect 252646 334568 252652 334620
rect 252704 334608 252710 334620
rect 253382 334608 253388 334620
rect 252704 334580 253388 334608
rect 252704 334568 252710 334580
rect 253382 334568 253388 334580
rect 253440 334568 253446 334620
rect 271414 334568 271420 334620
rect 271472 334608 271478 334620
rect 271690 334608 271696 334620
rect 271472 334580 271696 334608
rect 271472 334568 271478 334580
rect 271690 334568 271696 334580
rect 271748 334568 271754 334620
rect 276474 334568 276480 334620
rect 276532 334608 276538 334620
rect 276750 334608 276756 334620
rect 276532 334580 276756 334608
rect 276532 334568 276538 334580
rect 276750 334568 276756 334580
rect 276808 334568 276814 334620
rect 284754 334568 284760 334620
rect 284812 334608 284818 334620
rect 285398 334608 285404 334620
rect 284812 334580 285404 334608
rect 284812 334568 284818 334580
rect 285398 334568 285404 334580
rect 285456 334568 285462 334620
rect 525794 334608 525800 334620
rect 302206 334580 525800 334608
rect 239490 334540 239496 334552
rect 234586 334512 239496 334540
rect 239490 334500 239496 334512
rect 239548 334500 239554 334552
rect 251450 334500 251456 334552
rect 251508 334540 251514 334552
rect 251818 334540 251824 334552
rect 251508 334512 251824 334540
rect 251508 334500 251514 334512
rect 251818 334500 251824 334512
rect 251876 334500 251882 334552
rect 265066 334500 265072 334552
rect 265124 334540 265130 334552
rect 266078 334540 266084 334552
rect 265124 334512 266084 334540
rect 265124 334500 265130 334512
rect 266078 334500 266084 334512
rect 266136 334500 266142 334552
rect 284386 334500 284392 334552
rect 284444 334540 284450 334552
rect 285490 334540 285496 334552
rect 284444 334512 285496 334540
rect 284444 334500 284450 334512
rect 285490 334500 285496 334512
rect 285548 334500 285554 334552
rect 297450 334500 297456 334552
rect 297508 334540 297514 334552
rect 297818 334540 297824 334552
rect 297508 334512 297824 334540
rect 297508 334500 297514 334512
rect 297818 334500 297824 334512
rect 297876 334500 297882 334552
rect 298002 334500 298008 334552
rect 298060 334540 298066 334552
rect 302206 334540 302234 334580
rect 525794 334568 525800 334580
rect 525852 334568 525858 334620
rect 298060 334512 302234 334540
rect 298060 334500 298066 334512
rect 304074 334500 304080 334552
rect 304132 334540 304138 334552
rect 304442 334540 304448 334552
rect 304132 334512 304448 334540
rect 304132 334500 304138 334512
rect 304442 334500 304448 334512
rect 304500 334500 304506 334552
rect 296990 334432 296996 334484
rect 297048 334472 297054 334484
rect 297542 334472 297548 334484
rect 297048 334444 297548 334472
rect 297048 334432 297054 334444
rect 297542 334432 297548 334444
rect 297600 334432 297606 334484
rect 269206 334364 269212 334416
rect 269264 334404 269270 334416
rect 269942 334404 269948 334416
rect 269264 334376 269948 334404
rect 269264 334364 269270 334376
rect 269942 334364 269948 334376
rect 270000 334364 270006 334416
rect 284938 334364 284944 334416
rect 284996 334404 285002 334416
rect 285214 334404 285220 334416
rect 284996 334376 285220 334404
rect 284996 334364 285002 334376
rect 285214 334364 285220 334376
rect 285272 334364 285278 334416
rect 285861 334407 285919 334413
rect 285861 334373 285873 334407
rect 285907 334404 285919 334407
rect 285950 334404 285956 334416
rect 285907 334376 285956 334404
rect 285907 334373 285919 334376
rect 285861 334367 285919 334373
rect 285950 334364 285956 334376
rect 286008 334364 286014 334416
rect 291562 334364 291568 334416
rect 291620 334404 291626 334416
rect 292482 334404 292488 334416
rect 291620 334376 292488 334404
rect 291620 334364 291626 334376
rect 292482 334364 292488 334376
rect 292540 334364 292546 334416
rect 292850 334364 292856 334416
rect 292908 334404 292914 334416
rect 293218 334404 293224 334416
rect 292908 334376 293224 334404
rect 292908 334364 292914 334376
rect 293218 334364 293224 334376
rect 293276 334364 293282 334416
rect 297082 334364 297088 334416
rect 297140 334404 297146 334416
rect 297818 334404 297824 334416
rect 297140 334376 297824 334404
rect 297140 334364 297146 334376
rect 297818 334364 297824 334376
rect 297876 334364 297882 334416
rect 290274 334296 290280 334348
rect 290332 334336 290338 334348
rect 291010 334336 291016 334348
rect 290332 334308 291016 334336
rect 290332 334296 290338 334308
rect 291010 334296 291016 334308
rect 291068 334296 291074 334348
rect 292758 334228 292764 334280
rect 292816 334268 292822 334280
rect 293402 334268 293408 334280
rect 292816 334240 293408 334268
rect 292816 334228 292822 334240
rect 293402 334228 293408 334240
rect 293460 334228 293466 334280
rect 230382 333616 230388 333668
rect 230440 333656 230446 333668
rect 262306 333656 262312 333668
rect 230440 333628 262312 333656
rect 230440 333616 230446 333628
rect 262306 333616 262312 333628
rect 262364 333616 262370 333668
rect 272886 333616 272892 333668
rect 272944 333656 272950 333668
rect 316034 333656 316040 333668
rect 272944 333628 316040 333656
rect 272944 333616 272950 333628
rect 316034 333616 316040 333628
rect 316092 333616 316098 333668
rect 219250 333548 219256 333600
rect 219308 333588 219314 333600
rect 261110 333588 261116 333600
rect 219308 333560 261116 333588
rect 219308 333548 219314 333560
rect 261110 333548 261116 333560
rect 261168 333548 261174 333600
rect 288434 333548 288440 333600
rect 288492 333588 288498 333600
rect 338114 333588 338120 333600
rect 288492 333560 338120 333588
rect 288492 333548 288498 333560
rect 338114 333548 338120 333560
rect 338172 333548 338178 333600
rect 183462 333480 183468 333532
rect 183520 333520 183526 333532
rect 255314 333520 255320 333532
rect 183520 333492 255320 333520
rect 183520 333480 183526 333492
rect 255314 333480 255320 333492
rect 255372 333480 255378 333532
rect 273530 333480 273536 333532
rect 273588 333520 273594 333532
rect 324314 333520 324320 333532
rect 273588 333492 324320 333520
rect 273588 333480 273594 333492
rect 324314 333480 324320 333492
rect 324372 333480 324378 333532
rect 169662 333412 169668 333464
rect 169720 333452 169726 333464
rect 255130 333452 255136 333464
rect 169720 333424 255136 333452
rect 169720 333412 169726 333424
rect 255130 333412 255136 333424
rect 255188 333412 255194 333464
rect 279602 333412 279608 333464
rect 279660 333452 279666 333464
rect 372614 333452 372620 333464
rect 279660 333424 372620 333452
rect 279660 333412 279666 333424
rect 372614 333412 372620 333424
rect 372672 333412 372678 333464
rect 144822 333344 144828 333396
rect 144880 333384 144886 333396
rect 252094 333384 252100 333396
rect 144880 333356 252100 333384
rect 144880 333344 144886 333356
rect 252094 333344 252100 333356
rect 252152 333344 252158 333396
rect 268470 333344 268476 333396
rect 268528 333384 268534 333396
rect 269022 333384 269028 333396
rect 268528 333356 269028 333384
rect 268528 333344 268534 333356
rect 269022 333344 269028 333356
rect 269080 333344 269086 333396
rect 272702 333344 272708 333396
rect 272760 333384 272766 333396
rect 273070 333384 273076 333396
rect 272760 333356 273076 333384
rect 272760 333344 272766 333356
rect 273070 333344 273076 333356
rect 273128 333344 273134 333396
rect 282178 333344 282184 333396
rect 282236 333384 282242 333396
rect 282822 333384 282828 333396
rect 282236 333356 282828 333384
rect 282236 333344 282242 333356
rect 282822 333344 282828 333356
rect 282880 333344 282886 333396
rect 286410 333344 286416 333396
rect 286468 333384 286474 333396
rect 426434 333384 426440 333396
rect 286468 333356 426440 333384
rect 286468 333344 286474 333356
rect 426434 333344 426440 333356
rect 426492 333344 426498 333396
rect 95142 333276 95148 333328
rect 95200 333316 95206 333328
rect 246206 333316 246212 333328
rect 95200 333288 246212 333316
rect 95200 333276 95206 333288
rect 246206 333276 246212 333288
rect 246264 333276 246270 333328
rect 273714 333276 273720 333328
rect 273772 333316 273778 333328
rect 274082 333316 274088 333328
rect 273772 333288 274088 333316
rect 273772 333276 273778 333288
rect 274082 333276 274088 333288
rect 274140 333276 274146 333328
rect 277946 333276 277952 333328
rect 278004 333316 278010 333328
rect 278682 333316 278688 333328
rect 278004 333288 278688 333316
rect 278004 333276 278010 333288
rect 278682 333276 278688 333288
rect 278740 333276 278746 333328
rect 279234 333276 279240 333328
rect 279292 333316 279298 333328
rect 280062 333316 280068 333328
rect 279292 333288 280068 333316
rect 279292 333276 279298 333288
rect 280062 333276 280068 333288
rect 280120 333276 280126 333328
rect 287146 333276 287152 333328
rect 287204 333316 287210 333328
rect 434714 333316 434720 333328
rect 287204 333288 434720 333316
rect 287204 333276 287210 333288
rect 434714 333276 434720 333288
rect 434772 333276 434778 333328
rect 29638 333208 29644 333260
rect 29696 333248 29702 333260
rect 237742 333248 237748 333260
rect 29696 333220 237748 333248
rect 29696 333208 29702 333220
rect 237742 333208 237748 333220
rect 237800 333208 237806 333260
rect 241514 333208 241520 333260
rect 241572 333248 241578 333260
rect 242250 333248 242256 333260
rect 241572 333220 242256 333248
rect 241572 333208 241578 333220
rect 242250 333208 242256 333220
rect 242308 333208 242314 333260
rect 245930 333208 245936 333260
rect 245988 333248 245994 333260
rect 246390 333248 246396 333260
rect 245988 333220 246396 333248
rect 245988 333208 245994 333220
rect 246390 333208 246396 333220
rect 246448 333208 246454 333260
rect 251634 333208 251640 333260
rect 251692 333248 251698 333260
rect 252002 333248 252008 333260
rect 251692 333220 252008 333248
rect 251692 333208 251698 333220
rect 252002 333208 252008 333220
rect 252060 333208 252066 333260
rect 258350 333208 258356 333260
rect 258408 333248 258414 333260
rect 258718 333248 258724 333260
rect 258408 333220 258724 333248
rect 258408 333208 258414 333220
rect 258718 333208 258724 333220
rect 258776 333208 258782 333260
rect 266630 333208 266636 333260
rect 266688 333248 266694 333260
rect 266906 333248 266912 333260
rect 266688 333220 266912 333248
rect 266688 333208 266694 333220
rect 266906 333208 266912 333220
rect 266964 333208 266970 333260
rect 267182 333208 267188 333260
rect 267240 333248 267246 333260
rect 267458 333248 267464 333260
rect 267240 333220 267464 333248
rect 267240 333208 267246 333220
rect 267458 333208 267464 333220
rect 267516 333208 267522 333260
rect 268194 333208 268200 333260
rect 268252 333248 268258 333260
rect 269022 333248 269028 333260
rect 268252 333220 269028 333248
rect 268252 333208 268258 333220
rect 269022 333208 269028 333220
rect 269080 333208 269086 333260
rect 269574 333208 269580 333260
rect 269632 333248 269638 333260
rect 270126 333248 270132 333260
rect 269632 333220 270132 333248
rect 269632 333208 269638 333220
rect 270126 333208 270132 333220
rect 270184 333208 270190 333260
rect 270862 333208 270868 333260
rect 270920 333248 270926 333260
rect 271506 333248 271512 333260
rect 270920 333220 271512 333248
rect 270920 333208 270926 333220
rect 271506 333208 271512 333220
rect 271564 333208 271570 333260
rect 272426 333208 272432 333260
rect 272484 333248 272490 333260
rect 272702 333248 272708 333260
rect 272484 333220 272708 333248
rect 272484 333208 272490 333220
rect 272702 333208 272708 333220
rect 272760 333208 272766 333260
rect 273990 333208 273996 333260
rect 274048 333248 274054 333260
rect 274358 333248 274364 333260
rect 274048 333220 274364 333248
rect 274048 333208 274054 333220
rect 274358 333208 274364 333220
rect 274416 333208 274422 333260
rect 277670 333208 277676 333260
rect 277728 333248 277734 333260
rect 278498 333248 278504 333260
rect 277728 333220 278504 333248
rect 277728 333208 277734 333220
rect 278498 333208 278504 333220
rect 278556 333208 278562 333260
rect 279326 333208 279332 333260
rect 279384 333248 279390 333260
rect 279786 333248 279792 333260
rect 279384 333220 279792 333248
rect 279384 333208 279390 333220
rect 279786 333208 279792 333220
rect 279844 333208 279850 333260
rect 280614 333208 280620 333260
rect 280672 333248 280678 333260
rect 281074 333248 281080 333260
rect 280672 333220 281080 333248
rect 280672 333208 280678 333220
rect 281074 333208 281080 333220
rect 281132 333208 281138 333260
rect 282178 333208 282184 333260
rect 282236 333248 282242 333260
rect 282638 333248 282644 333260
rect 282236 333220 282644 333248
rect 282236 333208 282242 333220
rect 282638 333208 282644 333220
rect 282696 333208 282702 333260
rect 283742 333208 283748 333260
rect 283800 333248 283806 333260
rect 284018 333248 284024 333260
rect 283800 333220 284024 333248
rect 283800 333208 283806 333220
rect 284018 333208 284024 333220
rect 284076 333208 284082 333260
rect 284846 333208 284852 333260
rect 284904 333248 284910 333260
rect 285582 333248 285588 333260
rect 284904 333220 285588 333248
rect 284904 333208 284910 333220
rect 285582 333208 285588 333220
rect 285640 333208 285646 333260
rect 286134 333208 286140 333260
rect 286192 333248 286198 333260
rect 286870 333248 286876 333260
rect 286192 333220 286876 333248
rect 286192 333208 286198 333220
rect 286870 333208 286876 333220
rect 286928 333208 286934 333260
rect 287422 333208 287428 333260
rect 287480 333248 287486 333260
rect 288066 333248 288072 333260
rect 287480 333220 288072 333248
rect 287480 333208 287486 333220
rect 288066 333208 288072 333220
rect 288124 333208 288130 333260
rect 288986 333208 288992 333260
rect 289044 333248 289050 333260
rect 289630 333248 289636 333260
rect 289044 333220 289636 333248
rect 289044 333208 289050 333220
rect 289630 333208 289636 333220
rect 289688 333208 289694 333260
rect 291286 333208 291292 333260
rect 291344 333248 291350 333260
rect 292206 333248 292212 333260
rect 291344 333220 292212 333248
rect 291344 333208 291350 333220
rect 292206 333208 292212 333220
rect 292264 333208 292270 333260
rect 293126 333208 293132 333260
rect 293184 333248 293190 333260
rect 293678 333248 293684 333260
rect 293184 333220 293684 333248
rect 293184 333208 293190 333220
rect 293678 333208 293684 333220
rect 293736 333208 293742 333260
rect 295058 333208 295064 333260
rect 295116 333248 295122 333260
rect 500954 333248 500960 333260
rect 295116 333220 500960 333248
rect 295116 333208 295122 333220
rect 500954 333208 500960 333220
rect 501012 333208 501018 333260
rect 289446 333140 289452 333192
rect 289504 333180 289510 333192
rect 289722 333180 289728 333192
rect 289504 333152 289728 333180
rect 289504 333140 289510 333152
rect 289722 333140 289728 333152
rect 289780 333140 289786 333192
rect 295794 333140 295800 333192
rect 295852 333180 295858 333192
rect 296254 333180 296260 333192
rect 295852 333152 296260 333180
rect 295852 333140 295858 333152
rect 296254 333140 296260 333152
rect 296312 333140 296318 333192
rect 298646 333140 298652 333192
rect 298704 333180 298710 333192
rect 298922 333180 298928 333192
rect 298704 333152 298928 333180
rect 298704 333140 298710 333152
rect 298922 333140 298928 333152
rect 298980 333140 298986 333192
rect 299934 333140 299940 333192
rect 299992 333180 299998 333192
rect 300394 333180 300400 333192
rect 299992 333152 300400 333180
rect 299992 333140 299998 333152
rect 300394 333140 300400 333152
rect 300452 333140 300458 333192
rect 298370 333072 298376 333124
rect 298428 333112 298434 333124
rect 299014 333112 299020 333124
rect 298428 333084 299020 333112
rect 298428 333072 298434 333084
rect 299014 333072 299020 333084
rect 299072 333072 299078 333124
rect 300210 333072 300216 333124
rect 300268 333112 300274 333124
rect 300578 333112 300584 333124
rect 300268 333084 300584 333112
rect 300268 333072 300274 333084
rect 300578 333072 300584 333084
rect 300636 333072 300642 333124
rect 3050 332528 3056 332580
rect 3108 332568 3114 332580
rect 233142 332568 233148 332580
rect 3108 332540 233148 332568
rect 3108 332528 3114 332540
rect 233142 332528 233148 332540
rect 233200 332528 233206 332580
rect 234522 332188 234528 332240
rect 234580 332228 234586 332240
rect 262858 332228 262864 332240
rect 234580 332200 262864 332228
rect 234580 332188 234586 332200
rect 262858 332188 262864 332200
rect 262916 332188 262922 332240
rect 273346 332188 273352 332240
rect 273404 332228 273410 332240
rect 320174 332228 320180 332240
rect 273404 332200 320180 332228
rect 273404 332188 273410 332200
rect 320174 332188 320180 332200
rect 320232 332188 320238 332240
rect 223482 332120 223488 332172
rect 223540 332160 223546 332172
rect 261662 332160 261668 332172
rect 223540 332132 261668 332160
rect 223540 332120 223546 332132
rect 261662 332120 261668 332132
rect 261720 332120 261726 332172
rect 276566 332120 276572 332172
rect 276624 332120 276630 332172
rect 277949 332163 278007 332169
rect 277949 332129 277961 332163
rect 277995 332160 278007 332163
rect 342254 332160 342260 332172
rect 277995 332132 342260 332160
rect 277995 332129 278007 332132
rect 277949 332123 278007 332129
rect 342254 332120 342260 332132
rect 342312 332120 342318 332172
rect 162762 332052 162768 332104
rect 162820 332092 162826 332104
rect 254394 332092 254400 332104
rect 162820 332064 254400 332092
rect 162820 332052 162826 332064
rect 254394 332052 254400 332064
rect 254452 332052 254458 332104
rect 276584 332092 276612 332120
rect 347774 332092 347780 332104
rect 276584 332064 347780 332092
rect 347774 332052 347780 332064
rect 347832 332052 347838 332104
rect 136542 331984 136548 332036
rect 136600 332024 136606 332036
rect 251266 332024 251272 332036
rect 136600 331996 251272 332024
rect 136600 331984 136606 331996
rect 251266 331984 251272 331996
rect 251324 331984 251330 332036
rect 283374 331984 283380 332036
rect 283432 332024 283438 332036
rect 405734 332024 405740 332036
rect 283432 331996 405740 332024
rect 283432 331984 283438 331996
rect 405734 331984 405740 331996
rect 405792 331984 405798 332036
rect 108942 331916 108948 331968
rect 109000 331956 109006 331968
rect 247862 331956 247868 331968
rect 109000 331928 247868 331956
rect 109000 331916 109006 331928
rect 247862 331916 247868 331928
rect 247920 331916 247926 331968
rect 276566 331916 276572 331968
rect 276624 331956 276630 331968
rect 277118 331956 277124 331968
rect 276624 331928 277124 331956
rect 276624 331916 276630 331928
rect 277118 331916 277124 331928
rect 277176 331916 277182 331968
rect 290829 331959 290887 331965
rect 290829 331925 290841 331959
rect 290875 331956 290887 331959
rect 465166 331956 465172 331968
rect 290875 331928 465172 331956
rect 290875 331925 290887 331928
rect 290829 331919 290887 331925
rect 465166 331916 465172 331928
rect 465224 331916 465230 331968
rect 68922 331848 68928 331900
rect 68980 331888 68986 331900
rect 243078 331888 243084 331900
rect 68980 331860 243084 331888
rect 68980 331848 68986 331860
rect 243078 331848 243084 331860
rect 243136 331848 243142 331900
rect 296438 331848 296444 331900
rect 296496 331888 296502 331900
rect 507854 331888 507860 331900
rect 296496 331860 507860 331888
rect 296496 331848 296502 331860
rect 507854 331848 507860 331860
rect 507912 331848 507918 331900
rect 242986 331372 242992 331424
rect 243044 331412 243050 331424
rect 243354 331412 243360 331424
rect 243044 331384 243360 331412
rect 243044 331372 243050 331384
rect 243354 331372 243360 331384
rect 243412 331372 243418 331424
rect 239030 331168 239036 331220
rect 239088 331168 239094 331220
rect 239048 331140 239076 331168
rect 239214 331140 239220 331152
rect 239048 331112 239220 331140
rect 239214 331100 239220 331112
rect 239272 331100 239278 331152
rect 240686 331100 240692 331152
rect 240744 331140 240750 331152
rect 240962 331140 240968 331152
rect 240744 331112 240968 331140
rect 240744 331100 240750 331112
rect 240962 331100 240968 331112
rect 241020 331100 241026 331152
rect 301314 331100 301320 331152
rect 301372 331140 301378 331152
rect 301590 331140 301596 331152
rect 301372 331112 301596 331140
rect 301372 331100 301378 331112
rect 301590 331100 301596 331112
rect 301648 331100 301654 331152
rect 249705 331007 249763 331013
rect 249705 330973 249717 331007
rect 249751 331004 249763 331007
rect 257430 331004 257436 331016
rect 249751 330976 257436 331004
rect 249751 330973 249763 330976
rect 249705 330967 249763 330973
rect 257430 330964 257436 330976
rect 257488 330964 257494 331016
rect 244734 330896 244740 330948
rect 244792 330936 244798 330948
rect 244918 330936 244924 330948
rect 244792 330908 244924 330936
rect 244792 330896 244798 330908
rect 244918 330896 244924 330908
rect 244976 330896 244982 330948
rect 245010 330896 245016 330948
rect 245068 330936 245074 330948
rect 245194 330936 245200 330948
rect 245068 330908 245200 330936
rect 245068 330896 245074 330908
rect 245194 330896 245200 330908
rect 245252 330896 245258 330948
rect 249797 330939 249855 330945
rect 249797 330905 249809 330939
rect 249843 330936 249855 330939
rect 256418 330936 256424 330948
rect 249843 330908 256424 330936
rect 249843 330905 249855 330908
rect 249797 330899 249855 330905
rect 256418 330896 256424 330908
rect 256476 330896 256482 330948
rect 298833 330939 298891 330945
rect 298833 330905 298845 330939
rect 298879 330936 298891 330939
rect 299106 330936 299112 330948
rect 298879 330908 299112 330936
rect 298879 330905 298891 330908
rect 298833 330899 298891 330905
rect 299106 330896 299112 330908
rect 299164 330896 299170 330948
rect 213822 330828 213828 330880
rect 213880 330868 213886 330880
rect 260466 330868 260472 330880
rect 213880 330840 260472 330868
rect 213880 330828 213886 330840
rect 260466 330828 260472 330840
rect 260524 330828 260530 330880
rect 274266 330828 274272 330880
rect 274324 330868 274330 330880
rect 327074 330868 327080 330880
rect 274324 330840 327080 330868
rect 274324 330828 274330 330840
rect 327074 330828 327080 330840
rect 327132 330828 327138 330880
rect 187602 330760 187608 330812
rect 187660 330800 187666 330812
rect 249705 330803 249763 330809
rect 249705 330800 249717 330803
rect 187660 330772 249717 330800
rect 187660 330760 187666 330772
rect 249705 330769 249717 330772
rect 249751 330769 249763 330803
rect 252554 330800 252560 330812
rect 249705 330763 249763 330769
rect 249904 330772 252560 330800
rect 179322 330692 179328 330744
rect 179380 330732 179386 330744
rect 249797 330735 249855 330741
rect 249797 330732 249809 330735
rect 179380 330704 249809 330732
rect 179380 330692 179386 330704
rect 249797 330701 249809 330704
rect 249843 330701 249855 330735
rect 249797 330695 249855 330701
rect 147582 330624 147588 330676
rect 147640 330664 147646 330676
rect 249904 330664 249932 330772
rect 252554 330760 252560 330772
rect 252612 330760 252618 330812
rect 274818 330760 274824 330812
rect 274876 330800 274882 330812
rect 332594 330800 332600 330812
rect 274876 330772 332600 330800
rect 274876 330760 274882 330772
rect 332594 330760 332600 330772
rect 332652 330760 332658 330812
rect 250530 330732 250536 330744
rect 147640 330636 249932 330664
rect 249996 330704 250536 330732
rect 147640 330624 147646 330636
rect 102042 330556 102048 330608
rect 102100 330596 102106 330608
rect 246942 330596 246948 330608
rect 102100 330568 246948 330596
rect 102100 330556 102106 330568
rect 246942 330556 246948 330568
rect 247000 330556 247006 330608
rect 247678 330556 247684 330608
rect 247736 330596 247742 330608
rect 247862 330596 247868 330608
rect 247736 330568 247868 330596
rect 247736 330556 247742 330568
rect 247862 330556 247868 330568
rect 247920 330556 247926 330608
rect 35802 330488 35808 330540
rect 35860 330528 35866 330540
rect 35860 330500 219434 330528
rect 35860 330488 35866 330500
rect 219406 330256 219434 330500
rect 245010 330488 245016 330540
rect 245068 330528 245074 330540
rect 245562 330528 245568 330540
rect 245068 330500 245568 330528
rect 245068 330488 245074 330500
rect 245562 330488 245568 330500
rect 245620 330488 245626 330540
rect 246206 330488 246212 330540
rect 246264 330528 246270 330540
rect 246850 330528 246856 330540
rect 246264 330500 246856 330528
rect 246264 330488 246270 330500
rect 246850 330488 246856 330500
rect 246908 330488 246914 330540
rect 247310 330488 247316 330540
rect 247368 330528 247374 330540
rect 247954 330528 247960 330540
rect 247368 330500 247960 330528
rect 247368 330488 247374 330500
rect 247954 330488 247960 330500
rect 248012 330488 248018 330540
rect 249996 330472 250024 330704
rect 250530 330692 250536 330704
rect 250588 330692 250594 330744
rect 277762 330692 277768 330744
rect 277820 330732 277826 330744
rect 357434 330732 357440 330744
rect 277820 330704 357440 330732
rect 277820 330692 277826 330704
rect 357434 330692 357440 330704
rect 357492 330692 357498 330744
rect 250622 330664 250628 330676
rect 250088 330636 250628 330664
rect 250088 330472 250116 330636
rect 250622 330624 250628 330636
rect 250680 330624 250686 330676
rect 263778 330624 263784 330676
rect 263836 330664 263842 330676
rect 264422 330664 264428 330676
rect 263836 330636 264428 330664
rect 263836 330624 263842 330636
rect 264422 330624 264428 330636
rect 264480 330624 264486 330676
rect 270310 330624 270316 330676
rect 270368 330624 270374 330676
rect 271322 330624 271328 330676
rect 271380 330664 271386 330676
rect 271598 330664 271604 330676
rect 271380 330636 271604 330664
rect 271380 330624 271386 330636
rect 271598 330624 271604 330636
rect 271656 330624 271662 330676
rect 285766 330624 285772 330676
rect 285824 330664 285830 330676
rect 423674 330664 423680 330676
rect 285824 330636 423680 330664
rect 285824 330624 285830 330636
rect 423674 330624 423680 330636
rect 423732 330624 423738 330676
rect 265158 330556 265164 330608
rect 265216 330596 265222 330608
rect 265802 330596 265808 330608
rect 265216 330568 265808 330596
rect 265216 330556 265222 330568
rect 265802 330556 265808 330568
rect 265860 330556 265866 330608
rect 250254 330488 250260 330540
rect 250312 330528 250318 330540
rect 251082 330528 251088 330540
rect 250312 330500 251088 330528
rect 250312 330488 250318 330500
rect 251082 330488 251088 330500
rect 251140 330488 251146 330540
rect 252830 330488 252836 330540
rect 252888 330528 252894 330540
rect 253382 330528 253388 330540
rect 252888 330500 253388 330528
rect 252888 330488 252894 330500
rect 253382 330488 253388 330500
rect 253440 330488 253446 330540
rect 265526 330488 265532 330540
rect 265584 330528 265590 330540
rect 266262 330528 266268 330540
rect 265584 330500 266268 330528
rect 265584 330488 265590 330500
rect 266262 330488 266268 330500
rect 266320 330488 266326 330540
rect 244550 330420 244556 330472
rect 244608 330460 244614 330472
rect 245102 330460 245108 330472
rect 244608 330432 245108 330460
rect 244608 330420 244614 330432
rect 245102 330420 245108 330432
rect 245160 330420 245166 330472
rect 247218 330420 247224 330472
rect 247276 330460 247282 330472
rect 248138 330460 248144 330472
rect 247276 330432 248144 330460
rect 247276 330420 247282 330432
rect 248138 330420 248144 330432
rect 248196 330420 248202 330472
rect 249978 330420 249984 330472
rect 250036 330420 250042 330472
rect 250070 330420 250076 330472
rect 250128 330420 250134 330472
rect 251726 330420 251732 330472
rect 251784 330460 251790 330472
rect 252370 330460 252376 330472
rect 251784 330432 252376 330460
rect 251784 330420 251790 330432
rect 252370 330420 252376 330432
rect 252428 330420 252434 330472
rect 253106 330420 253112 330472
rect 253164 330460 253170 330472
rect 253290 330460 253296 330472
rect 253164 330432 253296 330460
rect 253164 330420 253170 330432
rect 253290 330420 253296 330432
rect 253348 330420 253354 330472
rect 265342 330420 265348 330472
rect 265400 330460 265406 330472
rect 265986 330460 265992 330472
rect 265400 330432 265992 330460
rect 265400 330420 265406 330432
rect 265986 330420 265992 330432
rect 266044 330420 266050 330472
rect 270328 330460 270356 330624
rect 305086 330556 305092 330608
rect 305144 330596 305150 330608
rect 514754 330596 514760 330608
rect 305144 330568 514760 330596
rect 305144 330556 305150 330568
rect 514754 330556 514760 330568
rect 514812 330556 514818 330608
rect 272886 330488 272892 330540
rect 272944 330528 272950 330540
rect 273162 330528 273168 330540
rect 272944 330500 273168 330528
rect 272944 330488 272950 330500
rect 273162 330488 273168 330500
rect 273220 330488 273226 330540
rect 282086 330488 282092 330540
rect 282144 330528 282150 330540
rect 282270 330528 282276 330540
rect 282144 330500 282276 330528
rect 282144 330488 282150 330500
rect 282270 330488 282276 330500
rect 282328 330488 282334 330540
rect 302510 330488 302516 330540
rect 302568 330528 302574 330540
rect 564434 330528 564440 330540
rect 302568 330500 564440 330528
rect 302568 330488 302574 330500
rect 564434 330488 564440 330500
rect 564492 330488 564498 330540
rect 270402 330460 270408 330472
rect 270328 330432 270408 330460
rect 270402 330420 270408 330432
rect 270460 330420 270466 330472
rect 270678 330420 270684 330472
rect 270736 330460 270742 330472
rect 271414 330460 271420 330472
rect 270736 330432 271420 330460
rect 270736 330420 270742 330432
rect 271414 330420 271420 330432
rect 271472 330420 271478 330472
rect 295702 330420 295708 330472
rect 295760 330460 295766 330472
rect 296622 330460 296628 330472
rect 295760 330432 296628 330460
rect 295760 330420 295766 330432
rect 296622 330420 296628 330432
rect 296680 330420 296686 330472
rect 298830 330460 298836 330472
rect 298791 330432 298836 330460
rect 298830 330420 298836 330432
rect 298888 330420 298894 330472
rect 301038 330420 301044 330472
rect 301096 330460 301102 330472
rect 301958 330460 301964 330472
rect 301096 330432 301964 330460
rect 301096 330420 301102 330432
rect 301958 330420 301964 330432
rect 302016 330420 302022 330472
rect 302878 330420 302884 330472
rect 302936 330460 302942 330472
rect 303154 330460 303160 330472
rect 302936 330432 303160 330460
rect 302936 330420 302942 330432
rect 303154 330420 303160 330432
rect 303212 330420 303218 330472
rect 303798 330420 303804 330472
rect 303856 330460 303862 330472
rect 304442 330460 304448 330472
rect 303856 330432 304448 330460
rect 303856 330420 303862 330432
rect 304442 330420 304448 330432
rect 304500 330420 304506 330472
rect 244826 330352 244832 330404
rect 244884 330392 244890 330404
rect 245286 330392 245292 330404
rect 244884 330364 245292 330392
rect 244884 330352 244890 330364
rect 245286 330352 245292 330364
rect 245344 330352 245350 330404
rect 245838 330352 245844 330404
rect 245896 330392 245902 330404
rect 246022 330392 246028 330404
rect 245896 330364 246028 330392
rect 245896 330352 245902 330364
rect 246022 330352 246028 330364
rect 246080 330352 246086 330404
rect 247494 330352 247500 330404
rect 247552 330392 247558 330404
rect 248230 330392 248236 330404
rect 247552 330364 248236 330392
rect 247552 330352 247558 330364
rect 248230 330352 248236 330364
rect 248288 330352 248294 330404
rect 263686 330352 263692 330404
rect 263744 330392 263750 330404
rect 264054 330392 264060 330404
rect 263744 330364 264060 330392
rect 263744 330352 263750 330364
rect 264054 330352 264060 330364
rect 264112 330352 264118 330404
rect 269298 330352 269304 330404
rect 269356 330392 269362 330404
rect 270310 330392 270316 330404
rect 269356 330364 270316 330392
rect 269356 330352 269362 330364
rect 270310 330352 270316 330364
rect 270368 330352 270374 330404
rect 274174 330352 274180 330404
rect 274232 330392 274238 330404
rect 274450 330392 274456 330404
rect 274232 330364 274456 330392
rect 274232 330352 274238 330364
rect 274450 330352 274456 330364
rect 274508 330352 274514 330404
rect 278406 330352 278412 330404
rect 278464 330392 278470 330404
rect 278590 330392 278596 330404
rect 278464 330364 278596 330392
rect 278464 330352 278470 330364
rect 278590 330352 278596 330364
rect 278648 330352 278654 330404
rect 279050 330352 279056 330404
rect 279108 330392 279114 330404
rect 279786 330392 279792 330404
rect 279108 330364 279792 330392
rect 279108 330352 279114 330364
rect 279786 330352 279792 330364
rect 279844 330352 279850 330404
rect 280798 330392 280804 330404
rect 280759 330364 280804 330392
rect 280798 330352 280804 330364
rect 280856 330352 280862 330404
rect 281902 330352 281908 330404
rect 281960 330392 281966 330404
rect 282730 330392 282736 330404
rect 281960 330364 282736 330392
rect 281960 330352 281966 330364
rect 282730 330352 282736 330364
rect 282788 330352 282794 330404
rect 299842 330352 299848 330404
rect 299900 330392 299906 330404
rect 300670 330392 300676 330404
rect 299900 330364 300676 330392
rect 299900 330352 299906 330364
rect 300670 330352 300676 330364
rect 300728 330352 300734 330404
rect 252738 330284 252744 330336
rect 252796 330324 252802 330336
rect 253290 330324 253296 330336
rect 252796 330296 253296 330324
rect 252796 330284 252802 330296
rect 253290 330284 253296 330296
rect 253348 330284 253354 330336
rect 280246 330284 280252 330336
rect 280304 330324 280310 330336
rect 281166 330324 281172 330336
rect 280304 330296 281172 330324
rect 280304 330284 280310 330296
rect 281166 330284 281172 330296
rect 281224 330284 281230 330336
rect 239033 330259 239091 330265
rect 239033 330256 239045 330259
rect 219406 330228 239045 330256
rect 239033 330225 239045 330228
rect 239079 330225 239091 330259
rect 239033 330219 239091 330225
rect 246022 330216 246028 330268
rect 246080 330256 246086 330268
rect 246666 330256 246672 330268
rect 246080 330228 246672 330256
rect 246080 330216 246086 330228
rect 246666 330216 246672 330228
rect 246724 330216 246730 330268
rect 248598 330216 248604 330268
rect 248656 330256 248662 330268
rect 249150 330256 249156 330268
rect 248656 330228 249156 330256
rect 248656 330216 248662 330228
rect 249150 330216 249156 330228
rect 249208 330216 249214 330268
rect 300302 330216 300308 330268
rect 300360 330256 300366 330268
rect 300673 330259 300731 330265
rect 300673 330256 300685 330259
rect 300360 330228 300685 330256
rect 300360 330216 300366 330228
rect 300673 330225 300685 330228
rect 300719 330225 300731 330259
rect 300673 330219 300731 330225
rect 280430 330148 280436 330200
rect 280488 330188 280494 330200
rect 281442 330188 281448 330200
rect 280488 330160 281448 330188
rect 280488 330148 280494 330160
rect 281442 330148 281448 330160
rect 281500 330148 281506 330200
rect 248874 329468 248880 329520
rect 248932 329508 248938 329520
rect 249242 329508 249248 329520
rect 248932 329480 249248 329508
rect 248932 329468 248938 329480
rect 249242 329468 249248 329480
rect 249300 329468 249306 329520
rect 227622 329400 227628 329452
rect 227680 329440 227686 329452
rect 262030 329440 262036 329452
rect 227680 329412 262036 329440
rect 227680 329400 227686 329412
rect 262030 329400 262036 329412
rect 262088 329400 262094 329452
rect 288618 329400 288624 329452
rect 288676 329440 288682 329452
rect 289538 329440 289544 329452
rect 288676 329412 289544 329440
rect 288676 329400 288682 329412
rect 289538 329400 289544 329412
rect 289596 329400 289602 329452
rect 188982 329332 188988 329384
rect 189040 329372 189046 329384
rect 257522 329372 257528 329384
rect 189040 329344 257528 329372
rect 189040 329332 189046 329344
rect 257522 329332 257528 329344
rect 257580 329332 257586 329384
rect 275646 329332 275652 329384
rect 275704 329372 275710 329384
rect 339494 329372 339500 329384
rect 275704 329344 339500 329372
rect 275704 329332 275710 329344
rect 339494 329332 339500 329344
rect 339552 329332 339558 329384
rect 166902 329264 166908 329316
rect 166960 329304 166966 329316
rect 254854 329304 254860 329316
rect 166960 329276 254860 329304
rect 166960 329264 166966 329276
rect 254854 329264 254860 329276
rect 254912 329264 254918 329316
rect 283926 329264 283932 329316
rect 283984 329304 283990 329316
rect 365714 329304 365720 329316
rect 283984 329276 365720 329304
rect 283984 329264 283990 329276
rect 365714 329264 365720 329276
rect 365772 329264 365778 329316
rect 140682 329196 140688 329248
rect 140740 329236 140746 329248
rect 251818 329236 251824 329248
rect 140740 329208 251824 329236
rect 140740 329196 140746 329208
rect 251818 329196 251824 329208
rect 251876 329196 251882 329248
rect 285306 329196 285312 329248
rect 285364 329236 285370 329248
rect 419534 329236 419540 329248
rect 285364 329208 419540 329236
rect 285364 329196 285370 329208
rect 419534 329196 419540 329208
rect 419592 329196 419598 329248
rect 115842 329128 115848 329180
rect 115900 329168 115906 329180
rect 248782 329168 248788 329180
rect 115900 329140 248788 329168
rect 115900 329128 115906 329140
rect 248782 329128 248788 329140
rect 248840 329128 248846 329180
rect 271782 329128 271788 329180
rect 271840 329168 271846 329180
rect 304994 329168 305000 329180
rect 271840 329140 305000 329168
rect 271840 329128 271846 329140
rect 304994 329128 305000 329140
rect 305052 329128 305058 329180
rect 305178 329128 305184 329180
rect 305236 329168 305242 329180
rect 518894 329168 518900 329180
rect 305236 329140 518900 329168
rect 305236 329128 305242 329140
rect 518894 329128 518900 329140
rect 518952 329128 518958 329180
rect 43438 329060 43444 329112
rect 43496 329100 43502 329112
rect 239858 329100 239864 329112
rect 43496 329072 239864 329100
rect 43496 329060 43502 329072
rect 239858 329060 239864 329072
rect 239916 329060 239922 329112
rect 298554 329060 298560 329112
rect 298612 329100 298618 329112
rect 529198 329100 529204 329112
rect 298612 329072 529204 329100
rect 298612 329060 298618 329072
rect 529198 329060 529204 329072
rect 529256 329060 529262 329112
rect 254578 329032 254584 329044
rect 254539 329004 254584 329032
rect 254578 328992 254584 329004
rect 254636 328992 254642 329044
rect 252830 328380 252836 328432
rect 252888 328420 252894 328432
rect 253474 328420 253480 328432
rect 252888 328392 253480 328420
rect 252888 328380 252894 328392
rect 253474 328380 253480 328392
rect 253532 328380 253538 328432
rect 253014 328312 253020 328364
rect 253072 328352 253078 328364
rect 253658 328352 253664 328364
rect 253072 328324 253664 328352
rect 253072 328312 253078 328324
rect 253658 328312 253664 328324
rect 253716 328312 253722 328364
rect 231762 328040 231768 328092
rect 231820 328080 231826 328092
rect 262674 328080 262680 328092
rect 231820 328052 262680 328080
rect 231820 328040 231826 328052
rect 262674 328040 262680 328052
rect 262732 328040 262738 328092
rect 184842 327972 184848 328024
rect 184900 328012 184906 328024
rect 256970 328012 256976 328024
rect 184900 327984 256976 328012
rect 184900 327972 184906 327984
rect 256970 327972 256976 327984
rect 257028 327972 257034 328024
rect 294138 327972 294144 328024
rect 294196 328012 294202 328024
rect 331214 328012 331220 328024
rect 294196 327984 331220 328012
rect 294196 327972 294202 327984
rect 331214 327972 331220 327984
rect 331272 327972 331278 328024
rect 160002 327904 160008 327956
rect 160060 327944 160066 327956
rect 254486 327944 254492 327956
rect 160060 327916 254492 327944
rect 160060 327904 160066 327916
rect 254486 327904 254492 327916
rect 254544 327904 254550 327956
rect 277210 327904 277216 327956
rect 277268 327944 277274 327956
rect 353294 327944 353300 327956
rect 277268 327916 353300 327944
rect 277268 327904 277274 327916
rect 353294 327904 353300 327916
rect 353352 327904 353358 327956
rect 151722 327836 151728 327888
rect 151780 327876 151786 327888
rect 252738 327876 252744 327888
rect 151780 327848 252744 327876
rect 151780 327836 151786 327848
rect 252738 327836 252744 327848
rect 252796 327836 252802 327888
rect 284570 327836 284576 327888
rect 284628 327876 284634 327888
rect 415486 327876 415492 327888
rect 284628 327848 415492 327876
rect 284628 327836 284634 327848
rect 415486 327836 415492 327848
rect 415544 327836 415550 327888
rect 85482 327768 85488 327820
rect 85540 327808 85546 327820
rect 245194 327808 245200 327820
rect 85540 327780 245200 327808
rect 85540 327768 85546 327780
rect 245194 327768 245200 327780
rect 245252 327768 245258 327820
rect 293586 327768 293592 327820
rect 293644 327808 293650 327820
rect 293644 327780 293724 327808
rect 293644 327768 293650 327780
rect 46198 327700 46204 327752
rect 46256 327740 46262 327752
rect 240318 327740 240324 327752
rect 46256 327712 240324 327740
rect 46256 327700 46262 327712
rect 240318 327700 240324 327712
rect 240376 327700 240382 327752
rect 293696 327616 293724 327780
rect 293770 327768 293776 327820
rect 293828 327808 293834 327820
rect 484394 327808 484400 327820
rect 293828 327780 484400 327808
rect 293828 327768 293834 327780
rect 484394 327768 484400 327780
rect 484452 327768 484458 327820
rect 303522 327700 303528 327752
rect 303580 327740 303586 327752
rect 566458 327740 566464 327752
rect 303580 327712 566464 327740
rect 303580 327700 303586 327712
rect 566458 327700 566464 327712
rect 566516 327700 566522 327752
rect 293678 327564 293684 327616
rect 293736 327564 293742 327616
rect 248782 327156 248788 327208
rect 248840 327196 248846 327208
rect 249702 327196 249708 327208
rect 248840 327168 249708 327196
rect 248840 327156 248846 327168
rect 249702 327156 249708 327168
rect 249760 327156 249766 327208
rect 302878 327088 302884 327140
rect 302936 327128 302942 327140
rect 303430 327128 303436 327140
rect 302936 327100 303436 327128
rect 302936 327088 302942 327100
rect 303430 327088 303436 327100
rect 303488 327088 303494 327140
rect 237558 326680 237564 326732
rect 237616 326720 237622 326732
rect 237742 326720 237748 326732
rect 237616 326692 237748 326720
rect 237616 326680 237622 326692
rect 237742 326680 237748 326692
rect 237800 326680 237806 326732
rect 217962 326612 217968 326664
rect 218020 326652 218026 326664
rect 261110 326652 261116 326664
rect 218020 326624 261116 326652
rect 218020 326612 218026 326624
rect 261110 326612 261116 326624
rect 261168 326612 261174 326664
rect 277302 326612 277308 326664
rect 277360 326652 277366 326664
rect 346394 326652 346400 326664
rect 277360 326624 346400 326652
rect 277360 326612 277366 326624
rect 346394 326612 346400 326624
rect 346452 326612 346458 326664
rect 191742 326544 191748 326596
rect 191800 326584 191806 326596
rect 257798 326584 257804 326596
rect 191800 326556 257804 326584
rect 191800 326544 191806 326556
rect 257798 326544 257804 326556
rect 257856 326544 257862 326596
rect 258442 326584 258448 326596
rect 258184 326556 258448 326584
rect 154482 326476 154488 326528
rect 154540 326516 154546 326528
rect 252646 326516 252652 326528
rect 154540 326488 252652 326516
rect 154540 326476 154546 326488
rect 252646 326476 252652 326488
rect 252704 326476 252710 326528
rect 113082 326408 113088 326460
rect 113140 326448 113146 326460
rect 248506 326448 248512 326460
rect 113140 326420 248512 326448
rect 113140 326408 113146 326420
rect 248506 326408 248512 326420
rect 248564 326408 248570 326460
rect 104802 326340 104808 326392
rect 104860 326380 104866 326392
rect 247126 326380 247132 326392
rect 104860 326352 247132 326380
rect 104860 326340 104866 326352
rect 247126 326340 247132 326352
rect 247184 326340 247190 326392
rect 254394 326340 254400 326392
rect 254452 326380 254458 326392
rect 254946 326380 254952 326392
rect 254452 326352 254952 326380
rect 254452 326340 254458 326352
rect 254946 326340 254952 326352
rect 255004 326340 255010 326392
rect 255406 326340 255412 326392
rect 255464 326380 255470 326392
rect 255774 326380 255780 326392
rect 255464 326352 255780 326380
rect 255464 326340 255470 326352
rect 255774 326340 255780 326352
rect 255832 326340 255838 326392
rect 257062 326340 257068 326392
rect 257120 326380 257126 326392
rect 257890 326380 257896 326392
rect 257120 326352 257896 326380
rect 257120 326340 257126 326352
rect 257890 326340 257896 326352
rect 257948 326340 257954 326392
rect 235166 326272 235172 326324
rect 235224 326312 235230 326324
rect 235902 326312 235908 326324
rect 235224 326284 235908 326312
rect 235224 326272 235230 326284
rect 235902 326272 235908 326284
rect 235960 326272 235966 326324
rect 236362 326272 236368 326324
rect 236420 326312 236426 326324
rect 237098 326312 237104 326324
rect 236420 326284 237104 326312
rect 236420 326272 236426 326284
rect 237098 326272 237104 326284
rect 237156 326272 237162 326324
rect 237834 326272 237840 326324
rect 237892 326312 237898 326324
rect 238478 326312 238484 326324
rect 237892 326284 238484 326312
rect 237892 326272 237898 326284
rect 238478 326272 238484 326284
rect 238536 326272 238542 326324
rect 243538 326272 243544 326324
rect 243596 326312 243602 326324
rect 244182 326312 244188 326324
rect 243596 326284 244188 326312
rect 243596 326272 243602 326284
rect 244182 326272 244188 326284
rect 244240 326272 244246 326324
rect 258184 326256 258212 326556
rect 258442 326544 258448 326556
rect 258500 326544 258506 326596
rect 279234 326544 279240 326596
rect 279292 326584 279298 326596
rect 375374 326584 375380 326596
rect 279292 326556 375380 326584
rect 279292 326544 279298 326556
rect 375374 326544 375380 326556
rect 375432 326544 375438 326596
rect 285030 326476 285036 326528
rect 285088 326516 285094 326528
rect 285214 326516 285220 326528
rect 285088 326488 285220 326516
rect 285088 326476 285094 326488
rect 285214 326476 285220 326488
rect 285272 326476 285278 326528
rect 292114 326516 292120 326528
rect 292075 326488 292120 326516
rect 292114 326476 292120 326488
rect 292172 326476 292178 326528
rect 294414 326476 294420 326528
rect 294472 326516 294478 326528
rect 412634 326516 412640 326528
rect 294472 326488 412640 326516
rect 294472 326476 294478 326488
rect 412634 326476 412640 326488
rect 412692 326476 412698 326528
rect 258902 326448 258908 326460
rect 258368 326420 258908 326448
rect 258368 326392 258396 326420
rect 258902 326408 258908 326420
rect 258960 326408 258966 326460
rect 259638 326408 259644 326460
rect 259696 326448 259702 326460
rect 260098 326448 260104 326460
rect 259696 326420 260104 326448
rect 259696 326408 259702 326420
rect 260098 326408 260104 326420
rect 260156 326408 260162 326460
rect 288342 326408 288348 326460
rect 288400 326448 288406 326460
rect 441614 326448 441620 326460
rect 288400 326420 441620 326448
rect 288400 326408 288406 326420
rect 441614 326408 441620 326420
rect 441672 326408 441678 326460
rect 258350 326340 258356 326392
rect 258408 326340 258414 326392
rect 258442 326340 258448 326392
rect 258500 326380 258506 326392
rect 258994 326380 259000 326392
rect 258500 326352 259000 326380
rect 258500 326340 258506 326352
rect 258994 326340 259000 326352
rect 259052 326340 259058 326392
rect 259546 326340 259552 326392
rect 259604 326380 259610 326392
rect 260006 326380 260012 326392
rect 259604 326352 260012 326380
rect 259604 326340 259610 326352
rect 260006 326340 260012 326352
rect 260064 326340 260070 326392
rect 262582 326340 262588 326392
rect 262640 326380 262646 326392
rect 263134 326380 263140 326392
rect 262640 326352 263140 326380
rect 262640 326340 262646 326352
rect 263134 326340 263140 326352
rect 263192 326340 263198 326392
rect 283558 326340 283564 326392
rect 283616 326380 283622 326392
rect 283742 326380 283748 326392
rect 283616 326352 283748 326380
rect 283616 326340 283622 326352
rect 283742 326340 283748 326352
rect 283800 326340 283806 326392
rect 283926 326340 283932 326392
rect 283984 326380 283990 326392
rect 284110 326380 284116 326392
rect 283984 326352 284116 326380
rect 283984 326340 283990 326352
rect 284110 326340 284116 326352
rect 284168 326340 284174 326392
rect 286318 326340 286324 326392
rect 286376 326380 286382 326392
rect 286686 326380 286692 326392
rect 286376 326352 286692 326380
rect 286376 326340 286382 326352
rect 286686 326340 286692 326352
rect 286744 326340 286750 326392
rect 287054 326340 287060 326392
rect 287112 326380 287118 326392
rect 287698 326380 287704 326392
rect 287112 326352 287704 326380
rect 287112 326340 287118 326352
rect 287698 326340 287704 326352
rect 287756 326340 287762 326392
rect 291010 326340 291016 326392
rect 291068 326380 291074 326392
rect 291068 326352 291148 326380
rect 291068 326340 291074 326352
rect 258810 326272 258816 326324
rect 258868 326312 258874 326324
rect 258868 326284 258948 326312
rect 258868 326272 258874 326284
rect 234706 326204 234712 326256
rect 234764 326244 234770 326256
rect 235810 326244 235816 326256
rect 234764 326216 235816 326244
rect 234764 326204 234770 326216
rect 235810 326204 235816 326216
rect 235868 326204 235874 326256
rect 237650 326204 237656 326256
rect 237708 326244 237714 326256
rect 238110 326244 238116 326256
rect 237708 326216 238116 326244
rect 237708 326204 237714 326216
rect 238110 326204 238116 326216
rect 238168 326204 238174 326256
rect 239122 326204 239128 326256
rect 239180 326244 239186 326256
rect 239766 326244 239772 326256
rect 239180 326216 239772 326244
rect 239180 326204 239186 326216
rect 239766 326204 239772 326216
rect 239824 326204 239830 326256
rect 240410 326204 240416 326256
rect 240468 326244 240474 326256
rect 241422 326244 241428 326256
rect 240468 326216 241428 326244
rect 240468 326204 240474 326216
rect 241422 326204 241428 326216
rect 241480 326204 241486 326256
rect 241790 326204 241796 326256
rect 241848 326244 241854 326256
rect 242434 326244 242440 326256
rect 241848 326216 242440 326244
rect 241848 326204 241854 326216
rect 242434 326204 242440 326216
rect 242492 326204 242498 326256
rect 243262 326204 243268 326256
rect 243320 326244 243326 326256
rect 243722 326244 243728 326256
rect 243320 326216 243728 326244
rect 243320 326204 243326 326216
rect 243722 326204 243728 326216
rect 243780 326204 243786 326256
rect 255406 326204 255412 326256
rect 255464 326244 255470 326256
rect 256050 326244 256056 326256
rect 255464 326216 256056 326244
rect 255464 326204 255470 326216
rect 256050 326204 256056 326216
rect 256108 326204 256114 326256
rect 258166 326204 258172 326256
rect 258224 326204 258230 326256
rect 237926 326136 237932 326188
rect 237984 326176 237990 326188
rect 238662 326176 238668 326188
rect 237984 326148 238668 326176
rect 237984 326136 237990 326148
rect 238662 326136 238668 326148
rect 238720 326136 238726 326188
rect 239030 326136 239036 326188
rect 239088 326176 239094 326188
rect 240042 326176 240048 326188
rect 239088 326148 240048 326176
rect 239088 326136 239094 326148
rect 240042 326136 240048 326148
rect 240100 326136 240106 326188
rect 240134 326136 240140 326188
rect 240192 326176 240198 326188
rect 241330 326176 241336 326188
rect 240192 326148 241336 326176
rect 240192 326136 240198 326148
rect 241330 326136 241336 326148
rect 241388 326136 241394 326188
rect 255682 326136 255688 326188
rect 255740 326176 255746 326188
rect 256602 326176 256608 326188
rect 255740 326148 256608 326176
rect 255740 326136 255746 326148
rect 256602 326136 256608 326148
rect 256660 326136 256666 326188
rect 258920 326120 258948 326284
rect 259822 326272 259828 326324
rect 259880 326312 259886 326324
rect 260742 326312 260748 326324
rect 259880 326284 260748 326312
rect 259880 326272 259886 326284
rect 260742 326272 260748 326284
rect 260800 326272 260806 326324
rect 259730 326204 259736 326256
rect 259788 326244 259794 326256
rect 260282 326244 260288 326256
rect 259788 326216 260288 326244
rect 259788 326204 259794 326216
rect 260282 326204 260288 326216
rect 260340 326204 260346 326256
rect 284662 326204 284668 326256
rect 284720 326244 284726 326256
rect 284938 326244 284944 326256
rect 284720 326216 284944 326244
rect 284720 326204 284726 326216
rect 284938 326204 284944 326216
rect 284996 326204 285002 326256
rect 259546 326136 259552 326188
rect 259604 326176 259610 326188
rect 260558 326176 260564 326188
rect 259604 326148 260564 326176
rect 259604 326136 259610 326148
rect 260558 326136 260564 326148
rect 260616 326136 260622 326188
rect 291120 326120 291148 326352
rect 292666 326340 292672 326392
rect 292724 326380 292730 326392
rect 481634 326380 481640 326392
rect 292724 326352 481640 326380
rect 292724 326340 292730 326352
rect 481634 326340 481640 326352
rect 481692 326340 481698 326392
rect 292117 326247 292175 326253
rect 292117 326213 292129 326247
rect 292163 326244 292175 326247
rect 292206 326244 292212 326256
rect 292163 326216 292212 326244
rect 292163 326213 292175 326216
rect 292117 326207 292175 326213
rect 292206 326204 292212 326216
rect 292264 326204 292270 326256
rect 237466 326068 237472 326120
rect 237524 326108 237530 326120
rect 238202 326108 238208 326120
rect 237524 326080 238208 326108
rect 237524 326068 237530 326080
rect 238202 326068 238208 326080
rect 238260 326068 238266 326120
rect 255498 326068 255504 326120
rect 255556 326108 255562 326120
rect 256510 326108 256516 326120
rect 255556 326080 256516 326108
rect 255556 326068 255562 326080
rect 256510 326068 256516 326080
rect 256568 326068 256574 326120
rect 258902 326068 258908 326120
rect 258960 326068 258966 326120
rect 285950 326068 285956 326120
rect 286008 326108 286014 326120
rect 286318 326108 286324 326120
rect 286008 326080 286324 326108
rect 286008 326068 286014 326080
rect 286318 326068 286324 326080
rect 286376 326068 286382 326120
rect 291102 326068 291108 326120
rect 291160 326068 291166 326120
rect 285858 326000 285864 326052
rect 285916 326040 285922 326052
rect 286594 326040 286600 326052
rect 285916 326012 286600 326040
rect 285916 326000 285922 326012
rect 286594 326000 286600 326012
rect 286652 326000 286658 326052
rect 242066 325864 242072 325916
rect 242124 325904 242130 325916
rect 242618 325904 242624 325916
rect 242124 325876 242624 325904
rect 242124 325864 242130 325876
rect 242618 325864 242624 325876
rect 242676 325864 242682 325916
rect 306374 325592 306380 325644
rect 306432 325632 306438 325644
rect 580166 325632 580172 325644
rect 306432 325604 580172 325632
rect 306432 325592 306438 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 289170 325184 289176 325236
rect 289228 325224 289234 325236
rect 289354 325224 289360 325236
rect 289228 325196 289360 325224
rect 289228 325184 289234 325196
rect 289354 325184 289360 325196
rect 289412 325184 289418 325236
rect 224862 325116 224868 325168
rect 224920 325156 224926 325168
rect 261754 325156 261760 325168
rect 224920 325128 261760 325156
rect 224920 325116 224926 325128
rect 261754 325116 261760 325128
rect 261812 325116 261818 325168
rect 272702 325116 272708 325168
rect 272760 325156 272766 325168
rect 311894 325156 311900 325168
rect 272760 325128 311900 325156
rect 272760 325116 272766 325128
rect 311894 325116 311900 325128
rect 311952 325116 311958 325168
rect 148962 325048 148968 325100
rect 149020 325088 149026 325100
rect 253290 325088 253296 325100
rect 149020 325060 253296 325088
rect 149020 325048 149026 325060
rect 253290 325048 253296 325060
rect 253348 325048 253354 325100
rect 276842 325048 276848 325100
rect 276900 325088 276906 325100
rect 349154 325088 349160 325100
rect 276900 325060 349160 325088
rect 276900 325048 276906 325060
rect 349154 325048 349160 325060
rect 349212 325048 349218 325100
rect 128262 324980 128268 325032
rect 128320 325020 128326 325032
rect 249886 325020 249892 325032
rect 128320 324992 249892 325020
rect 128320 324980 128326 324992
rect 249886 324980 249892 324992
rect 249944 324980 249950 325032
rect 278682 324980 278688 325032
rect 278740 325020 278746 325032
rect 357526 325020 357532 325032
rect 278740 324992 357532 325020
rect 278740 324980 278746 324992
rect 357526 324980 357532 324992
rect 357584 324980 357590 325032
rect 92382 324912 92388 324964
rect 92440 324952 92446 324964
rect 246390 324952 246396 324964
rect 92440 324924 246396 324952
rect 92440 324912 92446 324924
rect 246390 324912 246396 324924
rect 246448 324912 246454 324964
rect 288710 324912 288716 324964
rect 288768 324952 288774 324964
rect 289354 324952 289360 324964
rect 288768 324924 289360 324952
rect 288768 324912 288774 324924
rect 289354 324912 289360 324924
rect 289412 324912 289418 324964
rect 297542 324912 297548 324964
rect 297600 324952 297606 324964
rect 516134 324952 516140 324964
rect 297600 324924 516140 324952
rect 297600 324912 297606 324924
rect 516134 324912 516140 324924
rect 516192 324912 516198 324964
rect 240686 323960 240692 324012
rect 240744 324000 240750 324012
rect 241146 324000 241152 324012
rect 240744 323972 241152 324000
rect 240744 323960 240750 323972
rect 241146 323960 241152 323972
rect 241204 323960 241210 324012
rect 274082 323824 274088 323876
rect 274140 323864 274146 323876
rect 322934 323864 322940 323876
rect 274140 323836 322940 323864
rect 274140 323824 274146 323836
rect 322934 323824 322940 323836
rect 322992 323824 322998 323876
rect 169570 323756 169576 323808
rect 169628 323796 169634 323808
rect 255222 323796 255228 323808
rect 169628 323768 255228 323796
rect 169628 323756 169634 323768
rect 255222 323756 255228 323768
rect 255280 323756 255286 323808
rect 278130 323756 278136 323808
rect 278188 323796 278194 323808
rect 360194 323796 360200 323808
rect 278188 323768 360200 323796
rect 278188 323756 278194 323768
rect 360194 323756 360200 323768
rect 360252 323756 360258 323808
rect 144730 323688 144736 323740
rect 144788 323728 144794 323740
rect 252186 323728 252192 323740
rect 144788 323700 252192 323728
rect 144788 323688 144794 323700
rect 252186 323688 252192 323700
rect 252244 323688 252250 323740
rect 282822 323688 282828 323740
rect 282880 323728 282886 323740
rect 393314 323728 393320 323740
rect 282880 323700 393320 323728
rect 282880 323688 282886 323700
rect 393314 323688 393320 323700
rect 393372 323688 393378 323740
rect 50982 323620 50988 323672
rect 51040 323660 51046 323672
rect 240226 323660 240232 323672
rect 51040 323632 240232 323660
rect 51040 323620 51046 323632
rect 240226 323620 240232 323632
rect 240284 323620 240290 323672
rect 285674 323620 285680 323672
rect 285732 323660 285738 323672
rect 430574 323660 430580 323672
rect 285732 323632 430580 323660
rect 285732 323620 285738 323632
rect 430574 323620 430580 323632
rect 430632 323620 430638 323672
rect 14458 323552 14464 323604
rect 14516 323592 14522 323604
rect 236546 323592 236552 323604
rect 14516 323564 236552 323592
rect 14516 323552 14522 323564
rect 236546 323552 236552 323564
rect 236604 323552 236610 323604
rect 296622 323552 296628 323604
rect 296680 323592 296686 323604
rect 506474 323592 506480 323604
rect 296680 323564 506480 323592
rect 296680 323552 296686 323564
rect 506474 323552 506480 323564
rect 506532 323552 506538 323604
rect 257154 322504 257160 322516
rect 253906 322476 257160 322504
rect 186222 322396 186228 322448
rect 186280 322436 186286 322448
rect 253906 322436 253934 322476
rect 257154 322464 257160 322476
rect 257212 322464 257218 322516
rect 186280 322408 253934 322436
rect 186280 322396 186286 322408
rect 255866 322396 255872 322448
rect 255924 322436 255930 322448
rect 256234 322436 256240 322448
rect 255924 322408 256240 322436
rect 255924 322396 255930 322408
rect 256234 322396 256240 322408
rect 256292 322396 256298 322448
rect 281442 322396 281448 322448
rect 281500 322436 281506 322448
rect 379514 322436 379520 322448
rect 281500 322408 379520 322436
rect 281500 322396 281506 322408
rect 379514 322396 379520 322408
rect 379572 322396 379578 322448
rect 135162 322328 135168 322380
rect 135220 322368 135226 322380
rect 250990 322368 250996 322380
rect 135220 322340 250996 322368
rect 135220 322328 135226 322340
rect 250990 322328 250996 322340
rect 251048 322328 251054 322380
rect 286410 322328 286416 322380
rect 286468 322368 286474 322380
rect 433334 322368 433340 322380
rect 286468 322340 433340 322368
rect 286468 322328 286474 322340
rect 433334 322328 433340 322340
rect 433392 322328 433398 322380
rect 88242 322260 88248 322312
rect 88300 322300 88306 322312
rect 245378 322300 245384 322312
rect 88300 322272 245384 322300
rect 88300 322260 88306 322272
rect 245378 322260 245384 322272
rect 245436 322260 245442 322312
rect 290550 322260 290556 322312
rect 290608 322300 290614 322312
rect 463694 322300 463700 322312
rect 290608 322272 463700 322300
rect 290608 322260 290614 322272
rect 463694 322260 463700 322272
rect 463752 322260 463758 322312
rect 57882 322192 57888 322244
rect 57940 322232 57946 322244
rect 241606 322232 241612 322244
rect 57940 322204 241612 322232
rect 57940 322192 57946 322204
rect 241606 322192 241612 322204
rect 241664 322192 241670 322244
rect 297634 322192 297640 322244
rect 297692 322232 297698 322244
rect 520274 322232 520280 322244
rect 297692 322204 520280 322232
rect 297692 322192 297698 322204
rect 520274 322192 520280 322204
rect 520332 322192 520338 322244
rect 272794 321104 272800 321156
rect 272852 321144 272858 321156
rect 316126 321144 316132 321156
rect 272852 321116 316132 321144
rect 272852 321104 272858 321116
rect 316126 321104 316132 321116
rect 316184 321104 316190 321156
rect 227530 321036 227536 321088
rect 227588 321076 227594 321088
rect 261386 321076 261392 321088
rect 227588 321048 261392 321076
rect 227588 321036 227594 321048
rect 261386 321036 261392 321048
rect 261444 321036 261450 321088
rect 275554 321036 275560 321088
rect 275612 321076 275618 321088
rect 336734 321076 336740 321088
rect 275612 321048 336740 321076
rect 275612 321036 275618 321048
rect 336734 321036 336740 321048
rect 336792 321036 336798 321088
rect 137922 320968 137928 321020
rect 137980 321008 137986 321020
rect 251542 321008 251548 321020
rect 137980 320980 251548 321008
rect 137980 320968 137986 320980
rect 251542 320968 251548 320980
rect 251600 320968 251606 321020
rect 282178 320968 282184 321020
rect 282236 321008 282242 321020
rect 397454 321008 397460 321020
rect 282236 320980 397460 321008
rect 282236 320968 282242 320980
rect 397454 320968 397460 320980
rect 397512 320968 397518 321020
rect 111702 320900 111708 320952
rect 111760 320940 111766 320952
rect 247494 320940 247500 320952
rect 111760 320912 247500 320940
rect 111760 320900 111766 320912
rect 247494 320900 247500 320912
rect 247552 320900 247558 320952
rect 294598 320900 294604 320952
rect 294656 320940 294662 320952
rect 458174 320940 458180 320952
rect 294656 320912 458180 320940
rect 294656 320900 294662 320912
rect 458174 320900 458180 320912
rect 458232 320900 458238 320952
rect 33778 320832 33784 320884
rect 33836 320872 33842 320884
rect 33836 320844 219434 320872
rect 33836 320832 33842 320844
rect 219406 320804 219434 320844
rect 236086 320832 236092 320884
rect 236144 320872 236150 320884
rect 236270 320872 236276 320884
rect 236144 320844 236276 320872
rect 236144 320832 236150 320844
rect 236270 320832 236276 320844
rect 236328 320832 236334 320884
rect 242894 320832 242900 320884
rect 242952 320872 242958 320884
rect 243078 320872 243084 320884
rect 242952 320844 243084 320872
rect 242952 320832 242958 320844
rect 243078 320832 243084 320844
rect 243136 320832 243142 320884
rect 298738 320832 298744 320884
rect 298796 320872 298802 320884
rect 533338 320872 533344 320884
rect 298796 320844 533344 320872
rect 298796 320832 298802 320844
rect 533338 320832 533344 320844
rect 533396 320832 533402 320884
rect 238294 320804 238300 320816
rect 219406 320776 238300 320804
rect 238294 320764 238300 320776
rect 238352 320764 238358 320816
rect 3050 320084 3056 320136
rect 3108 320124 3114 320136
rect 233050 320124 233056 320136
rect 3108 320096 233056 320124
rect 3108 320084 3114 320096
rect 233050 320084 233056 320096
rect 233108 320084 233114 320136
rect 272886 319608 272892 319660
rect 272944 319648 272950 319660
rect 318794 319648 318800 319660
rect 272944 319620 318800 319648
rect 272944 319608 272950 319620
rect 318794 319608 318800 319620
rect 318852 319608 318858 319660
rect 280706 319540 280712 319592
rect 280764 319580 280770 319592
rect 382274 319580 382280 319592
rect 280764 319552 382280 319580
rect 280764 319540 280770 319552
rect 382274 319540 382280 319552
rect 382332 319540 382338 319592
rect 220722 319472 220728 319524
rect 220780 319512 220786 319524
rect 261294 319512 261300 319524
rect 220780 319484 261300 319512
rect 220780 319472 220786 319484
rect 261294 319472 261300 319484
rect 261352 319472 261358 319524
rect 287606 319472 287612 319524
rect 287664 319512 287670 319524
rect 438854 319512 438860 319524
rect 287664 319484 438860 319512
rect 287664 319472 287670 319484
rect 438854 319472 438860 319484
rect 438912 319472 438918 319524
rect 106182 319404 106188 319456
rect 106240 319444 106246 319456
rect 247770 319444 247776 319456
rect 106240 319416 247776 319444
rect 106240 319404 106246 319416
rect 247770 319404 247776 319416
rect 247828 319404 247834 319456
rect 293494 319404 293500 319456
rect 293552 319444 293558 319456
rect 488534 319444 488540 319456
rect 293552 319416 488540 319444
rect 293552 319404 293558 319416
rect 488534 319404 488540 319416
rect 488592 319404 488598 319456
rect 274174 318248 274180 318300
rect 274232 318288 274238 318300
rect 329834 318288 329840 318300
rect 274232 318260 329840 318288
rect 274232 318248 274238 318260
rect 329834 318248 329840 318260
rect 329892 318248 329898 318300
rect 142062 318180 142068 318232
rect 142120 318220 142126 318232
rect 251450 318220 251456 318232
rect 142120 318192 251456 318220
rect 142120 318180 142126 318192
rect 251450 318180 251456 318192
rect 251508 318180 251514 318232
rect 283650 318180 283656 318232
rect 283708 318220 283714 318232
rect 400214 318220 400220 318232
rect 283708 318192 400220 318220
rect 283708 318180 283714 318192
rect 400214 318180 400220 318192
rect 400272 318180 400278 318232
rect 95050 318112 95056 318164
rect 95108 318152 95114 318164
rect 246114 318152 246120 318164
rect 95108 318124 246120 318152
rect 95108 318112 95114 318124
rect 246114 318112 246120 318124
rect 246172 318112 246178 318164
rect 288894 318112 288900 318164
rect 288952 318152 288958 318164
rect 448514 318152 448520 318164
rect 288952 318124 448520 318152
rect 288952 318112 288958 318124
rect 448514 318112 448520 318124
rect 448572 318112 448578 318164
rect 53742 318044 53748 318096
rect 53800 318084 53806 318096
rect 240134 318084 240140 318096
rect 53800 318056 240140 318084
rect 53800 318044 53806 318056
rect 240134 318044 240140 318056
rect 240192 318044 240198 318096
rect 293586 318044 293592 318096
rect 293644 318084 293650 318096
rect 491294 318084 491300 318096
rect 293644 318056 491300 318084
rect 293644 318044 293650 318056
rect 491294 318044 491300 318056
rect 491352 318044 491358 318096
rect 153102 316820 153108 316872
rect 153160 316860 153166 316872
rect 252922 316860 252928 316872
rect 153160 316832 252928 316860
rect 153160 316820 153166 316832
rect 252922 316820 252928 316832
rect 252980 316820 252986 316872
rect 275738 316820 275744 316872
rect 275796 316860 275802 316872
rect 332686 316860 332692 316872
rect 275796 316832 332692 316860
rect 275796 316820 275802 316832
rect 332686 316820 332692 316832
rect 332744 316820 332750 316872
rect 99282 316752 99288 316804
rect 99340 316792 99346 316804
rect 246022 316792 246028 316804
rect 99340 316764 246028 316792
rect 99340 316752 99346 316764
rect 246022 316752 246028 316764
rect 246080 316752 246086 316804
rect 288158 316752 288164 316804
rect 288216 316752 288222 316804
rect 289078 316752 289084 316804
rect 289136 316792 289142 316804
rect 452654 316792 452660 316804
rect 289136 316764 452660 316792
rect 289136 316752 289142 316764
rect 452654 316752 452660 316764
rect 452712 316752 452718 316804
rect 62022 316684 62028 316736
rect 62080 316724 62086 316736
rect 241514 316724 241520 316736
rect 62080 316696 241520 316724
rect 62080 316684 62086 316696
rect 241514 316684 241520 316696
rect 241572 316684 241578 316736
rect 288176 316600 288204 316752
rect 296070 316684 296076 316736
rect 296128 316724 296134 316736
rect 509234 316724 509240 316736
rect 296128 316696 509240 316724
rect 296128 316684 296134 316696
rect 509234 316684 509240 316696
rect 509292 316684 509298 316736
rect 288158 316548 288164 316600
rect 288216 316548 288222 316600
rect 155862 315392 155868 315444
rect 155920 315432 155926 315444
rect 252830 315432 252836 315444
rect 155920 315404 252836 315432
rect 155920 315392 155926 315404
rect 252830 315392 252836 315404
rect 252888 315392 252894 315444
rect 280798 315392 280804 315444
rect 280856 315432 280862 315444
rect 386414 315432 386420 315444
rect 280856 315404 386420 315432
rect 280856 315392 280862 315404
rect 386414 315392 386420 315404
rect 386472 315392 386478 315444
rect 103422 315324 103428 315376
rect 103480 315364 103486 315376
rect 247402 315364 247408 315376
rect 103480 315336 247408 315364
rect 103480 315324 103486 315336
rect 247402 315324 247408 315336
rect 247460 315324 247466 315376
rect 290734 315324 290740 315376
rect 290792 315364 290798 315376
rect 466454 315364 466460 315376
rect 290792 315336 466460 315364
rect 290792 315324 290798 315336
rect 466454 315324 466460 315336
rect 466512 315324 466518 315376
rect 71682 315256 71688 315308
rect 71740 315296 71746 315308
rect 236638 315296 236644 315308
rect 71740 315268 236644 315296
rect 71740 315256 71746 315268
rect 236638 315256 236644 315268
rect 236696 315256 236702 315308
rect 296162 315256 296168 315308
rect 296220 315296 296226 315308
rect 513374 315296 513380 315308
rect 296220 315268 513380 315296
rect 296220 315256 296226 315268
rect 513374 315256 513380 315268
rect 513432 315256 513438 315308
rect 276934 314032 276940 314084
rect 276992 314072 276998 314084
rect 343634 314072 343640 314084
rect 276992 314044 343640 314072
rect 276992 314032 276998 314044
rect 343634 314032 343640 314044
rect 343692 314032 343698 314084
rect 164142 313964 164148 314016
rect 164200 314004 164206 314016
rect 254670 314004 254676 314016
rect 164200 313976 254676 314004
rect 164200 313964 164206 313976
rect 254670 313964 254676 313976
rect 254728 313964 254734 314016
rect 297726 313964 297732 314016
rect 297784 314004 297790 314016
rect 522298 314004 522304 314016
rect 297784 313976 522304 314004
rect 297784 313964 297790 313976
rect 522298 313964 522304 313976
rect 522356 313964 522362 314016
rect 117222 313896 117228 313948
rect 117280 313936 117286 313948
rect 248966 313936 248972 313948
rect 117280 313908 248972 313936
rect 117280 313896 117286 313908
rect 248966 313896 248972 313908
rect 249024 313896 249030 313948
rect 285306 313896 285312 313948
rect 285364 313936 285370 313948
rect 285490 313936 285496 313948
rect 285364 313908 285496 313936
rect 285364 313896 285370 313908
rect 285490 313896 285496 313908
rect 285548 313896 285554 313948
rect 304258 313896 304264 313948
rect 304316 313936 304322 313948
rect 576118 313936 576124 313948
rect 304316 313908 576124 313936
rect 304316 313896 304322 313908
rect 576118 313896 576124 313908
rect 576176 313896 576182 313948
rect 306466 313216 306472 313268
rect 306524 313256 306530 313268
rect 580166 313256 580172 313268
rect 306524 313228 580172 313256
rect 306524 313216 306530 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 168282 312604 168288 312656
rect 168340 312644 168346 312656
rect 254394 312644 254400 312656
rect 168340 312616 254400 312644
rect 168340 312604 168346 312616
rect 254394 312604 254400 312616
rect 254452 312604 254458 312656
rect 274266 312604 274272 312656
rect 274324 312644 274330 312656
rect 325694 312644 325700 312656
rect 274324 312616 325700 312644
rect 274324 312604 274330 312616
rect 325694 312604 325700 312616
rect 325752 312604 325758 312656
rect 119982 312536 119988 312588
rect 120040 312576 120046 312588
rect 248874 312576 248880 312588
rect 120040 312548 248880 312576
rect 120040 312536 120046 312548
rect 248874 312536 248880 312548
rect 248932 312536 248938 312588
rect 278222 312536 278228 312588
rect 278280 312576 278286 312588
rect 354674 312576 354680 312588
rect 278280 312548 354680 312576
rect 278280 312536 278286 312548
rect 354674 312536 354680 312548
rect 354732 312536 354738 312588
rect 193122 311176 193128 311228
rect 193180 311216 193186 311228
rect 257062 311216 257068 311228
rect 193180 311188 257068 311216
rect 193180 311176 193186 311188
rect 257062 311176 257068 311188
rect 257120 311176 257126 311228
rect 286502 311176 286508 311228
rect 286560 311216 286566 311228
rect 432046 311216 432052 311228
rect 286560 311188 432052 311216
rect 286560 311176 286566 311188
rect 432046 311176 432052 311188
rect 432104 311176 432110 311228
rect 22738 311108 22744 311160
rect 22796 311148 22802 311160
rect 236362 311148 236368 311160
rect 22796 311120 236368 311148
rect 22796 311108 22802 311120
rect 236362 311108 236368 311120
rect 236420 311108 236426 311160
rect 302878 311108 302884 311160
rect 302936 311148 302942 311160
rect 571334 311148 571340 311160
rect 302936 311120 571340 311148
rect 302936 311108 302942 311120
rect 571334 311108 571340 311120
rect 571392 311108 571398 311160
rect 136450 309816 136456 309868
rect 136508 309856 136514 309868
rect 250254 309856 250260 309868
rect 136508 309828 250260 309856
rect 136508 309816 136514 309828
rect 250254 309816 250260 309828
rect 250312 309816 250318 309868
rect 275830 309816 275836 309868
rect 275888 309856 275894 309868
rect 340874 309856 340880 309868
rect 275888 309828 340880 309856
rect 275888 309816 275894 309828
rect 340874 309816 340880 309828
rect 340932 309816 340938 309868
rect 36538 309748 36544 309800
rect 36596 309788 36602 309800
rect 237926 309788 237932 309800
rect 36596 309760 237932 309788
rect 36596 309748 36602 309760
rect 237926 309748 237932 309760
rect 237984 309748 237990 309800
rect 287790 309748 287796 309800
rect 287848 309788 287854 309800
rect 445754 309788 445760 309800
rect 287848 309760 445760 309788
rect 287848 309748 287854 309760
rect 445754 309748 445760 309760
rect 445812 309748 445818 309800
rect 161382 308456 161388 308508
rect 161440 308496 161446 308508
rect 254302 308496 254308 308508
rect 161440 308468 254308 308496
rect 161440 308456 161446 308468
rect 254302 308456 254308 308468
rect 254360 308456 254366 308508
rect 284938 308456 284944 308508
rect 284996 308496 285002 308508
rect 390554 308496 390560 308508
rect 284996 308468 390560 308496
rect 284996 308456 285002 308468
rect 390554 308456 390560 308468
rect 390612 308456 390618 308508
rect 64782 308388 64788 308440
rect 64840 308428 64846 308440
rect 242066 308428 242072 308440
rect 64840 308400 242072 308428
rect 64840 308388 64846 308400
rect 242066 308388 242072 308400
rect 242124 308388 242130 308440
rect 289170 308388 289176 308440
rect 289228 308428 289234 308440
rect 456886 308428 456892 308440
rect 289228 308400 456892 308428
rect 289228 308388 289234 308400
rect 456886 308388 456892 308400
rect 456944 308388 456950 308440
rect 283742 307096 283748 307148
rect 283800 307136 283806 307148
rect 404354 307136 404360 307148
rect 283800 307108 404360 307136
rect 283800 307096 283806 307108
rect 404354 307096 404360 307108
rect 404412 307096 404418 307148
rect 81342 307028 81348 307080
rect 81400 307068 81406 307080
rect 234062 307068 234068 307080
rect 81400 307040 234068 307068
rect 81400 307028 81406 307040
rect 234062 307028 234068 307040
rect 234120 307028 234126 307080
rect 293402 307028 293408 307080
rect 293460 307068 293466 307080
rect 459554 307068 459560 307080
rect 293460 307040 459560 307068
rect 293460 307028 293466 307040
rect 459554 307028 459560 307040
rect 459612 307028 459618 307080
rect 283834 305668 283840 305720
rect 283892 305708 283898 305720
rect 407114 305708 407120 305720
rect 283892 305680 407120 305708
rect 283892 305668 283898 305680
rect 407114 305668 407120 305680
rect 407172 305668 407178 305720
rect 110322 305600 110328 305652
rect 110380 305640 110386 305652
rect 247310 305640 247316 305652
rect 110380 305612 247316 305640
rect 110380 305600 110386 305612
rect 247310 305600 247316 305612
rect 247368 305600 247374 305652
rect 293678 305600 293684 305652
rect 293736 305640 293742 305652
rect 481726 305640 481732 305652
rect 293736 305612 481732 305640
rect 293736 305600 293742 305612
rect 481726 305600 481732 305612
rect 481784 305600 481790 305652
rect 124122 304240 124128 304292
rect 124180 304280 124186 304292
rect 248782 304280 248788 304292
rect 124180 304252 248788 304280
rect 124180 304240 124186 304252
rect 248782 304240 248788 304252
rect 248840 304240 248846 304292
rect 293034 304240 293040 304292
rect 293092 304280 293098 304292
rect 485774 304280 485780 304292
rect 293092 304252 485780 304280
rect 293092 304240 293098 304252
rect 485774 304240 485780 304252
rect 485832 304240 485838 304292
rect 293126 302880 293132 302932
rect 293184 302920 293190 302932
rect 490006 302920 490012 302932
rect 293184 302892 490012 302920
rect 293184 302880 293190 302892
rect 490006 302880 490012 302892
rect 490064 302880 490070 302932
rect 297818 301452 297824 301504
rect 297876 301492 297882 301504
rect 517514 301492 517520 301504
rect 297876 301464 517520 301492
rect 297876 301452 297882 301464
rect 517514 301452 517520 301464
rect 517572 301452 517578 301504
rect 297910 300092 297916 300144
rect 297968 300132 297974 300144
rect 521654 300132 521660 300144
rect 297968 300104 521660 300132
rect 297968 300092 297974 300104
rect 521654 300092 521660 300104
rect 521712 300092 521718 300144
rect 306558 299412 306564 299464
rect 306616 299452 306622 299464
rect 580166 299452 580172 299464
rect 306616 299424 580172 299452
rect 306616 299412 306622 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 297450 297372 297456 297424
rect 297508 297412 297514 297424
rect 524414 297412 524420 297424
rect 297508 297384 524420 297412
rect 297508 297372 297514 297384
rect 524414 297372 524420 297384
rect 524472 297372 524478 297424
rect 305914 295944 305920 295996
rect 305972 295984 305978 295996
rect 556154 295984 556160 295996
rect 305972 295956 556160 295984
rect 305972 295944 305978 295956
rect 556154 295944 556160 295956
rect 556212 295944 556218 295996
rect 305822 294584 305828 294636
rect 305880 294624 305886 294636
rect 574094 294624 574100 294636
rect 305880 294596 574100 294624
rect 305880 294584 305886 294596
rect 574094 294584 574100 294596
rect 574152 294584 574158 294636
rect 277026 293224 277032 293276
rect 277084 293264 277090 293276
rect 350534 293264 350540 293276
rect 277084 293236 350540 293264
rect 277084 293224 277090 293236
rect 350534 293224 350540 293236
rect 350592 293224 350598 293276
rect 3142 293156 3148 293208
rect 3200 293196 3206 293208
rect 7558 293196 7564 293208
rect 3200 293168 7564 293196
rect 3200 293156 3206 293168
rect 7558 293156 7564 293168
rect 7616 293156 7622 293208
rect 278314 291796 278320 291848
rect 278372 291836 278378 291848
rect 361574 291836 361580 291848
rect 278372 291808 361580 291836
rect 278372 291796 278378 291808
rect 361574 291796 361580 291808
rect 361632 291796 361638 291848
rect 461578 285608 461584 285660
rect 461636 285648 461642 285660
rect 580166 285648 580172 285660
rect 461636 285620 580172 285648
rect 461636 285608 461642 285620
rect 580166 285608 580172 285620
rect 580224 285608 580230 285660
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 232958 280140 232964 280152
rect 3200 280112 232964 280140
rect 3200 280100 3206 280112
rect 232958 280100 232964 280112
rect 233016 280100 233022 280152
rect 316678 273164 316684 273216
rect 316736 273204 316742 273216
rect 580166 273204 580172 273216
rect 316736 273176 580172 273204
rect 316736 273164 316742 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 232866 267696 232872 267708
rect 3016 267668 232872 267696
rect 3016 267656 3022 267668
rect 232866 267656 232872 267668
rect 232924 267656 232930 267708
rect 331858 259360 331864 259412
rect 331916 259400 331922 259412
rect 580166 259400 580172 259412
rect 331916 259372 580172 259400
rect 331916 259360 331922 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 22830 255252 22836 255264
rect 3200 255224 22836 255252
rect 3200 255212 3206 255224
rect 22830 255212 22836 255224
rect 22888 255212 22894 255264
rect 306650 245556 306656 245608
rect 306708 245596 306714 245608
rect 580166 245596 580172 245608
rect 306708 245568 580172 245596
rect 306708 245556 306714 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 306742 233180 306748 233232
rect 306800 233220 306806 233232
rect 579982 233220 579988 233232
rect 306800 233192 579988 233220
rect 306800 233180 306806 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3234 229032 3240 229084
rect 3292 229072 3298 229084
rect 232774 229072 232780 229084
rect 3292 229044 232780 229072
rect 3292 229032 3298 229044
rect 232774 229032 232780 229044
rect 232832 229032 232838 229084
rect 306834 219376 306840 219428
rect 306892 219416 306898 219428
rect 580166 219416 580172 219428
rect 306892 219388 580172 219416
rect 306892 219376 306898 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3234 215228 3240 215280
rect 3292 215268 3298 215280
rect 232682 215268 232688 215280
rect 3292 215240 232688 215268
rect 3292 215228 3298 215240
rect 232682 215228 232688 215240
rect 232740 215228 232746 215280
rect 306926 206932 306932 206984
rect 306984 206972 306990 206984
rect 579798 206972 579804 206984
rect 306984 206944 579804 206972
rect 306984 206932 306990 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 309778 193128 309784 193180
rect 309836 193168 309842 193180
rect 580166 193168 580172 193180
rect 309836 193140 580172 193168
rect 309836 193128 309842 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 14550 189020 14556 189032
rect 3384 188992 14556 189020
rect 3384 188980 3390 188992
rect 14550 188980 14556 188992
rect 14608 188980 14614 189032
rect 305730 181432 305736 181484
rect 305788 181472 305794 181484
rect 483014 181472 483020 181484
rect 305788 181444 483020 181472
rect 305788 181432 305794 181444
rect 483014 181432 483020 181444
rect 483072 181432 483078 181484
rect 324958 179324 324964 179376
rect 325016 179364 325022 179376
rect 580166 179364 580172 179376
rect 325016 179336 580172 179364
rect 325016 179324 325022 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 3326 176604 3332 176656
rect 3384 176644 3390 176656
rect 232590 176644 232596 176656
rect 3384 176616 232596 176644
rect 3384 176604 3390 176616
rect 232590 176604 232596 176616
rect 232648 176604 232654 176656
rect 307662 166948 307668 167000
rect 307720 166988 307726 167000
rect 580166 166988 580172 167000
rect 307720 166960 580172 166988
rect 307720 166948 307726 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 307570 153144 307576 153196
rect 307628 153184 307634 153196
rect 580166 153184 580172 153196
rect 307628 153156 580172 153184
rect 307628 153144 307634 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 25498 150396 25504 150408
rect 3384 150368 25504 150396
rect 3384 150356 3390 150368
rect 25498 150356 25504 150368
rect 25556 150356 25562 150408
rect 307478 139340 307484 139392
rect 307536 139380 307542 139392
rect 580166 139380 580172 139392
rect 307536 139352 580172 139380
rect 307536 139340 307542 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 307386 126896 307392 126948
rect 307444 126936 307450 126948
rect 580166 126936 580172 126948
rect 307444 126908 580172 126936
rect 307444 126896 307450 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3142 124108 3148 124160
rect 3200 124148 3206 124160
rect 232498 124148 232504 124160
rect 3200 124120 232504 124148
rect 3200 124108 3206 124120
rect 232498 124108 232504 124120
rect 232556 124108 232562 124160
rect 307294 113092 307300 113144
rect 307352 113132 307358 113144
rect 579798 113132 579804 113144
rect 307352 113104 579804 113132
rect 307352 113092 307358 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 323578 100648 323584 100700
rect 323636 100688 323642 100700
rect 580166 100688 580172 100700
rect 323636 100660 580172 100688
rect 323636 100648 323642 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 307202 86912 307208 86964
rect 307260 86952 307266 86964
rect 580166 86952 580172 86964
rect 307260 86924 580172 86952
rect 307260 86912 307266 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 15838 85524 15844 85536
rect 3200 85496 15844 85524
rect 3200 85484 3206 85496
rect 15838 85484 15844 85496
rect 15896 85484 15902 85536
rect 307110 73108 307116 73160
rect 307168 73148 307174 73160
rect 580166 73148 580172 73160
rect 307168 73120 580172 73148
rect 307168 73108 307174 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 307018 60664 307024 60716
rect 307076 60704 307082 60716
rect 580166 60704 580172 60716
rect 307076 60676 580172 60704
rect 307076 60664 307082 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 2866 59304 2872 59356
rect 2924 59344 2930 59356
rect 32398 59344 32404 59356
rect 2924 59316 32404 59344
rect 2924 59304 2930 59316
rect 32398 59304 32404 59316
rect 32456 59304 32462 59356
rect 460198 46860 460204 46912
rect 460256 46900 460262 46912
rect 580166 46900 580172 46912
rect 460256 46872 580172 46900
rect 460256 46860 460262 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 335998 22720 336004 22772
rect 336056 22760 336062 22772
rect 462314 22760 462320 22772
rect 336056 22732 462320 22760
rect 336056 22720 336062 22732
rect 462314 22720 462320 22732
rect 462372 22720 462378 22772
rect 327718 21360 327724 21412
rect 327776 21400 327782 21412
rect 523126 21400 523132 21412
rect 327776 21372 523132 21400
rect 327776 21360 327782 21372
rect 523126 21360 523132 21372
rect 523184 21360 523190 21412
rect 318058 20612 318064 20664
rect 318116 20652 318122 20664
rect 579982 20652 579988 20664
rect 318116 20624 579988 20652
rect 318116 20612 318122 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 139302 19932 139308 19984
rect 139360 19972 139366 19984
rect 251910 19972 251916 19984
rect 139360 19944 251916 19972
rect 139360 19932 139366 19944
rect 251910 19932 251916 19944
rect 251968 19932 251974 19984
rect 322198 18572 322204 18624
rect 322256 18612 322262 18624
rect 505094 18612 505100 18624
rect 322256 18584 505100 18612
rect 322256 18572 322262 18584
rect 505094 18572 505100 18584
rect 505152 18572 505158 18624
rect 190362 17212 190368 17264
rect 190420 17252 190426 17264
rect 233970 17252 233976 17264
rect 190420 17224 233976 17252
rect 190420 17212 190426 17224
rect 233970 17212 233976 17224
rect 234028 17212 234034 17264
rect 320818 17212 320824 17264
rect 320876 17252 320882 17264
rect 498194 17252 498200 17264
rect 320876 17224 498200 17252
rect 320876 17212 320882 17224
rect 498194 17212 498200 17224
rect 498252 17212 498258 17264
rect 186130 15852 186136 15904
rect 186188 15892 186194 15904
rect 226978 15892 226984 15904
rect 186188 15864 226984 15892
rect 186188 15852 186194 15864
rect 226978 15852 226984 15864
rect 227036 15852 227042 15904
rect 313918 15852 313924 15904
rect 313976 15892 313982 15904
rect 494698 15892 494704 15904
rect 313976 15864 494704 15892
rect 313976 15852 313982 15864
rect 494698 15852 494704 15864
rect 494756 15852 494762 15904
rect 305638 14560 305644 14612
rect 305696 14600 305702 14612
rect 306742 14600 306748 14612
rect 305696 14572 306748 14600
rect 305696 14560 305702 14572
rect 306742 14560 306748 14572
rect 306800 14560 306806 14612
rect 171962 14424 171968 14476
rect 172020 14464 172026 14476
rect 229738 14464 229744 14476
rect 172020 14436 229744 14464
rect 172020 14424 172026 14436
rect 229738 14424 229744 14436
rect 229796 14424 229802 14476
rect 312538 14424 312544 14476
rect 312596 14464 312602 14476
rect 487614 14464 487620 14476
rect 312596 14436 487620 14464
rect 312596 14424 312602 14436
rect 487614 14424 487620 14436
rect 487672 14424 487678 14476
rect 301314 13744 301320 13796
rect 301372 13784 301378 13796
rect 301682 13784 301688 13796
rect 301372 13756 301688 13784
rect 301372 13744 301378 13756
rect 301682 13744 301688 13756
rect 301740 13744 301746 13796
rect 301682 13608 301688 13660
rect 301740 13648 301746 13660
rect 301866 13648 301872 13660
rect 301740 13620 301872 13648
rect 301740 13608 301746 13620
rect 301866 13608 301872 13620
rect 301924 13608 301930 13660
rect 298922 13540 298928 13592
rect 298980 13580 298986 13592
rect 532510 13580 532516 13592
rect 298980 13552 532516 13580
rect 298980 13540 298986 13552
rect 532510 13540 532516 13552
rect 532568 13540 532574 13592
rect 298830 13472 298836 13524
rect 298888 13512 298894 13524
rect 536098 13512 536104 13524
rect 298888 13484 536104 13512
rect 298888 13472 298894 13484
rect 536098 13472 536104 13484
rect 536156 13472 536162 13524
rect 300210 13404 300216 13456
rect 300268 13444 300274 13456
rect 539594 13444 539600 13456
rect 300268 13416 539600 13444
rect 300268 13404 300274 13416
rect 539594 13404 539600 13416
rect 539652 13404 539658 13456
rect 300118 13336 300124 13388
rect 300176 13376 300182 13388
rect 543182 13376 543188 13388
rect 300176 13348 543188 13376
rect 300176 13336 300182 13348
rect 543182 13336 543188 13348
rect 543240 13336 543246 13388
rect 300026 13268 300032 13320
rect 300084 13308 300090 13320
rect 546678 13308 546684 13320
rect 300084 13280 546684 13308
rect 300084 13268 300090 13280
rect 546678 13268 546684 13280
rect 546736 13268 546742 13320
rect 301406 13200 301412 13252
rect 301464 13240 301470 13252
rect 550266 13240 550272 13252
rect 301464 13212 550272 13240
rect 301464 13200 301470 13212
rect 550266 13200 550272 13212
rect 550324 13200 550330 13252
rect 301590 13132 301596 13184
rect 301648 13172 301654 13184
rect 553762 13172 553768 13184
rect 301648 13144 553768 13172
rect 301648 13132 301654 13144
rect 553762 13132 553768 13144
rect 553820 13132 553826 13184
rect 164878 13064 164884 13116
rect 164936 13104 164942 13116
rect 231118 13104 231124 13116
rect 164936 13076 231124 13104
rect 164936 13064 164942 13076
rect 231118 13064 231124 13076
rect 231176 13064 231182 13116
rect 235810 13064 235816 13116
rect 235868 13104 235874 13116
rect 261570 13104 261576 13116
rect 235868 13076 261576 13104
rect 235868 13064 235874 13076
rect 261570 13064 261576 13076
rect 261628 13064 261634 13116
rect 268470 13064 268476 13116
rect 268528 13104 268534 13116
rect 284294 13104 284300 13116
rect 268528 13076 284300 13104
rect 268528 13064 268534 13076
rect 284294 13064 284300 13076
rect 284352 13064 284358 13116
rect 293310 13064 293316 13116
rect 293368 13104 293374 13116
rect 293368 13076 296714 13104
rect 293368 13064 293374 13076
rect 296686 13036 296714 13076
rect 301498 13064 301504 13116
rect 301556 13104 301562 13116
rect 560846 13104 560852 13116
rect 301556 13076 560852 13104
rect 301556 13064 301562 13076
rect 560846 13064 560852 13076
rect 560904 13064 560910 13116
rect 301866 13036 301872 13048
rect 296686 13008 301872 13036
rect 301866 12996 301872 13008
rect 301924 12996 301930 13048
rect 291746 12384 291752 12436
rect 291804 12424 291810 12436
rect 471054 12424 471060 12436
rect 291804 12396 471060 12424
rect 291804 12384 291810 12396
rect 471054 12384 471060 12396
rect 471112 12384 471118 12436
rect 294782 12316 294788 12368
rect 294840 12356 294846 12368
rect 295245 12359 295303 12365
rect 294840 12328 295104 12356
rect 294840 12316 294846 12328
rect 294874 12248 294880 12300
rect 294932 12288 294938 12300
rect 294932 12260 295012 12288
rect 294932 12248 294938 12260
rect 293218 12112 293224 12164
rect 293276 12152 293282 12164
rect 294874 12152 294880 12164
rect 293276 12124 294880 12152
rect 293276 12112 293282 12124
rect 294874 12112 294880 12124
rect 294932 12112 294938 12164
rect 294984 12152 295012 12260
rect 295076 12220 295104 12328
rect 295245 12325 295257 12359
rect 295291 12356 295303 12359
rect 473354 12356 473360 12368
rect 295291 12328 473360 12356
rect 295291 12325 295303 12328
rect 295245 12319 295303 12325
rect 473354 12316 473360 12328
rect 473412 12316 473418 12368
rect 295153 12291 295211 12297
rect 295153 12257 295165 12291
rect 295199 12288 295211 12291
rect 478138 12288 478144 12300
rect 295199 12260 478144 12288
rect 295199 12257 295211 12260
rect 295153 12251 295211 12257
rect 478138 12248 478144 12260
rect 478196 12248 478202 12300
rect 493502 12220 493508 12232
rect 295076 12192 493508 12220
rect 493502 12180 493508 12192
rect 493560 12180 493566 12232
rect 497090 12152 497096 12164
rect 294984 12124 497096 12152
rect 497090 12112 497096 12124
rect 497148 12112 497154 12164
rect 294966 12044 294972 12096
rect 295024 12084 295030 12096
rect 500586 12084 500592 12096
rect 295024 12056 500592 12084
rect 295024 12044 295030 12056
rect 500586 12044 500592 12056
rect 500644 12044 500650 12096
rect 291930 11976 291936 12028
rect 291988 12016 291994 12028
rect 295153 12019 295211 12025
rect 295153 12016 295165 12019
rect 291988 11988 295165 12016
rect 291988 11976 291994 11988
rect 295153 11985 295165 11988
rect 295199 11985 295211 12019
rect 295153 11979 295211 11985
rect 295886 11976 295892 12028
rect 295944 12016 295950 12028
rect 504174 12016 504180 12028
rect 295944 11988 504180 12016
rect 295944 11976 295950 11988
rect 504174 11976 504180 11988
rect 504232 11976 504238 12028
rect 287698 11908 287704 11960
rect 287756 11948 287762 11960
rect 291378 11948 291384 11960
rect 287756 11920 291384 11948
rect 287756 11908 287762 11920
rect 291378 11908 291384 11920
rect 291436 11908 291442 11960
rect 291562 11908 291568 11960
rect 291620 11948 291626 11960
rect 295245 11951 295303 11957
rect 295245 11948 295257 11951
rect 291620 11920 295257 11948
rect 291620 11908 291626 11920
rect 295245 11917 295257 11920
rect 295291 11917 295303 11951
rect 295245 11911 295303 11917
rect 296254 11908 296260 11960
rect 296312 11948 296318 11960
rect 507670 11948 507676 11960
rect 296312 11920 507676 11948
rect 296312 11908 296318 11920
rect 507670 11908 507676 11920
rect 507728 11908 507734 11960
rect 296346 11840 296352 11892
rect 296404 11880 296410 11892
rect 511258 11880 511264 11892
rect 296404 11852 511264 11880
rect 296404 11840 296410 11852
rect 511258 11840 511264 11852
rect 511316 11840 511322 11892
rect 241422 11772 241428 11824
rect 241480 11812 241486 11824
rect 254578 11812 254584 11824
rect 241480 11784 254584 11812
rect 241480 11772 241486 11784
rect 254578 11772 254584 11784
rect 254636 11772 254642 11824
rect 296438 11772 296444 11824
rect 296496 11812 296502 11824
rect 514846 11812 514852 11824
rect 296496 11784 514852 11812
rect 296496 11772 296502 11784
rect 514846 11772 514852 11784
rect 514904 11772 514910 11824
rect 161290 11704 161296 11756
rect 161348 11744 161354 11756
rect 233878 11744 233884 11756
rect 161348 11716 233884 11744
rect 161348 11704 161354 11716
rect 233878 11704 233884 11716
rect 233936 11704 233942 11756
rect 237006 11704 237012 11756
rect 237064 11744 237070 11756
rect 257338 11744 257344 11756
rect 237064 11716 257344 11744
rect 237064 11704 237070 11716
rect 257338 11704 257344 11716
rect 257396 11704 257402 11756
rect 299014 11704 299020 11756
rect 299072 11744 299078 11756
rect 529014 11744 529020 11756
rect 299072 11716 529020 11744
rect 299072 11704 299078 11716
rect 529014 11704 529020 11716
rect 529072 11704 529078 11756
rect 221550 11432 221556 11484
rect 221608 11472 221614 11484
rect 224218 11472 224224 11484
rect 221608 11444 224224 11472
rect 221608 11432 221614 11444
rect 224218 11432 224224 11444
rect 224276 11432 224282 11484
rect 56502 10956 56508 11008
rect 56560 10996 56566 11008
rect 241974 10996 241980 11008
rect 56560 10968 241980 10996
rect 56560 10956 56566 10968
rect 241974 10956 241980 10968
rect 242032 10956 242038 11008
rect 282270 10956 282276 11008
rect 282328 10996 282334 11008
rect 393038 10996 393044 11008
rect 282328 10968 393044 10996
rect 282328 10956 282334 10968
rect 393038 10956 393044 10968
rect 393096 10956 393102 11008
rect 53650 10888 53656 10940
rect 53708 10928 53714 10940
rect 240686 10928 240692 10940
rect 53708 10900 240692 10928
rect 53708 10888 53714 10900
rect 240686 10888 240692 10900
rect 240744 10888 240750 10940
rect 282454 10888 282460 10940
rect 282512 10928 282518 10940
rect 396534 10928 396540 10940
rect 282512 10900 396540 10928
rect 282512 10888 282518 10900
rect 396534 10888 396540 10900
rect 396592 10888 396598 10940
rect 49602 10820 49608 10872
rect 49660 10860 49666 10872
rect 240594 10860 240600 10872
rect 49660 10832 240600 10860
rect 49660 10820 49666 10832
rect 240594 10820 240600 10832
rect 240652 10820 240658 10872
rect 282362 10820 282368 10872
rect 282420 10860 282426 10872
rect 398834 10860 398840 10872
rect 282420 10832 398840 10860
rect 282420 10820 282426 10832
rect 398834 10820 398840 10832
rect 398892 10820 398898 10872
rect 45462 10752 45468 10804
rect 45520 10792 45526 10804
rect 240502 10792 240508 10804
rect 45520 10764 240508 10792
rect 45520 10752 45526 10764
rect 240502 10752 240508 10764
rect 240560 10752 240566 10804
rect 284110 10752 284116 10804
rect 284168 10792 284174 10804
rect 403618 10792 403624 10804
rect 284168 10764 403624 10792
rect 284168 10752 284174 10764
rect 403618 10752 403624 10764
rect 403676 10752 403682 10804
rect 41322 10684 41328 10736
rect 41380 10724 41386 10736
rect 239122 10724 239128 10736
rect 41380 10696 239128 10724
rect 41380 10684 41386 10696
rect 239122 10684 239128 10696
rect 239180 10684 239186 10736
rect 284018 10684 284024 10736
rect 284076 10724 284082 10736
rect 407206 10724 407212 10736
rect 284076 10696 407212 10724
rect 284076 10684 284082 10696
rect 407206 10684 407212 10696
rect 407264 10684 407270 10736
rect 37182 10616 37188 10668
rect 37240 10656 37246 10668
rect 239306 10656 239312 10668
rect 37240 10628 239312 10656
rect 37240 10616 37246 10628
rect 239306 10616 239312 10628
rect 239364 10616 239370 10668
rect 283926 10616 283932 10668
rect 283984 10656 283990 10668
rect 410794 10656 410800 10668
rect 283984 10628 410800 10656
rect 283984 10616 283990 10628
rect 410794 10616 410800 10628
rect 410852 10616 410858 10668
rect 34422 10548 34428 10600
rect 34480 10588 34486 10600
rect 239214 10588 239220 10600
rect 34480 10560 239220 10588
rect 34480 10548 34486 10560
rect 239214 10548 239220 10560
rect 239272 10548 239278 10600
rect 285122 10548 285128 10600
rect 285180 10588 285186 10600
rect 414290 10588 414296 10600
rect 285180 10560 414296 10588
rect 285180 10548 285186 10560
rect 414290 10548 414296 10560
rect 414348 10548 414354 10600
rect 30098 10480 30104 10532
rect 30156 10520 30162 10532
rect 237834 10520 237840 10532
rect 30156 10492 237840 10520
rect 30156 10480 30162 10492
rect 237834 10480 237840 10492
rect 237892 10480 237898 10532
rect 285214 10480 285220 10532
rect 285272 10520 285278 10532
rect 417878 10520 417884 10532
rect 285272 10492 417884 10520
rect 285272 10480 285278 10492
rect 417878 10480 417884 10492
rect 417936 10480 417942 10532
rect 27522 10412 27528 10464
rect 27580 10452 27586 10464
rect 237650 10452 237656 10464
rect 27580 10424 237656 10452
rect 27580 10412 27586 10424
rect 237650 10412 237656 10424
rect 237708 10412 237714 10464
rect 285030 10412 285036 10464
rect 285088 10452 285094 10464
rect 421374 10452 421380 10464
rect 285088 10424 421380 10452
rect 285088 10412 285094 10424
rect 421374 10412 421380 10424
rect 421432 10412 421438 10464
rect 21818 10344 21824 10396
rect 21876 10384 21882 10396
rect 237742 10384 237748 10396
rect 21876 10356 237748 10384
rect 21876 10344 21882 10356
rect 237742 10344 237748 10356
rect 237800 10344 237806 10396
rect 244090 10344 244096 10396
rect 244148 10384 244154 10396
rect 253198 10384 253204 10396
rect 244148 10356 253204 10384
rect 244148 10344 244154 10356
rect 253198 10344 253204 10356
rect 253256 10344 253262 10396
rect 286594 10344 286600 10396
rect 286652 10384 286658 10396
rect 423766 10384 423772 10396
rect 286652 10356 423772 10384
rect 286652 10344 286658 10356
rect 423766 10344 423772 10356
rect 423824 10344 423830 10396
rect 9582 10276 9588 10328
rect 9640 10316 9646 10328
rect 235166 10316 235172 10328
rect 9640 10288 235172 10316
rect 9640 10276 9646 10288
rect 235166 10276 235172 10288
rect 235224 10276 235230 10328
rect 242802 10276 242808 10328
rect 242860 10316 242866 10328
rect 261478 10316 261484 10328
rect 242860 10288 261484 10316
rect 242860 10276 242866 10288
rect 261478 10276 261484 10288
rect 261536 10276 261542 10328
rect 286686 10276 286692 10328
rect 286744 10316 286750 10328
rect 428458 10316 428464 10328
rect 286744 10288 428464 10316
rect 286744 10276 286750 10288
rect 428458 10276 428464 10288
rect 428516 10276 428522 10328
rect 60642 10208 60648 10260
rect 60700 10248 60706 10260
rect 241882 10248 241888 10260
rect 60700 10220 241888 10248
rect 60700 10208 60706 10220
rect 241882 10208 241888 10220
rect 241940 10208 241946 10260
rect 282546 10208 282552 10260
rect 282604 10248 282610 10260
rect 389450 10248 389456 10260
rect 282604 10220 389456 10248
rect 282604 10208 282610 10220
rect 389450 10208 389456 10220
rect 389508 10208 389514 10260
rect 63218 10140 63224 10192
rect 63276 10180 63282 10192
rect 241790 10180 241796 10192
rect 63276 10152 241796 10180
rect 63276 10140 63282 10152
rect 241790 10140 241796 10152
rect 241848 10140 241854 10192
rect 281074 10140 281080 10192
rect 281132 10180 281138 10192
rect 385954 10180 385960 10192
rect 281132 10152 385960 10180
rect 281132 10140 281138 10152
rect 385954 10140 385960 10152
rect 386012 10140 386018 10192
rect 67542 10072 67548 10124
rect 67600 10112 67606 10124
rect 243354 10112 243360 10124
rect 67600 10084 243360 10112
rect 67600 10072 67606 10084
rect 243354 10072 243360 10084
rect 243412 10072 243418 10124
rect 280890 10072 280896 10124
rect 280948 10112 280954 10124
rect 382366 10112 382372 10124
rect 280948 10084 382372 10112
rect 280948 10072 280954 10084
rect 382366 10072 382372 10084
rect 382424 10072 382430 10124
rect 70302 10004 70308 10056
rect 70360 10044 70366 10056
rect 243446 10044 243452 10056
rect 70360 10016 243452 10044
rect 70360 10004 70366 10016
rect 243446 10004 243452 10016
rect 243504 10004 243510 10056
rect 280982 10004 280988 10056
rect 281040 10044 281046 10056
rect 378870 10044 378876 10056
rect 281040 10016 378876 10044
rect 281040 10004 281046 10016
rect 378870 10004 378876 10016
rect 378928 10004 378934 10056
rect 74442 9936 74448 9988
rect 74500 9976 74506 9988
rect 243262 9976 243268 9988
rect 74500 9948 243268 9976
rect 74500 9936 74506 9948
rect 243262 9936 243268 9948
rect 243320 9936 243326 9988
rect 279694 9936 279700 9988
rect 279752 9976 279758 9988
rect 373994 9976 374000 9988
rect 279752 9948 374000 9976
rect 279752 9936 279758 9948
rect 373994 9936 374000 9948
rect 374052 9936 374058 9988
rect 78582 9868 78588 9920
rect 78640 9908 78646 9920
rect 243538 9908 243544 9920
rect 78640 9880 243544 9908
rect 78640 9868 78646 9880
rect 243538 9868 243544 9880
rect 243596 9868 243602 9920
rect 279602 9868 279608 9920
rect 279660 9908 279666 9920
rect 371694 9908 371700 9920
rect 279660 9880 371700 9908
rect 279660 9868 279666 9880
rect 371694 9868 371700 9880
rect 371752 9868 371758 9920
rect 119890 9800 119896 9852
rect 119948 9840 119954 9852
rect 248598 9840 248604 9852
rect 119948 9812 248604 9840
rect 119948 9800 119954 9812
rect 248598 9800 248604 9812
rect 248656 9800 248662 9852
rect 279786 9800 279792 9852
rect 279844 9840 279850 9852
rect 368198 9840 368204 9852
rect 279844 9812 368204 9840
rect 279844 9800 279850 9812
rect 368198 9800 368204 9812
rect 368256 9800 368262 9852
rect 122742 9732 122748 9784
rect 122800 9772 122806 9784
rect 248690 9772 248696 9784
rect 122800 9744 248696 9772
rect 122800 9732 122806 9744
rect 248690 9732 248696 9744
rect 248748 9732 248754 9784
rect 278406 9732 278412 9784
rect 278464 9772 278470 9784
rect 364610 9772 364616 9784
rect 278464 9744 364616 9772
rect 278464 9732 278470 9744
rect 364610 9732 364616 9744
rect 364668 9732 364674 9784
rect 83274 9596 83280 9648
rect 83332 9636 83338 9648
rect 244734 9636 244740 9648
rect 83332 9608 244740 9636
rect 83332 9596 83338 9608
rect 244734 9596 244740 9608
rect 244792 9596 244798 9648
rect 253474 9596 253480 9648
rect 253532 9636 253538 9648
rect 255958 9636 255964 9648
rect 253532 9608 255964 9636
rect 253532 9596 253538 9608
rect 255958 9596 255964 9608
rect 256016 9596 256022 9648
rect 300394 9596 300400 9648
rect 300452 9636 300458 9648
rect 541986 9636 541992 9648
rect 300452 9608 541992 9636
rect 300452 9596 300458 9608
rect 541986 9596 541992 9608
rect 542044 9596 542050 9648
rect 79686 9528 79692 9580
rect 79744 9568 79750 9580
rect 244642 9568 244648 9580
rect 79744 9540 244648 9568
rect 79744 9528 79750 9540
rect 244642 9528 244648 9540
rect 244700 9528 244706 9580
rect 300486 9528 300492 9580
rect 300544 9568 300550 9580
rect 545482 9568 545488 9580
rect 300544 9540 545488 9568
rect 300544 9528 300550 9540
rect 545482 9528 545488 9540
rect 545540 9528 545546 9580
rect 76190 9460 76196 9512
rect 76248 9500 76254 9512
rect 243078 9500 243084 9512
rect 76248 9472 243084 9500
rect 76248 9460 76254 9472
rect 243078 9460 243084 9472
rect 243136 9460 243142 9512
rect 300302 9460 300308 9512
rect 300360 9500 300366 9512
rect 549070 9500 549076 9512
rect 300360 9472 549076 9500
rect 300360 9460 300366 9472
rect 549070 9460 549076 9472
rect 549128 9460 549134 9512
rect 72602 9392 72608 9444
rect 72660 9432 72666 9444
rect 243170 9432 243176 9444
rect 72660 9404 243176 9432
rect 72660 9392 72666 9404
rect 243170 9392 243176 9404
rect 243228 9392 243234 9444
rect 301774 9392 301780 9444
rect 301832 9432 301838 9444
rect 552658 9432 552664 9444
rect 301832 9404 552664 9432
rect 301832 9392 301838 9404
rect 552658 9392 552664 9404
rect 552716 9392 552722 9444
rect 69106 9324 69112 9376
rect 69164 9364 69170 9376
rect 242986 9364 242992 9376
rect 69164 9336 242992 9364
rect 69164 9324 69170 9336
rect 242986 9324 242992 9336
rect 243044 9324 243050 9376
rect 301314 9324 301320 9376
rect 301372 9364 301378 9376
rect 556246 9364 556252 9376
rect 301372 9336 556252 9364
rect 301372 9324 301378 9336
rect 556246 9324 556252 9336
rect 556304 9324 556310 9376
rect 65518 9256 65524 9308
rect 65576 9296 65582 9308
rect 242434 9296 242440 9308
rect 65576 9268 242440 9296
rect 65576 9256 65582 9268
rect 242434 9256 242440 9268
rect 242492 9256 242498 9308
rect 301682 9256 301688 9308
rect 301740 9296 301746 9308
rect 559742 9296 559748 9308
rect 301740 9268 559748 9296
rect 301740 9256 301746 9268
rect 559742 9256 559748 9268
rect 559800 9256 559806 9308
rect 61930 9188 61936 9240
rect 61988 9228 61994 9240
rect 242342 9228 242348 9240
rect 61988 9200 242348 9228
rect 61988 9188 61994 9200
rect 242342 9188 242348 9200
rect 242400 9188 242406 9240
rect 303062 9188 303068 9240
rect 303120 9228 303126 9240
rect 563238 9228 563244 9240
rect 303120 9200 563244 9228
rect 303120 9188 303126 9200
rect 563238 9188 563244 9200
rect 563296 9188 563302 9240
rect 58434 9120 58440 9172
rect 58492 9160 58498 9172
rect 241698 9160 241704 9172
rect 58492 9132 241704 9160
rect 58492 9120 58498 9132
rect 241698 9120 241704 9132
rect 241756 9120 241762 9172
rect 303154 9120 303160 9172
rect 303212 9160 303218 9172
rect 566826 9160 566832 9172
rect 303212 9132 566832 9160
rect 303212 9120 303218 9132
rect 566826 9120 566832 9132
rect 566884 9120 566890 9172
rect 54938 9052 54944 9104
rect 54996 9092 55002 9104
rect 240410 9092 240416 9104
rect 54996 9064 240416 9092
rect 54996 9052 55002 9064
rect 240410 9052 240416 9064
rect 240468 9052 240474 9104
rect 302970 9052 302976 9104
rect 303028 9092 303034 9104
rect 570322 9092 570328 9104
rect 303028 9064 570328 9092
rect 303028 9052 303034 9064
rect 570322 9052 570328 9064
rect 570380 9052 570386 9104
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 236270 9024 236276 9036
rect 17092 8996 236276 9024
rect 17092 8984 17098 8996
rect 236270 8984 236276 8996
rect 236328 8984 236334 9036
rect 247586 8984 247592 9036
rect 247644 9024 247650 9036
rect 263962 9024 263968 9036
rect 247644 8996 263968 9024
rect 247644 8984 247650 8996
rect 263962 8984 263968 8996
rect 264020 8984 264026 9036
rect 304442 8984 304448 9036
rect 304500 9024 304506 9036
rect 573910 9024 573916 9036
rect 304500 8996 573916 9024
rect 304500 8984 304506 8996
rect 573910 8984 573916 8996
rect 573968 8984 573974 9036
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 235074 8956 235080 8968
rect 4120 8928 235080 8956
rect 4120 8916 4126 8928
rect 235074 8916 235080 8928
rect 235132 8916 235138 8968
rect 238110 8916 238116 8968
rect 238168 8956 238174 8968
rect 262490 8956 262496 8968
rect 238168 8928 262496 8956
rect 238168 8916 238174 8928
rect 262490 8916 262496 8928
rect 262548 8916 262554 8968
rect 304350 8916 304356 8968
rect 304408 8956 304414 8968
rect 577406 8956 577412 8968
rect 304408 8928 577412 8956
rect 304408 8916 304414 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 86862 8848 86868 8900
rect 86920 8888 86926 8900
rect 244826 8888 244832 8900
rect 86920 8860 244832 8888
rect 86920 8848 86926 8860
rect 244826 8848 244832 8860
rect 244884 8848 244890 8900
rect 299106 8848 299112 8900
rect 299164 8888 299170 8900
rect 538398 8888 538404 8900
rect 299164 8860 538404 8888
rect 299164 8848 299170 8860
rect 538398 8848 538404 8860
rect 538456 8848 538462 8900
rect 90358 8780 90364 8832
rect 90416 8820 90422 8832
rect 245930 8820 245936 8832
rect 90416 8792 245936 8820
rect 90416 8780 90422 8792
rect 245930 8780 245936 8792
rect 245988 8780 245994 8832
rect 273806 8780 273812 8832
rect 273864 8820 273870 8832
rect 329190 8820 329196 8832
rect 273864 8792 329196 8820
rect 273864 8780 273870 8792
rect 329190 8780 329196 8792
rect 329248 8780 329254 8832
rect 142430 8712 142436 8764
rect 142488 8752 142494 8764
rect 251634 8752 251640 8764
rect 142488 8724 251640 8752
rect 142488 8712 142494 8724
rect 251634 8712 251640 8724
rect 251692 8712 251698 8764
rect 274358 8712 274364 8764
rect 274416 8752 274422 8764
rect 325602 8752 325608 8764
rect 274416 8724 325608 8752
rect 274416 8712 274422 8724
rect 325602 8712 325608 8724
rect 325660 8712 325666 8764
rect 145926 8644 145932 8696
rect 145984 8684 145990 8696
rect 251726 8684 251732 8696
rect 145984 8656 251732 8684
rect 145984 8644 145990 8656
rect 251726 8644 251732 8656
rect 251784 8644 251790 8696
rect 273714 8644 273720 8696
rect 273772 8684 273778 8696
rect 322106 8684 322112 8696
rect 273772 8656 322112 8684
rect 273772 8644 273778 8656
rect 322106 8644 322112 8656
rect 322164 8644 322170 8696
rect 149514 8576 149520 8628
rect 149572 8616 149578 8628
rect 253382 8616 253388 8628
rect 149572 8588 253388 8616
rect 149572 8576 149578 8588
rect 253382 8576 253388 8588
rect 253440 8576 253446 8628
rect 272610 8576 272616 8628
rect 272668 8616 272674 8628
rect 318518 8616 318524 8628
rect 272668 8588 318524 8616
rect 272668 8576 272674 8588
rect 318518 8576 318524 8588
rect 318576 8576 318582 8628
rect 153010 8508 153016 8560
rect 153068 8548 153074 8560
rect 253106 8548 253112 8560
rect 153068 8520 253112 8548
rect 153068 8508 153074 8520
rect 253106 8508 253112 8520
rect 253164 8508 253170 8560
rect 273070 8508 273076 8560
rect 273128 8548 273134 8560
rect 315022 8548 315028 8560
rect 273128 8520 315028 8548
rect 273128 8508 273134 8520
rect 315022 8508 315028 8520
rect 315080 8508 315086 8560
rect 156598 8440 156604 8492
rect 156656 8480 156662 8492
rect 253014 8480 253020 8492
rect 156656 8452 253020 8480
rect 156656 8440 156662 8452
rect 253014 8440 253020 8452
rect 253072 8440 253078 8492
rect 272978 8440 272984 8492
rect 273036 8480 273042 8492
rect 311434 8480 311440 8492
rect 273036 8452 311440 8480
rect 273036 8440 273042 8452
rect 311434 8440 311440 8452
rect 311492 8440 311498 8492
rect 271322 8372 271328 8424
rect 271380 8412 271386 8424
rect 307938 8412 307944 8424
rect 271380 8384 307944 8412
rect 271380 8372 271386 8384
rect 307938 8372 307944 8384
rect 307996 8372 308002 8424
rect 199102 8236 199108 8288
rect 199160 8276 199166 8288
rect 258902 8276 258908 8288
rect 199160 8248 258908 8276
rect 199160 8236 199166 8248
rect 258902 8236 258908 8248
rect 258960 8236 258966 8288
rect 287882 8236 287888 8288
rect 287940 8276 287946 8288
rect 441522 8276 441528 8288
rect 287940 8248 441528 8276
rect 287940 8236 287946 8248
rect 441522 8236 441528 8248
rect 441580 8236 441586 8288
rect 195606 8168 195612 8220
rect 195664 8208 195670 8220
rect 258718 8208 258724 8220
rect 195664 8180 258724 8208
rect 195664 8168 195670 8180
rect 258718 8168 258724 8180
rect 258776 8168 258782 8220
rect 288066 8168 288072 8220
rect 288124 8208 288130 8220
rect 445018 8208 445024 8220
rect 288124 8180 445024 8208
rect 288124 8168 288130 8180
rect 445018 8168 445024 8180
rect 445076 8168 445082 8220
rect 181438 8100 181444 8152
rect 181496 8140 181502 8152
rect 255682 8140 255688 8152
rect 181496 8112 255688 8140
rect 181496 8100 181502 8112
rect 255682 8100 255688 8112
rect 255740 8100 255746 8152
rect 289354 8100 289360 8152
rect 289412 8140 289418 8152
rect 448606 8140 448612 8152
rect 289412 8112 448612 8140
rect 289412 8100 289418 8112
rect 448606 8100 448612 8112
rect 448664 8100 448670 8152
rect 177850 8032 177856 8084
rect 177908 8072 177914 8084
rect 255866 8072 255872 8084
rect 177908 8044 255872 8072
rect 177908 8032 177914 8044
rect 255866 8032 255872 8044
rect 255924 8032 255930 8084
rect 289262 8032 289268 8084
rect 289320 8072 289326 8084
rect 452102 8072 452108 8084
rect 289320 8044 452108 8072
rect 289320 8032 289326 8044
rect 452102 8032 452108 8044
rect 452160 8032 452166 8084
rect 174262 7964 174268 8016
rect 174320 8004 174326 8016
rect 255590 8004 255596 8016
rect 174320 7976 255596 8004
rect 174320 7964 174326 7976
rect 255590 7964 255596 7976
rect 255648 7964 255654 8016
rect 289446 7964 289452 8016
rect 289504 8004 289510 8016
rect 455690 8004 455696 8016
rect 289504 7976 455696 8004
rect 289504 7964 289510 7976
rect 455690 7964 455696 7976
rect 455748 7964 455754 8016
rect 170766 7896 170772 7948
rect 170824 7936 170830 7948
rect 255774 7936 255780 7948
rect 170824 7908 255780 7936
rect 170824 7896 170830 7908
rect 255774 7896 255780 7908
rect 255832 7896 255838 7948
rect 292114 7896 292120 7948
rect 292172 7936 292178 7948
rect 469858 7936 469864 7948
rect 292172 7908 469864 7936
rect 292172 7896 292178 7908
rect 469858 7896 469864 7908
rect 469916 7896 469922 7948
rect 131758 7828 131764 7880
rect 131816 7868 131822 7880
rect 250070 7868 250076 7880
rect 131816 7840 250076 7868
rect 131816 7828 131822 7840
rect 250070 7828 250076 7840
rect 250128 7828 250134 7880
rect 292022 7828 292028 7880
rect 292080 7868 292086 7880
rect 473446 7868 473452 7880
rect 292080 7840 473452 7868
rect 292080 7828 292086 7840
rect 473446 7828 473452 7840
rect 473504 7828 473510 7880
rect 128170 7760 128176 7812
rect 128228 7800 128234 7812
rect 250162 7800 250168 7812
rect 128228 7772 250168 7800
rect 128228 7760 128234 7772
rect 250162 7760 250168 7772
rect 250220 7760 250226 7812
rect 292206 7760 292212 7812
rect 292264 7800 292270 7812
rect 476942 7800 476948 7812
rect 292264 7772 476948 7800
rect 292264 7760 292270 7772
rect 476942 7760 476948 7772
rect 477000 7760 477006 7812
rect 51350 7692 51356 7744
rect 51408 7732 51414 7744
rect 240870 7732 240876 7744
rect 51408 7704 240876 7732
rect 51408 7692 51414 7704
rect 240870 7692 240876 7704
rect 240928 7692 240934 7744
rect 294138 7692 294144 7744
rect 294196 7732 294202 7744
rect 495894 7732 495900 7744
rect 294196 7704 495900 7732
rect 294196 7692 294202 7704
rect 495894 7692 495900 7704
rect 495952 7692 495958 7744
rect 47854 7624 47860 7676
rect 47912 7664 47918 7676
rect 240962 7664 240968 7676
rect 47912 7636 240968 7664
rect 47912 7624 47918 7636
rect 240962 7624 240968 7636
rect 241020 7624 241026 7676
rect 295150 7624 295156 7676
rect 295208 7664 295214 7676
rect 499390 7664 499396 7676
rect 295208 7636 499396 7664
rect 295208 7624 295214 7636
rect 499390 7624 499396 7636
rect 499448 7624 499454 7676
rect 12342 7556 12348 7608
rect 12400 7596 12406 7608
rect 236178 7596 236184 7608
rect 12400 7568 236184 7596
rect 12400 7556 12406 7568
rect 236178 7556 236184 7568
rect 236236 7556 236242 7608
rect 276658 7556 276664 7608
rect 276716 7596 276722 7608
rect 280706 7596 280712 7608
rect 276716 7568 280712 7596
rect 276716 7556 276722 7568
rect 280706 7556 280712 7568
rect 280764 7556 280770 7608
rect 295058 7556 295064 7608
rect 295116 7596 295122 7608
rect 502978 7596 502984 7608
rect 295116 7568 502984 7596
rect 295116 7556 295122 7568
rect 502978 7556 502984 7568
rect 503036 7556 503042 7608
rect 202690 7488 202696 7540
rect 202748 7528 202754 7540
rect 258810 7528 258816 7540
rect 202748 7500 258816 7528
rect 202748 7488 202754 7500
rect 258810 7488 258816 7500
rect 258868 7488 258874 7540
rect 287974 7488 287980 7540
rect 288032 7528 288038 7540
rect 437934 7528 437940 7540
rect 288032 7500 437940 7528
rect 288032 7488 288038 7500
rect 437934 7488 437940 7500
rect 437992 7488 437998 7540
rect 206186 7420 206192 7472
rect 206244 7460 206250 7472
rect 260098 7460 260104 7472
rect 206244 7432 260104 7460
rect 206244 7420 206250 7432
rect 260098 7420 260104 7432
rect 260156 7420 260162 7472
rect 286318 6876 286324 6928
rect 286376 6916 286382 6928
rect 287790 6916 287796 6928
rect 286376 6888 287796 6916
rect 286376 6876 286382 6888
rect 287790 6876 287796 6888
rect 287848 6876 287854 6928
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 17218 6848 17224 6860
rect 3476 6820 17224 6848
rect 3476 6808 3482 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 215662 6808 215668 6860
rect 215720 6848 215726 6860
rect 259822 6848 259828 6860
rect 215720 6820 259828 6848
rect 215720 6808 215726 6820
rect 259822 6808 259828 6820
rect 259880 6808 259886 6860
rect 279878 6808 279884 6860
rect 279936 6848 279942 6860
rect 367002 6848 367008 6860
rect 279936 6820 367008 6848
rect 279936 6808 279942 6820
rect 367002 6808 367008 6820
rect 367060 6808 367066 6860
rect 406378 6808 406384 6860
rect 406436 6848 406442 6860
rect 580166 6848 580172 6860
rect 406436 6820 580172 6848
rect 406436 6808 406442 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 212166 6740 212172 6792
rect 212224 6780 212230 6792
rect 259730 6780 259736 6792
rect 212224 6752 259736 6780
rect 212224 6740 212230 6752
rect 259730 6740 259736 6752
rect 259788 6740 259794 6792
rect 279510 6740 279516 6792
rect 279568 6780 279574 6792
rect 370590 6780 370596 6792
rect 279568 6752 370596 6780
rect 279568 6740 279574 6752
rect 370590 6740 370596 6752
rect 370648 6740 370654 6792
rect 208578 6672 208584 6724
rect 208636 6712 208642 6724
rect 259914 6712 259920 6724
rect 208636 6684 259920 6712
rect 208636 6672 208642 6684
rect 259914 6672 259920 6684
rect 259972 6672 259978 6724
rect 279418 6672 279424 6724
rect 279476 6712 279482 6724
rect 374086 6712 374092 6724
rect 279476 6684 374092 6712
rect 279476 6672 279482 6684
rect 374086 6672 374092 6684
rect 374144 6672 374150 6724
rect 205082 6604 205088 6656
rect 205140 6644 205146 6656
rect 260006 6644 260012 6656
rect 205140 6616 260012 6644
rect 205140 6604 205146 6616
rect 260006 6604 260012 6616
rect 260064 6604 260070 6656
rect 281166 6604 281172 6656
rect 281224 6644 281230 6656
rect 377674 6644 377680 6656
rect 281224 6616 377680 6644
rect 281224 6604 281230 6616
rect 377674 6604 377680 6616
rect 377732 6604 377738 6656
rect 201494 6536 201500 6588
rect 201552 6576 201558 6588
rect 258442 6576 258448 6588
rect 201552 6548 258448 6576
rect 201552 6536 201558 6548
rect 258442 6536 258448 6548
rect 258500 6536 258506 6588
rect 281258 6536 281264 6588
rect 281316 6576 281322 6588
rect 381170 6576 381176 6588
rect 281316 6548 381176 6576
rect 281316 6536 281322 6548
rect 381170 6536 381176 6548
rect 381228 6536 381234 6588
rect 197906 6468 197912 6520
rect 197964 6508 197970 6520
rect 258626 6508 258632 6520
rect 197964 6480 258632 6508
rect 197964 6468 197970 6480
rect 258626 6468 258632 6480
rect 258684 6468 258690 6520
rect 280614 6468 280620 6520
rect 280672 6508 280678 6520
rect 384758 6508 384764 6520
rect 280672 6480 384764 6508
rect 280672 6468 280678 6480
rect 384758 6468 384764 6480
rect 384816 6468 384822 6520
rect 194410 6400 194416 6452
rect 194468 6440 194474 6452
rect 258534 6440 258540 6452
rect 194468 6412 258540 6440
rect 194468 6400 194474 6412
rect 258534 6400 258540 6412
rect 258592 6400 258598 6452
rect 281350 6400 281356 6452
rect 281408 6440 281414 6452
rect 388254 6440 388260 6452
rect 281408 6412 388260 6440
rect 281408 6400 281414 6412
rect 388254 6400 388260 6412
rect 388312 6400 388318 6452
rect 180242 6332 180248 6384
rect 180300 6372 180306 6384
rect 255498 6372 255504 6384
rect 180300 6344 255504 6372
rect 180300 6332 180306 6344
rect 255498 6332 255504 6344
rect 255556 6332 255562 6384
rect 282730 6332 282736 6384
rect 282788 6372 282794 6384
rect 391842 6372 391848 6384
rect 282788 6344 391848 6372
rect 282788 6332 282794 6344
rect 391842 6332 391848 6344
rect 391900 6332 391906 6384
rect 176654 6264 176660 6316
rect 176712 6304 176718 6316
rect 255406 6304 255412 6316
rect 176712 6276 255412 6304
rect 176712 6264 176718 6276
rect 255406 6264 255412 6276
rect 255464 6264 255470 6316
rect 282086 6264 282092 6316
rect 282144 6304 282150 6316
rect 395338 6304 395344 6316
rect 282144 6276 395344 6304
rect 282144 6264 282150 6276
rect 395338 6264 395344 6276
rect 395396 6264 395402 6316
rect 173158 6196 173164 6248
rect 173216 6236 173222 6248
rect 256142 6236 256148 6248
rect 173216 6208 256148 6236
rect 173216 6196 173222 6208
rect 256142 6196 256148 6208
rect 256200 6196 256206 6248
rect 282638 6196 282644 6248
rect 282696 6236 282702 6248
rect 398926 6236 398932 6248
rect 282696 6208 398932 6236
rect 282696 6196 282702 6208
rect 398926 6196 398932 6208
rect 398984 6196 398990 6248
rect 400858 6196 400864 6248
rect 400916 6236 400922 6248
rect 409598 6236 409604 6248
rect 400916 6208 409604 6236
rect 400916 6196 400922 6208
rect 409598 6196 409604 6208
rect 409656 6196 409662 6248
rect 130562 6128 130568 6180
rect 130620 6168 130626 6180
rect 249978 6168 249984 6180
rect 130620 6140 249984 6168
rect 130620 6128 130626 6140
rect 249978 6128 249984 6140
rect 250036 6128 250042 6180
rect 283466 6128 283472 6180
rect 283524 6168 283530 6180
rect 402514 6168 402520 6180
rect 283524 6140 402520 6168
rect 283524 6128 283530 6140
rect 402514 6128 402520 6140
rect 402572 6128 402578 6180
rect 277854 6060 277860 6112
rect 277912 6100 277918 6112
rect 363506 6100 363512 6112
rect 277912 6072 363512 6100
rect 277912 6060 277918 6072
rect 363506 6060 363512 6072
rect 363564 6060 363570 6112
rect 277946 5992 277952 6044
rect 278004 6032 278010 6044
rect 359918 6032 359924 6044
rect 278004 6004 359924 6032
rect 278004 5992 278010 6004
rect 359918 5992 359924 6004
rect 359976 5992 359982 6044
rect 278498 5924 278504 5976
rect 278556 5964 278562 5976
rect 356330 5964 356336 5976
rect 278556 5936 356336 5964
rect 278556 5924 278562 5936
rect 356330 5924 356336 5936
rect 356388 5924 356394 5976
rect 276566 5856 276572 5908
rect 276624 5896 276630 5908
rect 352834 5896 352840 5908
rect 276624 5868 352840 5896
rect 276624 5856 276630 5868
rect 352834 5856 352840 5868
rect 352892 5856 352898 5908
rect 276474 5788 276480 5840
rect 276532 5828 276538 5840
rect 349246 5828 349252 5840
rect 276532 5800 349252 5828
rect 276532 5788 276538 5800
rect 349246 5788 349252 5800
rect 349304 5788 349310 5840
rect 276382 5720 276388 5772
rect 276440 5760 276446 5772
rect 345750 5760 345756 5772
rect 276440 5732 345756 5760
rect 276440 5720 276446 5732
rect 345750 5720 345756 5732
rect 345808 5720 345814 5772
rect 275462 5652 275468 5704
rect 275520 5692 275526 5704
rect 342162 5692 342168 5704
rect 275520 5664 342168 5692
rect 275520 5652 275526 5664
rect 342162 5652 342168 5664
rect 342220 5652 342226 5704
rect 268562 5584 268568 5636
rect 268620 5624 268626 5636
rect 274818 5624 274824 5636
rect 268620 5596 274824 5624
rect 268620 5584 268626 5596
rect 274818 5584 274824 5596
rect 274876 5584 274882 5636
rect 249245 5559 249303 5565
rect 249245 5525 249257 5559
rect 249291 5556 249303 5559
rect 250438 5556 250444 5568
rect 249291 5528 250444 5556
rect 249291 5525 249303 5528
rect 249245 5519 249303 5525
rect 250438 5516 250444 5528
rect 250496 5516 250502 5568
rect 273898 5516 273904 5568
rect 273956 5556 273962 5568
rect 279510 5556 279516 5568
rect 273956 5528 279516 5556
rect 273956 5516 273962 5528
rect 279510 5516 279516 5528
rect 279568 5516 279574 5568
rect 479518 5516 479524 5568
rect 479576 5556 479582 5568
rect 480530 5556 480536 5568
rect 479576 5528 480536 5556
rect 479576 5516 479582 5528
rect 480530 5516 480536 5528
rect 480588 5516 480594 5568
rect 207382 5448 207388 5500
rect 207440 5488 207446 5500
rect 259638 5488 259644 5500
rect 207440 5460 259644 5488
rect 207440 5448 207446 5460
rect 259638 5448 259644 5460
rect 259696 5448 259702 5500
rect 270310 5448 270316 5500
rect 270368 5488 270374 5500
rect 286594 5488 286600 5500
rect 270368 5460 286600 5488
rect 270368 5448 270374 5460
rect 286594 5448 286600 5460
rect 286652 5448 286658 5500
rect 300670 5448 300676 5500
rect 300728 5488 300734 5500
rect 540790 5488 540796 5500
rect 300728 5460 540796 5488
rect 300728 5448 300734 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 203886 5380 203892 5432
rect 203944 5420 203950 5432
rect 258258 5420 258264 5432
rect 203944 5392 258264 5420
rect 203944 5380 203950 5392
rect 258258 5380 258264 5392
rect 258316 5380 258322 5432
rect 270126 5380 270132 5432
rect 270184 5420 270190 5432
rect 288986 5420 288992 5432
rect 270184 5392 288992 5420
rect 270184 5380 270190 5392
rect 288986 5380 288992 5392
rect 289044 5380 289050 5432
rect 300578 5380 300584 5432
rect 300636 5420 300642 5432
rect 544378 5420 544384 5432
rect 300636 5392 544384 5420
rect 300636 5380 300642 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 200298 5312 200304 5364
rect 200356 5352 200362 5364
rect 258350 5352 258356 5364
rect 200356 5324 258356 5352
rect 200356 5312 200362 5324
rect 258350 5312 258356 5324
rect 258408 5312 258414 5364
rect 269850 5312 269856 5364
rect 269908 5352 269914 5364
rect 290182 5352 290188 5364
rect 269908 5324 290188 5352
rect 269908 5312 269914 5324
rect 290182 5312 290188 5324
rect 290240 5312 290246 5364
rect 300762 5312 300768 5364
rect 300820 5352 300826 5364
rect 547874 5352 547880 5364
rect 300820 5324 547880 5352
rect 300820 5312 300826 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 196802 5244 196808 5296
rect 196860 5284 196866 5296
rect 258166 5284 258172 5296
rect 196860 5256 258172 5284
rect 196860 5244 196866 5256
rect 258166 5244 258172 5256
rect 258224 5244 258230 5296
rect 270402 5244 270408 5296
rect 270460 5284 270466 5296
rect 293678 5284 293684 5296
rect 270460 5256 293684 5284
rect 270460 5244 270466 5256
rect 293678 5244 293684 5256
rect 293736 5244 293742 5296
rect 301958 5244 301964 5296
rect 302016 5284 302022 5296
rect 551462 5284 551468 5296
rect 302016 5256 551468 5284
rect 302016 5244 302022 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 193214 5176 193220 5228
rect 193272 5216 193278 5228
rect 258074 5216 258080 5228
rect 193272 5188 258080 5216
rect 193272 5176 193278 5188
rect 258074 5176 258080 5188
rect 258132 5176 258138 5228
rect 270218 5176 270224 5228
rect 270276 5216 270282 5228
rect 292574 5216 292580 5228
rect 270276 5188 292580 5216
rect 270276 5176 270282 5188
rect 292574 5176 292580 5188
rect 292632 5176 292638 5228
rect 302050 5176 302056 5228
rect 302108 5216 302114 5228
rect 554958 5216 554964 5228
rect 302108 5188 554964 5216
rect 302108 5176 302114 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 132954 5108 132960 5160
rect 133012 5148 133018 5160
rect 249245 5151 249303 5157
rect 249245 5148 249257 5151
rect 133012 5120 249257 5148
rect 133012 5108 133018 5120
rect 249245 5117 249257 5120
rect 249291 5117 249303 5151
rect 250346 5148 250352 5160
rect 249245 5111 249303 5117
rect 249352 5120 250352 5148
rect 129366 5040 129372 5092
rect 129424 5080 129430 5092
rect 249352 5080 249380 5120
rect 250346 5108 250352 5120
rect 250404 5108 250410 5160
rect 271414 5108 271420 5160
rect 271472 5148 271478 5160
rect 297266 5148 297272 5160
rect 271472 5120 297272 5148
rect 271472 5108 271478 5120
rect 297266 5108 297272 5120
rect 297324 5108 297330 5160
rect 302142 5108 302148 5160
rect 302200 5148 302206 5160
rect 558546 5148 558552 5160
rect 302200 5120 558552 5148
rect 302200 5108 302206 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 129424 5052 249380 5080
rect 129424 5040 129430 5052
rect 249978 5040 249984 5092
rect 250036 5080 250042 5092
rect 264422 5080 264428 5092
rect 250036 5052 264428 5080
rect 250036 5040 250042 5052
rect 264422 5040 264428 5052
rect 264480 5040 264486 5092
rect 270034 5040 270040 5092
rect 270092 5080 270098 5092
rect 296070 5080 296076 5092
rect 270092 5052 296076 5080
rect 270092 5040 270098 5052
rect 296070 5040 296076 5052
rect 296128 5040 296134 5092
rect 303338 5040 303344 5092
rect 303396 5080 303402 5092
rect 562042 5080 562048 5092
rect 303396 5052 562048 5080
rect 303396 5040 303402 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 234706 5012 234712 5024
rect 7708 4984 234712 5012
rect 7708 4972 7714 4984
rect 234706 4972 234712 4984
rect 234764 4972 234770 5024
rect 246390 4972 246396 5024
rect 246448 5012 246454 5024
rect 263778 5012 263784 5024
rect 246448 4984 263784 5012
rect 246448 4972 246454 4984
rect 263778 4972 263784 4984
rect 263836 4972 263842 5024
rect 271230 4972 271236 5024
rect 271288 5012 271294 5024
rect 300762 5012 300768 5024
rect 271288 4984 300768 5012
rect 271288 4972 271294 4984
rect 300762 4972 300768 4984
rect 300820 4972 300826 5024
rect 302786 4972 302792 5024
rect 302844 5012 302850 5024
rect 565630 5012 565636 5024
rect 302844 4984 565636 5012
rect 302844 4972 302850 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 234890 4944 234896 4956
rect 2924 4916 234896 4944
rect 2924 4904 2930 4916
rect 234890 4904 234896 4916
rect 234948 4904 234954 4956
rect 242894 4904 242900 4956
rect 242952 4944 242958 4956
rect 263870 4944 263876 4956
rect 242952 4916 263876 4944
rect 242952 4904 242958 4916
rect 263870 4904 263876 4916
rect 263928 4904 263934 4956
rect 271506 4904 271512 4956
rect 271564 4944 271570 4956
rect 299658 4944 299664 4956
rect 271564 4916 299664 4944
rect 271564 4904 271570 4916
rect 299658 4904 299664 4916
rect 299716 4904 299722 4956
rect 303246 4904 303252 4956
rect 303304 4944 303310 4956
rect 569126 4944 569132 4956
rect 303304 4916 569132 4944
rect 303304 4904 303310 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 234798 4876 234804 4888
rect 1728 4848 234804 4876
rect 1728 4836 1734 4848
rect 234798 4836 234804 4848
rect 234856 4836 234862 4888
rect 239306 4836 239312 4888
rect 239364 4876 239370 4888
rect 264054 4876 264060 4888
rect 239364 4848 264060 4876
rect 239364 4836 239370 4848
rect 264054 4836 264060 4848
rect 264112 4836 264118 4888
rect 271598 4836 271604 4888
rect 271656 4876 271662 4888
rect 303154 4876 303160 4888
rect 271656 4848 303160 4876
rect 271656 4836 271662 4848
rect 303154 4836 303160 4848
rect 303212 4836 303218 4888
rect 572714 4876 572720 4888
rect 304460 4848 572720 4876
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 234982 4808 234988 4820
rect 624 4780 234988 4808
rect 624 4768 630 4780
rect 234982 4768 234988 4780
rect 235040 4768 235046 4820
rect 235902 4768 235908 4820
rect 235960 4808 235966 4820
rect 262582 4808 262588 4820
rect 235960 4780 262588 4808
rect 235960 4768 235966 4780
rect 262582 4768 262588 4780
rect 262640 4768 262646 4820
rect 271690 4768 271696 4820
rect 271748 4808 271754 4820
rect 304350 4808 304356 4820
rect 271748 4780 304356 4808
rect 271748 4768 271754 4780
rect 304350 4768 304356 4780
rect 304408 4768 304414 4820
rect 211062 4700 211068 4752
rect 211120 4740 211126 4752
rect 260190 4740 260196 4752
rect 211120 4712 260196 4740
rect 211120 4700 211126 4712
rect 260190 4700 260196 4712
rect 260248 4700 260254 4752
rect 269942 4700 269948 4752
rect 270000 4740 270006 4752
rect 285398 4740 285404 4752
rect 270000 4712 285404 4740
rect 270000 4700 270006 4712
rect 285398 4700 285404 4712
rect 285456 4700 285462 4752
rect 302694 4700 302700 4752
rect 302752 4740 302758 4752
rect 304460 4740 304488 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 304534 4768 304540 4820
rect 304592 4808 304598 4820
rect 576302 4808 576308 4820
rect 304592 4780 576308 4808
rect 304592 4768 304598 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 537202 4740 537208 4752
rect 302752 4712 304488 4740
rect 304552 4712 537208 4740
rect 302752 4700 302758 4712
rect 259546 4672 259552 4684
rect 219406 4644 259552 4672
rect 214466 4564 214472 4616
rect 214524 4604 214530 4616
rect 219406 4604 219434 4644
rect 259546 4632 259552 4644
rect 259604 4632 259610 4684
rect 268838 4632 268844 4684
rect 268896 4672 268902 4684
rect 283098 4672 283104 4684
rect 268896 4644 283104 4672
rect 268896 4632 268902 4644
rect 283098 4632 283104 4644
rect 283156 4632 283162 4684
rect 299198 4632 299204 4684
rect 299256 4672 299262 4684
rect 304552 4672 304580 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 299256 4644 304580 4672
rect 304629 4675 304687 4681
rect 299256 4632 299262 4644
rect 304629 4641 304641 4675
rect 304675 4672 304687 4675
rect 533706 4672 533712 4684
rect 304675 4644 533712 4672
rect 304675 4641 304687 4644
rect 304629 4635 304687 4641
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 214524 4576 219434 4604
rect 214524 4564 214530 4576
rect 228726 4564 228732 4616
rect 228784 4604 228790 4616
rect 262398 4604 262404 4616
rect 228784 4576 262404 4604
rect 228784 4564 228790 4576
rect 262398 4564 262404 4576
rect 262456 4564 262462 4616
rect 268654 4564 268660 4616
rect 268712 4604 268718 4616
rect 281902 4604 281908 4616
rect 268712 4576 281908 4604
rect 268712 4564 268718 4576
rect 281902 4564 281908 4576
rect 281960 4564 281966 4616
rect 299290 4564 299296 4616
rect 299348 4604 299354 4616
rect 530118 4604 530124 4616
rect 299348 4576 530124 4604
rect 299348 4564 299354 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 232222 4496 232228 4548
rect 232280 4536 232286 4548
rect 262766 4536 262772 4548
rect 232280 4508 262772 4536
rect 232280 4496 232286 4508
rect 262766 4496 262772 4508
rect 262824 4496 262830 4548
rect 268746 4496 268752 4548
rect 268804 4536 268810 4548
rect 278314 4536 278320 4548
rect 268804 4508 278320 4536
rect 268804 4496 268810 4508
rect 278314 4496 278320 4508
rect 278372 4496 278378 4548
rect 295978 4496 295984 4548
rect 296036 4536 296042 4548
rect 512454 4536 512460 4548
rect 296036 4508 512460 4536
rect 296036 4496 296042 4508
rect 512454 4496 512460 4508
rect 512512 4496 512518 4548
rect 298646 4428 298652 4480
rect 298704 4468 298710 4480
rect 304629 4471 304687 4477
rect 304629 4468 304641 4471
rect 298704 4440 304641 4468
rect 298704 4428 298710 4440
rect 304629 4437 304641 4440
rect 304675 4437 304687 4471
rect 304629 4431 304687 4437
rect 126974 4156 126980 4208
rect 127032 4196 127038 4208
rect 128262 4196 128268 4208
rect 127032 4168 128268 4196
rect 127032 4156 127038 4168
rect 128262 4156 128268 4168
rect 128320 4156 128326 4208
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 144822 4196 144828 4208
rect 143592 4168 144828 4196
rect 143592 4156 143598 4168
rect 144822 4156 144828 4168
rect 144880 4156 144886 4208
rect 151814 4156 151820 4208
rect 151872 4196 151878 4208
rect 153102 4196 153108 4208
rect 151872 4168 153108 4196
rect 151872 4156 151878 4168
rect 153102 4156 153108 4168
rect 153160 4156 153166 4208
rect 160094 4156 160100 4208
rect 160152 4196 160158 4208
rect 161382 4196 161388 4208
rect 160152 4168 161388 4196
rect 160152 4156 160158 4168
rect 161382 4156 161388 4168
rect 161440 4156 161446 4208
rect 168374 4156 168380 4208
rect 168432 4196 168438 4208
rect 169662 4196 169668 4208
rect 168432 4168 169668 4196
rect 168432 4156 168438 4168
rect 169662 4156 169668 4168
rect 169720 4156 169726 4208
rect 184934 4156 184940 4208
rect 184992 4196 184998 4208
rect 186222 4196 186228 4208
rect 184992 4168 186228 4196
rect 184992 4156 184998 4168
rect 186222 4156 186228 4168
rect 186280 4156 186286 4208
rect 209774 4156 209780 4208
rect 209832 4196 209838 4208
rect 210970 4196 210976 4208
rect 209832 4168 210976 4196
rect 209832 4156 209838 4168
rect 210970 4156 210976 4168
rect 211028 4156 211034 4208
rect 218054 4156 218060 4208
rect 218112 4196 218118 4208
rect 219342 4196 219348 4208
rect 218112 4168 219348 4196
rect 218112 4156 218118 4168
rect 219342 4156 219348 4168
rect 219400 4156 219406 4208
rect 226334 4156 226340 4208
rect 226392 4196 226398 4208
rect 227622 4196 227628 4208
rect 226392 4168 227628 4196
rect 226392 4156 226398 4168
rect 227622 4156 227628 4168
rect 227680 4156 227686 4208
rect 229649 4199 229707 4205
rect 229649 4165 229661 4199
rect 229695 4196 229707 4199
rect 237558 4196 237564 4208
rect 229695 4168 237564 4196
rect 229695 4165 229707 4168
rect 229649 4159 229707 4165
rect 237558 4156 237564 4168
rect 237616 4156 237622 4208
rect 297358 4156 297364 4208
rect 297416 4196 297422 4208
rect 298462 4196 298468 4208
rect 297416 4168 298468 4196
rect 297416 4156 297422 4168
rect 298462 4156 298468 4168
rect 298520 4156 298526 4208
rect 307754 4156 307760 4208
rect 307812 4196 307818 4208
rect 309042 4196 309048 4208
rect 307812 4168 309048 4196
rect 307812 4156 307818 4168
rect 309042 4156 309048 4168
rect 309100 4156 309106 4208
rect 316034 4156 316040 4208
rect 316092 4196 316098 4208
rect 317322 4196 317328 4208
rect 316092 4168 317328 4196
rect 316092 4156 316098 4168
rect 317322 4156 317328 4168
rect 317380 4156 317386 4208
rect 332686 4156 332692 4208
rect 332744 4196 332750 4208
rect 333882 4196 333888 4208
rect 332744 4168 333888 4196
rect 332744 4156 332750 4168
rect 333882 4156 333888 4168
rect 333940 4156 333946 4208
rect 349154 4156 349160 4208
rect 349212 4196 349218 4208
rect 350442 4196 350448 4208
rect 349212 4168 350448 4196
rect 349212 4156 349218 4168
rect 350442 4156 350448 4168
rect 350500 4156 350506 4208
rect 357526 4156 357532 4208
rect 357584 4196 357590 4208
rect 358722 4196 358728 4208
rect 357584 4168 358728 4196
rect 357584 4156 357590 4168
rect 358722 4156 358728 4168
rect 358780 4156 358786 4208
rect 373994 4156 374000 4208
rect 374052 4196 374058 4208
rect 375282 4196 375288 4208
rect 374052 4168 375288 4196
rect 374052 4156 374058 4168
rect 375282 4156 375288 4168
rect 375340 4156 375346 4208
rect 382274 4156 382280 4208
rect 382332 4196 382338 4208
rect 383562 4196 383568 4208
rect 382332 4168 383568 4196
rect 382332 4156 382338 4168
rect 383562 4156 383568 4168
rect 383620 4156 383626 4208
rect 398834 4156 398840 4208
rect 398892 4196 398898 4208
rect 400122 4196 400128 4208
rect 398892 4168 400128 4196
rect 398892 4156 398898 4168
rect 400122 4156 400128 4168
rect 400180 4156 400186 4208
rect 423766 4156 423772 4208
rect 423824 4196 423830 4208
rect 424962 4196 424968 4208
rect 423824 4168 424968 4196
rect 423824 4156 423830 4168
rect 424962 4156 424968 4168
rect 425020 4156 425026 4208
rect 45370 4088 45376 4140
rect 45428 4128 45434 4140
rect 46198 4128 46204 4140
rect 45428 4100 46204 4128
rect 45428 4088 45434 4100
rect 46198 4088 46204 4100
rect 46256 4088 46262 4140
rect 85666 4088 85672 4140
rect 85724 4128 85730 4140
rect 244550 4128 244556 4140
rect 85724 4100 244556 4128
rect 85724 4088 85730 4100
rect 244550 4088 244556 4100
rect 244608 4088 244614 4140
rect 267366 4088 267372 4140
rect 267424 4128 267430 4140
rect 268838 4128 268844 4140
rect 267424 4100 268844 4128
rect 267424 4088 267430 4100
rect 268838 4088 268844 4100
rect 268896 4088 268902 4140
rect 287422 4088 287428 4140
rect 287480 4128 287486 4140
rect 443822 4128 443828 4140
rect 287480 4100 443828 4128
rect 287480 4088 287486 4100
rect 443822 4088 443828 4100
rect 443880 4088 443886 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 568022 4128 568028 4140
rect 566516 4100 568028 4128
rect 566516 4088 566522 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 18598 4060 18604 4072
rect 10008 4032 18604 4060
rect 10008 4020 10014 4032
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 244918 4060 244924 4072
rect 82136 4032 244924 4060
rect 82136 4020 82142 4032
rect 244918 4020 244924 4032
rect 244976 4020 244982 4072
rect 267458 4020 267464 4072
rect 267516 4060 267522 4072
rect 267642 4060 267648 4072
rect 267516 4032 267648 4060
rect 267516 4020 267522 4032
rect 267642 4020 267648 4032
rect 267700 4020 267706 4072
rect 289538 4020 289544 4072
rect 289596 4060 289602 4072
rect 447410 4060 447416 4072
rect 289596 4032 447416 4060
rect 289596 4020 289602 4032
rect 447410 4020 447416 4032
rect 447468 4020 447474 4072
rect 78490 3952 78496 4004
rect 78548 3992 78554 4004
rect 244458 3992 244464 4004
rect 78548 3964 244464 3992
rect 78548 3952 78554 3964
rect 244458 3952 244464 3964
rect 244516 3952 244522 4004
rect 289630 3952 289636 4004
rect 289688 3992 289694 4004
rect 450906 3992 450912 4004
rect 289688 3964 450912 3992
rect 289688 3952 289694 3964
rect 450906 3952 450912 3964
rect 450964 3952 450970 4004
rect 60826 3884 60832 3936
rect 60884 3924 60890 3936
rect 62022 3924 62028 3936
rect 60884 3896 62028 3924
rect 60884 3884 60890 3896
rect 62022 3884 62028 3896
rect 62080 3884 62086 3936
rect 74994 3884 75000 3936
rect 75052 3924 75058 3936
rect 243630 3924 243636 3936
rect 75052 3896 243636 3924
rect 75052 3884 75058 3896
rect 243630 3884 243636 3896
rect 243688 3884 243694 3936
rect 289722 3884 289728 3936
rect 289780 3924 289786 3936
rect 454494 3924 454500 3936
rect 289780 3896 454500 3924
rect 289780 3884 289786 3896
rect 454494 3884 454500 3896
rect 454552 3884 454558 3936
rect 576118 3884 576124 3936
rect 576176 3924 576182 3936
rect 578602 3924 578608 3936
rect 576176 3896 578608 3924
rect 576176 3884 576182 3896
rect 578602 3884 578608 3896
rect 578660 3884 578666 3936
rect 46658 3816 46664 3868
rect 46716 3856 46722 3868
rect 240778 3856 240784 3868
rect 46716 3828 240784 3856
rect 46716 3816 46722 3828
rect 240778 3816 240784 3828
rect 240836 3816 240842 3868
rect 260561 3859 260619 3865
rect 260561 3825 260573 3859
rect 260607 3856 260619 3859
rect 265434 3856 265440 3868
rect 260607 3828 265440 3856
rect 260607 3825 260619 3828
rect 260561 3819 260619 3825
rect 265434 3816 265440 3828
rect 265492 3816 265498 3868
rect 290826 3816 290832 3868
rect 290884 3856 290890 3868
rect 458082 3856 458088 3868
rect 290884 3828 458088 3856
rect 290884 3816 290890 3828
rect 458082 3816 458088 3828
rect 458140 3816 458146 3868
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 239030 3788 239036 3800
rect 43128 3760 239036 3788
rect 43128 3748 43134 3760
rect 239030 3748 239036 3760
rect 239088 3748 239094 3800
rect 262858 3788 262864 3800
rect 258046 3760 262864 3788
rect 28902 3680 28908 3732
rect 28960 3720 28966 3732
rect 35158 3720 35164 3732
rect 28960 3692 35164 3720
rect 28960 3680 28966 3692
rect 35158 3680 35164 3692
rect 35216 3680 35222 3732
rect 39574 3680 39580 3732
rect 39632 3720 39638 3732
rect 233789 3723 233847 3729
rect 233789 3720 233801 3723
rect 39632 3692 233801 3720
rect 39632 3680 39638 3692
rect 233789 3689 233801 3692
rect 233835 3689 233847 3723
rect 233789 3683 233847 3689
rect 233881 3723 233939 3729
rect 233881 3689 233893 3723
rect 233927 3720 233939 3723
rect 238846 3720 238852 3732
rect 233927 3692 238852 3720
rect 233927 3689 233939 3692
rect 233881 3683 233939 3689
rect 238846 3680 238852 3692
rect 238904 3680 238910 3732
rect 257062 3680 257068 3732
rect 257120 3720 257126 3732
rect 258046 3720 258074 3760
rect 262858 3748 262864 3760
rect 262916 3748 262922 3800
rect 263045 3791 263103 3797
rect 263045 3757 263057 3791
rect 263091 3788 263103 3791
rect 265618 3788 265624 3800
rect 263091 3760 265624 3788
rect 263091 3757 263103 3760
rect 263045 3751 263103 3757
rect 265618 3748 265624 3760
rect 265676 3748 265682 3800
rect 291102 3748 291108 3800
rect 291160 3788 291166 3800
rect 461578 3788 461584 3800
rect 291160 3760 461584 3788
rect 291160 3748 291166 3760
rect 461578 3748 461584 3760
rect 461636 3748 461642 3800
rect 257120 3692 258074 3720
rect 257120 3680 257126 3692
rect 259454 3680 259460 3732
rect 259512 3720 259518 3732
rect 265342 3720 265348 3732
rect 259512 3692 265348 3720
rect 259512 3680 259518 3692
rect 265342 3680 265348 3692
rect 265400 3680 265406 3732
rect 267550 3680 267556 3732
rect 267608 3720 267614 3732
rect 273622 3720 273628 3732
rect 267608 3692 273628 3720
rect 267608 3680 267614 3692
rect 273622 3680 273628 3692
rect 273680 3680 273686 3732
rect 290918 3680 290924 3732
rect 290976 3720 290982 3732
rect 465166 3720 465172 3732
rect 290976 3692 465172 3720
rect 290976 3680 290982 3692
rect 465166 3680 465172 3692
rect 465224 3680 465230 3732
rect 23014 3612 23020 3664
rect 23072 3652 23078 3664
rect 29638 3652 29644 3664
rect 23072 3624 29644 3652
rect 23072 3612 23078 3624
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 32398 3612 32404 3664
rect 32456 3652 32462 3664
rect 32456 3624 35894 3652
rect 32456 3612 32462 3624
rect 10318 3584 10324 3596
rect 6886 3556 10324 3584
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6886 3516 6914 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 28258 3584 28264 3596
rect 11204 3556 28264 3584
rect 11204 3544 11210 3556
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34422 3584 34428 3596
rect 33652 3556 34428 3584
rect 33652 3544 33658 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35866 3584 35894 3624
rect 35986 3612 35992 3664
rect 36044 3652 36050 3664
rect 238938 3652 238944 3664
rect 36044 3624 238944 3652
rect 36044 3612 36050 3624
rect 238938 3612 238944 3624
rect 238996 3612 239002 3664
rect 262950 3612 262956 3664
rect 263008 3652 263014 3664
rect 266538 3652 266544 3664
rect 263008 3624 266544 3652
rect 263008 3612 263014 3624
rect 266538 3612 266544 3624
rect 266596 3612 266602 3664
rect 291010 3612 291016 3664
rect 291068 3652 291074 3664
rect 468662 3652 468668 3664
rect 291068 3624 468668 3652
rect 291068 3612 291074 3624
rect 468662 3612 468668 3624
rect 468720 3612 468726 3664
rect 233881 3587 233939 3593
rect 233881 3584 233893 3587
rect 35866 3556 233893 3584
rect 233881 3553 233893 3556
rect 233927 3553 233939 3587
rect 233881 3547 233939 3553
rect 233973 3587 234031 3593
rect 233973 3553 233985 3587
rect 234019 3584 234031 3587
rect 238018 3584 238024 3596
rect 234019 3556 238024 3584
rect 234019 3553 234031 3556
rect 233973 3547 234031 3553
rect 238018 3544 238024 3556
rect 238076 3544 238082 3596
rect 255866 3544 255872 3596
rect 255924 3584 255930 3596
rect 263045 3587 263103 3593
rect 263045 3584 263057 3587
rect 255924 3556 263057 3584
rect 255924 3544 255930 3556
rect 263045 3553 263057 3556
rect 263091 3553 263103 3587
rect 263045 3547 263103 3553
rect 264146 3544 264152 3596
rect 264204 3584 264210 3596
rect 266906 3584 266912 3596
rect 264204 3556 266912 3584
rect 264204 3544 264210 3556
rect 266906 3544 266912 3556
rect 266964 3544 266970 3596
rect 292482 3544 292488 3596
rect 292540 3584 292546 3596
rect 472250 3584 472256 3596
rect 292540 3556 472256 3584
rect 292540 3544 292546 3556
rect 472250 3544 472256 3556
rect 472308 3544 472314 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 527818 3584 527824 3596
rect 525116 3556 527824 3584
rect 525116 3544 525122 3556
rect 527818 3544 527824 3556
rect 527876 3544 527882 3596
rect 5316 3488 6914 3516
rect 5316 3476 5322 3488
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 25372 3488 229784 3516
rect 25372 3476 25378 3488
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 229649 3451 229707 3457
rect 229649 3448 229661 3451
rect 24268 3420 229661 3448
rect 24268 3408 24274 3420
rect 229649 3417 229661 3420
rect 229695 3417 229707 3451
rect 229756 3448 229784 3488
rect 229830 3476 229836 3528
rect 229888 3516 229894 3528
rect 230382 3516 230388 3528
rect 229888 3488 230388 3516
rect 229888 3476 229894 3488
rect 230382 3476 230388 3488
rect 230440 3476 230446 3528
rect 231026 3476 231032 3528
rect 231084 3516 231090 3528
rect 231762 3516 231768 3528
rect 231084 3488 231768 3516
rect 231084 3476 231090 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 233418 3476 233424 3528
rect 233476 3516 233482 3528
rect 234522 3516 234528 3528
rect 233476 3488 234528 3516
rect 233476 3476 233482 3488
rect 234522 3476 234528 3488
rect 234580 3476 234586 3528
rect 234614 3476 234620 3528
rect 234672 3516 234678 3528
rect 235810 3516 235816 3528
rect 234672 3488 235816 3516
rect 234672 3476 234678 3488
rect 235810 3476 235816 3488
rect 235868 3476 235874 3528
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241422 3516 241428 3528
rect 240560 3488 241428 3516
rect 240560 3476 240566 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 241698 3476 241704 3528
rect 241756 3516 241762 3528
rect 242802 3516 242808 3528
rect 241756 3488 242808 3516
rect 241756 3476 241762 3488
rect 242802 3476 242808 3488
rect 242860 3476 242866 3528
rect 248782 3476 248788 3528
rect 248840 3516 248846 3528
rect 249702 3516 249708 3528
rect 248840 3488 249708 3516
rect 248840 3476 248846 3488
rect 249702 3476 249708 3488
rect 249760 3476 249766 3528
rect 254670 3476 254676 3528
rect 254728 3516 254734 3528
rect 260561 3519 260619 3525
rect 260561 3516 260573 3519
rect 254728 3488 260573 3516
rect 254728 3476 254734 3488
rect 260561 3485 260573 3488
rect 260607 3485 260619 3519
rect 260561 3479 260619 3485
rect 260650 3476 260656 3528
rect 260708 3516 260714 3528
rect 265066 3516 265072 3528
rect 260708 3488 265072 3516
rect 260708 3476 260714 3488
rect 265066 3476 265072 3488
rect 265124 3476 265130 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267090 3516 267096 3528
rect 266596 3488 267096 3516
rect 266596 3476 266602 3488
rect 267090 3476 267096 3488
rect 267148 3476 267154 3528
rect 268378 3476 268384 3528
rect 268436 3516 268442 3528
rect 272426 3516 272432 3528
rect 268436 3488 272432 3516
rect 268436 3476 268442 3488
rect 272426 3476 272432 3488
rect 272484 3476 272490 3528
rect 292298 3476 292304 3528
rect 292356 3516 292362 3528
rect 292356 3488 473216 3516
rect 292356 3476 292362 3488
rect 233697 3451 233755 3457
rect 233697 3448 233709 3451
rect 229756 3420 233709 3448
rect 229649 3411 229707 3417
rect 233697 3417 233709 3420
rect 233743 3417 233755 3451
rect 233697 3411 233755 3417
rect 233789 3451 233847 3457
rect 233789 3417 233801 3451
rect 233835 3448 233847 3451
rect 239398 3448 239404 3460
rect 233835 3420 239404 3448
rect 233835 3417 233847 3420
rect 233789 3411 233847 3417
rect 239398 3408 239404 3420
rect 239456 3408 239462 3460
rect 251174 3408 251180 3460
rect 251232 3448 251238 3460
rect 265250 3448 265256 3460
rect 251232 3420 265256 3448
rect 251232 3408 251238 3420
rect 265250 3408 265256 3420
rect 265308 3408 265314 3460
rect 265342 3408 265348 3460
rect 265400 3448 265406 3460
rect 266630 3448 266636 3460
rect 265400 3420 266636 3448
rect 265400 3408 265406 3420
rect 266630 3408 266636 3420
rect 266688 3408 266694 3460
rect 267274 3408 267280 3460
rect 267332 3448 267338 3460
rect 270034 3448 270040 3460
rect 267332 3420 270040 3448
rect 267332 3408 267338 3420
rect 270034 3408 270040 3420
rect 270092 3408 270098 3460
rect 292390 3408 292396 3460
rect 292448 3448 292454 3460
rect 473188 3448 473216 3488
rect 473354 3476 473360 3528
rect 473412 3516 473418 3528
rect 474550 3516 474556 3528
rect 473412 3488 474556 3516
rect 473412 3476 473418 3488
rect 474550 3476 474556 3488
rect 474608 3476 474614 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 491110 3516 491116 3528
rect 489972 3488 491116 3516
rect 489972 3476 489978 3488
rect 491110 3476 491116 3488
rect 491168 3476 491174 3528
rect 522298 3476 522304 3528
rect 522356 3516 522362 3528
rect 524230 3516 524236 3528
rect 522356 3488 524236 3516
rect 522356 3476 522362 3488
rect 524230 3476 524236 3488
rect 524288 3476 524294 3528
rect 533338 3476 533344 3528
rect 533396 3516 533402 3528
rect 534902 3516 534908 3528
rect 533396 3488 534908 3516
rect 533396 3476 533402 3488
rect 534902 3476 534908 3488
rect 534960 3476 534966 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 557350 3516 557356 3528
rect 556212 3488 557356 3516
rect 556212 3476 556218 3488
rect 557350 3476 557356 3488
rect 557408 3476 557414 3528
rect 475746 3448 475752 3460
rect 292448 3420 470594 3448
rect 473188 3420 475752 3448
rect 292448 3408 292454 3420
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 43438 3380 43444 3392
rect 41932 3352 43444 3380
rect 41932 3340 41938 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45462 3380 45468 3392
rect 44324 3352 45468 3380
rect 44324 3340 44330 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 48958 3340 48964 3392
rect 49016 3380 49022 3392
rect 49602 3380 49608 3392
rect 49016 3352 49608 3380
rect 49016 3340 49022 3352
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 50982 3380 50988 3392
rect 50212 3352 50988 3380
rect 50212 3340 50218 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 52546 3340 52552 3392
rect 52604 3380 52610 3392
rect 53650 3380 53656 3392
rect 52604 3352 53656 3380
rect 52604 3340 52610 3352
rect 53650 3340 53656 3352
rect 53708 3340 53714 3392
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 56502 3380 56508 3392
rect 56100 3352 56508 3380
rect 56100 3340 56106 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 57882 3380 57888 3392
rect 57296 3352 57888 3380
rect 57296 3340 57302 3352
rect 57882 3340 57888 3352
rect 57940 3340 57946 3392
rect 64322 3340 64328 3392
rect 64380 3380 64386 3392
rect 64782 3380 64788 3392
rect 64380 3352 64788 3380
rect 64380 3340 64386 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 67542 3380 67548 3392
rect 66772 3352 67548 3380
rect 66772 3340 66778 3352
rect 67542 3340 67548 3352
rect 67600 3340 67606 3392
rect 67910 3340 67916 3392
rect 67968 3380 67974 3392
rect 68922 3380 68928 3392
rect 67968 3352 68928 3380
rect 67968 3340 67974 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 73798 3340 73804 3392
rect 73856 3380 73862 3392
rect 74442 3380 74448 3392
rect 73856 3352 74448 3380
rect 73856 3340 73862 3352
rect 74442 3340 74448 3352
rect 74500 3340 74506 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 78582 3380 78588 3392
rect 77444 3352 78588 3380
rect 77444 3340 77450 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 85482 3380 85488 3392
rect 84528 3352 85488 3380
rect 84528 3340 84534 3352
rect 85482 3340 85488 3352
rect 85540 3340 85546 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 92382 3380 92388 3392
rect 91612 3352 92388 3380
rect 91612 3340 91618 3352
rect 92382 3340 92388 3352
rect 92440 3340 92446 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 95234 3380 95240 3392
rect 94004 3352 95240 3380
rect 94004 3340 94010 3352
rect 95234 3340 95240 3352
rect 95292 3340 95298 3392
rect 97442 3340 97448 3392
rect 97500 3380 97506 3392
rect 97902 3380 97908 3392
rect 97500 3352 97908 3380
rect 97500 3340 97506 3352
rect 97902 3340 97908 3352
rect 97960 3340 97966 3392
rect 98638 3340 98644 3392
rect 98696 3380 98702 3392
rect 99282 3380 99288 3392
rect 98696 3352 99288 3380
rect 98696 3340 98702 3352
rect 99282 3340 99288 3352
rect 99340 3340 99346 3392
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 102042 3380 102048 3392
rect 101088 3352 102048 3380
rect 101088 3340 101094 3352
rect 102042 3340 102048 3352
rect 102100 3340 102106 3392
rect 245010 3380 245016 3392
rect 102152 3352 245016 3380
rect 27706 3272 27712 3324
rect 27764 3312 27770 3324
rect 33778 3312 33784 3324
rect 27764 3284 33784 3312
rect 27764 3272 27770 3284
rect 33778 3272 33784 3284
rect 33836 3272 33842 3324
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 102152 3244 102180 3352
rect 245010 3340 245016 3352
rect 245068 3340 245074 3392
rect 287514 3340 287520 3392
rect 287572 3380 287578 3392
rect 440326 3380 440332 3392
rect 287572 3352 440332 3380
rect 287572 3340 287578 3352
rect 440326 3340 440332 3352
rect 440384 3340 440390 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 470566 3380 470594 3420
rect 475746 3408 475752 3420
rect 475804 3408 475810 3460
rect 514754 3408 514760 3460
rect 514812 3448 514818 3460
rect 515950 3448 515956 3460
rect 514812 3420 515956 3448
rect 514812 3408 514818 3420
rect 515950 3408 515956 3420
rect 516008 3408 516014 3460
rect 479334 3380 479340 3392
rect 470566 3352 479340 3380
rect 479334 3340 479340 3352
rect 479392 3340 479398 3392
rect 102229 3315 102287 3321
rect 102229 3281 102241 3315
rect 102275 3312 102287 3315
rect 245838 3312 245844 3324
rect 102275 3284 245844 3312
rect 102275 3281 102287 3284
rect 102229 3275 102287 3281
rect 245838 3272 245844 3284
rect 245896 3272 245902 3324
rect 269022 3272 269028 3324
rect 269080 3312 269086 3324
rect 277118 3312 277124 3324
rect 269080 3284 277124 3312
rect 269080 3272 269086 3284
rect 277118 3272 277124 3284
rect 277176 3272 277182 3324
rect 288158 3272 288164 3324
rect 288216 3312 288222 3324
rect 436738 3312 436744 3324
rect 288216 3284 436744 3312
rect 288216 3272 288222 3284
rect 436738 3272 436744 3284
rect 436796 3272 436802 3324
rect 246298 3244 246304 3256
rect 89220 3216 102180 3244
rect 102244 3216 246304 3244
rect 89220 3204 89226 3216
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 27522 3176 27528 3188
rect 26568 3148 27528 3176
rect 26568 3136 26574 3148
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 92750 3136 92756 3188
rect 92808 3176 92814 3188
rect 102137 3179 102195 3185
rect 102137 3176 102149 3179
rect 92808 3148 102149 3176
rect 92808 3136 92814 3148
rect 102137 3145 102149 3148
rect 102183 3145 102195 3179
rect 102137 3139 102195 3145
rect 31294 3068 31300 3120
rect 31352 3108 31358 3120
rect 36538 3108 36544 3120
rect 31352 3080 36544 3108
rect 31352 3068 31358 3080
rect 36538 3068 36544 3080
rect 36596 3068 36602 3120
rect 96246 3068 96252 3120
rect 96304 3108 96310 3120
rect 102244 3108 102272 3216
rect 246298 3204 246304 3216
rect 246356 3204 246362 3256
rect 261754 3204 261760 3256
rect 261812 3244 261818 3256
rect 265526 3244 265532 3256
rect 261812 3216 265532 3244
rect 261812 3204 261818 3216
rect 265526 3204 265532 3216
rect 265584 3204 265590 3256
rect 286134 3204 286140 3256
rect 286192 3244 286198 3256
rect 433242 3244 433248 3256
rect 286192 3216 433248 3244
rect 286192 3204 286198 3216
rect 433242 3204 433248 3216
rect 433300 3204 433306 3256
rect 105722 3136 105728 3188
rect 105780 3176 105786 3188
rect 106182 3176 106188 3188
rect 105780 3148 106188 3176
rect 105780 3136 105786 3148
rect 106182 3136 106188 3148
rect 106240 3136 106246 3188
rect 108114 3136 108120 3188
rect 108172 3176 108178 3188
rect 108942 3176 108948 3188
rect 108172 3148 108948 3176
rect 108172 3136 108178 3148
rect 108942 3136 108948 3148
rect 109000 3136 109006 3188
rect 109310 3136 109316 3188
rect 109368 3176 109374 3188
rect 110322 3176 110328 3188
rect 109368 3148 110328 3176
rect 109368 3136 109374 3148
rect 110322 3136 110328 3148
rect 110380 3136 110386 3188
rect 110417 3179 110475 3185
rect 110417 3145 110429 3179
rect 110463 3176 110475 3179
rect 246206 3176 246212 3188
rect 110463 3148 246212 3176
rect 110463 3145 110475 3148
rect 110417 3139 110475 3145
rect 246206 3136 246212 3148
rect 246264 3136 246270 3188
rect 268930 3136 268936 3188
rect 268988 3176 268994 3188
rect 276014 3176 276020 3188
rect 268988 3148 276020 3176
rect 268988 3136 268994 3148
rect 276014 3136 276020 3148
rect 276072 3136 276078 3188
rect 286778 3136 286784 3188
rect 286836 3176 286842 3188
rect 429654 3176 429660 3188
rect 286836 3148 429660 3176
rect 286836 3136 286842 3148
rect 429654 3136 429660 3148
rect 429712 3136 429718 3188
rect 96304 3080 102272 3108
rect 96304 3068 96310 3080
rect 103330 3068 103336 3120
rect 103388 3108 103394 3120
rect 247494 3108 247500 3120
rect 103388 3080 247500 3108
rect 103388 3068 103394 3080
rect 247494 3068 247500 3080
rect 247552 3068 247558 3120
rect 286226 3068 286232 3120
rect 286284 3108 286290 3120
rect 426158 3108 426164 3120
rect 286284 3080 426164 3108
rect 286284 3068 286290 3080
rect 426158 3068 426164 3080
rect 426216 3068 426222 3120
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 21358 3040 21364 3052
rect 19484 3012 21364 3040
rect 19484 3000 19490 3012
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 99834 3000 99840 3052
rect 99892 3040 99898 3052
rect 110417 3043 110475 3049
rect 110417 3040 110429 3043
rect 99892 3012 110429 3040
rect 99892 3000 99898 3012
rect 110417 3009 110429 3012
rect 110463 3009 110475 3043
rect 110417 3003 110475 3009
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 114462 3040 114468 3052
rect 114060 3012 114468 3040
rect 114060 3000 114066 3012
rect 114462 3000 114468 3012
rect 114520 3000 114526 3052
rect 115198 3000 115204 3052
rect 115256 3040 115262 3052
rect 115842 3040 115848 3052
rect 115256 3012 115848 3040
rect 115256 3000 115262 3012
rect 115842 3000 115848 3012
rect 115900 3000 115906 3052
rect 116394 3000 116400 3052
rect 116452 3040 116458 3052
rect 117222 3040 117228 3052
rect 116452 3012 117228 3040
rect 116452 3000 116458 3012
rect 117222 3000 117228 3012
rect 117280 3000 117286 3052
rect 118786 3000 118792 3052
rect 118844 3040 118850 3052
rect 119890 3040 119896 3052
rect 118844 3012 119896 3040
rect 118844 3000 118850 3012
rect 119890 3000 119896 3012
rect 119948 3000 119954 3052
rect 119985 3043 120043 3049
rect 119985 3009 119997 3043
rect 120031 3040 120043 3043
rect 247678 3040 247684 3052
rect 120031 3012 247684 3040
rect 120031 3009 120043 3012
rect 119985 3003 120043 3009
rect 247678 3000 247684 3012
rect 247736 3000 247742 3052
rect 284846 3000 284852 3052
rect 284904 3040 284910 3052
rect 422570 3040 422576 3052
rect 284904 3012 422576 3040
rect 284904 3000 284910 3012
rect 422570 3000 422576 3012
rect 422628 3000 422634 3052
rect 529198 3000 529204 3052
rect 529256 3040 529262 3052
rect 531314 3040 531320 3052
rect 529256 3012 531320 3040
rect 529256 3000 529262 3012
rect 531314 3000 531320 3012
rect 531372 3000 531378 3052
rect 59630 2932 59636 2984
rect 59688 2972 59694 2984
rect 60642 2972 60648 2984
rect 59688 2944 60648 2972
rect 59688 2932 59694 2944
rect 60642 2932 60648 2944
rect 60700 2932 60706 2984
rect 102226 2932 102232 2984
rect 102284 2972 102290 2984
rect 103422 2972 103428 2984
rect 102284 2944 103428 2972
rect 102284 2932 102290 2944
rect 103422 2932 103428 2944
rect 103480 2932 103486 2984
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 247218 2972 247224 2984
rect 110564 2944 247224 2972
rect 110564 2932 110570 2944
rect 247218 2932 247224 2944
rect 247276 2932 247282 2984
rect 258258 2932 258264 2984
rect 258316 2972 258322 2984
rect 265158 2972 265164 2984
rect 258316 2944 265164 2972
rect 258316 2932 258322 2944
rect 265158 2932 265164 2944
rect 265216 2932 265222 2984
rect 284754 2932 284760 2984
rect 284812 2972 284818 2984
rect 415397 2975 415455 2981
rect 415397 2972 415409 2975
rect 284812 2944 415409 2972
rect 284812 2932 284818 2944
rect 415397 2941 415409 2944
rect 415443 2941 415455 2975
rect 415397 2935 415455 2941
rect 415486 2932 415492 2984
rect 415544 2972 415550 2984
rect 416682 2972 416688 2984
rect 415544 2944 416688 2972
rect 415544 2932 415550 2944
rect 416682 2932 416688 2944
rect 416740 2932 416746 2984
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 22738 2904 22744 2916
rect 18288 2876 22744 2904
rect 18288 2864 18294 2876
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 106918 2864 106924 2916
rect 106976 2904 106982 2916
rect 119985 2907 120043 2913
rect 119985 2904 119997 2907
rect 106976 2876 119997 2904
rect 106976 2864 106982 2876
rect 119985 2873 119997 2876
rect 120031 2873 120043 2907
rect 122193 2907 122251 2913
rect 122193 2904 122205 2907
rect 119985 2867 120043 2873
rect 120092 2876 122205 2904
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 120092 2836 120120 2876
rect 122193 2873 122205 2876
rect 122239 2873 122251 2907
rect 122193 2867 122251 2873
rect 122282 2864 122288 2916
rect 122340 2904 122346 2916
rect 122742 2904 122748 2916
rect 122340 2876 122748 2904
rect 122340 2864 122346 2876
rect 122742 2864 122748 2876
rect 122800 2864 122806 2916
rect 123478 2864 123484 2916
rect 123536 2904 123542 2916
rect 124122 2904 124128 2916
rect 123536 2876 124128 2904
rect 123536 2864 123542 2876
rect 124122 2864 124128 2876
rect 124180 2864 124186 2916
rect 124674 2864 124680 2916
rect 124732 2904 124738 2916
rect 125502 2904 125508 2916
rect 124732 2876 125508 2904
rect 124732 2864 124738 2876
rect 125502 2864 125508 2876
rect 125560 2864 125566 2916
rect 125870 2864 125876 2916
rect 125928 2904 125934 2916
rect 126882 2904 126888 2916
rect 125928 2876 126888 2904
rect 125928 2864 125934 2876
rect 126882 2864 126888 2876
rect 126940 2864 126946 2916
rect 249058 2904 249064 2916
rect 127084 2876 249064 2904
rect 117648 2808 120120 2836
rect 117648 2796 117654 2808
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 126977 2839 127035 2845
rect 126977 2836 126989 2839
rect 121144 2808 122052 2836
rect 121144 2796 121150 2808
rect 122024 2700 122052 2808
rect 122300 2808 126989 2836
rect 122300 2700 122328 2808
rect 126977 2805 126989 2808
rect 127023 2805 127035 2839
rect 126977 2799 127035 2805
rect 122377 2771 122435 2777
rect 122377 2737 122389 2771
rect 122423 2768 122435 2771
rect 127084 2768 127112 2876
rect 249058 2864 249064 2876
rect 249116 2864 249122 2916
rect 285490 2864 285496 2916
rect 285548 2904 285554 2916
rect 415581 2907 415639 2913
rect 285548 2876 415532 2904
rect 285548 2864 285554 2876
rect 415504 2848 415532 2876
rect 415581 2873 415593 2907
rect 415627 2904 415639 2907
rect 418982 2904 418988 2916
rect 415627 2876 418988 2904
rect 415627 2873 415639 2876
rect 415581 2867 415639 2873
rect 418982 2864 418988 2876
rect 419040 2864 419046 2916
rect 127161 2839 127219 2845
rect 127161 2805 127173 2839
rect 127207 2836 127219 2839
rect 249150 2836 249156 2848
rect 127207 2808 249156 2836
rect 127207 2805 127219 2808
rect 127161 2799 127219 2805
rect 249150 2796 249156 2808
rect 249208 2796 249214 2848
rect 285306 2796 285312 2848
rect 285364 2836 285370 2848
rect 285364 2808 407068 2836
rect 285364 2796 285370 2808
rect 122423 2740 127112 2768
rect 407040 2768 407068 2808
rect 407114 2796 407120 2848
rect 407172 2836 407178 2848
rect 408402 2836 408408 2848
rect 407172 2808 408408 2836
rect 407172 2796 407178 2808
rect 408402 2796 408408 2808
rect 408460 2796 408466 2848
rect 411898 2836 411904 2848
rect 408512 2808 411904 2836
rect 408512 2768 408540 2808
rect 411898 2796 411904 2808
rect 411956 2796 411962 2848
rect 415486 2796 415492 2848
rect 415544 2796 415550 2848
rect 407040 2740 408540 2768
rect 122423 2737 122435 2740
rect 122377 2731 122435 2737
rect 122024 2672 122328 2700
<< via1 >>
rect 285588 700952 285640 701004
rect 413652 700952 413704 701004
rect 286968 700884 287020 700936
rect 429844 700884 429896 700936
rect 288348 700816 288400 700868
rect 446128 700816 446180 700868
rect 291108 700748 291160 700800
rect 462320 700748 462372 700800
rect 292488 700680 292540 700732
rect 478512 700680 478564 700732
rect 295248 700612 295300 700664
rect 494796 700612 494848 700664
rect 296628 700544 296680 700596
rect 510988 700544 511040 700596
rect 299388 700476 299440 700528
rect 527180 700476 527232 700528
rect 300768 700408 300820 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 235172 700340 235224 700392
rect 235908 700340 235960 700392
rect 269028 700340 269080 700392
rect 283840 700340 283892 700392
rect 302148 700340 302200 700392
rect 559656 700340 559708 700392
rect 271788 700272 271840 700324
rect 300124 700272 300176 700324
rect 304908 700272 304960 700324
rect 575848 700272 575900 700324
rect 282828 700204 282880 700256
rect 397460 700204 397512 700256
rect 56784 700136 56836 700188
rect 57888 700136 57940 700188
rect 186504 700136 186556 700188
rect 187608 700136 187660 700188
rect 281448 700136 281500 700188
rect 381176 700136 381228 700188
rect 251456 700068 251508 700120
rect 252468 700068 252520 700120
rect 278688 700068 278740 700120
rect 364984 700068 365036 700120
rect 277308 700000 277360 700052
rect 348792 700000 348844 700052
rect 275928 699932 275980 699984
rect 332508 699932 332560 699984
rect 273168 699864 273220 699916
rect 316316 699864 316368 699916
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 121644 699660 121696 699712
rect 122748 699660 122800 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 266360 699660 266412 699712
rect 267648 699660 267700 699712
rect 3424 696940 3476 696992
rect 184204 696940 184256 696992
rect 307024 696940 307076 696992
rect 580172 696940 580224 696992
rect 307116 683136 307168 683188
rect 580172 683136 580224 683188
rect 307208 670692 307260 670744
rect 580172 670692 580224 670744
rect 3332 644444 3384 644496
rect 195244 644444 195296 644496
rect 307300 643084 307352 643136
rect 580172 643084 580224 643136
rect 309784 630640 309836 630692
rect 579988 630640 580040 630692
rect 2780 619080 2832 619132
rect 4804 619080 4856 619132
rect 2964 592016 3016 592068
rect 198004 592016 198056 592068
rect 307392 590656 307444 590708
rect 580172 590656 580224 590708
rect 307484 576852 307536 576904
rect 579988 576852 580040 576904
rect 2872 539588 2924 539640
rect 220084 539588 220136 539640
rect 307576 536800 307628 536852
rect 580172 536800 580224 536852
rect 307668 524424 307720 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 10324 514768 10376 514820
rect 306932 484372 306984 484424
rect 580172 484372 580224 484424
rect 306840 470568 306892 470620
rect 579988 470568 580040 470620
rect 306748 430584 306800 430636
rect 580080 430584 580132 430636
rect 312544 418140 312596 418192
rect 580080 418140 580132 418192
rect 171048 411204 171100 411256
rect 255320 411204 255372 411256
rect 154488 411136 154540 411188
rect 253112 411136 253164 411188
rect 137928 411068 137980 411120
rect 251180 411068 251232 411120
rect 122748 411000 122800 411052
rect 249156 411000 249208 411052
rect 106188 410932 106240 410984
rect 247224 410932 247276 410984
rect 89628 410864 89680 410916
rect 245292 410864 245344 410916
rect 73068 410796 73120 410848
rect 243360 410796 243412 410848
rect 3516 410771 3568 410780
rect 3516 410737 3525 410771
rect 3525 410737 3559 410771
rect 3559 410737 3568 410771
rect 3516 410728 3568 410737
rect 57888 410728 57940 410780
rect 241520 410728 241572 410780
rect 41328 410660 41380 410712
rect 239496 410660 239548 410712
rect 24768 410592 24820 410644
rect 237564 410592 237616 410644
rect 252468 410592 252520 410644
rect 264980 410592 265032 410644
rect 8208 410524 8260 410576
rect 235632 410524 235684 410576
rect 235908 410524 235960 410576
rect 262772 410524 262824 410576
rect 3424 410456 3476 410508
rect 7564 410456 7616 410508
rect 187608 410456 187660 410508
rect 256976 410456 257028 410508
rect 202788 410388 202840 410440
rect 258908 410388 258960 410440
rect 3424 410320 3476 410372
rect 219348 410320 219400 410372
rect 260840 410320 260892 410372
rect 271236 409912 271288 409964
rect 271788 409912 271840 409964
rect 275100 409912 275152 409964
rect 275928 409912 275980 409964
rect 280988 409912 281040 409964
rect 281448 409912 281500 409964
rect 284852 409912 284904 409964
rect 285588 409912 285640 409964
rect 290648 409912 290700 409964
rect 291108 409912 291160 409964
rect 294604 409912 294656 409964
rect 295248 409912 295300 409964
rect 298468 409912 298520 409964
rect 299388 409912 299440 409964
rect 304264 409912 304316 409964
rect 304908 409912 304960 409964
rect 184204 408416 184256 408468
rect 232044 408416 232096 408468
rect 3516 405628 3568 405680
rect 232044 405628 232096 405680
rect 307024 404336 307076 404388
rect 580080 404336 580132 404388
rect 3424 404268 3476 404320
rect 232044 404268 232096 404320
rect 307208 404268 307260 404320
rect 580264 404268 580316 404320
rect 580080 404200 580132 404252
rect 580448 404200 580500 404252
rect 195244 402908 195296 402960
rect 232044 402908 232096 402960
rect 3608 401548 3660 401600
rect 232044 401548 232096 401600
rect 307300 401276 307352 401328
rect 309784 401276 309836 401328
rect 4804 400120 4856 400172
rect 232044 400120 232096 400172
rect 307208 400120 307260 400172
rect 580356 400120 580408 400172
rect 307300 398896 307352 398948
rect 307484 398896 307536 398948
rect 3700 398760 3752 398812
rect 232044 398760 232096 398812
rect 307484 398760 307536 398812
rect 580080 398760 580132 398812
rect 198004 397400 198056 397452
rect 232044 397400 232096 397452
rect 3792 395972 3844 396024
rect 232044 395972 232096 396024
rect 3884 394612 3936 394664
rect 231952 394612 232004 394664
rect 307484 394612 307536 394664
rect 580540 394612 580592 394664
rect 3976 393252 4028 393304
rect 232044 393252 232096 393304
rect 307484 393252 307536 393304
rect 580632 393252 580684 393304
rect 220084 391892 220136 391944
rect 232044 391892 232096 391944
rect 307116 390532 307168 390584
rect 580080 390532 580132 390584
rect 4068 390464 4120 390516
rect 232044 390464 232096 390516
rect 3332 389104 3384 389156
rect 231952 389104 232004 389156
rect 307668 389104 307720 389156
rect 580724 389104 580776 389156
rect 10324 389036 10376 389088
rect 232044 389036 232096 389088
rect 3240 387744 3292 387796
rect 232044 387744 232096 387796
rect 307668 387744 307720 387796
rect 580816 387744 580868 387796
rect 3148 386316 3200 386368
rect 232044 386316 232096 386368
rect 3056 384956 3108 385008
rect 232044 384956 232096 385008
rect 2964 383596 3016 383648
rect 231860 383596 231912 383648
rect 307668 383596 307720 383648
rect 580908 383596 580960 383648
rect 2872 382168 2924 382220
rect 232044 382168 232096 382220
rect 307668 382168 307720 382220
rect 580172 382168 580224 382220
rect 2780 380808 2832 380860
rect 232044 380808 232096 380860
rect 306840 380808 306892 380860
rect 312544 380808 312596 380860
rect 7564 379448 7616 379500
rect 232044 379448 232096 379500
rect 307668 378156 307720 378208
rect 580172 378156 580224 378208
rect 3424 378088 3476 378140
rect 232044 378088 232096 378140
rect 3516 376660 3568 376712
rect 232044 376660 232096 376712
rect 3516 374008 3568 374060
rect 232044 374008 232096 374060
rect 3608 372580 3660 372632
rect 232044 372580 232096 372632
rect 3424 371220 3476 371272
rect 232044 371220 232096 371272
rect 307668 371220 307720 371272
rect 320824 371220 320876 371272
rect 3148 367072 3200 367124
rect 232044 367072 232096 367124
rect 7564 365712 7616 365764
rect 232044 365712 232096 365764
rect 307668 365712 307720 365764
rect 461584 365712 461636 365764
rect 307116 365644 307168 365696
rect 580172 365644 580224 365696
rect 307668 364352 307720 364404
rect 316684 364352 316736 364404
rect 22836 362924 22888 362976
rect 232044 362924 232096 362976
rect 307300 362924 307352 362976
rect 331864 362924 331916 362976
rect 3240 361564 3292 361616
rect 232044 361564 232096 361616
rect 3332 357416 3384 357468
rect 232044 357416 232096 357468
rect 307668 356328 307720 356380
rect 309784 356328 309836 356380
rect 14556 356056 14608 356108
rect 232044 356056 232096 356108
rect 307668 354696 307720 354748
rect 324964 354696 325016 354748
rect 4068 353268 4120 353320
rect 232044 353268 232096 353320
rect 307116 353200 307168 353252
rect 580172 353200 580224 353252
rect 25504 351908 25556 351960
rect 232044 351908 232096 351960
rect 3976 350548 4028 350600
rect 232044 350548 232096 350600
rect 3884 347760 3936 347812
rect 232044 347760 232096 347812
rect 307668 347760 307720 347812
rect 323584 347760 323636 347812
rect 3792 346400 3844 346452
rect 232044 346400 232096 346452
rect 15844 345040 15896 345092
rect 232044 345040 232096 345092
rect 32404 343680 32456 343732
rect 232044 343680 232096 343732
rect 3700 343612 3752 343664
rect 231860 343612 231912 343664
rect 3608 342252 3660 342304
rect 232044 342252 232096 342304
rect 306288 342252 306340 342304
rect 460204 342252 460256 342304
rect 3516 340892 3568 340944
rect 232044 340892 232096 340944
rect 320824 340144 320876 340196
rect 580172 340144 580224 340196
rect 307208 339736 307260 339788
rect 3424 339464 3476 339516
rect 232044 339464 232096 339516
rect 307208 339464 307260 339516
rect 318064 339464 318116 339516
rect 17224 338104 17276 338156
rect 232044 338104 232096 338156
rect 307208 338104 307260 338156
rect 406384 338104 406436 338156
rect 234804 337900 234856 337952
rect 235126 337900 235178 337952
rect 236092 337943 236144 337952
rect 236092 337909 236101 337943
rect 236101 337909 236135 337943
rect 236135 337909 236144 337943
rect 236092 337900 236144 337909
rect 262450 337900 262502 337952
rect 303850 337900 303902 337952
rect 305828 337900 305880 337952
rect 235264 337832 235316 337884
rect 239082 337832 239134 337884
rect 241658 337832 241710 337884
rect 244602 337832 244654 337884
rect 246350 337832 246402 337884
rect 247454 337832 247506 337884
rect 257206 337832 257258 337884
rect 236092 337764 236144 337816
rect 236966 337764 237018 337816
rect 240140 337764 240192 337816
rect 240922 337764 240974 337816
rect 242164 337764 242216 337816
rect 243268 337764 243320 337816
rect 243590 337764 243642 337816
rect 246120 337764 246172 337816
rect 247132 337764 247184 337816
rect 251594 337764 251646 337816
rect 251916 337764 251968 337816
rect 253986 337764 254038 337816
rect 254492 337764 254544 337816
rect 255642 337764 255694 337816
rect 256148 337764 256200 337816
rect 258172 337764 258224 337816
rect 259322 337764 259374 337816
rect 261392 337764 261444 337816
rect 262174 337764 262226 337816
rect 234896 337696 234948 337748
rect 262312 337628 262364 337680
rect 275514 337832 275566 337884
rect 276066 337832 276118 337884
rect 280298 337832 280350 337884
rect 300446 337832 300498 337884
rect 300722 337832 300774 337884
rect 301734 337832 301786 337884
rect 305920 337832 305972 337884
rect 262496 337764 262548 337816
rect 263462 337764 263514 337816
rect 267970 337764 268022 337816
rect 268936 337764 268988 337816
rect 271650 337764 271702 337816
rect 278918 337764 278970 337816
rect 279976 337764 280028 337816
rect 281310 337764 281362 337816
rect 281586 337764 281638 337816
rect 282552 337764 282604 337816
rect 285680 337764 285732 337816
rect 286554 337764 286606 337816
rect 287336 337764 287388 337816
rect 288118 337764 288170 337816
rect 289360 337764 289412 337816
rect 289682 337764 289734 337816
rect 290786 337764 290838 337816
rect 292810 337764 292862 337816
rect 293592 337764 293644 337816
rect 296168 337764 296220 337816
rect 296490 337764 296542 337816
rect 280988 337696 281040 337748
rect 300032 337628 300084 337680
rect 302286 337764 302338 337816
rect 303344 337764 303396 337816
rect 304402 337764 304454 337816
rect 305000 337764 305052 337816
rect 277860 337152 277912 337204
rect 278412 337152 278464 337204
rect 231124 336608 231176 336660
rect 254676 336676 254728 336728
rect 262956 336676 263008 336728
rect 265716 336676 265768 336728
rect 293408 336676 293460 336728
rect 312544 336676 312596 336728
rect 272524 336608 272576 336660
rect 226984 336540 227036 336592
rect 274640 336608 274692 336660
rect 224224 336472 224276 336524
rect 261484 336472 261536 336524
rect 288440 336472 288492 336524
rect 294696 336472 294748 336524
rect 320824 336472 320876 336524
rect 125508 336404 125560 336456
rect 249800 336404 249852 336456
rect 263784 336404 263836 336456
rect 271144 336404 271196 336456
rect 295524 336404 295576 336456
rect 322204 336404 322256 336456
rect 114468 336336 114520 336388
rect 248604 336336 248656 336388
rect 255504 336336 255556 336388
rect 35164 336268 35216 336320
rect 238392 336268 238444 336320
rect 253204 336268 253256 336320
rect 28264 336200 28316 336252
rect 236276 336200 236328 336252
rect 261484 336268 261536 336320
rect 263968 336268 264020 336320
rect 270684 336268 270736 336320
rect 297272 336336 297324 336388
rect 307024 336336 307076 336388
rect 307208 336336 307260 336388
rect 290372 336268 290424 336320
rect 264152 336200 264204 336252
rect 21364 336132 21416 336184
rect 237196 336132 237248 336184
rect 249616 336132 249668 336184
rect 264704 336132 264756 336184
rect 270224 336132 270276 336184
rect 292948 336132 293000 336184
rect 297640 336200 297692 336252
rect 327724 336268 327776 336320
rect 336004 336132 336056 336184
rect 18604 336064 18656 336116
rect 252468 336064 252520 336116
rect 265256 336064 265308 336116
rect 269396 336064 269448 336116
rect 284024 336064 284076 336116
rect 400864 336064 400916 336116
rect 10324 335996 10376 336048
rect 235540 335996 235592 336048
rect 245476 335996 245528 336048
rect 233976 335928 234028 335980
rect 257620 335928 257672 335980
rect 264244 335996 264296 336048
rect 269948 335996 270000 336048
rect 287060 335996 287112 336048
rect 292580 335996 292632 336048
rect 479524 335996 479576 336048
rect 233884 335860 233936 335912
rect 254216 335860 254268 335912
rect 255872 335860 255924 335912
rect 234068 335792 234120 335844
rect 265164 335928 265216 335980
rect 294144 335928 294196 335980
rect 294236 335928 294288 335980
rect 313924 335928 313976 335980
rect 268476 335860 268528 335912
rect 273904 335860 273956 335912
rect 293040 335860 293092 335912
rect 305736 335860 305788 335912
rect 307024 335903 307076 335912
rect 307024 335869 307033 335903
rect 307033 335869 307067 335903
rect 307067 335869 307076 335903
rect 307024 335860 307076 335869
rect 268568 335792 268620 335844
rect 276664 335792 276716 335844
rect 282368 335792 282420 335844
rect 282828 335792 282880 335844
rect 284484 335792 284536 335844
rect 294420 335792 294472 335844
rect 301596 335792 301648 335844
rect 302148 335792 302200 335844
rect 305092 335792 305144 335844
rect 229744 335724 229796 335776
rect 267464 335724 267516 335776
rect 270500 335724 270552 335776
rect 278780 335724 278832 335776
rect 283012 335724 283064 335776
rect 283656 335724 283708 335776
rect 293776 335724 293828 335776
rect 306288 335724 306340 335776
rect 283380 335656 283432 335708
rect 283564 335656 283616 335708
rect 290096 335656 290148 335708
rect 292764 335656 292816 335708
rect 296812 335656 296864 335708
rect 305184 335656 305236 335708
rect 273536 335588 273588 335640
rect 273812 335588 273864 335640
rect 280620 335588 280672 335640
rect 281264 335588 281316 335640
rect 281724 335588 281776 335640
rect 284668 335588 284720 335640
rect 293408 335588 293460 335640
rect 302700 335588 302752 335640
rect 303528 335588 303580 335640
rect 267556 335520 267608 335572
rect 268384 335520 268436 335572
rect 294788 335520 294840 335572
rect 295248 335520 295300 335572
rect 297180 335520 297232 335572
rect 272616 335452 272668 335504
rect 273076 335452 273128 335504
rect 273812 335452 273864 335504
rect 274364 335452 274416 335504
rect 236736 335384 236788 335436
rect 243452 335384 243504 335436
rect 257344 335384 257396 335436
rect 263324 335384 263376 335436
rect 267004 335384 267056 335436
rect 267556 335384 267608 335436
rect 268292 335384 268344 335436
rect 268752 335384 268804 335436
rect 272248 335384 272300 335436
rect 272984 335384 273036 335436
rect 274916 335384 274968 335436
rect 275744 335384 275796 335436
rect 276480 335384 276532 335436
rect 277308 335384 277360 335436
rect 277492 335384 277544 335436
rect 278228 335384 278280 335436
rect 255320 335316 255372 335368
rect 256792 335316 256844 335368
rect 226248 335044 226300 335096
rect 219348 334976 219400 335028
rect 261024 335316 261076 335368
rect 261576 335316 261628 335368
rect 263048 335316 263100 335368
rect 267832 335316 267884 335368
rect 268568 335316 268620 335368
rect 269948 335316 270000 335368
rect 270408 335316 270460 335368
rect 271512 335316 271564 335368
rect 271788 335316 271840 335368
rect 275468 335316 275520 335368
rect 275928 335316 275980 335368
rect 276204 335316 276256 335368
rect 276940 335316 276992 335368
rect 280712 335316 280764 335368
rect 280896 335316 280948 335368
rect 282000 335316 282052 335368
rect 282276 335316 282328 335368
rect 283932 335452 283984 335504
rect 284484 335452 284536 335504
rect 284852 335452 284904 335504
rect 287796 335452 287848 335504
rect 288348 335452 288400 335504
rect 291936 335452 291988 335504
rect 292304 335452 292356 335504
rect 283288 335384 283340 335436
rect 284208 335384 284260 335436
rect 286508 335384 286560 335436
rect 286968 335384 287020 335436
rect 289820 335384 289872 335436
rect 290832 335384 290884 335436
rect 291660 335384 291712 335436
rect 292028 335384 292080 335436
rect 284576 335316 284628 335368
rect 284944 335316 284996 335368
rect 285128 335316 285180 335368
rect 285220 335316 285272 335368
rect 285404 335316 285456 335368
rect 286140 335316 286192 335368
rect 285128 335180 285180 335232
rect 286416 335316 286468 335368
rect 286784 335316 286836 335368
rect 287244 335316 287296 335368
rect 287520 335316 287572 335368
rect 287704 335316 287756 335368
rect 287980 335316 288032 335368
rect 288348 335316 288400 335368
rect 289084 335316 289136 335368
rect 289268 335316 289320 335368
rect 290648 335316 290700 335368
rect 291016 335316 291068 335368
rect 291384 335316 291436 335368
rect 291844 335316 291896 335368
rect 291936 335316 291988 335368
rect 292212 335316 292264 335368
rect 294052 335316 294104 335368
rect 294696 335316 294748 335368
rect 288164 335248 288216 335300
rect 295892 335452 295944 335504
rect 296444 335452 296496 335504
rect 298468 335452 298520 335504
rect 299480 335452 299532 335504
rect 299572 335452 299624 335504
rect 300308 335452 300360 335504
rect 295984 335384 296036 335436
rect 296352 335384 296404 335436
rect 298744 335384 298796 335436
rect 299020 335384 299072 335436
rect 301412 335520 301464 335572
rect 302056 335520 302108 335572
rect 301136 335452 301188 335504
rect 301780 335452 301832 335504
rect 302976 335452 303028 335504
rect 303528 335452 303580 335504
rect 302424 335384 302476 335436
rect 303068 335384 303120 335436
rect 304540 335384 304592 335436
rect 304908 335384 304960 335436
rect 295340 335316 295392 335368
rect 295892 335316 295944 335368
rect 297456 335316 297508 335368
rect 297916 335316 297968 335368
rect 299204 335316 299256 335368
rect 299388 335316 299440 335368
rect 300860 335316 300912 335368
rect 301412 335316 301464 335368
rect 301872 335316 301924 335368
rect 302148 335316 302200 335368
rect 302976 335316 303028 335368
rect 303252 335316 303304 335368
rect 304172 335316 304224 335368
rect 304356 335316 304408 335368
rect 286416 335180 286468 335232
rect 290004 335180 290056 335232
rect 294604 335180 294656 335232
rect 313280 335112 313332 335164
rect 271972 335044 272024 335096
rect 307760 335044 307812 335096
rect 272156 334976 272208 335028
rect 309140 334976 309192 335028
rect 210976 334908 211028 334960
rect 260012 334908 260064 334960
rect 275100 334908 275152 334960
rect 333980 334908 334032 334960
rect 176568 334840 176620 334892
rect 255964 334840 256016 334892
rect 261852 334840 261904 334892
rect 275284 334840 275336 334892
rect 335360 334840 335412 334892
rect 158628 334772 158680 334824
rect 253848 334772 253900 334824
rect 279148 334772 279200 334824
rect 368480 334772 368532 334824
rect 126888 334704 126940 334756
rect 249984 334704 250036 334756
rect 293132 334704 293184 334756
rect 293776 334704 293828 334756
rect 305644 334704 305696 334756
rect 306288 334704 306340 334756
rect 489920 334704 489972 334756
rect 97908 334636 97960 334688
rect 246580 334636 246632 334688
rect 298192 334636 298244 334688
rect 525064 334636 525116 334688
rect 39304 334568 39356 334620
rect 236460 334568 236512 334620
rect 236644 334568 236696 334620
rect 242900 334568 242952 334620
rect 244004 334568 244056 334620
rect 248696 334568 248748 334620
rect 249524 334568 249576 334620
rect 252652 334568 252704 334620
rect 253388 334568 253440 334620
rect 271420 334568 271472 334620
rect 271696 334568 271748 334620
rect 276480 334568 276532 334620
rect 276756 334568 276808 334620
rect 284760 334568 284812 334620
rect 285404 334568 285456 334620
rect 239496 334500 239548 334552
rect 251456 334500 251508 334552
rect 251824 334500 251876 334552
rect 265072 334500 265124 334552
rect 266084 334500 266136 334552
rect 284392 334500 284444 334552
rect 285496 334500 285548 334552
rect 297456 334500 297508 334552
rect 297824 334500 297876 334552
rect 298008 334500 298060 334552
rect 525800 334568 525852 334620
rect 304080 334500 304132 334552
rect 304448 334500 304500 334552
rect 296996 334432 297048 334484
rect 297548 334432 297600 334484
rect 269212 334364 269264 334416
rect 269948 334364 270000 334416
rect 284944 334364 284996 334416
rect 285220 334364 285272 334416
rect 285956 334364 286008 334416
rect 291568 334364 291620 334416
rect 292488 334364 292540 334416
rect 292856 334364 292908 334416
rect 293224 334364 293276 334416
rect 297088 334364 297140 334416
rect 297824 334364 297876 334416
rect 290280 334296 290332 334348
rect 291016 334296 291068 334348
rect 292764 334228 292816 334280
rect 293408 334228 293460 334280
rect 230388 333616 230440 333668
rect 262312 333616 262364 333668
rect 272892 333616 272944 333668
rect 316040 333616 316092 333668
rect 219256 333548 219308 333600
rect 261116 333548 261168 333600
rect 288440 333548 288492 333600
rect 338120 333548 338172 333600
rect 183468 333480 183520 333532
rect 255320 333480 255372 333532
rect 273536 333480 273588 333532
rect 324320 333480 324372 333532
rect 169668 333412 169720 333464
rect 255136 333412 255188 333464
rect 279608 333412 279660 333464
rect 372620 333412 372672 333464
rect 144828 333344 144880 333396
rect 252100 333344 252152 333396
rect 268476 333344 268528 333396
rect 269028 333344 269080 333396
rect 272708 333344 272760 333396
rect 273076 333344 273128 333396
rect 282184 333344 282236 333396
rect 282828 333344 282880 333396
rect 286416 333344 286468 333396
rect 426440 333344 426492 333396
rect 95148 333276 95200 333328
rect 246212 333276 246264 333328
rect 273720 333276 273772 333328
rect 274088 333276 274140 333328
rect 277952 333276 278004 333328
rect 278688 333276 278740 333328
rect 279240 333276 279292 333328
rect 280068 333276 280120 333328
rect 287152 333276 287204 333328
rect 434720 333276 434772 333328
rect 29644 333208 29696 333260
rect 237748 333208 237800 333260
rect 241520 333208 241572 333260
rect 242256 333208 242308 333260
rect 245936 333208 245988 333260
rect 246396 333208 246448 333260
rect 251640 333208 251692 333260
rect 252008 333208 252060 333260
rect 258356 333208 258408 333260
rect 258724 333208 258776 333260
rect 266636 333208 266688 333260
rect 266912 333208 266964 333260
rect 267188 333208 267240 333260
rect 267464 333208 267516 333260
rect 268200 333208 268252 333260
rect 269028 333208 269080 333260
rect 269580 333208 269632 333260
rect 270132 333208 270184 333260
rect 270868 333208 270920 333260
rect 271512 333208 271564 333260
rect 272432 333208 272484 333260
rect 272708 333208 272760 333260
rect 273996 333208 274048 333260
rect 274364 333208 274416 333260
rect 277676 333208 277728 333260
rect 278504 333208 278556 333260
rect 279332 333208 279384 333260
rect 279792 333208 279844 333260
rect 280620 333208 280672 333260
rect 281080 333208 281132 333260
rect 282184 333208 282236 333260
rect 282644 333208 282696 333260
rect 283748 333208 283800 333260
rect 284024 333208 284076 333260
rect 284852 333208 284904 333260
rect 285588 333208 285640 333260
rect 286140 333208 286192 333260
rect 286876 333208 286928 333260
rect 287428 333208 287480 333260
rect 288072 333208 288124 333260
rect 288992 333208 289044 333260
rect 289636 333208 289688 333260
rect 291292 333208 291344 333260
rect 292212 333208 292264 333260
rect 293132 333208 293184 333260
rect 293684 333208 293736 333260
rect 295064 333208 295116 333260
rect 500960 333208 501012 333260
rect 289452 333140 289504 333192
rect 289728 333140 289780 333192
rect 295800 333140 295852 333192
rect 296260 333140 296312 333192
rect 298652 333140 298704 333192
rect 298928 333140 298980 333192
rect 299940 333140 299992 333192
rect 300400 333140 300452 333192
rect 298376 333072 298428 333124
rect 299020 333072 299072 333124
rect 300216 333072 300268 333124
rect 300584 333072 300636 333124
rect 3056 332528 3108 332580
rect 233148 332528 233200 332580
rect 234528 332188 234580 332240
rect 262864 332188 262916 332240
rect 273352 332188 273404 332240
rect 320180 332188 320232 332240
rect 223488 332120 223540 332172
rect 261668 332120 261720 332172
rect 276572 332120 276624 332172
rect 342260 332120 342312 332172
rect 162768 332052 162820 332104
rect 254400 332052 254452 332104
rect 347780 332052 347832 332104
rect 136548 331984 136600 332036
rect 251272 331984 251324 332036
rect 283380 331984 283432 332036
rect 405740 331984 405792 332036
rect 108948 331916 109000 331968
rect 247868 331916 247920 331968
rect 276572 331916 276624 331968
rect 277124 331916 277176 331968
rect 465172 331916 465224 331968
rect 68928 331848 68980 331900
rect 243084 331848 243136 331900
rect 296444 331848 296496 331900
rect 507860 331848 507912 331900
rect 242992 331372 243044 331424
rect 243360 331372 243412 331424
rect 239036 331168 239088 331220
rect 239220 331100 239272 331152
rect 240692 331100 240744 331152
rect 240968 331100 241020 331152
rect 301320 331100 301372 331152
rect 301596 331100 301648 331152
rect 257436 330964 257488 331016
rect 244740 330896 244792 330948
rect 244924 330896 244976 330948
rect 245016 330896 245068 330948
rect 245200 330896 245252 330948
rect 256424 330896 256476 330948
rect 299112 330896 299164 330948
rect 213828 330828 213880 330880
rect 260472 330828 260524 330880
rect 274272 330828 274324 330880
rect 327080 330828 327132 330880
rect 187608 330760 187660 330812
rect 179328 330692 179380 330744
rect 147588 330624 147640 330676
rect 252560 330760 252612 330812
rect 274824 330760 274876 330812
rect 332600 330760 332652 330812
rect 102048 330556 102100 330608
rect 246948 330556 247000 330608
rect 247684 330556 247736 330608
rect 247868 330556 247920 330608
rect 35808 330488 35860 330540
rect 245016 330488 245068 330540
rect 245568 330488 245620 330540
rect 246212 330488 246264 330540
rect 246856 330488 246908 330540
rect 247316 330488 247368 330540
rect 247960 330488 248012 330540
rect 250536 330692 250588 330744
rect 277768 330692 277820 330744
rect 357440 330692 357492 330744
rect 250628 330624 250680 330676
rect 263784 330624 263836 330676
rect 264428 330624 264480 330676
rect 270316 330624 270368 330676
rect 271328 330624 271380 330676
rect 271604 330624 271656 330676
rect 285772 330624 285824 330676
rect 423680 330624 423732 330676
rect 265164 330556 265216 330608
rect 265808 330556 265860 330608
rect 250260 330488 250312 330540
rect 251088 330488 251140 330540
rect 252836 330488 252888 330540
rect 253388 330488 253440 330540
rect 265532 330488 265584 330540
rect 266268 330488 266320 330540
rect 244556 330420 244608 330472
rect 245108 330420 245160 330472
rect 247224 330420 247276 330472
rect 248144 330420 248196 330472
rect 249984 330420 250036 330472
rect 250076 330420 250128 330472
rect 251732 330420 251784 330472
rect 252376 330420 252428 330472
rect 253112 330420 253164 330472
rect 253296 330420 253348 330472
rect 265348 330420 265400 330472
rect 265992 330420 266044 330472
rect 305092 330556 305144 330608
rect 514760 330556 514812 330608
rect 272892 330488 272944 330540
rect 273168 330488 273220 330540
rect 282092 330488 282144 330540
rect 282276 330488 282328 330540
rect 302516 330488 302568 330540
rect 564440 330488 564492 330540
rect 270408 330420 270460 330472
rect 270684 330420 270736 330472
rect 271420 330420 271472 330472
rect 295708 330420 295760 330472
rect 296628 330420 296680 330472
rect 298836 330463 298888 330472
rect 298836 330429 298845 330463
rect 298845 330429 298879 330463
rect 298879 330429 298888 330463
rect 298836 330420 298888 330429
rect 301044 330420 301096 330472
rect 301964 330420 302016 330472
rect 302884 330420 302936 330472
rect 303160 330420 303212 330472
rect 303804 330420 303856 330472
rect 304448 330420 304500 330472
rect 244832 330352 244884 330404
rect 245292 330352 245344 330404
rect 245844 330352 245896 330404
rect 246028 330352 246080 330404
rect 247500 330352 247552 330404
rect 248236 330352 248288 330404
rect 263692 330352 263744 330404
rect 264060 330352 264112 330404
rect 269304 330352 269356 330404
rect 270316 330352 270368 330404
rect 274180 330352 274232 330404
rect 274456 330352 274508 330404
rect 278412 330352 278464 330404
rect 278596 330352 278648 330404
rect 279056 330352 279108 330404
rect 279792 330352 279844 330404
rect 280804 330395 280856 330404
rect 280804 330361 280813 330395
rect 280813 330361 280847 330395
rect 280847 330361 280856 330395
rect 280804 330352 280856 330361
rect 281908 330352 281960 330404
rect 282736 330352 282788 330404
rect 299848 330352 299900 330404
rect 300676 330352 300728 330404
rect 252744 330284 252796 330336
rect 253296 330284 253348 330336
rect 280252 330284 280304 330336
rect 281172 330284 281224 330336
rect 246028 330216 246080 330268
rect 246672 330216 246724 330268
rect 248604 330216 248656 330268
rect 249156 330216 249208 330268
rect 300308 330216 300360 330268
rect 280436 330148 280488 330200
rect 281448 330148 281500 330200
rect 248880 329468 248932 329520
rect 249248 329468 249300 329520
rect 227628 329400 227680 329452
rect 262036 329400 262088 329452
rect 288624 329400 288676 329452
rect 289544 329400 289596 329452
rect 188988 329332 189040 329384
rect 257528 329332 257580 329384
rect 275652 329332 275704 329384
rect 339500 329332 339552 329384
rect 166908 329264 166960 329316
rect 254860 329264 254912 329316
rect 283932 329264 283984 329316
rect 365720 329264 365772 329316
rect 140688 329196 140740 329248
rect 251824 329196 251876 329248
rect 285312 329196 285364 329248
rect 419540 329196 419592 329248
rect 115848 329128 115900 329180
rect 248788 329128 248840 329180
rect 271788 329128 271840 329180
rect 305000 329128 305052 329180
rect 305184 329128 305236 329180
rect 518900 329128 518952 329180
rect 43444 329060 43496 329112
rect 239864 329060 239916 329112
rect 298560 329060 298612 329112
rect 529204 329060 529256 329112
rect 254584 329035 254636 329044
rect 254584 329001 254593 329035
rect 254593 329001 254627 329035
rect 254627 329001 254636 329035
rect 254584 328992 254636 329001
rect 252836 328380 252888 328432
rect 253480 328380 253532 328432
rect 253020 328312 253072 328364
rect 253664 328312 253716 328364
rect 231768 328040 231820 328092
rect 262680 328040 262732 328092
rect 184848 327972 184900 328024
rect 256976 327972 257028 328024
rect 294144 327972 294196 328024
rect 331220 327972 331272 328024
rect 160008 327904 160060 327956
rect 254492 327904 254544 327956
rect 277216 327904 277268 327956
rect 353300 327904 353352 327956
rect 151728 327836 151780 327888
rect 252744 327836 252796 327888
rect 284576 327836 284628 327888
rect 415492 327836 415544 327888
rect 85488 327768 85540 327820
rect 245200 327768 245252 327820
rect 293592 327768 293644 327820
rect 46204 327700 46256 327752
rect 240324 327700 240376 327752
rect 293776 327768 293828 327820
rect 484400 327768 484452 327820
rect 303528 327700 303580 327752
rect 566464 327700 566516 327752
rect 293684 327564 293736 327616
rect 248788 327156 248840 327208
rect 249708 327156 249760 327208
rect 302884 327088 302936 327140
rect 303436 327088 303488 327140
rect 237564 326680 237616 326732
rect 237748 326680 237800 326732
rect 217968 326612 218020 326664
rect 261116 326612 261168 326664
rect 277308 326612 277360 326664
rect 346400 326612 346452 326664
rect 191748 326544 191800 326596
rect 257804 326544 257856 326596
rect 154488 326476 154540 326528
rect 252652 326476 252704 326528
rect 113088 326408 113140 326460
rect 248512 326408 248564 326460
rect 104808 326340 104860 326392
rect 247132 326340 247184 326392
rect 254400 326340 254452 326392
rect 254952 326340 255004 326392
rect 255412 326340 255464 326392
rect 255780 326340 255832 326392
rect 257068 326340 257120 326392
rect 257896 326340 257948 326392
rect 235172 326272 235224 326324
rect 235908 326272 235960 326324
rect 236368 326272 236420 326324
rect 237104 326272 237156 326324
rect 237840 326272 237892 326324
rect 238484 326272 238536 326324
rect 243544 326272 243596 326324
rect 244188 326272 244240 326324
rect 258448 326544 258500 326596
rect 279240 326544 279292 326596
rect 375380 326544 375432 326596
rect 285036 326476 285088 326528
rect 285220 326476 285272 326528
rect 292120 326519 292172 326528
rect 292120 326485 292129 326519
rect 292129 326485 292163 326519
rect 292163 326485 292172 326519
rect 292120 326476 292172 326485
rect 294420 326476 294472 326528
rect 412640 326476 412692 326528
rect 258908 326408 258960 326460
rect 259644 326408 259696 326460
rect 260104 326408 260156 326460
rect 288348 326408 288400 326460
rect 441620 326408 441672 326460
rect 258356 326340 258408 326392
rect 258448 326340 258500 326392
rect 259000 326340 259052 326392
rect 259552 326340 259604 326392
rect 260012 326340 260064 326392
rect 262588 326340 262640 326392
rect 263140 326340 263192 326392
rect 283564 326340 283616 326392
rect 283748 326340 283800 326392
rect 283932 326340 283984 326392
rect 284116 326340 284168 326392
rect 286324 326340 286376 326392
rect 286692 326340 286744 326392
rect 287060 326340 287112 326392
rect 287704 326340 287756 326392
rect 291016 326340 291068 326392
rect 258816 326272 258868 326324
rect 234712 326204 234764 326256
rect 235816 326204 235868 326256
rect 237656 326204 237708 326256
rect 238116 326204 238168 326256
rect 239128 326204 239180 326256
rect 239772 326204 239824 326256
rect 240416 326204 240468 326256
rect 241428 326204 241480 326256
rect 241796 326204 241848 326256
rect 242440 326204 242492 326256
rect 243268 326204 243320 326256
rect 243728 326204 243780 326256
rect 255412 326204 255464 326256
rect 256056 326204 256108 326256
rect 258172 326204 258224 326256
rect 237932 326136 237984 326188
rect 238668 326136 238720 326188
rect 239036 326136 239088 326188
rect 240048 326136 240100 326188
rect 240140 326136 240192 326188
rect 241336 326136 241388 326188
rect 255688 326136 255740 326188
rect 256608 326136 256660 326188
rect 259828 326272 259880 326324
rect 260748 326272 260800 326324
rect 259736 326204 259788 326256
rect 260288 326204 260340 326256
rect 284668 326204 284720 326256
rect 284944 326204 284996 326256
rect 259552 326136 259604 326188
rect 260564 326136 260616 326188
rect 292672 326340 292724 326392
rect 481640 326340 481692 326392
rect 292212 326204 292264 326256
rect 237472 326068 237524 326120
rect 238208 326068 238260 326120
rect 255504 326068 255556 326120
rect 256516 326068 256568 326120
rect 258908 326068 258960 326120
rect 285956 326068 286008 326120
rect 286324 326068 286376 326120
rect 291108 326068 291160 326120
rect 285864 326000 285916 326052
rect 286600 326000 286652 326052
rect 242072 325864 242124 325916
rect 242624 325864 242676 325916
rect 306380 325592 306432 325644
rect 580172 325592 580224 325644
rect 289176 325184 289228 325236
rect 289360 325184 289412 325236
rect 224868 325116 224920 325168
rect 261760 325116 261812 325168
rect 272708 325116 272760 325168
rect 311900 325116 311952 325168
rect 148968 325048 149020 325100
rect 253296 325048 253348 325100
rect 276848 325048 276900 325100
rect 349160 325048 349212 325100
rect 128268 324980 128320 325032
rect 249892 324980 249944 325032
rect 278688 324980 278740 325032
rect 357532 324980 357584 325032
rect 92388 324912 92440 324964
rect 246396 324912 246448 324964
rect 288716 324912 288768 324964
rect 289360 324912 289412 324964
rect 297548 324912 297600 324964
rect 516140 324912 516192 324964
rect 240692 323960 240744 324012
rect 241152 323960 241204 324012
rect 274088 323824 274140 323876
rect 322940 323824 322992 323876
rect 169576 323756 169628 323808
rect 255228 323756 255280 323808
rect 278136 323756 278188 323808
rect 360200 323756 360252 323808
rect 144736 323688 144788 323740
rect 252192 323688 252244 323740
rect 282828 323688 282880 323740
rect 393320 323688 393372 323740
rect 50988 323620 51040 323672
rect 240232 323620 240284 323672
rect 285680 323620 285732 323672
rect 430580 323620 430632 323672
rect 14464 323552 14516 323604
rect 236552 323552 236604 323604
rect 296628 323552 296680 323604
rect 506480 323552 506532 323604
rect 186228 322396 186280 322448
rect 257160 322464 257212 322516
rect 255872 322396 255924 322448
rect 256240 322396 256292 322448
rect 281448 322396 281500 322448
rect 379520 322396 379572 322448
rect 135168 322328 135220 322380
rect 250996 322328 251048 322380
rect 286416 322328 286468 322380
rect 433340 322328 433392 322380
rect 88248 322260 88300 322312
rect 245384 322260 245436 322312
rect 290556 322260 290608 322312
rect 463700 322260 463752 322312
rect 57888 322192 57940 322244
rect 241612 322192 241664 322244
rect 297640 322192 297692 322244
rect 520280 322192 520332 322244
rect 272800 321104 272852 321156
rect 316132 321104 316184 321156
rect 227536 321036 227588 321088
rect 261392 321036 261444 321088
rect 275560 321036 275612 321088
rect 336740 321036 336792 321088
rect 137928 320968 137980 321020
rect 251548 320968 251600 321020
rect 282184 320968 282236 321020
rect 397460 320968 397512 321020
rect 111708 320900 111760 320952
rect 247500 320900 247552 320952
rect 294604 320900 294656 320952
rect 458180 320900 458232 320952
rect 33784 320832 33836 320884
rect 236092 320832 236144 320884
rect 236276 320832 236328 320884
rect 242900 320832 242952 320884
rect 243084 320832 243136 320884
rect 298744 320832 298796 320884
rect 533344 320832 533396 320884
rect 238300 320764 238352 320816
rect 3056 320084 3108 320136
rect 233056 320084 233108 320136
rect 272892 319608 272944 319660
rect 318800 319608 318852 319660
rect 280712 319540 280764 319592
rect 382280 319540 382332 319592
rect 220728 319472 220780 319524
rect 261300 319472 261352 319524
rect 287612 319472 287664 319524
rect 438860 319472 438912 319524
rect 106188 319404 106240 319456
rect 247776 319404 247828 319456
rect 293500 319404 293552 319456
rect 488540 319404 488592 319456
rect 274180 318248 274232 318300
rect 329840 318248 329892 318300
rect 142068 318180 142120 318232
rect 251456 318180 251508 318232
rect 283656 318180 283708 318232
rect 400220 318180 400272 318232
rect 95056 318112 95108 318164
rect 246120 318112 246172 318164
rect 288900 318112 288952 318164
rect 448520 318112 448572 318164
rect 53748 318044 53800 318096
rect 240140 318044 240192 318096
rect 293592 318044 293644 318096
rect 491300 318044 491352 318096
rect 153108 316820 153160 316872
rect 252928 316820 252980 316872
rect 275744 316820 275796 316872
rect 332692 316820 332744 316872
rect 99288 316752 99340 316804
rect 246028 316752 246080 316804
rect 288164 316752 288216 316804
rect 289084 316752 289136 316804
rect 452660 316752 452712 316804
rect 62028 316684 62080 316736
rect 241520 316684 241572 316736
rect 296076 316684 296128 316736
rect 509240 316684 509292 316736
rect 288164 316548 288216 316600
rect 155868 315392 155920 315444
rect 252836 315392 252888 315444
rect 280804 315392 280856 315444
rect 386420 315392 386472 315444
rect 103428 315324 103480 315376
rect 247408 315324 247460 315376
rect 290740 315324 290792 315376
rect 466460 315324 466512 315376
rect 71688 315256 71740 315308
rect 236644 315256 236696 315308
rect 296168 315256 296220 315308
rect 513380 315256 513432 315308
rect 276940 314032 276992 314084
rect 343640 314032 343692 314084
rect 164148 313964 164200 314016
rect 254676 313964 254728 314016
rect 297732 313964 297784 314016
rect 522304 313964 522356 314016
rect 117228 313896 117280 313948
rect 248972 313896 249024 313948
rect 285312 313896 285364 313948
rect 285496 313896 285548 313948
rect 304264 313896 304316 313948
rect 576124 313896 576176 313948
rect 306472 313216 306524 313268
rect 580172 313216 580224 313268
rect 168288 312604 168340 312656
rect 254400 312604 254452 312656
rect 274272 312604 274324 312656
rect 325700 312604 325752 312656
rect 119988 312536 120040 312588
rect 248880 312536 248932 312588
rect 278228 312536 278280 312588
rect 354680 312536 354732 312588
rect 193128 311176 193180 311228
rect 257068 311176 257120 311228
rect 286508 311176 286560 311228
rect 432052 311176 432104 311228
rect 22744 311108 22796 311160
rect 236368 311108 236420 311160
rect 302884 311108 302936 311160
rect 571340 311108 571392 311160
rect 136456 309816 136508 309868
rect 250260 309816 250312 309868
rect 275836 309816 275888 309868
rect 340880 309816 340932 309868
rect 36544 309748 36596 309800
rect 237932 309748 237984 309800
rect 287796 309748 287848 309800
rect 445760 309748 445812 309800
rect 161388 308456 161440 308508
rect 254308 308456 254360 308508
rect 284944 308456 284996 308508
rect 390560 308456 390612 308508
rect 64788 308388 64840 308440
rect 242072 308388 242124 308440
rect 289176 308388 289228 308440
rect 456892 308388 456944 308440
rect 283748 307096 283800 307148
rect 404360 307096 404412 307148
rect 81348 307028 81400 307080
rect 234068 307028 234120 307080
rect 293408 307028 293460 307080
rect 459560 307028 459612 307080
rect 283840 305668 283892 305720
rect 407120 305668 407172 305720
rect 110328 305600 110380 305652
rect 247316 305600 247368 305652
rect 293684 305600 293736 305652
rect 481732 305600 481784 305652
rect 124128 304240 124180 304292
rect 248788 304240 248840 304292
rect 293040 304240 293092 304292
rect 485780 304240 485832 304292
rect 293132 302880 293184 302932
rect 490012 302880 490064 302932
rect 297824 301452 297876 301504
rect 517520 301452 517572 301504
rect 297916 300092 297968 300144
rect 521660 300092 521712 300144
rect 306564 299412 306616 299464
rect 580172 299412 580224 299464
rect 297456 297372 297508 297424
rect 524420 297372 524472 297424
rect 305920 295944 305972 295996
rect 556160 295944 556212 295996
rect 305828 294584 305880 294636
rect 574100 294584 574152 294636
rect 277032 293224 277084 293276
rect 350540 293224 350592 293276
rect 3148 293156 3200 293208
rect 7564 293156 7616 293208
rect 278320 291796 278372 291848
rect 361580 291796 361632 291848
rect 461584 285608 461636 285660
rect 580172 285608 580224 285660
rect 3148 280100 3200 280152
rect 232964 280100 233016 280152
rect 316684 273164 316736 273216
rect 580172 273164 580224 273216
rect 2964 267656 3016 267708
rect 232872 267656 232924 267708
rect 331864 259360 331916 259412
rect 580172 259360 580224 259412
rect 3148 255212 3200 255264
rect 22836 255212 22888 255264
rect 306656 245556 306708 245608
rect 580172 245556 580224 245608
rect 306748 233180 306800 233232
rect 579988 233180 580040 233232
rect 3240 229032 3292 229084
rect 232780 229032 232832 229084
rect 306840 219376 306892 219428
rect 580172 219376 580224 219428
rect 3240 215228 3292 215280
rect 232688 215228 232740 215280
rect 306932 206932 306984 206984
rect 579804 206932 579856 206984
rect 309784 193128 309836 193180
rect 580172 193128 580224 193180
rect 3332 188980 3384 189032
rect 14556 188980 14608 189032
rect 305736 181432 305788 181484
rect 483020 181432 483072 181484
rect 324964 179324 325016 179376
rect 580172 179324 580224 179376
rect 3332 176604 3384 176656
rect 232596 176604 232648 176656
rect 307668 166948 307720 167000
rect 580172 166948 580224 167000
rect 307576 153144 307628 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 25504 150356 25556 150408
rect 307484 139340 307536 139392
rect 580172 139340 580224 139392
rect 307392 126896 307444 126948
rect 580172 126896 580224 126948
rect 3148 124108 3200 124160
rect 232504 124108 232556 124160
rect 307300 113092 307352 113144
rect 579804 113092 579856 113144
rect 323584 100648 323636 100700
rect 580172 100648 580224 100700
rect 307208 86912 307260 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 15844 85484 15896 85536
rect 307116 73108 307168 73160
rect 580172 73108 580224 73160
rect 307024 60664 307076 60716
rect 580172 60664 580224 60716
rect 2872 59304 2924 59356
rect 32404 59304 32456 59356
rect 460204 46860 460256 46912
rect 580172 46860 580224 46912
rect 336004 22720 336056 22772
rect 462320 22720 462372 22772
rect 327724 21360 327776 21412
rect 523132 21360 523184 21412
rect 318064 20612 318116 20664
rect 579988 20612 580040 20664
rect 139308 19932 139360 19984
rect 251916 19932 251968 19984
rect 322204 18572 322256 18624
rect 505100 18572 505152 18624
rect 190368 17212 190420 17264
rect 233976 17212 234028 17264
rect 320824 17212 320876 17264
rect 498200 17212 498252 17264
rect 186136 15852 186188 15904
rect 226984 15852 227036 15904
rect 313924 15852 313976 15904
rect 494704 15852 494756 15904
rect 305644 14560 305696 14612
rect 306748 14560 306800 14612
rect 171968 14424 172020 14476
rect 229744 14424 229796 14476
rect 312544 14424 312596 14476
rect 487620 14424 487672 14476
rect 301320 13744 301372 13796
rect 301688 13744 301740 13796
rect 301688 13608 301740 13660
rect 301872 13608 301924 13660
rect 298928 13540 298980 13592
rect 532516 13540 532568 13592
rect 298836 13472 298888 13524
rect 536104 13472 536156 13524
rect 300216 13404 300268 13456
rect 539600 13404 539652 13456
rect 300124 13336 300176 13388
rect 543188 13336 543240 13388
rect 300032 13268 300084 13320
rect 546684 13268 546736 13320
rect 301412 13200 301464 13252
rect 550272 13200 550324 13252
rect 301596 13132 301648 13184
rect 553768 13132 553820 13184
rect 164884 13064 164936 13116
rect 231124 13064 231176 13116
rect 235816 13064 235868 13116
rect 261576 13064 261628 13116
rect 268476 13064 268528 13116
rect 284300 13064 284352 13116
rect 293316 13064 293368 13116
rect 301504 13064 301556 13116
rect 560852 13064 560904 13116
rect 301872 12996 301924 13048
rect 291752 12384 291804 12436
rect 471060 12384 471112 12436
rect 294788 12316 294840 12368
rect 294880 12248 294932 12300
rect 293224 12112 293276 12164
rect 294880 12112 294932 12164
rect 473360 12316 473412 12368
rect 478144 12248 478196 12300
rect 493508 12180 493560 12232
rect 497096 12112 497148 12164
rect 294972 12044 295024 12096
rect 500592 12044 500644 12096
rect 291936 11976 291988 12028
rect 295892 11976 295944 12028
rect 504180 11976 504232 12028
rect 287704 11908 287756 11960
rect 291384 11908 291436 11960
rect 291568 11908 291620 11960
rect 296260 11908 296312 11960
rect 507676 11908 507728 11960
rect 296352 11840 296404 11892
rect 511264 11840 511316 11892
rect 241428 11772 241480 11824
rect 254584 11772 254636 11824
rect 296444 11772 296496 11824
rect 514852 11772 514904 11824
rect 161296 11704 161348 11756
rect 233884 11704 233936 11756
rect 237012 11704 237064 11756
rect 257344 11704 257396 11756
rect 299020 11704 299072 11756
rect 529020 11704 529072 11756
rect 221556 11432 221608 11484
rect 224224 11432 224276 11484
rect 56508 10956 56560 11008
rect 241980 10956 242032 11008
rect 282276 10956 282328 11008
rect 393044 10956 393096 11008
rect 53656 10888 53708 10940
rect 240692 10888 240744 10940
rect 282460 10888 282512 10940
rect 396540 10888 396592 10940
rect 49608 10820 49660 10872
rect 240600 10820 240652 10872
rect 282368 10820 282420 10872
rect 398840 10820 398892 10872
rect 45468 10752 45520 10804
rect 240508 10752 240560 10804
rect 284116 10752 284168 10804
rect 403624 10752 403676 10804
rect 41328 10684 41380 10736
rect 239128 10684 239180 10736
rect 284024 10684 284076 10736
rect 407212 10684 407264 10736
rect 37188 10616 37240 10668
rect 239312 10616 239364 10668
rect 283932 10616 283984 10668
rect 410800 10616 410852 10668
rect 34428 10548 34480 10600
rect 239220 10548 239272 10600
rect 285128 10548 285180 10600
rect 414296 10548 414348 10600
rect 30104 10480 30156 10532
rect 237840 10480 237892 10532
rect 285220 10480 285272 10532
rect 417884 10480 417936 10532
rect 27528 10412 27580 10464
rect 237656 10412 237708 10464
rect 285036 10412 285088 10464
rect 421380 10412 421432 10464
rect 21824 10344 21876 10396
rect 237748 10344 237800 10396
rect 244096 10344 244148 10396
rect 253204 10344 253256 10396
rect 286600 10344 286652 10396
rect 423772 10344 423824 10396
rect 9588 10276 9640 10328
rect 235172 10276 235224 10328
rect 242808 10276 242860 10328
rect 261484 10276 261536 10328
rect 286692 10276 286744 10328
rect 428464 10276 428516 10328
rect 60648 10208 60700 10260
rect 241888 10208 241940 10260
rect 282552 10208 282604 10260
rect 389456 10208 389508 10260
rect 63224 10140 63276 10192
rect 241796 10140 241848 10192
rect 281080 10140 281132 10192
rect 385960 10140 386012 10192
rect 67548 10072 67600 10124
rect 243360 10072 243412 10124
rect 280896 10072 280948 10124
rect 382372 10072 382424 10124
rect 70308 10004 70360 10056
rect 243452 10004 243504 10056
rect 280988 10004 281040 10056
rect 378876 10004 378928 10056
rect 74448 9936 74500 9988
rect 243268 9936 243320 9988
rect 279700 9936 279752 9988
rect 374000 9936 374052 9988
rect 78588 9868 78640 9920
rect 243544 9868 243596 9920
rect 279608 9868 279660 9920
rect 371700 9868 371752 9920
rect 119896 9800 119948 9852
rect 248604 9800 248656 9852
rect 279792 9800 279844 9852
rect 368204 9800 368256 9852
rect 122748 9732 122800 9784
rect 248696 9732 248748 9784
rect 278412 9732 278464 9784
rect 364616 9732 364668 9784
rect 83280 9596 83332 9648
rect 244740 9596 244792 9648
rect 253480 9596 253532 9648
rect 255964 9596 256016 9648
rect 300400 9596 300452 9648
rect 541992 9596 542044 9648
rect 79692 9528 79744 9580
rect 244648 9528 244700 9580
rect 300492 9528 300544 9580
rect 545488 9528 545540 9580
rect 76196 9460 76248 9512
rect 243084 9460 243136 9512
rect 300308 9460 300360 9512
rect 549076 9460 549128 9512
rect 72608 9392 72660 9444
rect 243176 9392 243228 9444
rect 301780 9392 301832 9444
rect 552664 9392 552716 9444
rect 69112 9324 69164 9376
rect 242992 9324 243044 9376
rect 301320 9324 301372 9376
rect 556252 9324 556304 9376
rect 65524 9256 65576 9308
rect 242440 9256 242492 9308
rect 301688 9256 301740 9308
rect 559748 9256 559800 9308
rect 61936 9188 61988 9240
rect 242348 9188 242400 9240
rect 303068 9188 303120 9240
rect 563244 9188 563296 9240
rect 58440 9120 58492 9172
rect 241704 9120 241756 9172
rect 303160 9120 303212 9172
rect 566832 9120 566884 9172
rect 54944 9052 54996 9104
rect 240416 9052 240468 9104
rect 302976 9052 303028 9104
rect 570328 9052 570380 9104
rect 17040 8984 17092 9036
rect 236276 8984 236328 9036
rect 247592 8984 247644 9036
rect 263968 8984 264020 9036
rect 304448 8984 304500 9036
rect 573916 8984 573968 9036
rect 4068 8916 4120 8968
rect 235080 8916 235132 8968
rect 238116 8916 238168 8968
rect 262496 8916 262548 8968
rect 304356 8916 304408 8968
rect 577412 8916 577464 8968
rect 86868 8848 86920 8900
rect 244832 8848 244884 8900
rect 299112 8848 299164 8900
rect 538404 8848 538456 8900
rect 90364 8780 90416 8832
rect 245936 8780 245988 8832
rect 273812 8780 273864 8832
rect 329196 8780 329248 8832
rect 142436 8712 142488 8764
rect 251640 8712 251692 8764
rect 274364 8712 274416 8764
rect 325608 8712 325660 8764
rect 145932 8644 145984 8696
rect 251732 8644 251784 8696
rect 273720 8644 273772 8696
rect 322112 8644 322164 8696
rect 149520 8576 149572 8628
rect 253388 8576 253440 8628
rect 272616 8576 272668 8628
rect 318524 8576 318576 8628
rect 153016 8508 153068 8560
rect 253112 8508 253164 8560
rect 273076 8508 273128 8560
rect 315028 8508 315080 8560
rect 156604 8440 156656 8492
rect 253020 8440 253072 8492
rect 272984 8440 273036 8492
rect 311440 8440 311492 8492
rect 271328 8372 271380 8424
rect 307944 8372 307996 8424
rect 199108 8236 199160 8288
rect 258908 8236 258960 8288
rect 287888 8236 287940 8288
rect 441528 8236 441580 8288
rect 195612 8168 195664 8220
rect 258724 8168 258776 8220
rect 288072 8168 288124 8220
rect 445024 8168 445076 8220
rect 181444 8100 181496 8152
rect 255688 8100 255740 8152
rect 289360 8100 289412 8152
rect 448612 8100 448664 8152
rect 177856 8032 177908 8084
rect 255872 8032 255924 8084
rect 289268 8032 289320 8084
rect 452108 8032 452160 8084
rect 174268 7964 174320 8016
rect 255596 7964 255648 8016
rect 289452 7964 289504 8016
rect 455696 7964 455748 8016
rect 170772 7896 170824 7948
rect 255780 7896 255832 7948
rect 292120 7896 292172 7948
rect 469864 7896 469916 7948
rect 131764 7828 131816 7880
rect 250076 7828 250128 7880
rect 292028 7828 292080 7880
rect 473452 7828 473504 7880
rect 128176 7760 128228 7812
rect 250168 7760 250220 7812
rect 292212 7760 292264 7812
rect 476948 7760 477000 7812
rect 51356 7692 51408 7744
rect 240876 7692 240928 7744
rect 294144 7692 294196 7744
rect 495900 7692 495952 7744
rect 47860 7624 47912 7676
rect 240968 7624 241020 7676
rect 295156 7624 295208 7676
rect 499396 7624 499448 7676
rect 12348 7556 12400 7608
rect 236184 7556 236236 7608
rect 276664 7556 276716 7608
rect 280712 7556 280764 7608
rect 295064 7556 295116 7608
rect 502984 7556 503036 7608
rect 202696 7488 202748 7540
rect 258816 7488 258868 7540
rect 287980 7488 288032 7540
rect 437940 7488 437992 7540
rect 206192 7420 206244 7472
rect 260104 7420 260156 7472
rect 286324 6876 286376 6928
rect 287796 6876 287848 6928
rect 3424 6808 3476 6860
rect 17224 6808 17276 6860
rect 215668 6808 215720 6860
rect 259828 6808 259880 6860
rect 279884 6808 279936 6860
rect 367008 6808 367060 6860
rect 406384 6808 406436 6860
rect 580172 6808 580224 6860
rect 212172 6740 212224 6792
rect 259736 6740 259788 6792
rect 279516 6740 279568 6792
rect 370596 6740 370648 6792
rect 208584 6672 208636 6724
rect 259920 6672 259972 6724
rect 279424 6672 279476 6724
rect 374092 6672 374144 6724
rect 205088 6604 205140 6656
rect 260012 6604 260064 6656
rect 281172 6604 281224 6656
rect 377680 6604 377732 6656
rect 201500 6536 201552 6588
rect 258448 6536 258500 6588
rect 281264 6536 281316 6588
rect 381176 6536 381228 6588
rect 197912 6468 197964 6520
rect 258632 6468 258684 6520
rect 280620 6468 280672 6520
rect 384764 6468 384816 6520
rect 194416 6400 194468 6452
rect 258540 6400 258592 6452
rect 281356 6400 281408 6452
rect 388260 6400 388312 6452
rect 180248 6332 180300 6384
rect 255504 6332 255556 6384
rect 282736 6332 282788 6384
rect 391848 6332 391900 6384
rect 176660 6264 176712 6316
rect 255412 6264 255464 6316
rect 282092 6264 282144 6316
rect 395344 6264 395396 6316
rect 173164 6196 173216 6248
rect 256148 6196 256200 6248
rect 282644 6196 282696 6248
rect 398932 6196 398984 6248
rect 400864 6196 400916 6248
rect 409604 6196 409656 6248
rect 130568 6128 130620 6180
rect 249984 6128 250036 6180
rect 283472 6128 283524 6180
rect 402520 6128 402572 6180
rect 277860 6060 277912 6112
rect 363512 6060 363564 6112
rect 277952 5992 278004 6044
rect 359924 5992 359976 6044
rect 278504 5924 278556 5976
rect 356336 5924 356388 5976
rect 276572 5856 276624 5908
rect 352840 5856 352892 5908
rect 276480 5788 276532 5840
rect 349252 5788 349304 5840
rect 276388 5720 276440 5772
rect 345756 5720 345808 5772
rect 275468 5652 275520 5704
rect 342168 5652 342220 5704
rect 268568 5584 268620 5636
rect 274824 5584 274876 5636
rect 250444 5516 250496 5568
rect 273904 5516 273956 5568
rect 279516 5516 279568 5568
rect 479524 5516 479576 5568
rect 480536 5516 480588 5568
rect 207388 5448 207440 5500
rect 259644 5448 259696 5500
rect 270316 5448 270368 5500
rect 286600 5448 286652 5500
rect 300676 5448 300728 5500
rect 540796 5448 540848 5500
rect 203892 5380 203944 5432
rect 258264 5380 258316 5432
rect 270132 5380 270184 5432
rect 288992 5380 289044 5432
rect 300584 5380 300636 5432
rect 544384 5380 544436 5432
rect 200304 5312 200356 5364
rect 258356 5312 258408 5364
rect 269856 5312 269908 5364
rect 290188 5312 290240 5364
rect 300768 5312 300820 5364
rect 547880 5312 547932 5364
rect 196808 5244 196860 5296
rect 258172 5244 258224 5296
rect 270408 5244 270460 5296
rect 293684 5244 293736 5296
rect 301964 5244 302016 5296
rect 551468 5244 551520 5296
rect 193220 5176 193272 5228
rect 258080 5176 258132 5228
rect 270224 5176 270276 5228
rect 292580 5176 292632 5228
rect 302056 5176 302108 5228
rect 554964 5176 555016 5228
rect 132960 5108 133012 5160
rect 129372 5040 129424 5092
rect 250352 5108 250404 5160
rect 271420 5108 271472 5160
rect 297272 5108 297324 5160
rect 302148 5108 302200 5160
rect 558552 5108 558604 5160
rect 249984 5040 250036 5092
rect 264428 5040 264480 5092
rect 270040 5040 270092 5092
rect 296076 5040 296128 5092
rect 303344 5040 303396 5092
rect 562048 5040 562100 5092
rect 7656 4972 7708 5024
rect 234712 4972 234764 5024
rect 246396 4972 246448 5024
rect 263784 4972 263836 5024
rect 271236 4972 271288 5024
rect 300768 4972 300820 5024
rect 302792 4972 302844 5024
rect 565636 4972 565688 5024
rect 2872 4904 2924 4956
rect 234896 4904 234948 4956
rect 242900 4904 242952 4956
rect 263876 4904 263928 4956
rect 271512 4904 271564 4956
rect 299664 4904 299716 4956
rect 303252 4904 303304 4956
rect 569132 4904 569184 4956
rect 1676 4836 1728 4888
rect 234804 4836 234856 4888
rect 239312 4836 239364 4888
rect 264060 4836 264112 4888
rect 271604 4836 271656 4888
rect 303160 4836 303212 4888
rect 572 4768 624 4820
rect 234988 4768 235040 4820
rect 235908 4768 235960 4820
rect 262588 4768 262640 4820
rect 271696 4768 271748 4820
rect 304356 4768 304408 4820
rect 211068 4700 211120 4752
rect 260196 4700 260248 4752
rect 269948 4700 270000 4752
rect 285404 4700 285456 4752
rect 302700 4700 302752 4752
rect 572720 4836 572772 4888
rect 304540 4768 304592 4820
rect 576308 4768 576360 4820
rect 214472 4564 214524 4616
rect 259552 4632 259604 4684
rect 268844 4632 268896 4684
rect 283104 4632 283156 4684
rect 299204 4632 299256 4684
rect 537208 4700 537260 4752
rect 533712 4632 533764 4684
rect 228732 4564 228784 4616
rect 262404 4564 262456 4616
rect 268660 4564 268712 4616
rect 281908 4564 281960 4616
rect 299296 4564 299348 4616
rect 530124 4564 530176 4616
rect 232228 4496 232280 4548
rect 262772 4496 262824 4548
rect 268752 4496 268804 4548
rect 278320 4496 278372 4548
rect 295984 4496 296036 4548
rect 512460 4496 512512 4548
rect 298652 4428 298704 4480
rect 126980 4156 127032 4208
rect 128268 4156 128320 4208
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 143540 4156 143592 4208
rect 144828 4156 144880 4208
rect 151820 4156 151872 4208
rect 153108 4156 153160 4208
rect 160100 4156 160152 4208
rect 161388 4156 161440 4208
rect 168380 4156 168432 4208
rect 169668 4156 169720 4208
rect 184940 4156 184992 4208
rect 186228 4156 186280 4208
rect 209780 4156 209832 4208
rect 210976 4156 211028 4208
rect 218060 4156 218112 4208
rect 219348 4156 219400 4208
rect 226340 4156 226392 4208
rect 227628 4156 227680 4208
rect 237564 4156 237616 4208
rect 297364 4156 297416 4208
rect 298468 4156 298520 4208
rect 307760 4156 307812 4208
rect 309048 4156 309100 4208
rect 316040 4156 316092 4208
rect 317328 4156 317380 4208
rect 332692 4156 332744 4208
rect 333888 4156 333940 4208
rect 349160 4156 349212 4208
rect 350448 4156 350500 4208
rect 357532 4156 357584 4208
rect 358728 4156 358780 4208
rect 374000 4156 374052 4208
rect 375288 4156 375340 4208
rect 382280 4156 382332 4208
rect 383568 4156 383620 4208
rect 398840 4156 398892 4208
rect 400128 4156 400180 4208
rect 423772 4156 423824 4208
rect 424968 4156 425020 4208
rect 45376 4088 45428 4140
rect 46204 4088 46256 4140
rect 85672 4088 85724 4140
rect 244556 4088 244608 4140
rect 267372 4088 267424 4140
rect 268844 4088 268896 4140
rect 287428 4088 287480 4140
rect 443828 4088 443880 4140
rect 566464 4088 566516 4140
rect 568028 4088 568080 4140
rect 9956 4020 10008 4072
rect 18604 4020 18656 4072
rect 82084 4020 82136 4072
rect 244924 4020 244976 4072
rect 267464 4020 267516 4072
rect 267648 4020 267700 4072
rect 289544 4020 289596 4072
rect 447416 4020 447468 4072
rect 78496 3952 78548 4004
rect 244464 3952 244516 4004
rect 289636 3952 289688 4004
rect 450912 3952 450964 4004
rect 60832 3884 60884 3936
rect 62028 3884 62080 3936
rect 75000 3884 75052 3936
rect 243636 3884 243688 3936
rect 289728 3884 289780 3936
rect 454500 3884 454552 3936
rect 576124 3884 576176 3936
rect 578608 3884 578660 3936
rect 46664 3816 46716 3868
rect 240784 3816 240836 3868
rect 265440 3816 265492 3868
rect 290832 3816 290884 3868
rect 458088 3816 458140 3868
rect 43076 3748 43128 3800
rect 239036 3748 239088 3800
rect 28908 3680 28960 3732
rect 35164 3680 35216 3732
rect 39580 3680 39632 3732
rect 238852 3680 238904 3732
rect 257068 3680 257120 3732
rect 262864 3748 262916 3800
rect 265624 3748 265676 3800
rect 291108 3748 291160 3800
rect 461584 3748 461636 3800
rect 259460 3680 259512 3732
rect 265348 3680 265400 3732
rect 267556 3680 267608 3732
rect 273628 3680 273680 3732
rect 290924 3680 290976 3732
rect 465172 3680 465224 3732
rect 23020 3612 23072 3664
rect 29644 3612 29696 3664
rect 32404 3612 32456 3664
rect 5264 3476 5316 3528
rect 10324 3544 10376 3596
rect 11152 3544 11204 3596
rect 28264 3544 28316 3596
rect 33600 3544 33652 3596
rect 34428 3544 34480 3596
rect 35992 3612 36044 3664
rect 238944 3612 238996 3664
rect 262956 3612 263008 3664
rect 266544 3612 266596 3664
rect 291016 3612 291068 3664
rect 468668 3612 468720 3664
rect 238024 3544 238076 3596
rect 255872 3544 255924 3596
rect 264152 3544 264204 3596
rect 266912 3544 266964 3596
rect 292488 3544 292540 3596
rect 472256 3544 472308 3596
rect 525064 3544 525116 3596
rect 527824 3544 527876 3596
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 25320 3476 25372 3528
rect 24216 3408 24268 3460
rect 229836 3476 229888 3528
rect 230388 3476 230440 3528
rect 231032 3476 231084 3528
rect 231768 3476 231820 3528
rect 233424 3476 233476 3528
rect 234528 3476 234580 3528
rect 234620 3476 234672 3528
rect 235816 3476 235868 3528
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 241704 3476 241756 3528
rect 242808 3476 242860 3528
rect 248788 3476 248840 3528
rect 249708 3476 249760 3528
rect 254676 3476 254728 3528
rect 260656 3476 260708 3528
rect 265072 3476 265124 3528
rect 266544 3476 266596 3528
rect 267096 3476 267148 3528
rect 268384 3476 268436 3528
rect 272432 3476 272484 3528
rect 292304 3476 292356 3528
rect 239404 3408 239456 3460
rect 251180 3408 251232 3460
rect 265256 3408 265308 3460
rect 265348 3408 265400 3460
rect 266636 3408 266688 3460
rect 267280 3408 267332 3460
rect 270040 3408 270092 3460
rect 292396 3408 292448 3460
rect 473360 3476 473412 3528
rect 474556 3476 474608 3528
rect 489920 3476 489972 3528
rect 491116 3476 491168 3528
rect 522304 3476 522356 3528
rect 524236 3476 524288 3528
rect 533344 3476 533396 3528
rect 534908 3476 534960 3528
rect 556160 3476 556212 3528
rect 557356 3476 557408 3528
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 41880 3340 41932 3392
rect 43444 3340 43496 3392
rect 44272 3340 44324 3392
rect 45468 3340 45520 3392
rect 48964 3340 49016 3392
rect 49608 3340 49660 3392
rect 50160 3340 50212 3392
rect 50988 3340 51040 3392
rect 52552 3340 52604 3392
rect 53656 3340 53708 3392
rect 56048 3340 56100 3392
rect 56508 3340 56560 3392
rect 57244 3340 57296 3392
rect 57888 3340 57940 3392
rect 64328 3340 64380 3392
rect 64788 3340 64840 3392
rect 66720 3340 66772 3392
rect 67548 3340 67600 3392
rect 67916 3340 67968 3392
rect 68928 3340 68980 3392
rect 73804 3340 73856 3392
rect 74448 3340 74500 3392
rect 77392 3340 77444 3392
rect 78588 3340 78640 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 84476 3340 84528 3392
rect 85488 3340 85540 3392
rect 91560 3340 91612 3392
rect 92388 3340 92440 3392
rect 93952 3340 94004 3392
rect 95240 3340 95292 3392
rect 97448 3340 97500 3392
rect 97908 3340 97960 3392
rect 98644 3340 98696 3392
rect 99288 3340 99340 3392
rect 101036 3340 101088 3392
rect 102048 3340 102100 3392
rect 27712 3272 27764 3324
rect 33784 3272 33836 3324
rect 89168 3204 89220 3256
rect 245016 3340 245068 3392
rect 287520 3340 287572 3392
rect 440332 3340 440384 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 475752 3408 475804 3460
rect 514760 3408 514812 3460
rect 515956 3408 516008 3460
rect 479340 3340 479392 3392
rect 245844 3272 245896 3324
rect 269028 3272 269080 3324
rect 277124 3272 277176 3324
rect 288164 3272 288216 3324
rect 436744 3272 436796 3324
rect 26516 3136 26568 3188
rect 27528 3136 27580 3188
rect 92756 3136 92808 3188
rect 31300 3068 31352 3120
rect 36544 3068 36596 3120
rect 96252 3068 96304 3120
rect 246304 3204 246356 3256
rect 261760 3204 261812 3256
rect 265532 3204 265584 3256
rect 286140 3204 286192 3256
rect 433248 3204 433300 3256
rect 105728 3136 105780 3188
rect 106188 3136 106240 3188
rect 108120 3136 108172 3188
rect 108948 3136 109000 3188
rect 109316 3136 109368 3188
rect 110328 3136 110380 3188
rect 246212 3136 246264 3188
rect 268936 3136 268988 3188
rect 276020 3136 276072 3188
rect 286784 3136 286836 3188
rect 429660 3136 429712 3188
rect 103336 3068 103388 3120
rect 247500 3068 247552 3120
rect 286232 3068 286284 3120
rect 426164 3068 426216 3120
rect 19432 3000 19484 3052
rect 21364 3000 21416 3052
rect 99840 3000 99892 3052
rect 114008 3000 114060 3052
rect 114468 3000 114520 3052
rect 115204 3000 115256 3052
rect 115848 3000 115900 3052
rect 116400 3000 116452 3052
rect 117228 3000 117280 3052
rect 118792 3000 118844 3052
rect 119896 3000 119948 3052
rect 247684 3000 247736 3052
rect 284852 3000 284904 3052
rect 422576 3000 422628 3052
rect 529204 3000 529256 3052
rect 531320 3000 531372 3052
rect 59636 2932 59688 2984
rect 60648 2932 60700 2984
rect 102232 2932 102284 2984
rect 103428 2932 103480 2984
rect 110512 2932 110564 2984
rect 247224 2932 247276 2984
rect 258264 2932 258316 2984
rect 265164 2932 265216 2984
rect 284760 2932 284812 2984
rect 415492 2932 415544 2984
rect 416688 2932 416740 2984
rect 18236 2864 18288 2916
rect 22744 2864 22796 2916
rect 106924 2864 106976 2916
rect 117596 2796 117648 2848
rect 122288 2864 122340 2916
rect 122748 2864 122800 2916
rect 123484 2864 123536 2916
rect 124128 2864 124180 2916
rect 124680 2864 124732 2916
rect 125508 2864 125560 2916
rect 125876 2864 125928 2916
rect 126888 2864 126940 2916
rect 121092 2796 121144 2848
rect 249064 2864 249116 2916
rect 285496 2864 285548 2916
rect 418988 2864 419040 2916
rect 249156 2796 249208 2848
rect 285312 2796 285364 2848
rect 407120 2796 407172 2848
rect 408408 2796 408460 2848
rect 411904 2796 411956 2848
rect 415492 2796 415544 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 696998 3464 697303
rect 3424 696992 3476 696998
rect 3424 696934 3476 696940
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3330 645144 3386 645153
rect 3330 645079 3386 645088
rect 3344 644502 3372 645079
rect 3332 644496 3384 644502
rect 3332 644438 3384 644444
rect 2778 619168 2834 619177
rect 2778 619103 2780 619112
rect 2832 619103 2834 619112
rect 2780 619074 2832 619080
rect 2962 593056 3018 593065
rect 2962 592991 3018 593000
rect 2976 592074 3004 592991
rect 2964 592068 3016 592074
rect 2964 592010 3016 592016
rect 2870 540832 2926 540841
rect 2870 540767 2926 540776
rect 2884 539646 2912 540767
rect 2872 539640 2924 539646
rect 2872 539582 2924 539588
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3238 488744 3294 488753
rect 3238 488679 3294 488688
rect 3146 475688 3202 475697
rect 3146 475623 3202 475632
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 2962 449576 3018 449585
rect 2962 449511 3018 449520
rect 2870 436656 2926 436665
rect 2870 436591 2926 436600
rect 2778 423600 2834 423609
rect 2778 423535 2834 423544
rect 2792 380866 2820 423535
rect 2884 382226 2912 436591
rect 2976 383654 3004 449511
rect 3068 385014 3096 462567
rect 3160 386374 3188 475623
rect 3252 387802 3280 488679
rect 3344 389162 3372 501735
rect 3436 410666 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 410786 3556 658135
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3516 410780 3568 410786
rect 3516 410722 3568 410728
rect 3436 410638 3556 410666
rect 3422 410544 3478 410553
rect 3422 410479 3424 410488
rect 3476 410479 3478 410488
rect 3424 410450 3476 410456
rect 3424 410372 3476 410378
rect 3424 410314 3476 410320
rect 3436 404326 3464 410314
rect 3528 405686 3556 410638
rect 3516 405680 3568 405686
rect 3516 405622 3568 405628
rect 3424 404320 3476 404326
rect 3424 404262 3476 404268
rect 3620 401606 3648 632023
rect 4804 619132 4856 619138
rect 4804 619074 4856 619080
rect 3698 606112 3754 606121
rect 3698 606047 3754 606056
rect 3608 401600 3660 401606
rect 3608 401542 3660 401548
rect 3712 398818 3740 606047
rect 3790 580000 3846 580009
rect 3790 579935 3846 579944
rect 3700 398812 3752 398818
rect 3700 398754 3752 398760
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3332 389156 3384 389162
rect 3332 389098 3384 389104
rect 3240 387796 3292 387802
rect 3240 387738 3292 387744
rect 3148 386368 3200 386374
rect 3148 386310 3200 386316
rect 3056 385008 3108 385014
rect 3056 384950 3108 384956
rect 2964 383648 3016 383654
rect 2964 383590 3016 383596
rect 2872 382220 2924 382226
rect 2872 382162 2924 382168
rect 2780 380860 2832 380866
rect 2780 380802 2832 380808
rect 3436 378146 3464 397423
rect 3804 396030 3832 579935
rect 3882 566944 3938 566953
rect 3882 566879 3938 566888
rect 3792 396024 3844 396030
rect 3792 395966 3844 395972
rect 3896 394670 3924 566879
rect 3974 553888 4030 553897
rect 3974 553823 4030 553832
rect 3884 394664 3936 394670
rect 3884 394606 3936 394612
rect 3988 393310 4016 553823
rect 4066 527912 4122 527921
rect 4066 527847 4122 527856
rect 3976 393304 4028 393310
rect 3976 393246 4028 393252
rect 4080 390522 4108 527847
rect 4816 400178 4844 619074
rect 8220 410582 8248 702406
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 10324 514820 10376 514826
rect 10324 514762 10376 514768
rect 8208 410576 8260 410582
rect 8208 410518 8260 410524
rect 7564 410508 7616 410514
rect 7564 410450 7616 410456
rect 4804 400172 4856 400178
rect 4804 400114 4856 400120
rect 4068 390516 4120 390522
rect 4068 390458 4120 390464
rect 3514 384432 3570 384441
rect 3514 384367 3570 384376
rect 3424 378140 3476 378146
rect 3424 378082 3476 378088
rect 3528 376718 3556 384367
rect 7576 379506 7604 410450
rect 10336 389094 10364 514762
rect 24780 410650 24808 699654
rect 41340 410718 41368 700334
rect 56796 700194 56824 703520
rect 72988 702434 73016 703520
rect 72988 702406 73108 702434
rect 56784 700188 56836 700194
rect 56784 700130 56836 700136
rect 57888 700188 57940 700194
rect 57888 700130 57940 700136
rect 57900 410786 57928 700130
rect 73080 410854 73108 702406
rect 89180 699718 89208 703520
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 89640 410922 89668 699654
rect 106200 410990 106228 700334
rect 121656 699718 121684 703520
rect 137848 702434 137876 703520
rect 154132 702434 154160 703520
rect 137848 702406 137968 702434
rect 154132 702406 154528 702434
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 122748 699712 122800 699718
rect 122748 699654 122800 699660
rect 122760 411058 122788 699654
rect 137940 411126 137968 702406
rect 154500 411194 154528 702406
rect 170324 699718 170352 703520
rect 186516 700194 186544 703520
rect 186504 700188 186556 700194
rect 186504 700130 186556 700136
rect 187608 700188 187660 700194
rect 187608 700130 187660 700136
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 171060 411262 171088 699654
rect 184204 696992 184256 696998
rect 184204 696934 184256 696940
rect 171048 411256 171100 411262
rect 171048 411198 171100 411204
rect 154488 411188 154540 411194
rect 154488 411130 154540 411136
rect 137928 411120 137980 411126
rect 137928 411062 137980 411068
rect 122748 411052 122800 411058
rect 122748 410994 122800 411000
rect 106188 410984 106240 410990
rect 106188 410926 106240 410932
rect 89628 410916 89680 410922
rect 89628 410858 89680 410864
rect 73068 410848 73120 410854
rect 73068 410790 73120 410796
rect 57888 410780 57940 410786
rect 57888 410722 57940 410728
rect 41328 410712 41380 410718
rect 41328 410654 41380 410660
rect 24768 410644 24820 410650
rect 24768 410586 24820 410592
rect 184216 408474 184244 696934
rect 187620 410514 187648 700130
rect 195244 644496 195296 644502
rect 195244 644438 195296 644444
rect 187608 410508 187660 410514
rect 187608 410450 187660 410456
rect 184204 408468 184256 408474
rect 184204 408410 184256 408416
rect 195256 402966 195284 644438
rect 198004 592068 198056 592074
rect 198004 592010 198056 592016
rect 195244 402960 195296 402966
rect 195244 402902 195296 402908
rect 198016 397458 198044 592010
rect 202800 410446 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 410440 202840 410446
rect 202788 410382 202840 410388
rect 219360 410378 219388 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 235908 700392 235960 700398
rect 235908 700334 235960 700340
rect 220084 539640 220136 539646
rect 220084 539582 220136 539588
rect 219348 410372 219400 410378
rect 219348 410314 219400 410320
rect 198004 397452 198056 397458
rect 198004 397394 198056 397400
rect 220096 391950 220124 539582
rect 235920 410582 235948 700334
rect 251468 700126 251496 703520
rect 251456 700120 251508 700126
rect 251456 700062 251508 700068
rect 252468 700120 252520 700126
rect 252468 700062 252520 700068
rect 251180 411120 251232 411126
rect 251180 411062 251232 411068
rect 249156 411052 249208 411058
rect 249156 410994 249208 411000
rect 247224 410984 247276 410990
rect 247224 410926 247276 410932
rect 245292 410916 245344 410922
rect 245292 410858 245344 410864
rect 243360 410848 243412 410854
rect 243360 410790 243412 410796
rect 241520 410780 241572 410786
rect 241520 410722 241572 410728
rect 239496 410712 239548 410718
rect 239496 410654 239548 410660
rect 237564 410644 237616 410650
rect 237564 410586 237616 410592
rect 235632 410576 235684 410582
rect 235632 410518 235684 410524
rect 235908 410576 235960 410582
rect 235908 410518 235960 410524
rect 232044 408468 232096 408474
rect 232044 408410 232096 408416
rect 232056 407289 232084 408410
rect 235644 407946 235672 410518
rect 237576 407946 237604 410586
rect 239508 407946 239536 410654
rect 241532 407946 241560 410722
rect 243372 407946 243400 410790
rect 245304 407946 245332 410858
rect 247236 407946 247264 410926
rect 249168 407946 249196 410994
rect 251192 407946 251220 411062
rect 252480 410650 252508 700062
rect 267660 699718 267688 703520
rect 283852 700398 283880 703520
rect 285588 701004 285640 701010
rect 285588 700946 285640 700952
rect 269028 700392 269080 700398
rect 269028 700334 269080 700340
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 266360 699712 266412 699718
rect 266360 699654 266412 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 266372 422294 266400 699654
rect 266372 422266 266676 422294
rect 255320 411256 255372 411262
rect 255320 411198 255372 411204
rect 253112 411188 253164 411194
rect 253112 411130 253164 411136
rect 252468 410644 252520 410650
rect 252468 410586 252520 410592
rect 253124 407946 253152 411130
rect 255332 407946 255360 411198
rect 264980 410644 265032 410650
rect 264980 410586 265032 410592
rect 262772 410576 262824 410582
rect 262772 410518 262824 410524
rect 256976 410508 257028 410514
rect 256976 410450 257028 410456
rect 256988 407946 257016 410450
rect 258908 410440 258960 410446
rect 258908 410382 258960 410388
rect 258920 407946 258948 410382
rect 260840 410372 260892 410378
rect 260840 410314 260892 410320
rect 260852 407946 260880 410314
rect 262784 407946 262812 410518
rect 264992 407946 265020 410586
rect 266648 407946 266676 422266
rect 269040 408218 269068 700334
rect 271788 700324 271840 700330
rect 271788 700266 271840 700272
rect 271800 409970 271828 700266
rect 282828 700256 282880 700262
rect 282828 700198 282880 700204
rect 281448 700188 281500 700194
rect 281448 700130 281500 700136
rect 278688 700120 278740 700126
rect 278688 700062 278740 700068
rect 277308 700052 277360 700058
rect 277308 699994 277360 700000
rect 275928 699984 275980 699990
rect 275928 699926 275980 699932
rect 273168 699916 273220 699922
rect 273168 699858 273220 699864
rect 271236 409964 271288 409970
rect 271236 409906 271288 409912
rect 271788 409964 271840 409970
rect 271788 409906 271840 409912
rect 268994 408190 269068 408218
rect 235644 407918 235980 407946
rect 237576 407918 237912 407946
rect 239508 407918 239844 407946
rect 241532 407918 241776 407946
rect 243372 407918 243708 407946
rect 245304 407918 245640 407946
rect 247236 407918 247572 407946
rect 249168 407918 249504 407946
rect 251192 407918 251528 407946
rect 253124 407918 253460 407946
rect 255332 407918 255392 407946
rect 256988 407918 257324 407946
rect 258920 407918 259256 407946
rect 260852 407918 261188 407946
rect 262784 407918 263120 407946
rect 264992 407918 265144 407946
rect 266648 407918 267076 407946
rect 268994 407932 269022 408190
rect 271248 407946 271276 409906
rect 273180 407946 273208 699858
rect 275940 409970 275968 699926
rect 277320 412634 277348 699994
rect 277136 412606 277348 412634
rect 275100 409964 275152 409970
rect 275100 409906 275152 409912
rect 275928 409964 275980 409970
rect 275928 409906 275980 409912
rect 275112 407946 275140 409906
rect 277136 407946 277164 412606
rect 270940 407918 271276 407946
rect 272872 407918 273208 407946
rect 274804 407918 275140 407946
rect 276736 407918 277164 407946
rect 278700 407946 278728 700062
rect 281460 409970 281488 700130
rect 280988 409964 281040 409970
rect 280988 409906 281040 409912
rect 281448 409964 281500 409970
rect 281448 409906 281500 409912
rect 281000 407946 281028 409906
rect 282840 407946 282868 700198
rect 285600 409970 285628 700946
rect 286968 700936 287020 700942
rect 286968 700878 287020 700884
rect 286980 412634 287008 700878
rect 288348 700868 288400 700874
rect 288348 700810 288400 700816
rect 286888 412606 287008 412634
rect 284852 409964 284904 409970
rect 284852 409906 284904 409912
rect 285588 409964 285640 409970
rect 285588 409906 285640 409912
rect 284864 407946 284892 409906
rect 286888 407946 286916 412606
rect 278700 407918 278760 407946
rect 280692 407918 281028 407946
rect 282624 407918 282868 407946
rect 284556 407918 284892 407946
rect 286488 407918 286916 407946
rect 288360 407946 288388 700810
rect 291108 700800 291160 700806
rect 291108 700742 291160 700748
rect 291120 409970 291148 700742
rect 292488 700732 292540 700738
rect 292488 700674 292540 700680
rect 290648 409964 290700 409970
rect 290648 409906 290700 409912
rect 291108 409964 291160 409970
rect 291108 409906 291160 409912
rect 290660 407946 290688 409906
rect 292500 407946 292528 700674
rect 295248 700664 295300 700670
rect 295248 700606 295300 700612
rect 295260 409970 295288 700606
rect 296628 700596 296680 700602
rect 296628 700538 296680 700544
rect 294604 409964 294656 409970
rect 294604 409906 294656 409912
rect 295248 409964 295300 409970
rect 295248 409906 295300 409912
rect 294616 407946 294644 409906
rect 296640 407946 296668 700538
rect 299388 700528 299440 700534
rect 299388 700470 299440 700476
rect 299400 409970 299428 700470
rect 300136 700330 300164 703520
rect 300768 700460 300820 700466
rect 300768 700402 300820 700408
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 300780 412634 300808 700402
rect 302148 700392 302200 700398
rect 302148 700334 302200 700340
rect 300504 412606 300808 412634
rect 298468 409964 298520 409970
rect 298468 409906 298520 409912
rect 299388 409964 299440 409970
rect 299388 409906 299440 409912
rect 298480 407946 298508 409906
rect 300504 407946 300532 412606
rect 302160 407946 302188 700334
rect 304908 700324 304960 700330
rect 304908 700266 304960 700272
rect 304920 409970 304948 700266
rect 316328 699922 316356 703520
rect 332520 699990 332548 703520
rect 348804 700058 348832 703520
rect 364996 700126 365024 703520
rect 381188 700194 381216 703520
rect 397472 700262 397500 703520
rect 413664 701010 413692 703520
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 429856 700942 429884 703520
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 446140 700874 446168 703520
rect 446128 700868 446180 700874
rect 446128 700810 446180 700816
rect 462332 700806 462360 703520
rect 462320 700800 462372 700806
rect 462320 700742 462372 700748
rect 478524 700738 478552 703520
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 511000 700602 511028 703520
rect 510988 700596 511040 700602
rect 510988 700538 511040 700544
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 575860 700330 575888 703520
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 381176 700188 381228 700194
rect 381176 700130 381228 700136
rect 364984 700120 365036 700126
rect 364984 700062 365036 700068
rect 348792 700052 348844 700058
rect 348792 699994 348844 700000
rect 332508 699984 332560 699990
rect 332508 699926 332560 699932
rect 316316 699916 316368 699922
rect 316316 699858 316368 699864
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 307024 696992 307076 696998
rect 307024 696934 307076 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 306932 484424 306984 484430
rect 306932 484366 306984 484372
rect 306840 470620 306892 470626
rect 306840 470562 306892 470568
rect 306748 430636 306800 430642
rect 306748 430578 306800 430584
rect 304264 409964 304316 409970
rect 304264 409906 304316 409912
rect 304908 409964 304960 409970
rect 304908 409906 304960 409912
rect 304276 407946 304304 409906
rect 288360 407918 288420 407946
rect 290352 407918 290688 407946
rect 292376 407918 292528 407946
rect 294308 407918 294644 407946
rect 296240 407918 296668 407946
rect 298172 407918 298508 407946
rect 300104 407918 300532 407946
rect 302036 407918 302188 407946
rect 303968 407918 304304 407946
rect 232042 407280 232098 407289
rect 232042 407215 232098 407224
rect 232044 405680 232096 405686
rect 232044 405622 232096 405628
rect 232056 404705 232084 405622
rect 232042 404696 232098 404705
rect 232042 404631 232098 404640
rect 232044 404320 232096 404326
rect 232044 404262 232096 404268
rect 232056 403345 232084 404262
rect 232042 403336 232098 403345
rect 232042 403271 232098 403280
rect 232044 402960 232096 402966
rect 232044 402902 232096 402908
rect 232056 402121 232084 402902
rect 232042 402112 232098 402121
rect 232042 402047 232098 402056
rect 232044 401600 232096 401606
rect 232044 401542 232096 401548
rect 232056 400761 232084 401542
rect 232042 400752 232098 400761
rect 232042 400687 232098 400696
rect 232044 400172 232096 400178
rect 232044 400114 232096 400120
rect 232056 399537 232084 400114
rect 232042 399528 232098 399537
rect 232042 399463 232098 399472
rect 232044 398812 232096 398818
rect 232044 398754 232096 398760
rect 232056 398177 232084 398754
rect 232042 398168 232098 398177
rect 232042 398103 232098 398112
rect 232044 397452 232096 397458
rect 232044 397394 232096 397400
rect 232056 396953 232084 397394
rect 232042 396944 232098 396953
rect 232042 396879 232098 396888
rect 232044 396024 232096 396030
rect 232044 395966 232096 395972
rect 232056 395593 232084 395966
rect 232042 395584 232098 395593
rect 232042 395519 232098 395528
rect 231952 394664 232004 394670
rect 231952 394606 232004 394612
rect 231964 394369 231992 394606
rect 231950 394360 232006 394369
rect 231950 394295 232006 394304
rect 232044 393304 232096 393310
rect 232044 393246 232096 393252
rect 232056 393009 232084 393246
rect 232042 393000 232098 393009
rect 232042 392935 232098 392944
rect 220084 391944 220136 391950
rect 220084 391886 220136 391892
rect 232044 391944 232096 391950
rect 232044 391886 232096 391892
rect 232056 391785 232084 391886
rect 232042 391776 232098 391785
rect 232042 391711 232098 391720
rect 232044 390516 232096 390522
rect 232044 390458 232096 390464
rect 232056 390425 232084 390458
rect 232042 390416 232098 390425
rect 232042 390351 232098 390360
rect 231952 389156 232004 389162
rect 231952 389098 232004 389104
rect 10324 389088 10376 389094
rect 10324 389030 10376 389036
rect 231964 387841 231992 389098
rect 232044 389088 232096 389094
rect 232042 389056 232044 389065
rect 232096 389056 232098 389065
rect 232042 388991 232098 389000
rect 231950 387832 232006 387841
rect 231950 387767 232006 387776
rect 232044 387796 232096 387802
rect 232044 387738 232096 387744
rect 232056 386481 232084 387738
rect 232042 386472 232098 386481
rect 232042 386407 232098 386416
rect 232044 386368 232096 386374
rect 232044 386310 232096 386316
rect 232056 385257 232084 386310
rect 232042 385248 232098 385257
rect 232042 385183 232098 385192
rect 232044 385008 232096 385014
rect 232044 384950 232096 384956
rect 232056 383897 232084 384950
rect 232042 383888 232098 383897
rect 232042 383823 232098 383832
rect 231860 383648 231912 383654
rect 231860 383590 231912 383596
rect 231872 382673 231900 383590
rect 231858 382664 231914 382673
rect 231858 382599 231914 382608
rect 232044 382220 232096 382226
rect 232044 382162 232096 382168
rect 232056 381313 232084 382162
rect 232042 381304 232098 381313
rect 232042 381239 232098 381248
rect 306760 380905 306788 430578
rect 306852 384985 306880 470562
rect 306944 386209 306972 484366
rect 307036 407833 307064 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 307116 683188 307168 683194
rect 307116 683130 307168 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 307022 407824 307078 407833
rect 307022 407759 307078 407768
rect 307128 406473 307156 683130
rect 307208 670744 307260 670750
rect 580172 670744 580224 670750
rect 307208 670686 307260 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 307114 406464 307170 406473
rect 307114 406399 307170 406408
rect 307220 405113 307248 670686
rect 580170 670647 580226 670656
rect 580262 657384 580318 657393
rect 580262 657319 580318 657328
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 307300 643136 307352 643142
rect 307300 643078 307352 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 307206 405104 307262 405113
rect 307206 405039 307262 405048
rect 307024 404388 307076 404394
rect 307024 404330 307076 404336
rect 306930 386200 306986 386209
rect 306930 386135 306986 386144
rect 306838 384976 306894 384985
rect 306838 384911 306894 384920
rect 306746 380896 306802 380905
rect 232044 380860 232096 380866
rect 306746 380831 306802 380840
rect 306840 380860 306892 380866
rect 232044 380802 232096 380808
rect 306840 380802 306892 380808
rect 232056 380089 232084 380802
rect 306852 380089 306880 380802
rect 232042 380080 232098 380089
rect 232042 380015 232098 380024
rect 306838 380080 306894 380089
rect 306838 380015 306894 380024
rect 7564 379500 7616 379506
rect 7564 379442 7616 379448
rect 232044 379500 232096 379506
rect 232044 379442 232096 379448
rect 232056 378729 232084 379442
rect 307036 378729 307064 404330
rect 307208 404320 307260 404326
rect 307208 404262 307260 404268
rect 307220 403889 307248 404262
rect 307206 403880 307262 403889
rect 307206 403815 307262 403824
rect 307312 402529 307340 643078
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 309784 630692 309836 630698
rect 309784 630634 309836 630640
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 307392 590708 307444 590714
rect 307392 590650 307444 590656
rect 307298 402520 307354 402529
rect 307298 402455 307354 402464
rect 307300 401328 307352 401334
rect 307300 401270 307352 401276
rect 307312 401169 307340 401270
rect 307298 401160 307354 401169
rect 307298 401095 307354 401104
rect 307208 400172 307260 400178
rect 307208 400114 307260 400120
rect 307220 399673 307248 400114
rect 307206 399664 307262 399673
rect 307206 399599 307262 399608
rect 307300 398948 307352 398954
rect 307300 398890 307352 398896
rect 307312 395729 307340 398890
rect 307404 397225 307432 590650
rect 307484 576904 307536 576910
rect 307484 576846 307536 576852
rect 307496 398954 307524 576846
rect 307576 536852 307628 536858
rect 307576 536794 307628 536800
rect 307484 398948 307536 398954
rect 307484 398890 307536 398896
rect 307484 398812 307536 398818
rect 307484 398754 307536 398760
rect 307496 398449 307524 398754
rect 307482 398440 307538 398449
rect 307482 398375 307538 398384
rect 307390 397216 307446 397225
rect 307390 397151 307446 397160
rect 307298 395720 307354 395729
rect 307298 395655 307354 395664
rect 307484 394664 307536 394670
rect 307484 394606 307536 394612
rect 307496 394369 307524 394606
rect 307482 394360 307538 394369
rect 307482 394295 307538 394304
rect 307484 393304 307536 393310
rect 307484 393246 307536 393252
rect 307496 393009 307524 393246
rect 307482 393000 307538 393009
rect 307482 392935 307538 392944
rect 307588 391921 307616 536794
rect 307668 524476 307720 524482
rect 307668 524418 307720 524424
rect 307574 391912 307630 391921
rect 307574 391847 307630 391856
rect 307116 390584 307168 390590
rect 307680 390561 307708 524418
rect 309796 401334 309824 630634
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579986 577688 580042 577697
rect 579986 577623 580042 577632
rect 580000 576910 580028 577623
rect 579988 576904 580040 576910
rect 579988 576846 580040 576852
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580078 431624 580134 431633
rect 580078 431559 580134 431568
rect 580092 430642 580120 431559
rect 580080 430636 580132 430642
rect 580080 430578 580132 430584
rect 580078 418296 580134 418305
rect 580078 418231 580134 418240
rect 580092 418198 580120 418231
rect 312544 418192 312596 418198
rect 312544 418134 312596 418140
rect 580080 418192 580132 418198
rect 580080 418134 580132 418140
rect 309784 401328 309836 401334
rect 309784 401270 309836 401276
rect 307116 390526 307168 390532
rect 307666 390552 307722 390561
rect 232042 378720 232098 378729
rect 232042 378655 232098 378664
rect 307022 378720 307078 378729
rect 307022 378655 307078 378664
rect 232044 378140 232096 378146
rect 232044 378082 232096 378088
rect 232056 377505 232084 378082
rect 232042 377496 232098 377505
rect 232042 377431 232098 377440
rect 307128 377369 307156 390526
rect 307666 390487 307722 390496
rect 307668 389156 307720 389162
rect 307668 389098 307720 389104
rect 307680 388929 307708 389098
rect 307666 388920 307722 388929
rect 307666 388855 307722 388864
rect 307668 387796 307720 387802
rect 307668 387738 307720 387744
rect 307680 387569 307708 387738
rect 307666 387560 307722 387569
rect 307666 387495 307722 387504
rect 307668 383648 307720 383654
rect 307666 383616 307668 383625
rect 307720 383616 307722 383625
rect 307666 383551 307722 383560
rect 307666 382256 307722 382265
rect 307666 382191 307668 382200
rect 307720 382191 307722 382200
rect 307668 382162 307720 382168
rect 312556 380866 312584 418134
rect 580078 404968 580134 404977
rect 580078 404903 580134 404912
rect 580092 404394 580120 404903
rect 580080 404388 580132 404394
rect 580080 404330 580132 404336
rect 580080 404252 580132 404258
rect 580080 404194 580132 404200
rect 580092 398818 580120 404194
rect 580080 398812 580132 398818
rect 580080 398754 580132 398760
rect 580078 391776 580134 391785
rect 580078 391711 580134 391720
rect 580092 390590 580120 391711
rect 580080 390584 580132 390590
rect 580080 390526 580132 390532
rect 580184 382226 580212 444751
rect 580276 404326 580304 657319
rect 580354 617536 580410 617545
rect 580354 617471 580410 617480
rect 580264 404320 580316 404326
rect 580264 404262 580316 404268
rect 580368 400178 580396 617471
rect 580446 604208 580502 604217
rect 580446 604143 580502 604152
rect 580460 404258 580488 604143
rect 580538 564360 580594 564369
rect 580538 564295 580594 564304
rect 580448 404252 580500 404258
rect 580448 404194 580500 404200
rect 580356 400172 580408 400178
rect 580356 400114 580408 400120
rect 580552 394670 580580 564295
rect 580630 551168 580686 551177
rect 580630 551103 580686 551112
rect 580540 394664 580592 394670
rect 580540 394606 580592 394612
rect 580644 393310 580672 551103
rect 580722 511320 580778 511329
rect 580722 511255 580778 511264
rect 580632 393304 580684 393310
rect 580632 393246 580684 393252
rect 580736 389162 580764 511255
rect 580814 497992 580870 498001
rect 580814 497927 580870 497936
rect 580724 389156 580776 389162
rect 580724 389098 580776 389104
rect 580828 387802 580856 497927
rect 580906 458144 580962 458153
rect 580906 458079 580962 458088
rect 580816 387796 580868 387802
rect 580816 387738 580868 387744
rect 580920 383654 580948 458079
rect 580908 383648 580960 383654
rect 580908 383590 580960 383596
rect 580172 382220 580224 382226
rect 580172 382162 580224 382168
rect 312544 380860 312596 380866
rect 312544 380802 312596 380808
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 307668 378208 307720 378214
rect 307668 378150 307720 378156
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 307114 377360 307170 377369
rect 307114 377295 307170 377304
rect 3516 376712 3568 376718
rect 3516 376654 3568 376660
rect 232044 376712 232096 376718
rect 232044 376654 232096 376660
rect 232056 376145 232084 376654
rect 307680 376145 307708 378150
rect 232042 376136 232098 376145
rect 232042 376071 232098 376080
rect 307666 376136 307722 376145
rect 307666 376071 307722 376080
rect 232042 374912 232098 374921
rect 232042 374847 232098 374856
rect 232056 374066 232084 374847
rect 307114 374096 307170 374105
rect 3516 374060 3568 374066
rect 3516 374002 3568 374008
rect 232044 374060 232096 374066
rect 307114 374031 307170 374040
rect 232044 374002 232096 374008
rect 3528 371385 3556 374002
rect 232042 373552 232098 373561
rect 232042 373487 232098 373496
rect 232056 372638 232084 373487
rect 307022 372736 307078 372745
rect 307022 372671 307078 372680
rect 3608 372632 3660 372638
rect 3608 372574 3660 372580
rect 232044 372632 232096 372638
rect 232044 372574 232096 372580
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3148 367124 3200 367130
rect 3148 367066 3200 367072
rect 3056 332580 3108 332586
rect 3056 332522 3108 332528
rect 3068 332353 3096 332522
rect 3054 332344 3110 332353
rect 3054 332279 3110 332288
rect 3056 320136 3108 320142
rect 3056 320078 3108 320084
rect 3068 319297 3096 320078
rect 3054 319288 3110 319297
rect 3054 319223 3110 319232
rect 3160 306241 3188 367066
rect 3240 361616 3292 361622
rect 3240 361558 3292 361564
rect 3146 306232 3202 306241
rect 3146 306167 3202 306176
rect 3148 293208 3200 293214
rect 3146 293176 3148 293185
rect 3200 293176 3202 293185
rect 3146 293111 3202 293120
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3252 241097 3280 361558
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3240 229084 3292 229090
rect 3240 229026 3292 229032
rect 3252 228041 3280 229026
rect 3238 228032 3294 228041
rect 3238 227967 3294 227976
rect 3240 215280 3292 215286
rect 3240 215222 3292 215228
rect 3252 214985 3280 215222
rect 3238 214976 3294 214985
rect 3238 214911 3294 214920
rect 3344 201929 3372 357410
rect 3436 345409 3464 371214
rect 3620 358465 3648 372574
rect 232042 372192 232098 372201
rect 232042 372127 232098 372136
rect 232056 371278 232084 372127
rect 232044 371272 232096 371278
rect 232044 371214 232096 371220
rect 233146 370968 233202 370977
rect 233146 370903 233202 370912
rect 233054 369608 233110 369617
rect 233054 369543 233110 369552
rect 232042 368384 232098 368393
rect 232042 368319 232098 368328
rect 232056 367130 232084 368319
rect 232044 367124 232096 367130
rect 232044 367066 232096 367072
rect 232042 367024 232098 367033
rect 232042 366959 232098 366968
rect 232056 365770 232084 366959
rect 232778 365800 232834 365809
rect 7564 365764 7616 365770
rect 7564 365706 7616 365712
rect 232044 365764 232096 365770
rect 232778 365735 232834 365744
rect 232044 365706 232096 365712
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 4068 353320 4120 353326
rect 4068 353262 4120 353268
rect 3976 350600 4028 350606
rect 3976 350542 4028 350548
rect 3884 347812 3936 347818
rect 3884 347754 3936 347760
rect 3792 346452 3844 346458
rect 3792 346394 3844 346400
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3700 343664 3752 343670
rect 3700 343606 3752 343612
rect 3608 342304 3660 342310
rect 3608 342246 3660 342252
rect 3516 340944 3568 340950
rect 3516 340886 3568 340892
rect 3424 339516 3476 339522
rect 3424 339458 3476 339464
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3332 176656 3384 176662
rect 3332 176598 3384 176604
rect 3344 175953 3372 176598
rect 3330 175944 3386 175953
rect 3330 175879 3386 175888
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3148 124160 3200 124166
rect 3148 124102 3200 124108
rect 3160 123729 3188 124102
rect 3146 123720 3202 123729
rect 3146 123655 3202 123664
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 2872 59356 2924 59362
rect 2872 59298 2924 59304
rect 2884 58585 2912 59298
rect 2870 58576 2926 58585
rect 2870 58511 2926 58520
rect 3436 19417 3464 339458
rect 3528 32473 3556 340886
rect 3620 45529 3648 342246
rect 3712 71641 3740 343606
rect 3804 97617 3832 346394
rect 3896 110673 3924 347754
rect 3988 136785 4016 350542
rect 4080 162897 4108 353262
rect 7576 293214 7604 365706
rect 232686 364440 232742 364449
rect 232686 364375 232742 364384
rect 232042 363216 232098 363225
rect 232042 363151 232098 363160
rect 232056 362982 232084 363151
rect 22836 362976 22888 362982
rect 22836 362918 22888 362924
rect 232044 362976 232096 362982
rect 232044 362918 232096 362924
rect 14556 356108 14608 356114
rect 14556 356050 14608 356056
rect 10324 336048 10376 336054
rect 10324 335990 10376 335996
rect 7564 293208 7616 293214
rect 7564 293150 7616 293156
rect 4066 162888 4122 162897
rect 4066 162823 4122 162832
rect 3974 136776 4030 136785
rect 3974 136711 4030 136720
rect 3882 110664 3938 110673
rect 3882 110599 3938 110608
rect 3790 97608 3846 97617
rect 3790 97543 3846 97552
rect 3698 71632 3754 71641
rect 3698 71567 3754 71576
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 9588 10328 9640 10334
rect 9588 10270 9640 10276
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 8910
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 480 5304 3470
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 9600 3534 9628 10270
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 8772 480 8800 3470
rect 9968 480 9996 4014
rect 10336 3602 10364 335990
rect 14464 323604 14516 323610
rect 14464 323546 14516 323552
rect 12348 7608 12400 7614
rect 12348 7550 12400 7556
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 480 11192 3538
rect 12360 480 12388 7550
rect 14476 3534 14504 323546
rect 14568 189038 14596 356050
rect 15844 345092 15896 345098
rect 15844 345034 15896 345040
rect 14556 189032 14608 189038
rect 14556 188974 14608 188980
rect 15856 85542 15884 345034
rect 17224 338156 17276 338162
rect 17224 338098 17276 338104
rect 15844 85536 15896 85542
rect 15844 85478 15896 85484
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14738 3496 14794 3505
rect 13556 480 13584 3470
rect 14738 3431 14794 3440
rect 14752 480 14780 3431
rect 15948 480 15976 3567
rect 17052 480 17080 8978
rect 17236 6866 17264 338098
rect 21364 336184 21416 336190
rect 21364 336126 21416 336132
rect 18604 336116 18656 336122
rect 18604 336058 18656 336064
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 18616 4078 18644 336058
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 20626 3768 20682 3777
rect 20626 3703 20682 3712
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18248 480 18276 2858
rect 19444 480 19472 2994
rect 20640 480 20668 3703
rect 21376 3058 21404 336126
rect 22744 311160 22796 311166
rect 22744 311102 22796 311108
rect 21824 10396 21876 10402
rect 21824 10338 21876 10344
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21836 480 21864 10338
rect 22756 2922 22784 311102
rect 22848 255270 22876 362918
rect 232042 361856 232098 361865
rect 232042 361791 232098 361800
rect 232056 361622 232084 361791
rect 232044 361616 232096 361622
rect 232044 361558 232096 361564
rect 232594 360632 232650 360641
rect 232594 360567 232650 360576
rect 232608 359394 232636 360567
rect 232700 359530 232728 364375
rect 232792 364334 232820 365735
rect 232792 364306 233004 364334
rect 232700 359502 232912 359530
rect 232608 359366 232820 359394
rect 232686 359272 232742 359281
rect 232686 359207 232742 359216
rect 232042 358048 232098 358057
rect 232042 357983 232098 357992
rect 232056 357474 232084 357983
rect 232044 357468 232096 357474
rect 232044 357410 232096 357416
rect 232042 356688 232098 356697
rect 232042 356623 232098 356632
rect 232056 356114 232084 356623
rect 232044 356108 232096 356114
rect 232044 356050 232096 356056
rect 232594 355328 232650 355337
rect 232594 355263 232650 355272
rect 232042 354104 232098 354113
rect 232042 354039 232098 354048
rect 232056 353326 232084 354039
rect 232044 353320 232096 353326
rect 232044 353262 232096 353268
rect 232042 352744 232098 352753
rect 232042 352679 232098 352688
rect 232056 351966 232084 352679
rect 25504 351960 25556 351966
rect 25504 351902 25556 351908
rect 232044 351960 232096 351966
rect 232044 351902 232096 351908
rect 22836 255264 22888 255270
rect 22836 255206 22888 255212
rect 25516 150414 25544 351902
rect 232042 351520 232098 351529
rect 232042 351455 232098 351464
rect 232056 350606 232084 351455
rect 232044 350600 232096 350606
rect 232044 350542 232096 350548
rect 232502 350160 232558 350169
rect 232502 350095 232558 350104
rect 232042 348936 232098 348945
rect 232042 348871 232098 348880
rect 232056 347818 232084 348871
rect 232044 347812 232096 347818
rect 232044 347754 232096 347760
rect 232042 347576 232098 347585
rect 232042 347511 232098 347520
rect 232056 346458 232084 347511
rect 232044 346452 232096 346458
rect 232044 346394 232096 346400
rect 232042 346352 232098 346361
rect 232042 346287 232098 346296
rect 232056 345098 232084 346287
rect 232044 345092 232096 345098
rect 232044 345034 232096 345040
rect 231858 344992 231914 345001
rect 231858 344927 231914 344936
rect 32404 343732 32456 343738
rect 32404 343674 32456 343680
rect 28264 336252 28316 336258
rect 28264 336194 28316 336200
rect 25504 150408 25556 150414
rect 25504 150350 25556 150356
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 23032 480 23060 3606
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3470
rect 27540 3194 27568 10406
rect 28276 3602 28304 336194
rect 29644 333260 29696 333266
rect 29644 333202 29696 333208
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 27712 3324 27764 3330
rect 27712 3266 27764 3272
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 26528 480 26556 3130
rect 27724 480 27752 3266
rect 28920 480 28948 3674
rect 29656 3670 29684 333202
rect 32416 59362 32444 343674
rect 231872 343670 231900 344927
rect 232042 343768 232098 343777
rect 232042 343703 232044 343712
rect 232096 343703 232098 343712
rect 232044 343674 232096 343680
rect 231860 343664 231912 343670
rect 231860 343606 231912 343612
rect 232042 342408 232098 342417
rect 232042 342343 232098 342352
rect 232056 342310 232084 342343
rect 232044 342304 232096 342310
rect 232044 342246 232096 342252
rect 232042 341184 232098 341193
rect 232042 341119 232098 341128
rect 232056 340950 232084 341119
rect 232044 340944 232096 340950
rect 232044 340886 232096 340892
rect 232042 339824 232098 339833
rect 232042 339759 232098 339768
rect 232056 339522 232084 339759
rect 232044 339516 232096 339522
rect 232044 339458 232096 339464
rect 232042 338600 232098 338609
rect 232042 338535 232098 338544
rect 232056 338162 232084 338535
rect 232044 338156 232096 338162
rect 232044 338098 232096 338104
rect 231124 336660 231176 336666
rect 231124 336602 231176 336608
rect 226984 336592 227036 336598
rect 226984 336534 227036 336540
rect 224224 336524 224276 336530
rect 224224 336466 224276 336472
rect 125508 336456 125560 336462
rect 125508 336398 125560 336404
rect 114468 336388 114520 336394
rect 114468 336330 114520 336336
rect 35164 336320 35216 336326
rect 35164 336262 35216 336268
rect 33784 320884 33836 320890
rect 33784 320826 33836 320832
rect 32404 59356 32456 59362
rect 32404 59298 32456 59304
rect 30104 10532 30156 10538
rect 30104 10474 30156 10480
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 30116 480 30144 10474
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 31312 480 31340 3062
rect 32416 480 32444 3606
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 33612 480 33640 3538
rect 33796 3330 33824 320826
rect 34428 10600 34480 10606
rect 34428 10542 34480 10548
rect 34440 3602 34468 10542
rect 35176 3738 35204 336262
rect 97908 334688 97960 334694
rect 97908 334630 97960 334636
rect 39304 334620 39356 334626
rect 39304 334562 39356 334568
rect 35808 330540 35860 330546
rect 35808 330482 35860 330488
rect 35164 3732 35216 3738
rect 35164 3674 35216 3680
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 35820 3398 35848 330482
rect 36544 309800 36596 309806
rect 36544 309742 36596 309748
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 33784 3324 33836 3330
rect 33784 3266 33836 3272
rect 34808 480 34836 3334
rect 36004 480 36032 3606
rect 36556 3126 36584 309742
rect 37188 10668 37240 10674
rect 37188 10610 37240 10616
rect 36544 3120 36596 3126
rect 36544 3062 36596 3068
rect 37200 480 37228 10610
rect 39316 3398 39344 334562
rect 95148 333328 95200 333334
rect 95148 333270 95200 333276
rect 68928 331900 68980 331906
rect 68928 331842 68980 331848
rect 43444 329112 43496 329118
rect 43444 329054 43496 329060
rect 41328 10736 41380 10742
rect 41328 10678 41380 10684
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 38396 480 38424 3334
rect 39592 480 39620 3674
rect 41340 3398 41368 10678
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 40696 480 40724 3334
rect 41892 480 41920 3334
rect 43088 480 43116 3742
rect 43456 3398 43484 329054
rect 46204 327752 46256 327758
rect 46204 327694 46256 327700
rect 45468 10804 45520 10810
rect 45468 10746 45520 10752
rect 45376 4140 45428 4146
rect 45376 4082 45428 4088
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 44284 480 44312 3334
rect 45388 2122 45416 4082
rect 45480 3398 45508 10746
rect 46216 4146 46244 327694
rect 50988 323672 51040 323678
rect 50988 323614 51040 323620
rect 49608 10872 49660 10878
rect 49608 10814 49660 10820
rect 47860 7676 47912 7682
rect 47860 7618 47912 7624
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 46664 3868 46716 3874
rect 46664 3810 46716 3816
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45388 2094 45508 2122
rect 45480 480 45508 2094
rect 46676 480 46704 3810
rect 47872 480 47900 7618
rect 49620 3398 49648 10814
rect 51000 3398 51028 323614
rect 57888 322244 57940 322250
rect 57888 322186 57940 322192
rect 53748 318096 53800 318102
rect 53748 318038 53800 318044
rect 53656 10940 53708 10946
rect 53656 10882 53708 10888
rect 51356 7744 51408 7750
rect 51356 7686 51408 7692
rect 48964 3392 49016 3398
rect 48964 3334 49016 3340
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 48976 480 49004 3334
rect 50172 480 50200 3334
rect 51368 480 51396 7686
rect 53668 3398 53696 10882
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 53656 3392 53708 3398
rect 53656 3334 53708 3340
rect 52564 480 52592 3334
rect 53760 480 53788 318038
rect 56508 11008 56560 11014
rect 56508 10950 56560 10956
rect 54944 9104 54996 9110
rect 54944 9046 54996 9052
rect 54956 480 54984 9046
rect 56520 3398 56548 10950
rect 57900 3398 57928 322186
rect 62028 316736 62080 316742
rect 62028 316678 62080 316684
rect 60648 10260 60700 10266
rect 60648 10202 60700 10208
rect 58440 9172 58492 9178
rect 58440 9114 58492 9120
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56508 3392 56560 3398
rect 56508 3334 56560 3340
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 57888 3392 57940 3398
rect 57888 3334 57940 3340
rect 56060 480 56088 3334
rect 57256 480 57284 3334
rect 58452 480 58480 9114
rect 60660 2990 60688 10202
rect 61936 9240 61988 9246
rect 61936 9182 61988 9188
rect 60832 3936 60884 3942
rect 60832 3878 60884 3884
rect 59636 2984 59688 2990
rect 59636 2926 59688 2932
rect 60648 2984 60700 2990
rect 60648 2926 60700 2932
rect 59648 480 59676 2926
rect 60844 480 60872 3878
rect 61948 3482 61976 9182
rect 62040 3942 62068 316678
rect 64788 308440 64840 308446
rect 64788 308382 64840 308388
rect 63224 10192 63276 10198
rect 63224 10134 63276 10140
rect 62028 3936 62080 3942
rect 62028 3878 62080 3884
rect 61948 3454 62068 3482
rect 62040 480 62068 3454
rect 63236 480 63264 10134
rect 64800 3398 64828 308382
rect 67548 10124 67600 10130
rect 67548 10066 67600 10072
rect 65524 9308 65576 9314
rect 65524 9250 65576 9256
rect 64328 3392 64380 3398
rect 64328 3334 64380 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64340 480 64368 3334
rect 65536 480 65564 9250
rect 67560 3398 67588 10066
rect 68940 3398 68968 331842
rect 85488 327820 85540 327826
rect 85488 327762 85540 327768
rect 71688 315308 71740 315314
rect 71688 315250 71740 315256
rect 70308 10056 70360 10062
rect 70308 9998 70360 10004
rect 69112 9376 69164 9382
rect 69112 9318 69164 9324
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 67548 3392 67600 3398
rect 67548 3334 67600 3340
rect 67916 3392 67968 3398
rect 67916 3334 67968 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 66732 480 66760 3334
rect 67928 480 67956 3334
rect 69124 480 69152 9318
rect 70320 480 70348 9998
rect 71700 6914 71728 315250
rect 81348 307080 81400 307086
rect 81348 307022 81400 307028
rect 74448 9988 74500 9994
rect 74448 9930 74500 9936
rect 72608 9444 72660 9450
rect 72608 9386 72660 9392
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 72620 480 72648 9386
rect 74460 3398 74488 9930
rect 78588 9920 78640 9926
rect 78588 9862 78640 9868
rect 76196 9512 76248 9518
rect 76196 9454 76248 9460
rect 75000 3936 75052 3942
rect 75000 3878 75052 3884
rect 73804 3392 73856 3398
rect 73804 3334 73856 3340
rect 74448 3392 74500 3398
rect 74448 3334 74500 3340
rect 73816 480 73844 3334
rect 75012 480 75040 3878
rect 76208 480 76236 9454
rect 78496 4004 78548 4010
rect 78496 3946 78548 3952
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 77404 480 77432 3334
rect 78508 1986 78536 3946
rect 78600 3398 78628 9862
rect 79692 9580 79744 9586
rect 79692 9522 79744 9528
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78508 1958 78628 1986
rect 78600 480 78628 1958
rect 79704 480 79732 9522
rect 81360 3398 81388 307022
rect 83280 9648 83332 9654
rect 83280 9590 83332 9596
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82096 480 82124 4014
rect 83292 480 83320 9590
rect 85500 3398 85528 327762
rect 92388 324964 92440 324970
rect 92388 324906 92440 324912
rect 88248 322312 88300 322318
rect 88248 322254 88300 322260
rect 86868 8900 86920 8906
rect 86868 8842 86920 8848
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 85488 3392 85540 3398
rect 85488 3334 85540 3340
rect 84488 480 84516 3334
rect 85684 480 85712 4082
rect 86880 480 86908 8842
rect 88260 6914 88288 322254
rect 90364 8832 90416 8838
rect 90364 8774 90416 8780
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 8774
rect 92400 3398 92428 324906
rect 95056 318164 95108 318170
rect 95056 318106 95108 318112
rect 95068 3482 95096 318106
rect 95160 3618 95188 333270
rect 95160 3590 95280 3618
rect 95068 3454 95188 3482
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 92388 3392 92440 3398
rect 92388 3334 92440 3340
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 91572 480 91600 3334
rect 92756 3188 92808 3194
rect 92756 3130 92808 3136
rect 92768 480 92796 3130
rect 93964 480 93992 3334
rect 95160 480 95188 3454
rect 95252 3398 95280 3590
rect 97920 3398 97948 334630
rect 108948 331968 109000 331974
rect 108948 331910 109000 331916
rect 102048 330608 102100 330614
rect 102048 330550 102100 330556
rect 99288 316804 99340 316810
rect 99288 316746 99340 316752
rect 99300 3398 99328 316746
rect 102060 3398 102088 330550
rect 104808 326392 104860 326398
rect 104808 326334 104860 326340
rect 103428 315376 103480 315382
rect 103428 315318 103480 315324
rect 95240 3392 95292 3398
rect 95240 3334 95292 3340
rect 97448 3392 97500 3398
rect 97448 3334 97500 3340
rect 97908 3392 97960 3398
rect 97908 3334 97960 3340
rect 98644 3392 98696 3398
rect 98644 3334 98696 3340
rect 99288 3392 99340 3398
rect 99288 3334 99340 3340
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 102048 3392 102100 3398
rect 102048 3334 102100 3340
rect 96252 3120 96304 3126
rect 96252 3062 96304 3068
rect 96264 480 96292 3062
rect 97460 480 97488 3334
rect 98656 480 98684 3334
rect 99840 3052 99892 3058
rect 99840 2994 99892 3000
rect 99852 480 99880 2994
rect 101048 480 101076 3334
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 102232 2984 102284 2990
rect 102232 2926 102284 2932
rect 102244 480 102272 2926
rect 103348 480 103376 3062
rect 103440 2990 103468 315318
rect 104820 6914 104848 326334
rect 106188 319456 106240 319462
rect 106188 319398 106240 319404
rect 104544 6886 104848 6914
rect 103428 2984 103480 2990
rect 103428 2926 103480 2932
rect 104544 480 104572 6886
rect 106200 3194 106228 319398
rect 108960 3194 108988 331910
rect 113088 326460 113140 326466
rect 113088 326402 113140 326408
rect 111708 320952 111760 320958
rect 111708 320894 111760 320900
rect 110328 305652 110380 305658
rect 110328 305594 110380 305600
rect 110340 3194 110368 305594
rect 111720 6914 111748 320894
rect 113100 6914 113128 326402
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 105728 3188 105780 3194
rect 105728 3130 105780 3136
rect 106188 3188 106240 3194
rect 106188 3130 106240 3136
rect 108120 3188 108172 3194
rect 108120 3130 108172 3136
rect 108948 3188 109000 3194
rect 108948 3130 109000 3136
rect 109316 3188 109368 3194
rect 109316 3130 109368 3136
rect 110328 3188 110380 3194
rect 110328 3130 110380 3136
rect 105740 480 105768 3130
rect 106924 2916 106976 2922
rect 106924 2858 106976 2864
rect 106936 480 106964 2858
rect 108132 480 108160 3130
rect 109328 480 109356 3130
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110524 480 110552 2926
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114480 3058 114508 336330
rect 115848 329180 115900 329186
rect 115848 329122 115900 329128
rect 115860 3058 115888 329122
rect 117228 313948 117280 313954
rect 117228 313890 117280 313896
rect 117240 3058 117268 313890
rect 119988 312588 120040 312594
rect 119988 312530 120040 312536
rect 119896 9852 119948 9858
rect 119896 9794 119948 9800
rect 119908 3058 119936 9794
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 114468 3052 114520 3058
rect 114468 2994 114520 3000
rect 115204 3052 115256 3058
rect 115204 2994 115256 3000
rect 115848 3052 115900 3058
rect 115848 2994 115900 3000
rect 116400 3052 116452 3058
rect 116400 2994 116452 3000
rect 117228 3052 117280 3058
rect 117228 2994 117280 3000
rect 118792 3052 118844 3058
rect 118792 2994 118844 3000
rect 119896 3052 119948 3058
rect 119896 2994 119948 3000
rect 114020 480 114048 2994
rect 115216 480 115244 2994
rect 116412 480 116440 2994
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 117608 480 117636 2790
rect 118804 480 118832 2994
rect 120000 1442 120028 312530
rect 124128 304292 124180 304298
rect 124128 304234 124180 304240
rect 122748 9784 122800 9790
rect 122748 9726 122800 9732
rect 122760 2922 122788 9726
rect 124140 2922 124168 304234
rect 125520 2922 125548 336398
rect 219348 335028 219400 335034
rect 219348 334970 219400 334976
rect 210976 334960 211028 334966
rect 210976 334902 211028 334908
rect 176568 334892 176620 334898
rect 176568 334834 176620 334840
rect 158628 334824 158680 334830
rect 158628 334766 158680 334772
rect 126888 334756 126940 334762
rect 126888 334698 126940 334704
rect 126900 2922 126928 334698
rect 144828 333396 144880 333402
rect 144828 333338 144880 333344
rect 136548 332036 136600 332042
rect 136548 331978 136600 331984
rect 128268 325032 128320 325038
rect 128268 324974 128320 324980
rect 128176 7812 128228 7818
rect 128176 7754 128228 7760
rect 126980 4208 127032 4214
rect 126980 4150 127032 4156
rect 122288 2916 122340 2922
rect 122288 2858 122340 2864
rect 122748 2916 122800 2922
rect 122748 2858 122800 2864
rect 123484 2916 123536 2922
rect 123484 2858 123536 2864
rect 124128 2916 124180 2922
rect 124128 2858 124180 2864
rect 124680 2916 124732 2922
rect 124680 2858 124732 2864
rect 125508 2916 125560 2922
rect 125508 2858 125560 2864
rect 125876 2916 125928 2922
rect 125876 2858 125928 2864
rect 126888 2916 126940 2922
rect 126888 2858 126940 2864
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 119908 1414 120028 1442
rect 119908 480 119936 1414
rect 121104 480 121132 2790
rect 122300 480 122328 2858
rect 123496 480 123524 2858
rect 124692 480 124720 2858
rect 125888 480 125916 2858
rect 126992 480 127020 4150
rect 128188 480 128216 7754
rect 128280 4214 128308 324974
rect 135168 322380 135220 322386
rect 135168 322322 135220 322328
rect 131764 7880 131816 7886
rect 131764 7822 131816 7828
rect 130568 6180 130620 6186
rect 130568 6122 130620 6128
rect 129372 5092 129424 5098
rect 129372 5034 129424 5040
rect 128268 4208 128320 4214
rect 128268 4150 128320 4156
rect 129384 480 129412 5034
rect 130580 480 130608 6122
rect 131776 480 131804 7822
rect 135180 6914 135208 322322
rect 136456 309868 136508 309874
rect 136456 309810 136508 309816
rect 134168 6886 135208 6914
rect 132960 5160 133012 5166
rect 132960 5102 133012 5108
rect 132972 480 133000 5102
rect 134168 480 134196 6886
rect 136468 4214 136496 309810
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 480 135300 4150
rect 136560 1442 136588 331978
rect 140688 329248 140740 329254
rect 140688 329190 140740 329196
rect 137928 321020 137980 321026
rect 137928 320962 137980 320968
rect 137940 6914 137968 320962
rect 139308 19984 139360 19990
rect 139308 19926 139360 19932
rect 139320 6914 139348 19926
rect 140700 6914 140728 329190
rect 144736 323740 144788 323746
rect 144736 323682 144788 323688
rect 142068 318232 142120 318238
rect 142068 318174 142120 318180
rect 142080 6914 142108 318174
rect 142436 8764 142488 8770
rect 142436 8706 142488 8712
rect 136468 1414 136588 1442
rect 137664 6886 137968 6914
rect 138860 6886 139348 6914
rect 140056 6886 140728 6914
rect 141252 6886 142108 6914
rect 136468 480 136496 1414
rect 137664 480 137692 6886
rect 138860 480 138888 6886
rect 140056 480 140084 6886
rect 141252 480 141280 6886
rect 142448 480 142476 8706
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 144748 480 144776 323682
rect 144840 4214 144868 333338
rect 147588 330676 147640 330682
rect 147588 330618 147640 330624
rect 145932 8696 145984 8702
rect 145932 8638 145984 8644
rect 144828 4208 144880 4214
rect 144828 4150 144880 4156
rect 145944 480 145972 8638
rect 147600 6914 147628 330618
rect 151728 327888 151780 327894
rect 151728 327830 151780 327836
rect 148968 325100 149020 325106
rect 148968 325042 149020 325048
rect 148980 6914 149008 325042
rect 149520 8628 149572 8634
rect 149520 8570 149572 8576
rect 147140 6886 147628 6914
rect 148336 6886 149008 6914
rect 147140 480 147168 6886
rect 148336 480 148364 6886
rect 149532 480 149560 8570
rect 151740 6914 151768 327830
rect 154488 326528 154540 326534
rect 154488 326470 154540 326476
rect 153108 316872 153160 316878
rect 153108 316814 153160 316820
rect 153016 8560 153068 8566
rect 153016 8502 153068 8508
rect 150636 6886 151768 6914
rect 150636 480 150664 6886
rect 151820 4208 151872 4214
rect 151820 4150 151872 4156
rect 151832 480 151860 4150
rect 153028 480 153056 8502
rect 153120 4214 153148 316814
rect 154500 6914 154528 326470
rect 155868 315444 155920 315450
rect 155868 315386 155920 315392
rect 155880 6914 155908 315386
rect 156604 8492 156656 8498
rect 156604 8434 156656 8440
rect 154224 6886 154528 6914
rect 155420 6886 155908 6914
rect 153108 4208 153160 4214
rect 153108 4150 153160 4156
rect 154224 480 154252 6886
rect 155420 480 155448 6886
rect 156616 480 156644 8434
rect 158640 6914 158668 334766
rect 169668 333464 169720 333470
rect 169668 333406 169720 333412
rect 162768 332104 162820 332110
rect 162768 332046 162820 332052
rect 160008 327956 160060 327962
rect 160008 327898 160060 327904
rect 160020 6914 160048 327898
rect 161388 308508 161440 308514
rect 161388 308450 161440 308456
rect 161296 11756 161348 11762
rect 161296 11698 161348 11704
rect 157812 6886 158668 6914
rect 158916 6886 160048 6914
rect 157812 480 157840 6886
rect 158916 480 158944 6886
rect 160100 4208 160152 4214
rect 160100 4150 160152 4156
rect 160112 480 160140 4150
rect 161308 480 161336 11698
rect 161400 4214 161428 308450
rect 162780 6914 162808 332046
rect 166908 329316 166960 329322
rect 166908 329258 166960 329264
rect 164148 314016 164200 314022
rect 164148 313958 164200 313964
rect 164160 6914 164188 313958
rect 164884 13116 164936 13122
rect 164884 13058 164936 13064
rect 162504 6886 162808 6914
rect 163700 6886 164188 6914
rect 161388 4208 161440 4214
rect 161388 4150 161440 4156
rect 162504 480 162532 6886
rect 163700 480 163728 6886
rect 164896 480 164924 13058
rect 166920 6914 166948 329258
rect 169576 323808 169628 323814
rect 169576 323750 169628 323756
rect 168288 312656 168340 312662
rect 168288 312598 168340 312604
rect 168300 6914 168328 312598
rect 166092 6886 166948 6914
rect 167196 6886 168328 6914
rect 166092 480 166120 6886
rect 167196 480 167224 6886
rect 168380 4208 168432 4214
rect 168380 4150 168432 4156
rect 168392 480 168420 4150
rect 169588 480 169616 323750
rect 169680 4214 169708 333406
rect 171968 14476 172020 14482
rect 171968 14418 172020 14424
rect 170772 7948 170824 7954
rect 170772 7890 170824 7896
rect 169668 4208 169720 4214
rect 169668 4150 169720 4156
rect 170784 480 170812 7890
rect 171980 480 172008 14418
rect 174268 8016 174320 8022
rect 174268 7958 174320 7964
rect 173164 6248 173216 6254
rect 173164 6190 173216 6196
rect 173176 480 173204 6190
rect 174280 480 174308 7958
rect 176580 6914 176608 334834
rect 183468 333532 183520 333538
rect 183468 333474 183520 333480
rect 179328 330744 179380 330750
rect 179328 330686 179380 330692
rect 177856 8084 177908 8090
rect 177856 8026 177908 8032
rect 175476 6886 176608 6914
rect 175476 480 175504 6886
rect 176660 6316 176712 6322
rect 176660 6258 176712 6264
rect 176672 480 176700 6258
rect 177868 480 177896 8026
rect 179340 6914 179368 330686
rect 181444 8152 181496 8158
rect 181444 8094 181496 8100
rect 179064 6886 179368 6914
rect 179064 480 179092 6886
rect 180248 6384 180300 6390
rect 180248 6326 180300 6332
rect 180260 480 180288 6326
rect 181456 480 181484 8094
rect 183480 6914 183508 333474
rect 187608 330812 187660 330818
rect 187608 330754 187660 330760
rect 184848 328024 184900 328030
rect 184848 327966 184900 327972
rect 184860 6914 184888 327966
rect 186228 322448 186280 322454
rect 186228 322390 186280 322396
rect 186136 15904 186188 15910
rect 186136 15846 186188 15852
rect 182560 6886 183508 6914
rect 183756 6886 184888 6914
rect 182560 480 182588 6886
rect 183756 480 183784 6886
rect 184940 4208 184992 4214
rect 184940 4150 184992 4156
rect 184952 480 184980 4150
rect 186148 480 186176 15846
rect 186240 4214 186268 322390
rect 187620 6914 187648 330754
rect 188988 329384 189040 329390
rect 188988 329326 189040 329332
rect 189000 6914 189028 329326
rect 191748 326596 191800 326602
rect 191748 326538 191800 326544
rect 190368 17264 190420 17270
rect 190368 17206 190420 17212
rect 190380 6914 190408 17206
rect 191760 6914 191788 326538
rect 193128 311228 193180 311234
rect 193128 311170 193180 311176
rect 193140 6914 193168 311170
rect 199108 8288 199160 8294
rect 199108 8230 199160 8236
rect 195612 8220 195664 8226
rect 195612 8162 195664 8168
rect 187344 6886 187648 6914
rect 188540 6886 189028 6914
rect 189736 6886 190408 6914
rect 190840 6886 191788 6914
rect 192036 6886 193168 6914
rect 186228 4208 186280 4214
rect 186228 4150 186280 4156
rect 187344 480 187372 6886
rect 188540 480 188568 6886
rect 189736 480 189764 6886
rect 190840 480 190868 6886
rect 192036 480 192064 6886
rect 194416 6452 194468 6458
rect 194416 6394 194468 6400
rect 193220 5228 193272 5234
rect 193220 5170 193272 5176
rect 193232 480 193260 5170
rect 194428 480 194456 6394
rect 195624 480 195652 8162
rect 197912 6520 197964 6526
rect 197912 6462 197964 6468
rect 196808 5296 196860 5302
rect 196808 5238 196860 5244
rect 196820 480 196848 5238
rect 197924 480 197952 6462
rect 199120 480 199148 8230
rect 202696 7540 202748 7546
rect 202696 7482 202748 7488
rect 201500 6588 201552 6594
rect 201500 6530 201552 6536
rect 200304 5364 200356 5370
rect 200304 5306 200356 5312
rect 200316 480 200344 5306
rect 201512 480 201540 6530
rect 202708 480 202736 7482
rect 206192 7472 206244 7478
rect 206192 7414 206244 7420
rect 205088 6656 205140 6662
rect 205088 6598 205140 6604
rect 203892 5432 203944 5438
rect 203892 5374 203944 5380
rect 203904 480 203932 5374
rect 205100 480 205128 6598
rect 206204 480 206232 7414
rect 208584 6724 208636 6730
rect 208584 6666 208636 6672
rect 207388 5500 207440 5506
rect 207388 5442 207440 5448
rect 207400 480 207428 5442
rect 208596 480 208624 6666
rect 210988 4214 211016 334902
rect 219256 333600 219308 333606
rect 219256 333542 219308 333548
rect 213828 330880 213880 330886
rect 213828 330822 213880 330828
rect 213840 6914 213868 330822
rect 217968 326664 218020 326670
rect 217968 326606 218020 326612
rect 217980 6914 218008 326606
rect 213380 6886 213868 6914
rect 216876 6886 218008 6914
rect 212172 6792 212224 6798
rect 212172 6734 212224 6740
rect 211068 4752 211120 4758
rect 211068 4694 211120 4700
rect 209780 4208 209832 4214
rect 209780 4150 209832 4156
rect 210976 4208 211028 4214
rect 210976 4150 211028 4156
rect 209792 480 209820 4150
rect 211080 2394 211108 4694
rect 210988 2366 211108 2394
rect 210988 480 211016 2366
rect 212184 480 212212 6734
rect 213380 480 213408 6886
rect 215668 6860 215720 6866
rect 215668 6802 215720 6808
rect 214472 4616 214524 4622
rect 214472 4558 214524 4564
rect 214484 480 214512 4558
rect 215680 480 215708 6802
rect 216876 480 216904 6886
rect 218060 4208 218112 4214
rect 218060 4150 218112 4156
rect 218072 480 218100 4150
rect 219268 480 219296 333542
rect 219360 4214 219388 334970
rect 223488 332172 223540 332178
rect 223488 332114 223540 332120
rect 220728 319524 220780 319530
rect 220728 319466 220780 319472
rect 220740 6914 220768 319466
rect 221556 11484 221608 11490
rect 221556 11426 221608 11432
rect 220464 6886 220768 6914
rect 219348 4208 219400 4214
rect 219348 4150 219400 4156
rect 220464 480 220492 6886
rect 221568 480 221596 11426
rect 223500 6914 223528 332114
rect 224236 11490 224264 336466
rect 226248 335096 226300 335102
rect 226248 335038 226300 335044
rect 224868 325168 224920 325174
rect 224868 325110 224920 325116
rect 224224 11484 224276 11490
rect 224224 11426 224276 11432
rect 224880 6914 224908 325110
rect 226260 6914 226288 335038
rect 226996 15910 227024 336534
rect 229744 335776 229796 335782
rect 229744 335718 229796 335724
rect 227628 329452 227680 329458
rect 227628 329394 227680 329400
rect 227536 321088 227588 321094
rect 227536 321030 227588 321036
rect 226984 15904 227036 15910
rect 226984 15846 227036 15852
rect 222764 6886 223528 6914
rect 223960 6886 224908 6914
rect 225156 6886 226288 6914
rect 222764 480 222792 6886
rect 223960 480 223988 6886
rect 225156 480 225184 6886
rect 226340 4208 226392 4214
rect 226340 4150 226392 4156
rect 226352 480 226380 4150
rect 227548 480 227576 321030
rect 227640 4214 227668 329394
rect 229756 14482 229784 335718
rect 230388 333668 230440 333674
rect 230388 333610 230440 333616
rect 229744 14476 229796 14482
rect 229744 14418 229796 14424
rect 228732 4616 228784 4622
rect 228732 4558 228784 4564
rect 227628 4208 227680 4214
rect 227628 4150 227680 4156
rect 228744 480 228772 4558
rect 230400 3534 230428 333610
rect 231136 13122 231164 336602
rect 231768 328092 231820 328098
rect 231768 328034 231820 328040
rect 231124 13116 231176 13122
rect 231124 13058 231176 13064
rect 231780 3534 231808 328034
rect 232516 124166 232544 350095
rect 232608 176662 232636 355263
rect 232700 215286 232728 359207
rect 232792 229090 232820 359366
rect 232884 267714 232912 359502
rect 232976 280158 233004 364306
rect 233068 320142 233096 369543
rect 233160 332586 233188 370903
rect 306378 369880 306434 369889
rect 306378 369815 306434 369824
rect 306286 342408 306342 342417
rect 306286 342343 306342 342352
rect 306300 342310 306328 342343
rect 306288 342304 306340 342310
rect 306288 342246 306340 342252
rect 235000 338014 235060 338042
rect 234804 337952 234856 337958
rect 234804 337894 234856 337900
rect 233976 335980 234028 335986
rect 233976 335922 234028 335928
rect 233884 335912 233936 335918
rect 233884 335854 233936 335860
rect 233148 332580 233200 332586
rect 233148 332522 233200 332528
rect 233056 320136 233108 320142
rect 233056 320078 233108 320084
rect 232964 280152 233016 280158
rect 232964 280094 233016 280100
rect 232872 267708 232924 267714
rect 232872 267650 232924 267656
rect 232780 229084 232832 229090
rect 232780 229026 232832 229032
rect 232688 215280 232740 215286
rect 232688 215222 232740 215228
rect 232596 176656 232648 176662
rect 232596 176598 232648 176604
rect 232504 124160 232556 124166
rect 232504 124102 232556 124108
rect 233896 11762 233924 335854
rect 233988 17270 234016 335922
rect 234068 335844 234120 335850
rect 234068 335786 234120 335792
rect 234080 307086 234108 335786
rect 234528 332240 234580 332246
rect 234528 332182 234580 332188
rect 234068 307080 234120 307086
rect 234068 307022 234120 307028
rect 233976 17264 234028 17270
rect 233976 17206 234028 17212
rect 233884 11756 233936 11762
rect 233884 11698 233936 11704
rect 232228 4548 232280 4554
rect 232228 4490 232280 4496
rect 229836 3528 229888 3534
rect 229836 3470 229888 3476
rect 230388 3528 230440 3534
rect 230388 3470 230440 3476
rect 231032 3528 231084 3534
rect 231032 3470 231084 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 229848 480 229876 3470
rect 231044 480 231072 3470
rect 232240 480 232268 4490
rect 234540 3534 234568 332182
rect 234712 326256 234764 326262
rect 234712 326198 234764 326204
rect 234724 5030 234752 326198
rect 234712 5024 234764 5030
rect 234712 4966 234764 4972
rect 234816 4894 234844 337894
rect 234896 337748 234948 337754
rect 234896 337690 234948 337696
rect 234908 4962 234936 337690
rect 234896 4956 234948 4962
rect 234896 4898 234948 4904
rect 234804 4888 234856 4894
rect 234804 4830 234856 4836
rect 235000 4826 235028 338014
rect 235138 337958 235166 338028
rect 235276 338014 235336 338042
rect 235126 337952 235178 337958
rect 235126 337894 235178 337900
rect 235276 337890 235304 338014
rect 235264 337884 235316 337890
rect 235264 337826 235316 337832
rect 235414 337770 235442 338028
rect 235092 337742 235442 337770
rect 235552 338014 235612 338042
rect 235092 8974 235120 337742
rect 235552 336054 235580 338014
rect 235690 337770 235718 338028
rect 235644 337742 235718 337770
rect 235828 338014 235888 338042
rect 235540 336048 235592 336054
rect 235540 335990 235592 335996
rect 235172 326324 235224 326330
rect 235172 326266 235224 326272
rect 235184 10334 235212 326266
rect 235644 316034 235672 337742
rect 235828 326262 235856 338014
rect 235966 337770 235994 338028
rect 236104 338014 236164 338042
rect 236104 337958 236132 338014
rect 236092 337952 236144 337958
rect 236242 337940 236270 338028
rect 236380 338014 236440 338042
rect 236242 337912 236316 337940
rect 236092 337894 236144 337900
rect 235920 337742 235994 337770
rect 236092 337816 236144 337822
rect 236092 337758 236144 337764
rect 235920 326330 235948 337742
rect 235908 326324 235960 326330
rect 235908 326266 235960 326272
rect 235816 326256 235868 326262
rect 235816 326198 235868 326204
rect 236104 320890 236132 337758
rect 236288 336258 236316 337912
rect 236276 336252 236328 336258
rect 236276 336194 236328 336200
rect 236380 331214 236408 338014
rect 236518 337736 236546 338028
rect 236656 338014 236716 338042
rect 236840 338014 236900 338042
rect 236518 337708 236592 337736
rect 236460 334620 236512 334626
rect 236460 334562 236512 334568
rect 236196 331186 236408 331214
rect 236092 320884 236144 320890
rect 236092 320826 236144 320832
rect 235276 316006 235672 316034
rect 235172 10328 235224 10334
rect 235172 10270 235224 10276
rect 235080 8968 235132 8974
rect 235080 8910 235132 8916
rect 234988 4820 235040 4826
rect 234988 4762 235040 4768
rect 233424 3528 233476 3534
rect 233424 3470 233476 3476
rect 234528 3528 234580 3534
rect 234528 3470 234580 3476
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 233436 480 233464 3470
rect 234632 480 234660 3470
rect 235276 3369 235304 316006
rect 235816 13116 235868 13122
rect 235816 13058 235868 13064
rect 235828 3534 235856 13058
rect 236196 7614 236224 331186
rect 236368 326324 236420 326330
rect 236368 326266 236420 326272
rect 236276 320884 236328 320890
rect 236276 320826 236328 320832
rect 236288 9042 236316 320826
rect 236380 311166 236408 326266
rect 236368 311160 236420 311166
rect 236368 311102 236420 311108
rect 236276 9036 236328 9042
rect 236276 8978 236328 8984
rect 236184 7608 236236 7614
rect 236184 7550 236236 7556
rect 235908 4820 235960 4826
rect 235908 4762 235960 4768
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 235262 3360 235318 3369
rect 235262 3295 235318 3304
rect 235920 2394 235948 4762
rect 236472 3505 236500 334562
rect 236564 323610 236592 337708
rect 236656 334626 236684 338014
rect 236736 335436 236788 335442
rect 236736 335378 236788 335384
rect 236644 334620 236696 334626
rect 236644 334562 236696 334568
rect 236748 331214 236776 335378
rect 236656 331186 236776 331214
rect 236552 323604 236604 323610
rect 236552 323546 236604 323552
rect 236656 315314 236684 331186
rect 236840 316034 236868 338014
rect 236978 337822 237006 338028
rect 237116 338014 237176 338042
rect 236966 337816 237018 337822
rect 236966 337758 237018 337764
rect 237116 326330 237144 338014
rect 237254 337770 237282 338028
rect 237208 337742 237282 337770
rect 237438 337770 237466 338028
rect 237530 337872 237558 338028
rect 237714 337872 237742 338028
rect 237806 337940 237834 338028
rect 237806 337912 237880 337940
rect 237530 337844 237604 337872
rect 237714 337844 237788 337872
rect 237438 337742 237512 337770
rect 237208 336190 237236 337742
rect 237196 336184 237248 336190
rect 237196 336126 237248 336132
rect 237104 326324 237156 326330
rect 237104 326266 237156 326272
rect 237484 326126 237512 337742
rect 237576 326738 237604 337844
rect 237760 333266 237788 337844
rect 237748 333260 237800 333266
rect 237748 333202 237800 333208
rect 237852 328454 237880 337912
rect 237990 337770 238018 338028
rect 238082 337872 238110 338028
rect 238082 337844 238156 337872
rect 237990 337742 238064 337770
rect 237668 328426 237880 328454
rect 237564 326732 237616 326738
rect 237564 326674 237616 326680
rect 237668 326346 237696 328426
rect 237748 326732 237800 326738
rect 237748 326674 237800 326680
rect 237576 326318 237696 326346
rect 237472 326120 237524 326126
rect 237472 326062 237524 326068
rect 236748 316006 236868 316034
rect 236644 315308 236696 315314
rect 236644 315250 236696 315256
rect 236748 3641 236776 316006
rect 237012 11756 237064 11762
rect 237012 11698 237064 11704
rect 236734 3632 236790 3641
rect 236734 3567 236790 3576
rect 236458 3496 236514 3505
rect 236458 3431 236514 3440
rect 235828 2366 235948 2394
rect 235828 480 235856 2366
rect 237024 480 237052 11698
rect 237576 4214 237604 326318
rect 237656 326256 237708 326262
rect 237656 326198 237708 326204
rect 237668 10470 237696 326198
rect 237656 10464 237708 10470
rect 237656 10406 237708 10412
rect 237760 10402 237788 326674
rect 237840 326324 237892 326330
rect 237840 326266 237892 326272
rect 237852 10538 237880 326266
rect 237932 326188 237984 326194
rect 237932 326130 237984 326136
rect 237944 309806 237972 326130
rect 238036 321554 238064 337742
rect 238128 326262 238156 337844
rect 238266 337770 238294 338028
rect 238358 337906 238386 338028
rect 238496 338014 238556 338042
rect 238680 338014 238740 338042
rect 238358 337878 238432 337906
rect 238266 337742 238340 337770
rect 238116 326256 238168 326262
rect 238116 326198 238168 326204
rect 238208 326120 238260 326126
rect 238208 326062 238260 326068
rect 238036 321526 238156 321554
rect 237932 309800 237984 309806
rect 237932 309742 237984 309748
rect 238128 16574 238156 321526
rect 238036 16546 238156 16574
rect 237840 10532 237892 10538
rect 237840 10474 237892 10480
rect 237748 10396 237800 10402
rect 237748 10338 237800 10344
rect 237564 4208 237616 4214
rect 237564 4150 237616 4156
rect 238036 3602 238064 16546
rect 238116 8968 238168 8974
rect 238116 8910 238168 8916
rect 238024 3596 238076 3602
rect 238024 3538 238076 3544
rect 238128 480 238156 8910
rect 238220 3777 238248 326062
rect 238312 320822 238340 337742
rect 238404 336326 238432 337878
rect 238392 336320 238444 336326
rect 238392 336262 238444 336268
rect 238496 326330 238524 338014
rect 238484 326324 238536 326330
rect 238484 326266 238536 326272
rect 238680 326194 238708 338014
rect 238818 337736 238846 338028
rect 239002 337770 239030 338028
rect 239094 337890 239122 338028
rect 239232 338014 239292 338042
rect 239082 337884 239134 337890
rect 239082 337826 239134 337832
rect 239002 337742 239076 337770
rect 238818 337708 238892 337736
rect 238668 326188 238720 326194
rect 238668 326130 238720 326136
rect 238300 320816 238352 320822
rect 238300 320758 238352 320764
rect 238206 3768 238262 3777
rect 238864 3738 238892 337708
rect 239048 331226 239076 337742
rect 239036 331220 239088 331226
rect 239232 331214 239260 338014
rect 239370 337770 239398 338028
rect 239036 331162 239088 331168
rect 239140 331186 239260 331214
rect 239324 337742 239398 337770
rect 239508 338014 239568 338042
rect 239140 326346 239168 331186
rect 239220 331152 239272 331158
rect 239220 331094 239272 331100
rect 238956 326318 239168 326346
rect 238206 3703 238262 3712
rect 238852 3732 238904 3738
rect 238852 3674 238904 3680
rect 238956 3670 238984 326318
rect 239128 326256 239180 326262
rect 239128 326198 239180 326204
rect 239036 326188 239088 326194
rect 239036 326130 239088 326136
rect 239048 3806 239076 326130
rect 239140 10742 239168 326198
rect 239128 10736 239180 10742
rect 239128 10678 239180 10684
rect 239232 10606 239260 331094
rect 239324 10674 239352 337742
rect 239508 334558 239536 338014
rect 239646 337770 239674 338028
rect 239600 337742 239674 337770
rect 239784 338014 239844 338042
rect 239496 334552 239548 334558
rect 239496 334494 239548 334500
rect 239600 316034 239628 337742
rect 239784 326262 239812 338014
rect 239922 337906 239950 338028
rect 239876 337878 239950 337906
rect 240060 338014 240120 338042
rect 239876 329118 239904 337878
rect 239864 329112 239916 329118
rect 239864 329054 239916 329060
rect 239772 326256 239824 326262
rect 239772 326198 239824 326204
rect 240060 326194 240088 338014
rect 240198 337906 240226 338028
rect 240336 338014 240396 338042
rect 240198 337878 240272 337906
rect 240140 337816 240192 337822
rect 240140 337758 240192 337764
rect 240152 326346 240180 337758
rect 240244 326482 240272 337878
rect 240336 327758 240364 338014
rect 240566 337770 240594 338028
rect 240658 337906 240686 338028
rect 240796 338014 240856 338042
rect 240658 337878 240732 337906
rect 240566 337742 240640 337770
rect 240324 327752 240376 327758
rect 240324 327694 240376 327700
rect 240244 326454 240548 326482
rect 240152 326318 240272 326346
rect 240048 326188 240100 326194
rect 240048 326130 240100 326136
rect 240140 326188 240192 326194
rect 240140 326130 240192 326136
rect 240152 318102 240180 326130
rect 240244 323678 240272 326318
rect 240416 326256 240468 326262
rect 240416 326198 240468 326204
rect 240232 323672 240284 323678
rect 240232 323614 240284 323620
rect 240140 318096 240192 318102
rect 240140 318038 240192 318044
rect 239416 316006 239628 316034
rect 239312 10668 239364 10674
rect 239312 10610 239364 10616
rect 239220 10600 239272 10606
rect 239220 10542 239272 10548
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 239036 3800 239088 3806
rect 239036 3742 239088 3748
rect 238944 3664 238996 3670
rect 238944 3606 238996 3612
rect 239324 480 239352 4830
rect 239416 3466 239444 316006
rect 240428 9110 240456 326198
rect 240520 10810 240548 326454
rect 240612 326369 240640 337742
rect 240704 331158 240732 337878
rect 240692 331152 240744 331158
rect 240692 331094 240744 331100
rect 240598 326360 240654 326369
rect 240598 326295 240654 326304
rect 240796 326210 240824 338014
rect 240934 337822 240962 338028
rect 241072 338014 241132 338042
rect 240922 337816 240974 337822
rect 240922 337758 240974 337764
rect 241072 331214 241100 338014
rect 241210 337770 241238 338028
rect 240704 326182 240824 326210
rect 240888 331186 241100 331214
rect 241164 337742 241238 337770
rect 241348 338014 241408 338042
rect 240704 326074 240732 326182
rect 240612 326046 240732 326074
rect 240782 326088 240838 326097
rect 240612 10878 240640 326046
rect 240782 326023 240838 326032
rect 240692 324012 240744 324018
rect 240692 323954 240744 323960
rect 240704 10946 240732 323954
rect 240692 10940 240744 10946
rect 240692 10882 240744 10888
rect 240600 10872 240652 10878
rect 240600 10814 240652 10820
rect 240508 10804 240560 10810
rect 240508 10746 240560 10752
rect 240416 9104 240468 9110
rect 240416 9046 240468 9052
rect 240796 3874 240824 326023
rect 240888 7750 240916 331186
rect 240968 331152 241020 331158
rect 240968 331094 241020 331100
rect 240876 7744 240928 7750
rect 240876 7686 240928 7692
rect 240980 7682 241008 331094
rect 241164 324018 241192 337742
rect 241348 326194 241376 338014
rect 241486 337770 241514 338028
rect 241670 337890 241698 338028
rect 241658 337884 241710 337890
rect 241658 337826 241710 337832
rect 241762 337770 241790 338028
rect 241440 337742 241514 337770
rect 241624 337742 241790 337770
rect 241900 338014 241960 338042
rect 242084 338014 242144 338042
rect 241440 326262 241468 337742
rect 241520 333260 241572 333266
rect 241520 333202 241572 333208
rect 241428 326256 241480 326262
rect 241428 326198 241480 326204
rect 241336 326188 241388 326194
rect 241336 326130 241388 326136
rect 241152 324012 241204 324018
rect 241152 323954 241204 323960
rect 241532 316742 241560 333202
rect 241624 322250 241652 337742
rect 241900 333010 241928 338014
rect 241808 332982 241928 333010
rect 241808 326346 241836 332982
rect 242084 331214 242112 338014
rect 242222 337906 242250 338028
rect 242360 338014 242420 338042
rect 242222 337878 242296 337906
rect 242164 337816 242216 337822
rect 242164 337758 242216 337764
rect 241716 326318 241836 326346
rect 241900 331186 242112 331214
rect 241612 322244 241664 322250
rect 241612 322186 241664 322192
rect 241520 316736 241572 316742
rect 241520 316678 241572 316684
rect 241428 11824 241480 11830
rect 241428 11766 241480 11772
rect 240968 7676 241020 7682
rect 240968 7618 241020 7624
rect 240784 3868 240836 3874
rect 240784 3810 240836 3816
rect 241440 3534 241468 11766
rect 241716 9178 241744 326318
rect 241796 326256 241848 326262
rect 241796 326198 241848 326204
rect 241808 10198 241836 326198
rect 241900 10266 241928 331186
rect 242176 326346 242204 337758
rect 242268 333266 242296 337878
rect 242256 333260 242308 333266
rect 242256 333202 242308 333208
rect 241992 326318 242204 326346
rect 241992 11014 242020 326318
rect 242072 325916 242124 325922
rect 242072 325858 242124 325864
rect 242084 308446 242112 325858
rect 242072 308440 242124 308446
rect 242072 308382 242124 308388
rect 241980 11008 242032 11014
rect 241980 10950 242032 10956
rect 241888 10260 241940 10266
rect 241888 10202 241940 10208
rect 241796 10192 241848 10198
rect 241796 10134 241848 10140
rect 242360 9246 242388 338014
rect 242498 337770 242526 338028
rect 242452 337742 242526 337770
rect 242636 338014 242696 338042
rect 242452 326262 242480 337742
rect 242440 326256 242492 326262
rect 242440 326198 242492 326204
rect 242636 325922 242664 338014
rect 242774 337770 242802 338028
rect 242728 337742 242802 337770
rect 242958 337770 242986 338028
rect 243050 337906 243078 338028
rect 243188 338014 243248 338042
rect 243050 337878 243124 337906
rect 242958 337742 243032 337770
rect 242624 325916 242676 325922
rect 242624 325858 242676 325864
rect 242728 316034 242756 337742
rect 242900 334620 242952 334626
rect 242900 334562 242952 334568
rect 242912 320890 242940 334562
rect 243004 331430 243032 337742
rect 243096 331906 243124 337878
rect 243084 331900 243136 331906
rect 243084 331842 243136 331848
rect 242992 331424 243044 331430
rect 242992 331366 243044 331372
rect 243188 326482 243216 338014
rect 243326 337906 243354 338028
rect 243464 338014 243524 338042
rect 243326 337878 243400 337906
rect 243268 337816 243320 337822
rect 243268 337758 243320 337764
rect 243004 326454 243216 326482
rect 242900 320884 242952 320890
rect 242900 320826 242952 320832
rect 242452 316006 242756 316034
rect 242452 9314 242480 316006
rect 242808 10328 242860 10334
rect 242808 10270 242860 10276
rect 242440 9308 242492 9314
rect 242440 9250 242492 9256
rect 242348 9240 242400 9246
rect 242348 9182 242400 9188
rect 241704 9172 241756 9178
rect 241704 9114 241756 9120
rect 242820 3534 242848 10270
rect 243004 9382 243032 326454
rect 243280 326346 243308 337758
rect 243372 333146 243400 337878
rect 243464 335442 243492 338014
rect 243602 337822 243630 338028
rect 243740 338014 243800 338042
rect 243924 338014 243984 338042
rect 243590 337816 243642 337822
rect 243590 337758 243642 337764
rect 243452 335436 243504 335442
rect 243452 335378 243504 335384
rect 243372 333118 243492 333146
rect 243360 331424 243412 331430
rect 243360 331366 243412 331372
rect 243188 326318 243308 326346
rect 243084 320884 243136 320890
rect 243084 320826 243136 320832
rect 243096 9518 243124 320826
rect 243084 9512 243136 9518
rect 243084 9454 243136 9460
rect 243188 9450 243216 326318
rect 243268 326256 243320 326262
rect 243268 326198 243320 326204
rect 243280 9994 243308 326198
rect 243372 10130 243400 331366
rect 243360 10124 243412 10130
rect 243360 10066 243412 10072
rect 243464 10062 243492 333118
rect 243544 326324 243596 326330
rect 243544 326266 243596 326272
rect 243452 10056 243504 10062
rect 243452 9998 243504 10004
rect 243268 9988 243320 9994
rect 243268 9930 243320 9936
rect 243556 9926 243584 326266
rect 243740 326262 243768 338014
rect 243728 326256 243780 326262
rect 243728 326198 243780 326204
rect 243924 316034 243952 338014
rect 244062 337770 244090 338028
rect 244016 337742 244090 337770
rect 244200 338014 244260 338042
rect 244016 334626 244044 337742
rect 244004 334620 244056 334626
rect 244004 334562 244056 334568
rect 244200 326330 244228 338014
rect 244338 337906 244366 338028
rect 244338 337878 244412 337906
rect 244384 328454 244412 337878
rect 244522 337770 244550 338028
rect 244614 337890 244642 338028
rect 244752 338014 244812 338042
rect 244602 337884 244654 337890
rect 244602 337826 244654 337832
rect 244522 337742 244688 337770
rect 244556 330472 244608 330478
rect 244556 330414 244608 330420
rect 244384 328426 244504 328454
rect 244188 326324 244240 326330
rect 244188 326266 244240 326272
rect 243648 316006 243952 316034
rect 243544 9920 243596 9926
rect 243544 9862 243596 9868
rect 243176 9444 243228 9450
rect 243176 9386 243228 9392
rect 242992 9376 243044 9382
rect 242992 9318 243044 9324
rect 242900 4956 242952 4962
rect 242900 4898 242952 4904
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 241704 3528 241756 3534
rect 241704 3470 241756 3476
rect 242808 3528 242860 3534
rect 242808 3470 242860 3476
rect 239404 3460 239456 3466
rect 239404 3402 239456 3408
rect 240520 480 240548 3470
rect 241716 480 241744 3470
rect 242912 480 242940 4898
rect 243648 3942 243676 316006
rect 244096 10396 244148 10402
rect 244096 10338 244148 10344
rect 243636 3936 243688 3942
rect 243636 3878 243688 3884
rect 244108 480 244136 10338
rect 244476 4010 244504 328426
rect 244568 4146 244596 330414
rect 244660 9586 244688 337742
rect 244752 330954 244780 338014
rect 244890 337770 244918 338028
rect 244844 337742 244918 337770
rect 245028 338014 245088 338042
rect 244740 330948 244792 330954
rect 244740 330890 244792 330896
rect 244844 330528 244872 337742
rect 245028 330954 245056 338014
rect 245166 337770 245194 338028
rect 245120 337742 245194 337770
rect 245304 338014 245364 338042
rect 244924 330948 244976 330954
rect 244924 330890 244976 330896
rect 245016 330948 245068 330954
rect 245016 330890 245068 330896
rect 244752 330500 244872 330528
rect 244752 9654 244780 330500
rect 244832 330404 244884 330410
rect 244832 330346 244884 330352
rect 244740 9648 244792 9654
rect 244740 9590 244792 9596
rect 244648 9580 244700 9586
rect 244648 9522 244700 9528
rect 244844 8906 244872 330346
rect 244832 8900 244884 8906
rect 244832 8842 244884 8848
rect 244556 4140 244608 4146
rect 244556 4082 244608 4088
rect 244936 4078 244964 330890
rect 245016 330540 245068 330546
rect 245016 330482 245068 330488
rect 244924 4072 244976 4078
rect 244924 4014 244976 4020
rect 244464 4004 244516 4010
rect 244464 3946 244516 3952
rect 245028 3398 245056 330482
rect 245120 330478 245148 337742
rect 245200 330948 245252 330954
rect 245200 330890 245252 330896
rect 245108 330472 245160 330478
rect 245108 330414 245160 330420
rect 245212 327826 245240 330890
rect 245304 330410 245332 338014
rect 245442 337770 245470 338028
rect 245396 337742 245470 337770
rect 245580 338014 245640 338042
rect 245292 330404 245344 330410
rect 245292 330346 245344 330352
rect 245200 327820 245252 327826
rect 245200 327762 245252 327768
rect 245396 322318 245424 337742
rect 245476 336048 245528 336054
rect 245476 335990 245528 335996
rect 245488 325694 245516 335990
rect 245580 330546 245608 338014
rect 245810 337770 245838 338028
rect 245902 337906 245930 338028
rect 246040 338014 246100 338042
rect 245902 337878 245976 337906
rect 245810 337742 245884 337770
rect 245568 330540 245620 330546
rect 245856 330528 245884 337742
rect 245948 333266 245976 337878
rect 245936 333260 245988 333266
rect 245936 333202 245988 333208
rect 245856 330500 245976 330528
rect 245568 330482 245620 330488
rect 245844 330404 245896 330410
rect 245844 330346 245896 330352
rect 245488 325666 245608 325694
rect 245384 322312 245436 322318
rect 245384 322254 245436 322260
rect 245580 6914 245608 325666
rect 245212 6886 245608 6914
rect 245016 3392 245068 3398
rect 245016 3334 245068 3340
rect 245212 480 245240 6886
rect 245856 3330 245884 330346
rect 245948 8838 245976 330500
rect 246040 330410 246068 338014
rect 246178 337906 246206 338028
rect 246178 337878 246252 337906
rect 246362 337890 246390 338028
rect 246120 337816 246172 337822
rect 246120 337758 246172 337764
rect 246028 330404 246080 330410
rect 246028 330346 246080 330352
rect 246028 330268 246080 330274
rect 246028 330210 246080 330216
rect 246040 316810 246068 330210
rect 246132 318170 246160 337758
rect 246224 333334 246252 337878
rect 246350 337884 246402 337890
rect 246350 337826 246402 337832
rect 246454 337770 246482 338028
rect 246316 337742 246482 337770
rect 246592 338014 246652 338042
rect 246212 333328 246264 333334
rect 246212 333270 246264 333276
rect 246212 330540 246264 330546
rect 246212 330482 246264 330488
rect 246120 318164 246172 318170
rect 246120 318106 246172 318112
rect 246028 316804 246080 316810
rect 246028 316746 246080 316752
rect 245936 8832 245988 8838
rect 245936 8774 245988 8780
rect 245844 3324 245896 3330
rect 245844 3266 245896 3272
rect 246224 3194 246252 330482
rect 246316 3262 246344 337742
rect 246592 334694 246620 338014
rect 246730 337770 246758 338028
rect 246684 337742 246758 337770
rect 246868 338014 246928 338042
rect 246580 334688 246632 334694
rect 246580 334630 246632 334636
rect 246396 333260 246448 333266
rect 246396 333202 246448 333208
rect 246408 324970 246436 333202
rect 246684 330274 246712 337742
rect 246868 330546 246896 338014
rect 247006 337770 247034 338028
rect 247190 337906 247218 338028
rect 247190 337878 247264 337906
rect 246960 337742 247034 337770
rect 247132 337816 247184 337822
rect 247132 337758 247184 337764
rect 246960 330614 246988 337742
rect 246948 330608 247000 330614
rect 246948 330550 247000 330556
rect 246856 330540 246908 330546
rect 246856 330482 246908 330488
rect 246672 330268 246724 330274
rect 246672 330210 246724 330216
rect 247144 326398 247172 337758
rect 247236 337634 247264 337878
rect 247374 337770 247402 338028
rect 247466 337890 247494 338028
rect 247604 338014 247664 338042
rect 247454 337884 247506 337890
rect 247454 337826 247506 337832
rect 247374 337742 247540 337770
rect 247236 337606 247448 337634
rect 247316 330540 247368 330546
rect 247316 330482 247368 330488
rect 247224 330472 247276 330478
rect 247224 330414 247276 330420
rect 247132 326392 247184 326398
rect 247132 326334 247184 326340
rect 246396 324964 246448 324970
rect 246396 324906 246448 324912
rect 246396 5024 246448 5030
rect 246396 4966 246448 4972
rect 246304 3256 246356 3262
rect 246304 3198 246356 3204
rect 246212 3188 246264 3194
rect 246212 3130 246264 3136
rect 246408 480 246436 4966
rect 247236 2990 247264 330414
rect 247328 305658 247356 330482
rect 247420 315382 247448 337606
rect 247512 330528 247540 337742
rect 247604 330698 247632 338014
rect 247742 337770 247770 338028
rect 247696 337742 247770 337770
rect 247880 338014 247940 338042
rect 247696 330834 247724 337742
rect 247880 331974 247908 338014
rect 248018 337770 248046 338028
rect 247972 337742 248046 337770
rect 248156 338014 248216 338042
rect 247868 331968 247920 331974
rect 247868 331910 247920 331916
rect 247696 330806 247908 330834
rect 247604 330670 247816 330698
rect 247684 330608 247736 330614
rect 247684 330550 247736 330556
rect 247512 330500 247632 330528
rect 247500 330404 247552 330410
rect 247500 330346 247552 330352
rect 247512 320958 247540 330346
rect 247500 320952 247552 320958
rect 247500 320894 247552 320900
rect 247408 315376 247460 315382
rect 247408 315318 247460 315324
rect 247316 305652 247368 305658
rect 247316 305594 247368 305600
rect 247604 16574 247632 330500
rect 247512 16546 247632 16574
rect 247512 3126 247540 16546
rect 247592 9036 247644 9042
rect 247592 8978 247644 8984
rect 247500 3120 247552 3126
rect 247500 3062 247552 3068
rect 247224 2984 247276 2990
rect 247224 2926 247276 2932
rect 247604 480 247632 8978
rect 247696 3058 247724 330550
rect 247788 319462 247816 330670
rect 247880 330614 247908 330806
rect 247868 330608 247920 330614
rect 247868 330550 247920 330556
rect 247972 330546 248000 337742
rect 247960 330540 248012 330546
rect 247960 330482 248012 330488
rect 248156 330478 248184 338014
rect 248294 337770 248322 338028
rect 248248 337742 248322 337770
rect 248478 337770 248506 338028
rect 248570 337906 248598 338028
rect 248708 338014 248768 338042
rect 248570 337878 248644 337906
rect 248478 337742 248552 337770
rect 248144 330472 248196 330478
rect 248144 330414 248196 330420
rect 248248 330410 248276 337742
rect 248236 330404 248288 330410
rect 248236 330346 248288 330352
rect 248524 326466 248552 337742
rect 248616 336394 248644 337878
rect 248708 337634 248736 338014
rect 248846 337770 248874 338028
rect 249030 337906 249058 338028
rect 249168 338014 249228 338042
rect 249030 337878 249104 337906
rect 248846 337742 249012 337770
rect 248708 337606 248828 337634
rect 248604 336388 248656 336394
rect 248604 336330 248656 336336
rect 248696 334620 248748 334626
rect 248696 334562 248748 334568
rect 248604 330268 248656 330274
rect 248604 330210 248656 330216
rect 248512 326460 248564 326466
rect 248512 326402 248564 326408
rect 247776 319456 247828 319462
rect 247776 319398 247828 319404
rect 248616 9858 248644 330210
rect 248604 9852 248656 9858
rect 248604 9794 248656 9800
rect 248708 9790 248736 334562
rect 248800 329186 248828 337606
rect 248880 329520 248932 329526
rect 248880 329462 248932 329468
rect 248788 329180 248840 329186
rect 248788 329122 248840 329128
rect 248788 327208 248840 327214
rect 248788 327150 248840 327156
rect 248800 304298 248828 327150
rect 248892 312594 248920 329462
rect 248984 313954 249012 337742
rect 248972 313948 249024 313954
rect 248972 313890 249024 313896
rect 248880 312588 248932 312594
rect 248880 312530 248932 312536
rect 248788 304292 248840 304298
rect 248788 304234 248840 304240
rect 248696 9784 248748 9790
rect 248696 9726 248748 9732
rect 248788 3528 248840 3534
rect 248788 3470 248840 3476
rect 247684 3052 247736 3058
rect 247684 2994 247736 3000
rect 248800 480 248828 3470
rect 249076 2922 249104 337878
rect 249168 330274 249196 338014
rect 249306 337770 249334 338028
rect 249260 337742 249334 337770
rect 249444 338014 249504 338042
rect 249156 330268 249208 330274
rect 249156 330210 249208 330216
rect 249260 329526 249288 337742
rect 249248 329520 249300 329526
rect 249248 329462 249300 329468
rect 249444 316034 249472 338014
rect 249582 337770 249610 338028
rect 249536 337742 249610 337770
rect 249720 338014 249780 338042
rect 249536 334626 249564 337742
rect 249616 336184 249668 336190
rect 249616 336126 249668 336132
rect 249524 334620 249576 334626
rect 249524 334562 249576 334568
rect 249628 325694 249656 336126
rect 249720 327214 249748 338014
rect 249858 337906 249886 338028
rect 249812 337878 249886 337906
rect 249996 338014 250056 338042
rect 249812 336462 249840 337878
rect 249800 336456 249852 336462
rect 249800 336398 249852 336404
rect 249996 334762 250024 338014
rect 250134 337770 250162 338028
rect 250088 337742 250162 337770
rect 250272 338014 250332 338042
rect 249984 334756 250036 334762
rect 249984 334698 250036 334704
rect 250088 330562 250116 337742
rect 250272 331214 250300 338014
rect 250410 337770 250438 338028
rect 249904 330534 250116 330562
rect 250180 331186 250300 331214
rect 250364 337742 250438 337770
rect 250548 338014 250608 338042
rect 249708 327208 249760 327214
rect 249708 327150 249760 327156
rect 249628 325666 249748 325694
rect 249168 316006 249472 316034
rect 249064 2916 249116 2922
rect 249064 2858 249116 2864
rect 249168 2854 249196 316006
rect 249720 3534 249748 325666
rect 249904 325038 249932 330534
rect 249984 330472 250036 330478
rect 249984 330414 250036 330420
rect 250076 330472 250128 330478
rect 250076 330414 250128 330420
rect 249892 325032 249944 325038
rect 249892 324974 249944 324980
rect 249996 6186 250024 330414
rect 250088 7886 250116 330414
rect 250076 7880 250128 7886
rect 250076 7822 250128 7828
rect 250180 7818 250208 331186
rect 250260 330540 250312 330546
rect 250260 330482 250312 330488
rect 250272 309874 250300 330482
rect 250260 309868 250312 309874
rect 250260 309810 250312 309816
rect 250168 7812 250220 7818
rect 250168 7754 250220 7760
rect 249984 6180 250036 6186
rect 249984 6122 250036 6128
rect 250364 5166 250392 337742
rect 250548 330750 250576 338014
rect 250686 337770 250714 338028
rect 250640 337742 250714 337770
rect 250824 338014 250884 338042
rect 251008 338014 251068 338042
rect 250536 330744 250588 330750
rect 250536 330686 250588 330692
rect 250640 330682 250668 337742
rect 250824 331214 250852 338014
rect 250732 331186 250852 331214
rect 250628 330676 250680 330682
rect 250628 330618 250680 330624
rect 250732 330562 250760 331186
rect 250456 330534 250760 330562
rect 250456 5574 250484 330534
rect 251008 322386 251036 338014
rect 251146 337770 251174 338028
rect 251100 337742 251174 337770
rect 251284 338014 251344 338042
rect 251100 330546 251128 337742
rect 251284 332042 251312 338014
rect 251422 337770 251450 338028
rect 251606 337822 251634 338028
rect 251594 337816 251646 337822
rect 251422 337742 251496 337770
rect 251594 337758 251646 337764
rect 251698 337770 251726 338028
rect 251836 338014 251896 338042
rect 251698 337742 251772 337770
rect 251468 337634 251496 337742
rect 251468 337606 251588 337634
rect 251456 334552 251508 334558
rect 251456 334494 251508 334500
rect 251272 332036 251324 332042
rect 251272 331978 251324 331984
rect 251088 330540 251140 330546
rect 251088 330482 251140 330488
rect 250996 322380 251048 322386
rect 250996 322322 251048 322328
rect 251468 318238 251496 334494
rect 251560 321026 251588 337606
rect 251744 334370 251772 337742
rect 251836 334558 251864 338014
rect 251974 337906 252002 338028
rect 252112 338014 252172 338042
rect 251974 337878 252048 337906
rect 251916 337816 251968 337822
rect 251916 337758 251968 337764
rect 251824 334552 251876 334558
rect 251824 334494 251876 334500
rect 251744 334342 251864 334370
rect 251640 333260 251692 333266
rect 251640 333202 251692 333208
rect 251548 321020 251600 321026
rect 251548 320962 251600 320968
rect 251456 318232 251508 318238
rect 251456 318174 251508 318180
rect 251652 8770 251680 333202
rect 251732 330472 251784 330478
rect 251732 330414 251784 330420
rect 251640 8764 251692 8770
rect 251640 8706 251692 8712
rect 251744 8702 251772 330414
rect 251836 329254 251864 334342
rect 251824 329248 251876 329254
rect 251824 329190 251876 329196
rect 251928 329202 251956 337758
rect 252020 333266 252048 337878
rect 252112 333402 252140 338014
rect 252250 337770 252278 338028
rect 252204 337742 252278 337770
rect 252388 338014 252448 338042
rect 252572 338014 252632 338042
rect 252100 333396 252152 333402
rect 252100 333338 252152 333344
rect 252008 333260 252060 333266
rect 252008 333202 252060 333208
rect 251928 329174 252048 329202
rect 252020 328930 252048 329174
rect 251928 328902 252048 328930
rect 251928 19990 251956 328902
rect 252204 323746 252232 337742
rect 252388 330478 252416 338014
rect 252468 336116 252520 336122
rect 252468 336058 252520 336064
rect 252376 330472 252428 330478
rect 252376 330414 252428 330420
rect 252192 323740 252244 323746
rect 252192 323682 252244 323688
rect 251916 19984 251968 19990
rect 251916 19926 251968 19932
rect 251732 8696 251784 8702
rect 251732 8638 251784 8644
rect 252480 6914 252508 336058
rect 252572 330818 252600 338014
rect 252710 337770 252738 338028
rect 252848 338014 252908 338042
rect 252710 337742 252784 337770
rect 252652 334620 252704 334626
rect 252652 334562 252704 334568
rect 252560 330812 252612 330818
rect 252560 330754 252612 330760
rect 252664 326534 252692 334562
rect 252756 330342 252784 337742
rect 252848 330546 252876 338014
rect 252986 337770 253014 338028
rect 252940 337742 253014 337770
rect 253124 338014 253184 338042
rect 252836 330540 252888 330546
rect 252836 330482 252888 330488
rect 252744 330336 252796 330342
rect 252744 330278 252796 330284
rect 252940 328522 252968 337742
rect 253124 334642 253152 338014
rect 253262 337770 253290 338028
rect 253400 338014 253460 338042
rect 253262 337742 253336 337770
rect 253204 336320 253256 336326
rect 253204 336262 253256 336268
rect 252756 328494 252968 328522
rect 253032 334614 253152 334642
rect 252756 327894 252784 328494
rect 253032 328454 253060 334614
rect 253216 331214 253244 336262
rect 253124 331186 253244 331214
rect 253124 330562 253152 331186
rect 253124 330534 253244 330562
rect 253112 330472 253164 330478
rect 253112 330414 253164 330420
rect 252836 328432 252888 328438
rect 252836 328374 252888 328380
rect 252940 328426 253060 328454
rect 252744 327888 252796 327894
rect 252744 327830 252796 327836
rect 252652 326528 252704 326534
rect 252652 326470 252704 326476
rect 252848 315450 252876 328374
rect 252940 316878 252968 328426
rect 253020 328364 253072 328370
rect 253020 328306 253072 328312
rect 252928 316872 252980 316878
rect 252928 316814 252980 316820
rect 252836 315444 252888 315450
rect 252836 315386 252888 315392
rect 253032 8498 253060 328306
rect 253124 8566 253152 330414
rect 253216 10402 253244 330534
rect 253308 330478 253336 337742
rect 253400 334626 253428 338014
rect 253538 337770 253566 338028
rect 253492 337742 253566 337770
rect 253676 338014 253736 338042
rect 253388 334620 253440 334626
rect 253388 334562 253440 334568
rect 253388 330540 253440 330546
rect 253388 330482 253440 330488
rect 253296 330472 253348 330478
rect 253296 330414 253348 330420
rect 253296 330336 253348 330342
rect 253296 330278 253348 330284
rect 253308 325106 253336 330278
rect 253296 325100 253348 325106
rect 253296 325042 253348 325048
rect 253204 10396 253256 10402
rect 253204 10338 253256 10344
rect 253400 8634 253428 330482
rect 253492 328438 253520 337742
rect 253480 328432 253532 328438
rect 253480 328374 253532 328380
rect 253676 328370 253704 338014
rect 253814 337770 253842 338028
rect 253998 337822 254026 338028
rect 253986 337816 254038 337822
rect 253814 337742 253888 337770
rect 253986 337758 254038 337764
rect 254090 337770 254118 338028
rect 254228 338014 254288 338042
rect 254412 338014 254472 338042
rect 254090 337742 254164 337770
rect 253860 334830 253888 337742
rect 253848 334824 253900 334830
rect 253848 334766 253900 334772
rect 254136 328454 254164 337742
rect 254228 335918 254256 338014
rect 254216 335912 254268 335918
rect 254216 335854 254268 335860
rect 254412 332110 254440 338014
rect 254550 337906 254578 338028
rect 254688 338014 254748 338042
rect 254550 337878 254624 337906
rect 254492 337816 254544 337822
rect 254492 337758 254544 337764
rect 254400 332104 254452 332110
rect 254400 332046 254452 332052
rect 254136 328426 254348 328454
rect 253664 328364 253716 328370
rect 253664 328306 253716 328312
rect 254320 308514 254348 328426
rect 254504 327962 254532 337758
rect 254596 331106 254624 337878
rect 254688 336734 254716 338014
rect 254826 337770 254854 338028
rect 254964 338014 255024 338042
rect 254826 337742 254900 337770
rect 254676 336728 254728 336734
rect 254676 336670 254728 336676
rect 254596 331078 254716 331106
rect 254584 329044 254636 329050
rect 254584 328986 254636 328992
rect 254492 327956 254544 327962
rect 254492 327898 254544 327904
rect 254400 326392 254452 326398
rect 254400 326334 254452 326340
rect 254412 312662 254440 326334
rect 254400 312656 254452 312662
rect 254400 312598 254452 312604
rect 254308 308508 254360 308514
rect 254308 308450 254360 308456
rect 254596 11830 254624 328986
rect 254688 314022 254716 331078
rect 254872 329322 254900 337742
rect 254860 329316 254912 329322
rect 254860 329258 254912 329264
rect 254964 326398 254992 338014
rect 255102 337770 255130 338028
rect 255240 338014 255300 338042
rect 255102 337742 255176 337770
rect 255148 333470 255176 337742
rect 255136 333464 255188 333470
rect 255136 333406 255188 333412
rect 254952 326392 255004 326398
rect 254952 326334 255004 326340
rect 255240 323814 255268 338014
rect 255378 337770 255406 338028
rect 255516 338014 255576 338042
rect 255378 337742 255452 337770
rect 255320 335368 255372 335374
rect 255320 335310 255372 335316
rect 255332 333538 255360 335310
rect 255320 333532 255372 333538
rect 255320 333474 255372 333480
rect 255424 326398 255452 337742
rect 255516 336394 255544 338014
rect 255654 337822 255682 338028
rect 255792 338014 255852 338042
rect 255642 337816 255694 337822
rect 255642 337758 255694 337764
rect 255504 336388 255556 336394
rect 255504 336330 255556 336336
rect 255792 331214 255820 338014
rect 255930 337770 255958 338028
rect 256068 338014 256128 338042
rect 256252 338014 256312 338042
rect 255930 337742 256004 337770
rect 255872 335912 255924 335918
rect 255872 335854 255924 335860
rect 255516 331186 255820 331214
rect 255884 331214 255912 335854
rect 255976 334898 256004 337742
rect 255964 334892 256016 334898
rect 255964 334834 256016 334840
rect 255884 331186 256004 331214
rect 255412 326392 255464 326398
rect 255412 326334 255464 326340
rect 255412 326256 255464 326262
rect 255412 326198 255464 326204
rect 255516 326210 255544 331186
rect 255780 326392 255832 326398
rect 255780 326334 255832 326340
rect 255228 323808 255280 323814
rect 255228 323750 255280 323756
rect 254676 314016 254728 314022
rect 254676 313958 254728 313964
rect 254584 11824 254636 11830
rect 254584 11766 254636 11772
rect 253480 9648 253532 9654
rect 253480 9590 253532 9596
rect 253388 8628 253440 8634
rect 253388 8570 253440 8576
rect 253112 8560 253164 8566
rect 253112 8502 253164 8508
rect 253020 8492 253072 8498
rect 253020 8434 253072 8440
rect 252388 6886 252508 6914
rect 250444 5568 250496 5574
rect 250444 5510 250496 5516
rect 250352 5160 250404 5166
rect 250352 5102 250404 5108
rect 249984 5092 250036 5098
rect 249984 5034 250036 5040
rect 249708 3528 249760 3534
rect 249708 3470 249760 3476
rect 249156 2848 249208 2854
rect 249156 2790 249208 2796
rect 249996 480 250024 5034
rect 251180 3460 251232 3466
rect 251180 3402 251232 3408
rect 251192 480 251220 3402
rect 252388 480 252416 6886
rect 253492 480 253520 9590
rect 255424 6322 255452 326198
rect 255516 326182 255636 326210
rect 255504 326120 255556 326126
rect 255504 326062 255556 326068
rect 255516 6390 255544 326062
rect 255608 8022 255636 326182
rect 255688 326188 255740 326194
rect 255688 326130 255740 326136
rect 255700 8158 255728 326130
rect 255688 8152 255740 8158
rect 255688 8094 255740 8100
rect 255596 8016 255648 8022
rect 255596 7958 255648 7964
rect 255792 7954 255820 326334
rect 255872 322448 255924 322454
rect 255872 322390 255924 322396
rect 255884 8090 255912 322390
rect 255976 9654 256004 331186
rect 256068 326262 256096 338014
rect 256148 337816 256200 337822
rect 256148 337758 256200 337764
rect 256056 326256 256108 326262
rect 256056 326198 256108 326204
rect 255964 9648 256016 9654
rect 255964 9590 256016 9596
rect 255872 8084 255924 8090
rect 255872 8026 255924 8032
rect 255780 7948 255832 7954
rect 255780 7890 255832 7896
rect 255504 6384 255556 6390
rect 255504 6326 255556 6332
rect 255412 6316 255464 6322
rect 255412 6258 255464 6264
rect 256160 6254 256188 337758
rect 256252 322454 256280 338014
rect 256390 337770 256418 338028
rect 256528 338014 256588 338042
rect 256390 337742 256464 337770
rect 256436 330954 256464 337742
rect 256424 330948 256476 330954
rect 256424 330890 256476 330896
rect 256528 326126 256556 338014
rect 256666 337770 256694 338028
rect 256620 337742 256694 337770
rect 256804 338014 256864 338042
rect 256620 326194 256648 337742
rect 256804 335374 256832 338014
rect 256942 337770 256970 338028
rect 257126 337770 257154 338028
rect 257218 337890 257246 338028
rect 257206 337884 257258 337890
rect 257206 337826 257258 337832
rect 257402 337770 257430 338028
rect 257494 337906 257522 338028
rect 257632 338014 257692 338042
rect 257816 338014 257876 338042
rect 257494 337878 257568 337906
rect 256942 337742 257016 337770
rect 257126 337742 257200 337770
rect 257402 337742 257476 337770
rect 256792 335368 256844 335374
rect 256792 335310 256844 335316
rect 256988 328030 257016 337742
rect 256976 328024 257028 328030
rect 256976 327966 257028 327972
rect 257068 326392 257120 326398
rect 257068 326334 257120 326340
rect 256608 326188 256660 326194
rect 256608 326130 256660 326136
rect 256516 326120 256568 326126
rect 256516 326062 256568 326068
rect 256240 322448 256292 322454
rect 256240 322390 256292 322396
rect 257080 311234 257108 326334
rect 257172 322522 257200 337742
rect 257344 335436 257396 335442
rect 257344 335378 257396 335384
rect 257160 322516 257212 322522
rect 257160 322458 257212 322464
rect 257068 311228 257120 311234
rect 257068 311170 257120 311176
rect 257356 11762 257384 335378
rect 257448 331022 257476 337742
rect 257436 331016 257488 331022
rect 257436 330958 257488 330964
rect 257540 329390 257568 337878
rect 257632 335986 257660 338014
rect 257620 335980 257672 335986
rect 257620 335922 257672 335928
rect 257528 329384 257580 329390
rect 257528 329326 257580 329332
rect 257816 326602 257844 338014
rect 257954 337770 257982 338028
rect 257908 337742 257982 337770
rect 258092 338014 258152 338042
rect 257804 326596 257856 326602
rect 257804 326538 257856 326544
rect 257908 326398 257936 337742
rect 257896 326392 257948 326398
rect 257896 326334 257948 326340
rect 257344 11756 257396 11762
rect 257344 11698 257396 11704
rect 256148 6248 256200 6254
rect 256148 6190 256200 6196
rect 258092 5234 258120 338014
rect 258230 337906 258258 338028
rect 258368 338014 258428 338042
rect 258230 337878 258304 337906
rect 258172 337816 258224 337822
rect 258172 337758 258224 337764
rect 258184 326346 258212 337758
rect 258276 326482 258304 337878
rect 258368 333266 258396 338014
rect 258506 337770 258534 338028
rect 258460 337742 258534 337770
rect 258644 338014 258704 338042
rect 258356 333260 258408 333266
rect 258356 333202 258408 333208
rect 258460 326602 258488 337742
rect 258448 326596 258500 326602
rect 258448 326538 258500 326544
rect 258276 326454 258580 326482
rect 258356 326392 258408 326398
rect 258184 326318 258304 326346
rect 258356 326334 258408 326340
rect 258448 326392 258500 326398
rect 258448 326334 258500 326340
rect 258172 326256 258224 326262
rect 258172 326198 258224 326204
rect 258184 5302 258212 326198
rect 258276 5438 258304 326318
rect 258264 5432 258316 5438
rect 258264 5374 258316 5380
rect 258368 5370 258396 326334
rect 258460 6594 258488 326334
rect 258448 6588 258500 6594
rect 258448 6530 258500 6536
rect 258552 6458 258580 326454
rect 258644 6526 258672 338014
rect 258782 337906 258810 338028
rect 258920 338014 258980 338042
rect 258782 337878 258856 337906
rect 258724 333260 258776 333266
rect 258724 333202 258776 333208
rect 258736 8226 258764 333202
rect 258828 326330 258856 337878
rect 258920 326466 258948 338014
rect 259058 337770 259086 338028
rect 259012 337742 259086 337770
rect 259196 338014 259256 338042
rect 258908 326460 258960 326466
rect 258908 326402 258960 326408
rect 259012 326398 259040 337742
rect 259196 331214 259224 338014
rect 259334 337822 259362 338028
rect 259322 337816 259374 337822
rect 259322 337758 259374 337764
rect 259518 337770 259546 338028
rect 259656 338014 259716 338042
rect 259518 337742 259592 337770
rect 259104 331186 259224 331214
rect 259000 326392 259052 326398
rect 259000 326334 259052 326340
rect 258816 326324 258868 326330
rect 258816 326266 258868 326272
rect 259104 326210 259132 331186
rect 259564 326398 259592 337742
rect 259656 326466 259684 338014
rect 259794 337770 259822 338028
rect 259748 337742 259822 337770
rect 259932 338014 259992 338042
rect 259644 326460 259696 326466
rect 259644 326402 259696 326408
rect 259552 326392 259604 326398
rect 259748 326346 259776 337742
rect 259552 326334 259604 326340
rect 258828 326182 259132 326210
rect 259656 326318 259776 326346
rect 259828 326324 259880 326330
rect 259552 326188 259604 326194
rect 258724 8220 258776 8226
rect 258724 8162 258776 8168
rect 258828 7546 258856 326182
rect 259552 326130 259604 326136
rect 258908 326120 258960 326126
rect 258908 326062 258960 326068
rect 258920 8294 258948 326062
rect 258908 8288 258960 8294
rect 258908 8230 258960 8236
rect 258816 7540 258868 7546
rect 258816 7482 258868 7488
rect 258632 6520 258684 6526
rect 258632 6462 258684 6468
rect 258540 6452 258592 6458
rect 258540 6394 258592 6400
rect 258356 5364 258408 5370
rect 258356 5306 258408 5312
rect 258172 5296 258224 5302
rect 258172 5238 258224 5244
rect 258080 5228 258132 5234
rect 258080 5170 258132 5176
rect 259564 4690 259592 326130
rect 259656 5506 259684 326318
rect 259828 326266 259880 326272
rect 259736 326256 259788 326262
rect 259736 326198 259788 326204
rect 259748 6798 259776 326198
rect 259840 6866 259868 326266
rect 259828 6860 259880 6866
rect 259828 6802 259880 6808
rect 259736 6792 259788 6798
rect 259736 6734 259788 6740
rect 259932 6730 259960 338014
rect 260070 337872 260098 338028
rect 260024 337844 260098 337872
rect 260208 338014 260268 338042
rect 260024 334966 260052 337844
rect 260012 334960 260064 334966
rect 260012 334902 260064 334908
rect 260104 326460 260156 326466
rect 260104 326402 260156 326408
rect 260012 326392 260064 326398
rect 260012 326334 260064 326340
rect 259920 6724 259972 6730
rect 259920 6666 259972 6672
rect 260024 6662 260052 326334
rect 260116 7478 260144 326402
rect 260104 7472 260156 7478
rect 260104 7414 260156 7420
rect 260012 6656 260064 6662
rect 260012 6598 260064 6604
rect 259644 5500 259696 5506
rect 259644 5442 259696 5448
rect 260208 4758 260236 338014
rect 260346 337770 260374 338028
rect 260300 337742 260374 337770
rect 260484 338014 260544 338042
rect 260300 326262 260328 337742
rect 260484 330886 260512 338014
rect 260622 337770 260650 338028
rect 260576 337742 260650 337770
rect 260760 338014 260820 338042
rect 260472 330880 260524 330886
rect 260472 330822 260524 330828
rect 260288 326256 260340 326262
rect 260288 326198 260340 326204
rect 260576 326194 260604 337742
rect 260760 326330 260788 338014
rect 260898 337770 260926 338028
rect 261036 338014 261096 338042
rect 260898 337742 260972 337770
rect 260944 328454 260972 337742
rect 261036 335374 261064 338014
rect 261174 337906 261202 338028
rect 261128 337878 261202 337906
rect 261312 338014 261372 338042
rect 261496 338014 261556 338042
rect 261024 335368 261076 335374
rect 261024 335310 261076 335316
rect 261128 333606 261156 337878
rect 261116 333600 261168 333606
rect 261116 333542 261168 333548
rect 260944 328426 261156 328454
rect 261128 326670 261156 328426
rect 261116 326664 261168 326670
rect 261116 326606 261168 326612
rect 260748 326324 260800 326330
rect 260748 326266 260800 326272
rect 260564 326188 260616 326194
rect 260564 326130 260616 326136
rect 261312 319530 261340 338014
rect 261392 337816 261444 337822
rect 261392 337758 261444 337764
rect 261404 321094 261432 337758
rect 261496 336530 261524 338014
rect 261634 337940 261662 338028
rect 261772 338014 261832 338042
rect 261634 337912 261708 337940
rect 261484 336524 261536 336530
rect 261484 336466 261536 336472
rect 261484 336320 261536 336326
rect 261484 336262 261536 336268
rect 261392 321088 261444 321094
rect 261392 321030 261444 321036
rect 261300 319524 261352 319530
rect 261300 319466 261352 319472
rect 261496 10334 261524 336262
rect 261576 335368 261628 335374
rect 261576 335310 261628 335316
rect 261588 13122 261616 335310
rect 261680 332178 261708 337912
rect 261668 332172 261720 332178
rect 261668 332114 261720 332120
rect 261772 325174 261800 338014
rect 261910 337906 261938 338028
rect 261864 337878 261938 337906
rect 262048 338014 262108 338042
rect 261864 334898 261892 337878
rect 261852 334892 261904 334898
rect 261852 334834 261904 334840
rect 262048 329458 262076 338014
rect 262186 337822 262214 338028
rect 262174 337816 262226 337822
rect 262174 337758 262226 337764
rect 262370 337770 262398 338028
rect 262462 337958 262490 338028
rect 262450 337952 262502 337958
rect 262450 337894 262502 337900
rect 262496 337816 262548 337822
rect 262370 337742 262444 337770
rect 262496 337758 262548 337764
rect 262646 337770 262674 338028
rect 262738 337872 262766 338028
rect 262876 338014 262936 338042
rect 263060 338014 263120 338042
rect 262738 337844 262812 337872
rect 262312 337680 262364 337686
rect 262312 337622 262364 337628
rect 262324 333674 262352 337622
rect 262312 333668 262364 333674
rect 262312 333610 262364 333616
rect 262036 329452 262088 329458
rect 262036 329394 262088 329400
rect 261760 325168 261812 325174
rect 261760 325110 261812 325116
rect 261576 13116 261628 13122
rect 261576 13058 261628 13064
rect 261484 10328 261536 10334
rect 261484 10270 261536 10276
rect 260196 4752 260248 4758
rect 260196 4694 260248 4700
rect 259552 4684 259604 4690
rect 259552 4626 259604 4632
rect 262416 4622 262444 337742
rect 262508 8974 262536 337758
rect 262646 337742 262720 337770
rect 262692 328098 262720 337742
rect 262680 328092 262732 328098
rect 262680 328034 262732 328040
rect 262588 326392 262640 326398
rect 262588 326334 262640 326340
rect 262496 8968 262548 8974
rect 262496 8910 262548 8916
rect 262600 4826 262628 326334
rect 262588 4820 262640 4826
rect 262588 4762 262640 4768
rect 262404 4616 262456 4622
rect 262404 4558 262456 4564
rect 262784 4554 262812 337844
rect 262876 332246 262904 338014
rect 262956 336728 263008 336734
rect 262956 336670 263008 336676
rect 262864 332240 262916 332246
rect 262864 332182 262916 332188
rect 262968 316034 262996 336670
rect 263060 335374 263088 338014
rect 263198 337770 263226 338028
rect 263152 337742 263226 337770
rect 263336 338014 263396 338042
rect 263048 335368 263100 335374
rect 263048 335310 263100 335316
rect 263152 326398 263180 337742
rect 263336 335442 263364 338014
rect 263474 337822 263502 338028
rect 263462 337816 263514 337822
rect 263462 337758 263514 337764
rect 263658 337770 263686 338028
rect 263750 337906 263778 338028
rect 263750 337878 263824 337906
rect 263658 337742 263732 337770
rect 263324 335436 263376 335442
rect 263324 335378 263376 335384
rect 263704 330410 263732 337742
rect 263796 336462 263824 337878
rect 263934 337770 263962 338028
rect 264026 337872 264054 338028
rect 264164 338014 264224 338042
rect 264026 337844 264100 337872
rect 263934 337742 264008 337770
rect 263784 336456 263836 336462
rect 263784 336398 263836 336404
rect 263980 336326 264008 337742
rect 263968 336320 264020 336326
rect 263968 336262 264020 336268
rect 264072 336172 264100 337844
rect 264164 336258 264192 338014
rect 264302 337906 264330 338028
rect 264256 337878 264330 337906
rect 264440 338014 264500 338042
rect 264152 336252 264204 336258
rect 264152 336194 264204 336200
rect 263888 336144 264100 336172
rect 263784 330676 263836 330682
rect 263784 330618 263836 330624
rect 263692 330404 263744 330410
rect 263692 330346 263744 330352
rect 263140 326392 263192 326398
rect 263140 326334 263192 326340
rect 262876 316006 262996 316034
rect 262772 4548 262824 4554
rect 262772 4490 262824 4496
rect 262876 3806 262904 316006
rect 263796 5030 263824 330618
rect 263784 5024 263836 5030
rect 263784 4966 263836 4972
rect 263888 4962 263916 336144
rect 264256 336054 264284 337878
rect 264244 336048 264296 336054
rect 264244 335990 264296 335996
rect 264440 330682 264468 338014
rect 264578 337770 264606 338028
rect 264532 337742 264606 337770
rect 264716 338014 264776 338042
rect 264900 338014 264960 338042
rect 264428 330676 264480 330682
rect 264428 330618 264480 330624
rect 264532 330528 264560 337742
rect 264716 336190 264744 338014
rect 264704 336184 264756 336190
rect 264704 336126 264756 336132
rect 263980 330500 264560 330528
rect 263980 9042 264008 330500
rect 264060 330404 264112 330410
rect 264060 330346 264112 330352
rect 263968 9036 264020 9042
rect 263968 8978 264020 8984
rect 263876 4956 263928 4962
rect 263876 4898 263928 4904
rect 264072 4894 264100 330346
rect 264900 316034 264928 338014
rect 265038 337770 265066 338028
rect 265176 338014 265236 338042
rect 265038 337742 265112 337770
rect 265084 335322 265112 337742
rect 265176 335986 265204 338014
rect 265314 337872 265342 338028
rect 265268 337844 265342 337872
rect 265452 338014 265512 338042
rect 265268 336122 265296 337844
rect 265256 336116 265308 336122
rect 265256 336058 265308 336064
rect 265164 335980 265216 335986
rect 265164 335922 265216 335928
rect 265084 335294 265296 335322
rect 265072 334552 265124 334558
rect 265072 334494 265124 334500
rect 264440 316006 264928 316034
rect 264440 5098 264468 316006
rect 264428 5092 264480 5098
rect 264428 5034 264480 5040
rect 264060 4888 264112 4894
rect 264060 4830 264112 4836
rect 262864 3800 262916 3806
rect 262864 3742 262916 3748
rect 257068 3732 257120 3738
rect 257068 3674 257120 3680
rect 259460 3732 259512 3738
rect 259460 3674 259512 3680
rect 255872 3596 255924 3602
rect 255872 3538 255924 3544
rect 254676 3528 254728 3534
rect 254676 3470 254728 3476
rect 254688 480 254716 3470
rect 255884 480 255912 3538
rect 257080 480 257108 3674
rect 258264 2984 258316 2990
rect 258264 2926 258316 2932
rect 258276 480 258304 2926
rect 259472 480 259500 3674
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 260668 480 260696 3470
rect 261760 3256 261812 3262
rect 261760 3198 261812 3204
rect 261772 480 261800 3198
rect 262968 480 262996 3606
rect 264152 3596 264204 3602
rect 264152 3538 264204 3544
rect 264164 480 264192 3538
rect 265084 3534 265112 334494
rect 265164 330608 265216 330614
rect 265164 330550 265216 330556
rect 265072 3528 265124 3534
rect 265072 3470 265124 3476
rect 265176 2990 265204 330550
rect 265268 3466 265296 335294
rect 265348 330472 265400 330478
rect 265348 330414 265400 330420
rect 265360 3738 265388 330414
rect 265452 3874 265480 338014
rect 265590 337770 265618 338028
rect 265728 338014 265788 338042
rect 265590 337742 265664 337770
rect 265532 330540 265584 330546
rect 265532 330482 265584 330488
rect 265440 3868 265492 3874
rect 265440 3810 265492 3816
rect 265348 3732 265400 3738
rect 265348 3674 265400 3680
rect 265256 3460 265308 3466
rect 265256 3402 265308 3408
rect 265348 3460 265400 3466
rect 265348 3402 265400 3408
rect 265164 2984 265216 2990
rect 265164 2926 265216 2932
rect 265360 480 265388 3402
rect 265544 3262 265572 330482
rect 265636 3806 265664 337742
rect 265728 336734 265756 338014
rect 265866 337770 265894 338028
rect 265820 337742 265894 337770
rect 266004 338014 266064 338042
rect 265716 336728 265768 336734
rect 265716 336670 265768 336676
rect 265820 330614 265848 337742
rect 265808 330608 265860 330614
rect 265808 330550 265860 330556
rect 266004 330478 266032 338014
rect 266142 337770 266170 338028
rect 266096 337742 266170 337770
rect 266280 338014 266340 338042
rect 266096 334558 266124 337742
rect 266084 334552 266136 334558
rect 266084 334494 266136 334500
rect 266280 330546 266308 338014
rect 266418 337770 266446 338028
rect 266602 337770 266630 338028
rect 266740 338014 266800 338042
rect 266418 337742 266492 337770
rect 266602 337742 266676 337770
rect 266268 330540 266320 330546
rect 266268 330482 266320 330488
rect 265992 330472 266044 330478
rect 265992 330414 266044 330420
rect 266464 328454 266492 337742
rect 266648 333266 266676 337742
rect 266636 333260 266688 333266
rect 266636 333202 266688 333208
rect 266464 328426 266584 328454
rect 265624 3800 265676 3806
rect 265624 3742 265676 3748
rect 266556 3670 266584 328426
rect 266740 316034 266768 338014
rect 266878 337770 266906 338028
rect 267016 338014 267076 338042
rect 266878 337742 266952 337770
rect 266924 335322 266952 337742
rect 267016 335442 267044 338014
rect 267154 337770 267182 338028
rect 267338 337770 267366 338028
rect 267430 337872 267458 338028
rect 267568 338014 267628 338042
rect 267430 337844 267504 337872
rect 267154 337742 267228 337770
rect 267338 337742 267412 337770
rect 267004 335436 267056 335442
rect 267004 335378 267056 335384
rect 266924 335294 267136 335322
rect 266912 333260 266964 333266
rect 266912 333202 266964 333208
rect 266648 316006 266768 316034
rect 266544 3664 266596 3670
rect 266544 3606 266596 3612
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 265532 3256 265584 3262
rect 265532 3198 265584 3204
rect 266556 480 266584 3470
rect 266648 3466 266676 316006
rect 266924 3602 266952 333202
rect 266912 3596 266964 3602
rect 266912 3538 266964 3544
rect 267108 3534 267136 335294
rect 267200 333266 267228 337742
rect 267188 333260 267240 333266
rect 267188 333202 267240 333208
rect 267384 6914 267412 337742
rect 267476 335782 267504 337844
rect 267464 335776 267516 335782
rect 267464 335718 267516 335724
rect 267568 335578 267596 338014
rect 267706 337770 267734 338028
rect 267660 337742 267734 337770
rect 267844 338014 267904 338042
rect 267556 335572 267608 335578
rect 267556 335514 267608 335520
rect 267556 335436 267608 335442
rect 267556 335378 267608 335384
rect 267464 333260 267516 333266
rect 267464 333202 267516 333208
rect 267292 6886 267412 6914
rect 267096 3528 267148 3534
rect 267096 3470 267148 3476
rect 267292 3466 267320 6886
rect 267476 5658 267504 333202
rect 267384 5630 267504 5658
rect 267384 4146 267412 5630
rect 267568 5522 267596 335378
rect 267476 5494 267596 5522
rect 267372 4140 267424 4146
rect 267372 4082 267424 4088
rect 267476 4078 267504 5494
rect 267660 5250 267688 337742
rect 267844 335374 267872 338014
rect 267982 337822 268010 338028
rect 267970 337816 268022 337822
rect 267970 337758 268022 337764
rect 268166 337770 268194 338028
rect 268304 338014 268364 338042
rect 268166 337742 268240 337770
rect 267832 335368 267884 335374
rect 267832 335310 267884 335316
rect 268212 333266 268240 337742
rect 268304 335442 268332 338014
rect 268442 337770 268470 338028
rect 268580 338014 268640 338042
rect 268442 337742 268516 337770
rect 268488 335918 268516 337742
rect 268476 335912 268528 335918
rect 268476 335854 268528 335860
rect 268580 335850 268608 338014
rect 268718 337770 268746 338028
rect 268672 337742 268746 337770
rect 268856 338014 268916 338042
rect 268568 335844 268620 335850
rect 268568 335786 268620 335792
rect 268384 335572 268436 335578
rect 268384 335514 268436 335520
rect 268292 335436 268344 335442
rect 268292 335378 268344 335384
rect 268200 333260 268252 333266
rect 268200 333202 268252 333208
rect 267568 5222 267688 5250
rect 267464 4072 267516 4078
rect 267464 4014 267516 4020
rect 267568 3738 267596 5222
rect 267648 4072 267700 4078
rect 267700 4020 267780 4026
rect 267648 4014 267780 4020
rect 267660 3998 267780 4014
rect 267556 3732 267608 3738
rect 267556 3674 267608 3680
rect 266636 3460 266688 3466
rect 266636 3402 266688 3408
rect 267280 3460 267332 3466
rect 267280 3402 267332 3408
rect 267752 480 267780 3998
rect 268396 3534 268424 335514
rect 268568 335368 268620 335374
rect 268568 335310 268620 335316
rect 268476 333396 268528 333402
rect 268476 333338 268528 333344
rect 268488 13122 268516 333338
rect 268476 13116 268528 13122
rect 268476 13058 268528 13064
rect 268580 5642 268608 335310
rect 268568 5636 268620 5642
rect 268568 5578 268620 5584
rect 268672 4622 268700 337742
rect 268752 335436 268804 335442
rect 268752 335378 268804 335384
rect 268660 4616 268712 4622
rect 268660 4558 268712 4564
rect 268764 4554 268792 335378
rect 268856 4690 268884 338014
rect 268994 337906 269022 338028
rect 268994 337878 269068 337906
rect 268936 337816 268988 337822
rect 268936 337758 268988 337764
rect 268844 4684 268896 4690
rect 268844 4626 268896 4632
rect 268752 4548 268804 4554
rect 268752 4490 268804 4496
rect 268844 4140 268896 4146
rect 268844 4082 268896 4088
rect 268384 3528 268436 3534
rect 268384 3470 268436 3476
rect 268856 480 268884 4082
rect 268948 3194 268976 337758
rect 269040 333402 269068 337878
rect 269178 337770 269206 338028
rect 269270 337872 269298 338028
rect 269408 338014 269468 338042
rect 269270 337844 269344 337872
rect 269178 337742 269252 337770
rect 269224 334422 269252 337742
rect 269212 334416 269264 334422
rect 269212 334358 269264 334364
rect 269028 333396 269080 333402
rect 269028 333338 269080 333344
rect 269028 333260 269080 333266
rect 269028 333202 269080 333208
rect 269040 3330 269068 333202
rect 269316 330410 269344 337844
rect 269408 336122 269436 338014
rect 269546 337770 269574 338028
rect 269730 337770 269758 338028
rect 269822 337872 269850 338028
rect 270006 337940 270034 338028
rect 270144 338014 270204 338042
rect 270006 337912 270080 337940
rect 269822 337844 269988 337872
rect 269546 337742 269620 337770
rect 269730 337742 269896 337770
rect 269396 336116 269448 336122
rect 269396 336058 269448 336064
rect 269592 333266 269620 337742
rect 269580 333260 269632 333266
rect 269580 333202 269632 333208
rect 269304 330404 269356 330410
rect 269304 330346 269356 330352
rect 269868 5370 269896 337742
rect 269960 336054 269988 337844
rect 269948 336048 270000 336054
rect 269948 335990 270000 335996
rect 269948 335368 270000 335374
rect 269948 335310 270000 335316
rect 269960 334506 269988 335310
rect 270052 334642 270080 337912
rect 270144 334778 270172 338014
rect 270282 337770 270310 338028
rect 270236 337742 270310 337770
rect 270420 338014 270480 338042
rect 270236 336190 270264 337742
rect 270224 336184 270276 336190
rect 270224 336126 270276 336132
rect 270420 335374 270448 338014
rect 270558 337770 270586 338028
rect 270696 338014 270756 338042
rect 270558 337742 270632 337770
rect 270604 336172 270632 337742
rect 270696 336326 270724 338014
rect 270834 337872 270862 338028
rect 270834 337844 270908 337872
rect 270684 336320 270736 336326
rect 270684 336262 270736 336268
rect 270604 336144 270724 336172
rect 270500 335776 270552 335782
rect 270500 335718 270552 335724
rect 270408 335368 270460 335374
rect 270408 335310 270460 335316
rect 270144 334750 270356 334778
rect 270052 334614 270264 334642
rect 269960 334478 270080 334506
rect 269948 334416 270000 334422
rect 269948 334358 270000 334364
rect 269856 5364 269908 5370
rect 269856 5306 269908 5312
rect 269960 4758 269988 334358
rect 270052 5098 270080 334478
rect 270132 333260 270184 333266
rect 270132 333202 270184 333208
rect 270144 5438 270172 333202
rect 270132 5432 270184 5438
rect 270132 5374 270184 5380
rect 270236 5234 270264 334614
rect 270328 330682 270356 334750
rect 270512 331214 270540 335718
rect 270512 331186 270632 331214
rect 270316 330676 270368 330682
rect 270316 330618 270368 330624
rect 270408 330472 270460 330478
rect 270408 330414 270460 330420
rect 270316 330404 270368 330410
rect 270316 330346 270368 330352
rect 270328 5506 270356 330346
rect 270316 5500 270368 5506
rect 270316 5442 270368 5448
rect 270420 5302 270448 330414
rect 270604 16574 270632 331186
rect 270696 330478 270724 336144
rect 270880 333266 270908 337844
rect 271018 337770 271046 338028
rect 271110 337906 271138 338028
rect 271110 337878 271184 337906
rect 271018 337742 271092 337770
rect 270868 333260 270920 333266
rect 270868 333202 270920 333208
rect 270684 330472 270736 330478
rect 270684 330414 270736 330420
rect 271064 325694 271092 337742
rect 271156 336462 271184 337878
rect 271294 337770 271322 338028
rect 271386 337906 271414 338028
rect 271524 338014 271584 338042
rect 271386 337878 271460 337906
rect 271294 337742 271368 337770
rect 271144 336456 271196 336462
rect 271144 336398 271196 336404
rect 271340 330682 271368 337742
rect 271432 334626 271460 337878
rect 271524 335374 271552 338014
rect 271662 337822 271690 338028
rect 271800 338014 271860 338042
rect 271984 338014 272044 338042
rect 271650 337816 271702 337822
rect 271650 337758 271702 337764
rect 271800 335458 271828 338014
rect 271616 335430 271828 335458
rect 271512 335368 271564 335374
rect 271512 335310 271564 335316
rect 271420 334620 271472 334626
rect 271420 334562 271472 334568
rect 271616 334506 271644 335430
rect 271788 335368 271840 335374
rect 271788 335310 271840 335316
rect 271696 334620 271748 334626
rect 271696 334562 271748 334568
rect 271432 334478 271644 334506
rect 271328 330676 271380 330682
rect 271328 330618 271380 330624
rect 271432 330562 271460 334478
rect 271512 333260 271564 333266
rect 271512 333202 271564 333208
rect 271340 330534 271460 330562
rect 271064 325666 271276 325694
rect 270604 16546 271184 16574
rect 270408 5296 270460 5302
rect 270408 5238 270460 5244
rect 270224 5228 270276 5234
rect 270224 5170 270276 5176
rect 270040 5092 270092 5098
rect 270040 5034 270092 5040
rect 269948 4752 270000 4758
rect 269948 4694 270000 4700
rect 271156 3482 271184 16546
rect 271248 5030 271276 325666
rect 271340 8430 271368 330534
rect 271420 330472 271472 330478
rect 271420 330414 271472 330420
rect 271328 8424 271380 8430
rect 271328 8366 271380 8372
rect 271432 5166 271460 330414
rect 271420 5160 271472 5166
rect 271420 5102 271472 5108
rect 271236 5024 271288 5030
rect 271236 4966 271288 4972
rect 271524 4962 271552 333202
rect 271604 330676 271656 330682
rect 271604 330618 271656 330624
rect 271512 4956 271564 4962
rect 271512 4898 271564 4904
rect 271616 4894 271644 330618
rect 271604 4888 271656 4894
rect 271604 4830 271656 4836
rect 271708 4826 271736 334562
rect 271800 329186 271828 335310
rect 271984 335102 272012 338014
rect 272122 337906 272150 338028
rect 272260 338014 272320 338042
rect 272122 337878 272196 337906
rect 271972 335096 272024 335102
rect 271972 335038 272024 335044
rect 272168 335034 272196 337878
rect 272260 335442 272288 338014
rect 272398 337906 272426 338028
rect 272536 338014 272596 338042
rect 272398 337878 272472 337906
rect 272248 335436 272300 335442
rect 272248 335378 272300 335384
rect 272156 335028 272208 335034
rect 272156 334970 272208 334976
rect 272444 333266 272472 337878
rect 272536 336666 272564 338014
rect 272674 337906 272702 338028
rect 272812 338014 272872 338042
rect 272674 337878 272748 337906
rect 272524 336660 272576 336666
rect 272524 336602 272576 336608
rect 272616 335504 272668 335510
rect 272616 335446 272668 335452
rect 272432 333260 272484 333266
rect 272432 333202 272484 333208
rect 271788 329180 271840 329186
rect 271788 329122 271840 329128
rect 272628 8634 272656 335446
rect 272720 333402 272748 337878
rect 272708 333396 272760 333402
rect 272708 333338 272760 333344
rect 272708 333260 272760 333266
rect 272708 333202 272760 333208
rect 272720 325174 272748 333202
rect 272708 325168 272760 325174
rect 272708 325110 272760 325116
rect 272812 321162 272840 338014
rect 272950 337770 272978 338028
rect 272904 337742 272978 337770
rect 273088 338014 273148 338042
rect 272904 333674 272932 337742
rect 273088 335510 273116 338014
rect 273226 337770 273254 338028
rect 273180 337742 273254 337770
rect 273364 338014 273424 338042
rect 273076 335504 273128 335510
rect 273076 335446 273128 335452
rect 272984 335436 273036 335442
rect 272984 335378 273036 335384
rect 272892 333668 272944 333674
rect 272892 333610 272944 333616
rect 272892 330540 272944 330546
rect 272892 330482 272944 330488
rect 272800 321156 272852 321162
rect 272800 321098 272852 321104
rect 272904 319666 272932 330482
rect 272892 319660 272944 319666
rect 272892 319602 272944 319608
rect 272616 8628 272668 8634
rect 272616 8570 272668 8576
rect 272996 8498 273024 335378
rect 273076 333396 273128 333402
rect 273076 333338 273128 333344
rect 273088 8566 273116 333338
rect 273180 330546 273208 337742
rect 273364 332246 273392 338014
rect 273594 337770 273622 338028
rect 273686 337872 273714 338028
rect 273824 338014 273884 338042
rect 273686 337844 273760 337872
rect 273594 337742 273668 337770
rect 273536 335640 273588 335646
rect 273536 335582 273588 335588
rect 273548 333538 273576 335582
rect 273536 333532 273588 333538
rect 273536 333474 273588 333480
rect 273352 332240 273404 332246
rect 273352 332182 273404 332188
rect 273168 330540 273220 330546
rect 273168 330482 273220 330488
rect 273640 325694 273668 337742
rect 273732 333334 273760 337844
rect 273824 335646 273852 338014
rect 273962 337770 273990 338028
rect 274146 337770 274174 338028
rect 274238 337872 274266 338028
rect 274376 338014 274436 338042
rect 274238 337844 274312 337872
rect 273962 337742 274036 337770
rect 274146 337742 274220 337770
rect 273904 335912 273956 335918
rect 273904 335854 273956 335860
rect 273812 335640 273864 335646
rect 273812 335582 273864 335588
rect 273812 335504 273864 335510
rect 273812 335446 273864 335452
rect 273720 333328 273772 333334
rect 273720 333270 273772 333276
rect 273824 331214 273852 335446
rect 273732 331186 273852 331214
rect 273732 330562 273760 331186
rect 273732 330534 273852 330562
rect 273640 325666 273760 325694
rect 273732 8702 273760 325666
rect 273824 8838 273852 330534
rect 273812 8832 273864 8838
rect 273812 8774 273864 8780
rect 273720 8696 273772 8702
rect 273720 8638 273772 8644
rect 273076 8560 273128 8566
rect 273076 8502 273128 8508
rect 272984 8492 273036 8498
rect 272984 8434 273036 8440
rect 273916 5574 273944 335854
rect 274008 333266 274036 337742
rect 274088 333328 274140 333334
rect 274088 333270 274140 333276
rect 273996 333260 274048 333266
rect 273996 333202 274048 333208
rect 274100 323882 274128 333270
rect 274192 330562 274220 337742
rect 274284 330886 274312 337844
rect 274376 335510 274404 338014
rect 274514 337770 274542 338028
rect 274468 337742 274542 337770
rect 274652 338014 274712 338042
rect 274364 335504 274416 335510
rect 274364 335446 274416 335452
rect 274364 333260 274416 333266
rect 274364 333202 274416 333208
rect 274272 330880 274324 330886
rect 274272 330822 274324 330828
rect 274192 330534 274312 330562
rect 274180 330404 274232 330410
rect 274180 330346 274232 330352
rect 274088 323876 274140 323882
rect 274088 323818 274140 323824
rect 274192 318306 274220 330346
rect 274180 318300 274232 318306
rect 274180 318242 274232 318248
rect 274284 312662 274312 330534
rect 274272 312656 274324 312662
rect 274272 312598 274324 312604
rect 274376 8770 274404 333202
rect 274468 330410 274496 337742
rect 274652 336666 274680 338014
rect 274790 337770 274818 338028
rect 274928 338014 274988 338042
rect 274790 337742 274864 337770
rect 274640 336660 274692 336666
rect 274640 336602 274692 336608
rect 274836 330818 274864 337742
rect 274928 335442 274956 338014
rect 275066 337770 275094 338028
rect 275250 337770 275278 338028
rect 275434 337770 275462 338028
rect 275526 337890 275554 338028
rect 275664 338014 275724 338042
rect 275514 337884 275566 337890
rect 275514 337826 275566 337832
rect 275066 337742 275140 337770
rect 275250 337742 275324 337770
rect 275434 337742 275600 337770
rect 274916 335436 274968 335442
rect 274916 335378 274968 335384
rect 275112 334966 275140 337742
rect 275100 334960 275152 334966
rect 275100 334902 275152 334908
rect 275296 334898 275324 337742
rect 275468 335368 275520 335374
rect 275468 335310 275520 335316
rect 275284 334892 275336 334898
rect 275284 334834 275336 334840
rect 274824 330812 274876 330818
rect 274824 330754 274876 330760
rect 274456 330404 274508 330410
rect 274456 330346 274508 330352
rect 274364 8764 274416 8770
rect 274364 8706 274416 8712
rect 275480 5710 275508 335310
rect 275572 321094 275600 337742
rect 275664 329390 275692 338014
rect 275802 337770 275830 338028
rect 275940 338014 276000 338042
rect 275802 337742 275876 337770
rect 275744 335436 275796 335442
rect 275744 335378 275796 335384
rect 275652 329384 275704 329390
rect 275652 329326 275704 329332
rect 275560 321088 275612 321094
rect 275560 321030 275612 321036
rect 275756 316878 275784 335378
rect 275744 316872 275796 316878
rect 275744 316814 275796 316820
rect 275848 309874 275876 337742
rect 275940 335374 275968 338014
rect 276078 337890 276106 338028
rect 276216 338014 276276 338042
rect 276066 337884 276118 337890
rect 276066 337826 276118 337832
rect 276216 335374 276244 338014
rect 276354 337770 276382 338028
rect 276492 338014 276552 338042
rect 276354 337742 276428 337770
rect 275928 335368 275980 335374
rect 275928 335310 275980 335316
rect 276204 335368 276256 335374
rect 276204 335310 276256 335316
rect 275836 309868 275888 309874
rect 275836 309810 275888 309816
rect 276400 5778 276428 337742
rect 276492 335442 276520 338014
rect 276630 337770 276658 338028
rect 276584 337742 276658 337770
rect 276768 338014 276828 338042
rect 276480 335436 276532 335442
rect 276480 335378 276532 335384
rect 276480 334620 276532 334626
rect 276480 334562 276532 334568
rect 276492 5846 276520 334562
rect 276584 332178 276612 337742
rect 276664 335844 276716 335850
rect 276664 335786 276716 335792
rect 276572 332172 276624 332178
rect 276572 332114 276624 332120
rect 276572 331968 276624 331974
rect 276572 331910 276624 331916
rect 276584 5914 276612 331910
rect 276676 7614 276704 335786
rect 276768 334626 276796 338014
rect 276906 337770 276934 338028
rect 276860 337742 276934 337770
rect 277044 338014 277104 338042
rect 277228 338014 277288 338042
rect 276756 334620 276808 334626
rect 276756 334562 276808 334568
rect 276860 325106 276888 337742
rect 276940 335368 276992 335374
rect 276940 335310 276992 335316
rect 276848 325100 276900 325106
rect 276848 325042 276900 325048
rect 276952 314090 276980 335310
rect 276940 314084 276992 314090
rect 276940 314026 276992 314032
rect 277044 293282 277072 338014
rect 277228 337906 277256 338014
rect 277136 337878 277256 337906
rect 277136 331974 277164 337878
rect 277366 337770 277394 338028
rect 277228 337742 277394 337770
rect 277504 338014 277564 338042
rect 277124 331968 277176 331974
rect 277124 331910 277176 331916
rect 277228 327962 277256 337742
rect 277504 335442 277532 338014
rect 277642 337770 277670 338028
rect 277780 338014 277840 338042
rect 277642 337742 277716 337770
rect 277308 335436 277360 335442
rect 277308 335378 277360 335384
rect 277492 335436 277544 335442
rect 277492 335378 277544 335384
rect 277216 327956 277268 327962
rect 277216 327898 277268 327904
rect 277320 326670 277348 335378
rect 277688 333266 277716 337742
rect 277676 333260 277728 333266
rect 277676 333202 277728 333208
rect 277780 330750 277808 338014
rect 277918 337940 277946 338028
rect 278056 338014 278116 338042
rect 277918 337912 277992 337940
rect 277860 337204 277912 337210
rect 277860 337146 277912 337152
rect 277768 330744 277820 330750
rect 277768 330686 277820 330692
rect 277308 326664 277360 326670
rect 277308 326606 277360 326612
rect 277032 293276 277084 293282
rect 277032 293218 277084 293224
rect 276664 7608 276716 7614
rect 276664 7550 276716 7556
rect 277872 6118 277900 337146
rect 277964 333334 277992 337912
rect 277952 333328 278004 333334
rect 277952 333270 278004 333276
rect 278056 316034 278084 338014
rect 278194 337770 278222 338028
rect 278148 337742 278222 337770
rect 278332 338014 278392 338042
rect 278148 323814 278176 337742
rect 278228 335436 278280 335442
rect 278228 335378 278280 335384
rect 278136 323808 278188 323814
rect 278136 323750 278188 323756
rect 277964 316006 278084 316034
rect 277860 6112 277912 6118
rect 277860 6054 277912 6060
rect 277964 6050 277992 316006
rect 278240 312594 278268 335378
rect 278228 312588 278280 312594
rect 278228 312530 278280 312536
rect 278332 291854 278360 338014
rect 278470 337770 278498 338028
rect 278424 337742 278498 337770
rect 278608 338014 278668 338042
rect 278792 338014 278852 338042
rect 278424 337210 278452 337742
rect 278412 337204 278464 337210
rect 278412 337146 278464 337152
rect 278504 333260 278556 333266
rect 278504 333202 278556 333208
rect 278412 330404 278464 330410
rect 278412 330346 278464 330352
rect 278320 291848 278372 291854
rect 278320 291790 278372 291796
rect 278424 9790 278452 330346
rect 278412 9784 278464 9790
rect 278412 9726 278464 9732
rect 277952 6044 278004 6050
rect 277952 5986 278004 5992
rect 278516 5982 278544 333202
rect 278608 330410 278636 338014
rect 278792 335782 278820 338014
rect 278930 337822 278958 338028
rect 279068 338014 279128 338042
rect 278918 337816 278970 337822
rect 278918 337758 278970 337764
rect 278780 335776 278832 335782
rect 278780 335718 278832 335724
rect 278688 333328 278740 333334
rect 278688 333270 278740 333276
rect 278596 330404 278648 330410
rect 278596 330346 278648 330352
rect 278700 325038 278728 333270
rect 279068 330410 279096 338014
rect 279206 337770 279234 338028
rect 279160 337742 279234 337770
rect 279390 337770 279418 338028
rect 279482 337872 279510 338028
rect 279620 338014 279680 338042
rect 279482 337844 279556 337872
rect 279390 337742 279464 337770
rect 279160 334830 279188 337742
rect 279148 334824 279200 334830
rect 279148 334766 279200 334772
rect 279240 333328 279292 333334
rect 279240 333270 279292 333276
rect 279056 330404 279108 330410
rect 279056 330346 279108 330352
rect 279252 326602 279280 333270
rect 279332 333260 279384 333266
rect 279332 333202 279384 333208
rect 279240 326596 279292 326602
rect 279240 326538 279292 326544
rect 279344 325694 279372 333202
rect 279436 330528 279464 337742
rect 279528 333282 279556 337844
rect 279620 333470 279648 338014
rect 279758 337736 279786 338028
rect 279896 338014 279956 338042
rect 279758 337708 279832 337736
rect 279608 333464 279660 333470
rect 279608 333406 279660 333412
rect 279528 333254 279648 333282
rect 279804 333266 279832 337708
rect 279436 330500 279556 330528
rect 279344 325666 279464 325694
rect 278688 325032 278740 325038
rect 278688 324974 278740 324980
rect 279436 6730 279464 325666
rect 279528 6798 279556 330500
rect 279620 9926 279648 333254
rect 279792 333260 279844 333266
rect 279792 333202 279844 333208
rect 279896 330528 279924 338014
rect 280034 337906 280062 338028
rect 280034 337878 280108 337906
rect 279976 337816 280028 337822
rect 279976 337758 280028 337764
rect 279712 330500 279924 330528
rect 279712 9994 279740 330500
rect 279792 330404 279844 330410
rect 279792 330346 279844 330352
rect 279700 9988 279752 9994
rect 279700 9930 279752 9936
rect 279608 9920 279660 9926
rect 279608 9862 279660 9868
rect 279804 9858 279832 330346
rect 279988 316034 280016 337758
rect 280080 333334 280108 337878
rect 280218 337770 280246 338028
rect 280310 337890 280338 338028
rect 280448 338014 280508 338042
rect 280632 338014 280692 338042
rect 280298 337884 280350 337890
rect 280298 337826 280350 337832
rect 280218 337742 280292 337770
rect 280068 333328 280120 333334
rect 280068 333270 280120 333276
rect 280264 330342 280292 337742
rect 280252 330336 280304 330342
rect 280252 330278 280304 330284
rect 280448 330206 280476 338014
rect 280632 335646 280660 338014
rect 280770 337906 280798 338028
rect 280908 338014 280968 338042
rect 280770 337878 280844 337906
rect 280620 335640 280672 335646
rect 280620 335582 280672 335588
rect 280712 335368 280764 335374
rect 280712 335310 280764 335316
rect 280620 333260 280672 333266
rect 280620 333202 280672 333208
rect 280436 330200 280488 330206
rect 280436 330142 280488 330148
rect 279896 316006 280016 316034
rect 279792 9852 279844 9858
rect 279792 9794 279844 9800
rect 279896 6866 279924 316006
rect 279884 6860 279936 6866
rect 279884 6802 279936 6808
rect 279516 6792 279568 6798
rect 279516 6734 279568 6740
rect 279424 6724 279476 6730
rect 279424 6666 279476 6672
rect 280632 6526 280660 333202
rect 280724 319598 280752 335310
rect 280816 335186 280844 337878
rect 280908 335374 280936 338014
rect 281046 337872 281074 338028
rect 281184 338014 281244 338042
rect 281046 337844 281120 337872
rect 280988 337748 281040 337754
rect 280988 337690 281040 337696
rect 280896 335368 280948 335374
rect 280896 335310 280948 335316
rect 280816 335158 280936 335186
rect 280804 330404 280856 330410
rect 280804 330346 280856 330352
rect 280712 319592 280764 319598
rect 280712 319534 280764 319540
rect 280816 315450 280844 330346
rect 280804 315444 280856 315450
rect 280804 315386 280856 315392
rect 280908 10130 280936 335158
rect 280896 10124 280948 10130
rect 280896 10066 280948 10072
rect 281000 10062 281028 337690
rect 281092 333266 281120 337844
rect 281080 333260 281132 333266
rect 281080 333202 281132 333208
rect 281184 330528 281212 338014
rect 281322 337822 281350 338028
rect 281460 338014 281520 338042
rect 281310 337816 281362 337822
rect 281310 337758 281362 337764
rect 281264 335640 281316 335646
rect 281264 335582 281316 335588
rect 281092 330500 281212 330528
rect 281092 10198 281120 330500
rect 281172 330336 281224 330342
rect 281172 330278 281224 330284
rect 281080 10192 281132 10198
rect 281080 10134 281132 10140
rect 280988 10056 281040 10062
rect 280988 9998 281040 10004
rect 280712 7608 280764 7614
rect 280712 7550 280764 7556
rect 280620 6520 280672 6526
rect 280620 6462 280672 6468
rect 278504 5976 278556 5982
rect 278504 5918 278556 5924
rect 276572 5908 276624 5914
rect 276572 5850 276624 5856
rect 276480 5840 276532 5846
rect 276480 5782 276532 5788
rect 276388 5772 276440 5778
rect 276388 5714 276440 5720
rect 275468 5704 275520 5710
rect 275468 5646 275520 5652
rect 274824 5636 274876 5642
rect 274824 5578 274876 5584
rect 273904 5568 273956 5574
rect 273904 5510 273956 5516
rect 271696 4820 271748 4826
rect 271696 4762 271748 4768
rect 273628 3732 273680 3738
rect 273628 3674 273680 3680
rect 272432 3528 272484 3534
rect 270040 3460 270092 3466
rect 271156 3454 271276 3482
rect 272432 3470 272484 3476
rect 270040 3402 270092 3408
rect 269028 3324 269080 3330
rect 269028 3266 269080 3272
rect 268936 3188 268988 3194
rect 268936 3130 268988 3136
rect 270052 480 270080 3402
rect 271248 480 271276 3454
rect 272444 480 272472 3470
rect 273640 480 273668 3674
rect 274836 480 274864 5578
rect 279516 5568 279568 5574
rect 279516 5510 279568 5516
rect 278320 4548 278372 4554
rect 278320 4490 278372 4496
rect 277124 3324 277176 3330
rect 277124 3266 277176 3272
rect 276020 3188 276072 3194
rect 276020 3130 276072 3136
rect 276032 480 276060 3130
rect 277136 480 277164 3266
rect 278332 480 278360 4490
rect 279528 480 279556 5510
rect 280724 480 280752 7550
rect 281184 6662 281212 330278
rect 281172 6656 281224 6662
rect 281172 6598 281224 6604
rect 281276 6594 281304 335582
rect 281460 330528 281488 338014
rect 281598 337822 281626 338028
rect 281736 338014 281796 338042
rect 281586 337816 281638 337822
rect 281586 337758 281638 337764
rect 281736 335646 281764 338014
rect 281874 337906 281902 338028
rect 281874 337878 281948 337906
rect 281724 335640 281776 335646
rect 281724 335582 281776 335588
rect 281368 330500 281488 330528
rect 281264 6588 281316 6594
rect 281264 6530 281316 6536
rect 281368 6458 281396 330500
rect 281920 330410 281948 337878
rect 282058 337770 282086 338028
rect 282150 337906 282178 338028
rect 282288 338014 282348 338042
rect 282472 338014 282532 338042
rect 282150 337878 282224 337906
rect 282058 337742 282132 337770
rect 282000 335368 282052 335374
rect 282000 335310 282052 335316
rect 281908 330404 281960 330410
rect 281908 330346 281960 330352
rect 281448 330200 281500 330206
rect 281448 330142 281500 330148
rect 281460 322454 281488 330142
rect 282012 325694 282040 335310
rect 282104 330546 282132 337742
rect 282196 333402 282224 337878
rect 282288 335374 282316 338014
rect 282368 335844 282420 335850
rect 282368 335786 282420 335792
rect 282276 335368 282328 335374
rect 282276 335310 282328 335316
rect 282184 333396 282236 333402
rect 282184 333338 282236 333344
rect 282184 333260 282236 333266
rect 282184 333202 282236 333208
rect 282092 330540 282144 330546
rect 282092 330482 282144 330488
rect 282012 325666 282132 325694
rect 281448 322448 281500 322454
rect 281448 322390 281500 322396
rect 281356 6452 281408 6458
rect 281356 6394 281408 6400
rect 282104 6322 282132 325666
rect 282196 321026 282224 333202
rect 282276 330540 282328 330546
rect 282276 330482 282328 330488
rect 282184 321020 282236 321026
rect 282184 320962 282236 320968
rect 282288 11014 282316 330482
rect 282276 11008 282328 11014
rect 282276 10950 282328 10956
rect 282380 10878 282408 335786
rect 282472 10946 282500 338014
rect 282610 337906 282638 338028
rect 282748 338014 282808 338042
rect 282610 337878 282684 337906
rect 282552 337816 282604 337822
rect 282552 337758 282604 337764
rect 282460 10940 282512 10946
rect 282460 10882 282512 10888
rect 282368 10872 282420 10878
rect 282368 10814 282420 10820
rect 282564 10266 282592 337758
rect 282656 333266 282684 337878
rect 282644 333260 282696 333266
rect 282644 333202 282696 333208
rect 282748 330528 282776 338014
rect 282886 337770 282914 338028
rect 282840 337742 282914 337770
rect 283024 338014 283084 338042
rect 282840 335850 282868 337742
rect 282828 335844 282880 335850
rect 282828 335786 282880 335792
rect 283024 335782 283052 338014
rect 283162 337736 283190 338028
rect 283300 338014 283360 338042
rect 283162 337708 283236 337736
rect 283012 335776 283064 335782
rect 283012 335718 283064 335724
rect 282828 333396 282880 333402
rect 282828 333338 282880 333344
rect 282656 330500 282776 330528
rect 282552 10260 282604 10266
rect 282552 10202 282604 10208
rect 282092 6316 282144 6322
rect 282092 6258 282144 6264
rect 282656 6254 282684 330500
rect 282736 330404 282788 330410
rect 282736 330346 282788 330352
rect 282748 6390 282776 330346
rect 282840 323746 282868 333338
rect 283208 328454 283236 337708
rect 283300 335442 283328 338014
rect 283438 337736 283466 338028
rect 283576 338014 283636 338042
rect 283438 337708 283512 337736
rect 283380 335708 283432 335714
rect 283380 335650 283432 335656
rect 283288 335436 283340 335442
rect 283288 335378 283340 335384
rect 283392 332042 283420 335650
rect 283484 335594 283512 337708
rect 283576 335714 283604 338014
rect 283714 337736 283742 338028
rect 283852 338014 283912 338042
rect 284036 338014 284096 338042
rect 283714 337708 283788 337736
rect 283656 335776 283708 335782
rect 283656 335718 283708 335724
rect 283564 335708 283616 335714
rect 283564 335650 283616 335656
rect 283484 335566 283604 335594
rect 283380 332036 283432 332042
rect 283380 331978 283432 331984
rect 283208 328426 283512 328454
rect 282828 323740 282880 323746
rect 282828 323682 282880 323688
rect 282736 6384 282788 6390
rect 282736 6326 282788 6332
rect 282644 6248 282696 6254
rect 282644 6190 282696 6196
rect 283484 6186 283512 328426
rect 283576 326398 283604 335566
rect 283564 326392 283616 326398
rect 283564 326334 283616 326340
rect 283668 318238 283696 335718
rect 283760 333266 283788 337708
rect 283748 333260 283800 333266
rect 283748 333202 283800 333208
rect 283748 326392 283800 326398
rect 283748 326334 283800 326340
rect 283656 318232 283708 318238
rect 283656 318174 283708 318180
rect 283760 307154 283788 326334
rect 283748 307148 283800 307154
rect 283748 307090 283800 307096
rect 283852 305726 283880 338014
rect 284036 336122 284064 338014
rect 284174 337770 284202 338028
rect 284128 337742 284202 337770
rect 284358 337770 284386 338028
rect 284450 337872 284478 338028
rect 284588 338014 284648 338042
rect 284450 337844 284524 337872
rect 284358 337742 284432 337770
rect 284024 336116 284076 336122
rect 284024 336058 284076 336064
rect 283932 335504 283984 335510
rect 283932 335446 283984 335452
rect 283944 329322 283972 335446
rect 284024 333260 284076 333266
rect 284024 333202 284076 333208
rect 283932 329316 283984 329322
rect 283932 329258 283984 329264
rect 283932 326392 283984 326398
rect 283932 326334 283984 326340
rect 283840 305720 283892 305726
rect 283840 305662 283892 305668
rect 283944 10674 283972 326334
rect 284036 10742 284064 333202
rect 284128 326398 284156 337742
rect 284208 335436 284260 335442
rect 284208 335378 284260 335384
rect 284116 326392 284168 326398
rect 284116 326334 284168 326340
rect 284220 311894 284248 335378
rect 284404 334558 284432 337742
rect 284496 335850 284524 337844
rect 284484 335844 284536 335850
rect 284484 335786 284536 335792
rect 284484 335504 284536 335510
rect 284484 335446 284536 335452
rect 284392 334552 284444 334558
rect 284392 334494 284444 334500
rect 284496 331214 284524 335446
rect 284588 335374 284616 338014
rect 284726 337736 284754 338028
rect 284864 338014 284924 338042
rect 284726 337708 284800 337736
rect 284668 335640 284720 335646
rect 284668 335582 284720 335588
rect 284576 335368 284628 335374
rect 284576 335310 284628 335316
rect 284496 331186 284616 331214
rect 284588 327894 284616 331186
rect 284576 327888 284628 327894
rect 284576 327830 284628 327836
rect 284680 326262 284708 335582
rect 284772 334626 284800 337708
rect 284864 335510 284892 338014
rect 285002 337736 285030 338028
rect 285140 338014 285200 338042
rect 285002 337708 285076 337736
rect 284852 335504 284904 335510
rect 284852 335446 284904 335452
rect 284944 335368 284996 335374
rect 284944 335310 284996 335316
rect 284760 334620 284812 334626
rect 284760 334562 284812 334568
rect 284956 334506 284984 335310
rect 284772 334478 284984 334506
rect 284668 326256 284720 326262
rect 284668 326198 284720 326204
rect 284128 311866 284248 311894
rect 284128 10810 284156 311866
rect 284300 13116 284352 13122
rect 284300 13058 284352 13064
rect 284116 10804 284168 10810
rect 284116 10746 284168 10752
rect 284024 10736 284076 10742
rect 284024 10678 284076 10684
rect 283932 10668 283984 10674
rect 283932 10610 283984 10616
rect 283472 6180 283524 6186
rect 283472 6122 283524 6128
rect 283104 4684 283156 4690
rect 283104 4626 283156 4632
rect 281908 4616 281960 4622
rect 281908 4558 281960 4564
rect 281920 480 281948 4558
rect 283116 480 283144 4626
rect 284312 480 284340 13058
rect 284772 2990 284800 334478
rect 284944 334416 284996 334422
rect 284944 334358 284996 334364
rect 284852 333260 284904 333266
rect 284852 333202 284904 333208
rect 284864 3058 284892 333202
rect 284956 326380 284984 334358
rect 285048 326534 285076 337708
rect 285140 335374 285168 338014
rect 285278 337736 285306 338028
rect 285416 338014 285476 338042
rect 285278 337708 285352 337736
rect 285128 335368 285180 335374
rect 285128 335310 285180 335316
rect 285220 335368 285272 335374
rect 285220 335310 285272 335316
rect 285128 335232 285180 335238
rect 285128 335174 285180 335180
rect 285036 326528 285088 326534
rect 285036 326470 285088 326476
rect 284956 326352 285076 326380
rect 284944 326256 284996 326262
rect 284944 326198 284996 326204
rect 284956 308514 284984 326198
rect 284944 308508 284996 308514
rect 284944 308450 284996 308456
rect 285048 10470 285076 326352
rect 285140 10606 285168 335174
rect 285232 334422 285260 335310
rect 285220 334416 285272 334422
rect 285220 334358 285272 334364
rect 285324 329254 285352 337708
rect 285416 335374 285444 338014
rect 285554 337736 285582 338028
rect 285738 337906 285766 338028
rect 285876 338014 285936 338042
rect 285738 337878 285812 337906
rect 285680 337816 285732 337822
rect 285680 337758 285732 337764
rect 285554 337708 285628 337736
rect 285404 335368 285456 335374
rect 285404 335310 285456 335316
rect 285404 334620 285456 334626
rect 285404 334562 285456 334568
rect 285312 329248 285364 329254
rect 285312 329190 285364 329196
rect 285220 326528 285272 326534
rect 285220 326470 285272 326476
rect 285128 10600 285180 10606
rect 285128 10542 285180 10548
rect 285232 10538 285260 326470
rect 285416 318794 285444 334562
rect 285496 334552 285548 334558
rect 285496 334494 285548 334500
rect 285324 318766 285444 318794
rect 285324 314106 285352 318766
rect 285324 314078 285444 314106
rect 285312 313948 285364 313954
rect 285312 313890 285364 313896
rect 285220 10532 285272 10538
rect 285220 10474 285272 10480
rect 285036 10464 285088 10470
rect 285036 10406 285088 10412
rect 284852 3052 284904 3058
rect 284852 2994 284904 3000
rect 284760 2984 284812 2990
rect 284760 2926 284812 2932
rect 285324 2854 285352 313890
rect 285416 16574 285444 314078
rect 285508 313954 285536 334494
rect 285600 333266 285628 337708
rect 285588 333260 285640 333266
rect 285588 333202 285640 333208
rect 285692 323678 285720 337758
rect 285784 330682 285812 337878
rect 285772 330676 285824 330682
rect 285772 330618 285824 330624
rect 285876 326058 285904 338014
rect 286014 337736 286042 338028
rect 286152 338014 286212 338042
rect 286014 337708 286088 337736
rect 286060 335220 286088 337708
rect 286152 335374 286180 338014
rect 286290 337736 286318 338028
rect 286428 338014 286488 338042
rect 286290 337708 286364 337736
rect 286140 335368 286192 335374
rect 286140 335310 286192 335316
rect 286060 335192 286272 335220
rect 285956 334416 286008 334422
rect 285956 334358 286008 334364
rect 285968 326126 285996 334358
rect 286140 333260 286192 333266
rect 286140 333202 286192 333208
rect 285956 326120 286008 326126
rect 285956 326062 286008 326068
rect 285864 326052 285916 326058
rect 285864 325994 285916 326000
rect 285680 323672 285732 323678
rect 285680 323614 285732 323620
rect 285496 313948 285548 313954
rect 285496 313890 285548 313896
rect 285416 16546 285536 16574
rect 285404 4752 285456 4758
rect 285404 4694 285456 4700
rect 285312 2848 285364 2854
rect 285312 2790 285364 2796
rect 285416 480 285444 4694
rect 285508 2922 285536 16546
rect 286152 3262 286180 333202
rect 286140 3256 286192 3262
rect 286140 3198 286192 3204
rect 286244 3126 286272 335192
rect 286336 326398 286364 337708
rect 286428 335374 286456 338014
rect 286566 337822 286594 338028
rect 286704 338014 286764 338042
rect 286554 337816 286606 337822
rect 286554 337758 286606 337764
rect 286508 335436 286560 335442
rect 286508 335378 286560 335384
rect 286416 335368 286468 335374
rect 286416 335310 286468 335316
rect 286416 335232 286468 335238
rect 286416 335174 286468 335180
rect 286428 333402 286456 335174
rect 286416 333396 286468 333402
rect 286416 333338 286468 333344
rect 286520 331214 286548 335378
rect 286704 331214 286732 338014
rect 286842 337736 286870 338028
rect 286980 338014 287040 338042
rect 286842 337708 286916 337736
rect 286784 335368 286836 335374
rect 286784 335310 286836 335316
rect 286428 331186 286548 331214
rect 286612 331186 286732 331214
rect 286324 326392 286376 326398
rect 286324 326334 286376 326340
rect 286324 326120 286376 326126
rect 286324 326062 286376 326068
rect 286336 6934 286364 326062
rect 286428 322386 286456 331186
rect 286612 326380 286640 331186
rect 286520 326352 286640 326380
rect 286692 326392 286744 326398
rect 286416 322380 286468 322386
rect 286416 322322 286468 322328
rect 286520 311234 286548 326352
rect 286692 326334 286744 326340
rect 286600 326052 286652 326058
rect 286600 325994 286652 326000
rect 286508 311228 286560 311234
rect 286508 311170 286560 311176
rect 286612 10402 286640 325994
rect 286600 10396 286652 10402
rect 286600 10338 286652 10344
rect 286704 10334 286732 326334
rect 286692 10328 286744 10334
rect 286692 10270 286744 10276
rect 286324 6928 286376 6934
rect 286324 6870 286376 6876
rect 286600 5500 286652 5506
rect 286600 5442 286652 5448
rect 286232 3120 286284 3126
rect 286232 3062 286284 3068
rect 285496 2916 285548 2922
rect 285496 2858 285548 2864
rect 286612 480 286640 5442
rect 286796 3194 286824 335310
rect 286888 333266 286916 337708
rect 286980 335442 287008 338014
rect 287118 337736 287146 338028
rect 287256 338014 287316 338042
rect 287118 337708 287192 337736
rect 287060 336048 287112 336054
rect 287060 335990 287112 335996
rect 286968 335436 287020 335442
rect 286968 335378 287020 335384
rect 286876 333260 286928 333266
rect 286876 333202 286928 333208
rect 287072 326398 287100 335990
rect 287164 333334 287192 337708
rect 287256 335374 287284 338014
rect 287394 337906 287422 338028
rect 287394 337878 287468 337906
rect 287336 337816 287388 337822
rect 287336 337758 287388 337764
rect 287244 335368 287296 335374
rect 287244 335310 287296 335316
rect 287152 333328 287204 333334
rect 287152 333270 287204 333276
rect 287348 328454 287376 337758
rect 287440 333266 287468 337878
rect 287578 337736 287606 338028
rect 287716 338014 287776 338042
rect 287578 337708 287652 337736
rect 287520 335368 287572 335374
rect 287520 335310 287572 335316
rect 287428 333260 287480 333266
rect 287428 333202 287480 333208
rect 287348 328426 287468 328454
rect 287060 326392 287112 326398
rect 287060 326334 287112 326340
rect 287440 4146 287468 328426
rect 287428 4140 287480 4146
rect 287428 4082 287480 4088
rect 287532 3398 287560 335310
rect 287624 319530 287652 337708
rect 287716 335374 287744 338014
rect 287854 337736 287882 338028
rect 287992 338014 288052 338042
rect 287854 337708 287928 337736
rect 287796 335504 287848 335510
rect 287796 335446 287848 335452
rect 287704 335368 287756 335374
rect 287704 335310 287756 335316
rect 287704 326392 287756 326398
rect 287704 326334 287756 326340
rect 287612 319524 287664 319530
rect 287612 319466 287664 319472
rect 287716 11966 287744 326334
rect 287808 309806 287836 335446
rect 287796 309800 287848 309806
rect 287796 309742 287848 309748
rect 287704 11960 287756 11966
rect 287704 11902 287756 11908
rect 287900 8294 287928 337708
rect 287992 335374 288020 338014
rect 288130 337822 288158 338028
rect 288268 338014 288328 338042
rect 288118 337816 288170 337822
rect 288118 337758 288170 337764
rect 287980 335368 288032 335374
rect 287980 335310 288032 335316
rect 288164 335300 288216 335306
rect 288164 335242 288216 335248
rect 288072 333260 288124 333266
rect 288072 333202 288124 333208
rect 288084 321554 288112 333202
rect 287992 321526 288112 321554
rect 287888 8288 287940 8294
rect 287888 8230 287940 8236
rect 287992 7546 288020 321526
rect 288176 316810 288204 335242
rect 288164 316804 288216 316810
rect 288164 316746 288216 316752
rect 288268 316690 288296 338014
rect 288406 337770 288434 338028
rect 288360 337742 288434 337770
rect 288590 337770 288618 338028
rect 288682 337906 288710 338028
rect 288682 337878 288756 337906
rect 288590 337742 288664 337770
rect 288360 335510 288388 337742
rect 288440 336524 288492 336530
rect 288440 336466 288492 336472
rect 288348 335504 288400 335510
rect 288348 335446 288400 335452
rect 288348 335368 288400 335374
rect 288348 335310 288400 335316
rect 288360 326466 288388 335310
rect 288452 333606 288480 336466
rect 288440 333600 288492 333606
rect 288440 333542 288492 333548
rect 288636 329458 288664 337742
rect 288624 329452 288676 329458
rect 288624 329394 288676 329400
rect 288348 326460 288400 326466
rect 288348 326402 288400 326408
rect 288728 324970 288756 337878
rect 288866 337770 288894 338028
rect 288958 337906 288986 338028
rect 288958 337878 289032 337906
rect 288866 337742 288940 337770
rect 288716 324964 288768 324970
rect 288716 324906 288768 324912
rect 288912 318170 288940 337742
rect 289004 333266 289032 337878
rect 289142 337770 289170 338028
rect 289280 338014 289340 338042
rect 289142 337742 289216 337770
rect 289084 335368 289136 335374
rect 289084 335310 289136 335316
rect 288992 333260 289044 333266
rect 288992 333202 289044 333208
rect 288900 318164 288952 318170
rect 288900 318106 288952 318112
rect 289096 316810 289124 335310
rect 289188 325394 289216 337742
rect 289280 335374 289308 338014
rect 289418 337906 289446 338028
rect 289556 338014 289616 338042
rect 289418 337878 289492 337906
rect 289360 337816 289412 337822
rect 289360 337758 289412 337764
rect 289268 335368 289320 335374
rect 289268 335310 289320 335316
rect 289188 325366 289308 325394
rect 289176 325236 289228 325242
rect 289176 325178 289228 325184
rect 289084 316804 289136 316810
rect 289084 316746 289136 316752
rect 288084 316662 288296 316690
rect 288084 8226 288112 316662
rect 288164 316600 288216 316606
rect 288164 316542 288216 316548
rect 288072 8220 288124 8226
rect 288072 8162 288124 8168
rect 287980 7540 288032 7546
rect 287980 7482 288032 7488
rect 287796 6928 287848 6934
rect 287796 6870 287848 6876
rect 287520 3392 287572 3398
rect 287520 3334 287572 3340
rect 286784 3188 286836 3194
rect 286784 3130 286836 3136
rect 287808 480 287836 6870
rect 288176 3330 288204 316542
rect 289188 308446 289216 325178
rect 289176 308440 289228 308446
rect 289176 308382 289228 308388
rect 289280 8090 289308 325366
rect 289372 325242 289400 337758
rect 289464 333198 289492 337878
rect 289452 333192 289504 333198
rect 289452 333134 289504 333140
rect 289556 331214 289584 338014
rect 289694 337822 289722 338028
rect 289832 338014 289892 338042
rect 289682 337816 289734 337822
rect 289682 337758 289734 337764
rect 289832 335442 289860 338014
rect 289970 337770 289998 338028
rect 290108 338014 290168 338042
rect 289970 337742 290044 337770
rect 289820 335436 289872 335442
rect 289820 335378 289872 335384
rect 290016 335238 290044 337742
rect 290108 335714 290136 338014
rect 290246 337906 290274 338028
rect 290384 338014 290444 338042
rect 290246 337878 290320 337906
rect 290096 335708 290148 335714
rect 290096 335650 290148 335656
rect 290004 335232 290056 335238
rect 290004 335174 290056 335180
rect 290292 334354 290320 337878
rect 290384 336326 290412 338014
rect 290522 337770 290550 338028
rect 290660 338014 290720 338042
rect 290522 337742 290596 337770
rect 290372 336320 290424 336326
rect 290372 336262 290424 336268
rect 290280 334348 290332 334354
rect 290280 334290 290332 334296
rect 289636 333260 289688 333266
rect 289636 333202 289688 333208
rect 289464 331186 289584 331214
rect 289360 325236 289412 325242
rect 289360 325178 289412 325184
rect 289360 324964 289412 324970
rect 289360 324906 289412 324912
rect 289372 8158 289400 324906
rect 289360 8152 289412 8158
rect 289360 8094 289412 8100
rect 289268 8084 289320 8090
rect 289268 8026 289320 8032
rect 289464 8022 289492 331186
rect 289544 329452 289596 329458
rect 289544 329394 289596 329400
rect 289452 8016 289504 8022
rect 289452 7958 289504 7964
rect 288992 5432 289044 5438
rect 288992 5374 289044 5380
rect 288164 3324 288216 3330
rect 288164 3266 288216 3272
rect 289004 480 289032 5374
rect 289556 4078 289584 329394
rect 289544 4072 289596 4078
rect 289544 4014 289596 4020
rect 289648 4010 289676 333202
rect 289728 333192 289780 333198
rect 289728 333134 289780 333140
rect 289636 4004 289688 4010
rect 289636 3946 289688 3952
rect 289740 3942 289768 333134
rect 290568 322318 290596 337742
rect 290660 335374 290688 338014
rect 290798 337822 290826 338028
rect 290936 338014 290996 338042
rect 291120 338014 291180 338042
rect 290786 337816 290838 337822
rect 290786 337758 290838 337764
rect 290936 335594 290964 338014
rect 290752 335566 290964 335594
rect 290648 335368 290700 335374
rect 290648 335310 290700 335316
rect 290556 322312 290608 322318
rect 290556 322254 290608 322260
rect 290752 315382 290780 335566
rect 290832 335436 290884 335442
rect 290832 335378 290884 335384
rect 290740 315376 290792 315382
rect 290740 315318 290792 315324
rect 290188 5364 290240 5370
rect 290188 5306 290240 5312
rect 289728 3936 289780 3942
rect 289728 3878 289780 3884
rect 290200 480 290228 5306
rect 290844 3874 290872 335378
rect 291016 335368 291068 335374
rect 291016 335310 291068 335316
rect 291028 334506 291056 335310
rect 290936 334478 291056 334506
rect 290832 3868 290884 3874
rect 290832 3810 290884 3816
rect 290936 3738 290964 334478
rect 291016 334348 291068 334354
rect 291016 334290 291068 334296
rect 291028 326398 291056 334290
rect 291120 326482 291148 338014
rect 291258 337906 291286 338028
rect 291396 338014 291456 338042
rect 291258 337878 291332 337906
rect 291304 333266 291332 337878
rect 291396 335374 291424 338014
rect 291534 337906 291562 338028
rect 291672 338014 291732 338042
rect 291534 337878 291608 337906
rect 291384 335368 291436 335374
rect 291384 335310 291436 335316
rect 291580 334422 291608 337878
rect 291672 335442 291700 338014
rect 291810 337770 291838 338028
rect 291764 337742 291838 337770
rect 291948 338014 292008 338042
rect 291660 335436 291712 335442
rect 291660 335378 291712 335384
rect 291568 334416 291620 334422
rect 291568 334358 291620 334364
rect 291292 333260 291344 333266
rect 291292 333202 291344 333208
rect 291120 326454 291240 326482
rect 291016 326392 291068 326398
rect 291016 326334 291068 326340
rect 291212 326210 291240 326454
rect 291028 326182 291240 326210
rect 290924 3732 290976 3738
rect 290924 3674 290976 3680
rect 291028 3670 291056 326182
rect 291108 326120 291160 326126
rect 291108 326062 291160 326068
rect 291120 3806 291148 326062
rect 291764 321554 291792 337742
rect 291948 335510 291976 338014
rect 292086 337770 292114 338028
rect 292224 338014 292284 338042
rect 292086 337742 292160 337770
rect 291936 335504 291988 335510
rect 291936 335446 291988 335452
rect 292028 335436 292080 335442
rect 292028 335378 292080 335384
rect 291844 335368 291896 335374
rect 291844 335310 291896 335316
rect 291936 335368 291988 335374
rect 291936 335310 291988 335316
rect 291580 321526 291792 321554
rect 291580 11966 291608 321526
rect 291856 311894 291884 335310
rect 291764 311866 291884 311894
rect 291764 12442 291792 311866
rect 291752 12436 291804 12442
rect 291752 12378 291804 12384
rect 291948 12034 291976 335310
rect 291936 12028 291988 12034
rect 291936 11970 291988 11976
rect 291384 11960 291436 11966
rect 291384 11902 291436 11908
rect 291568 11960 291620 11966
rect 291568 11902 291620 11908
rect 291108 3800 291160 3806
rect 291108 3742 291160 3748
rect 291016 3664 291068 3670
rect 291016 3606 291068 3612
rect 291396 480 291424 11902
rect 292040 7886 292068 335378
rect 292132 326534 292160 337742
rect 292224 335374 292252 338014
rect 292362 337770 292390 338028
rect 292500 338014 292560 338042
rect 292362 337742 292436 337770
rect 292304 335504 292356 335510
rect 292304 335446 292356 335452
rect 292212 335368 292264 335374
rect 292212 335310 292264 335316
rect 292212 333260 292264 333266
rect 292212 333202 292264 333208
rect 292120 326528 292172 326534
rect 292120 326470 292172 326476
rect 292224 326346 292252 333202
rect 292132 326318 292252 326346
rect 292132 7954 292160 326318
rect 292212 326256 292264 326262
rect 292212 326198 292264 326204
rect 292120 7948 292172 7954
rect 292120 7890 292172 7896
rect 292028 7880 292080 7886
rect 292028 7822 292080 7828
rect 292224 7818 292252 326198
rect 292212 7812 292264 7818
rect 292212 7754 292264 7760
rect 292316 3534 292344 335446
rect 292304 3528 292356 3534
rect 292304 3470 292356 3476
rect 292408 3466 292436 337742
rect 292500 336648 292528 338014
rect 292638 337770 292666 338028
rect 292822 337822 292850 338028
rect 292810 337816 292862 337822
rect 292638 337742 292712 337770
rect 292810 337758 292862 337764
rect 293006 337770 293034 338028
rect 293098 337906 293126 338028
rect 293236 338014 293296 338042
rect 293098 337878 293172 337906
rect 293006 337742 293080 337770
rect 292500 336620 292620 336648
rect 292592 336054 292620 336620
rect 292580 336048 292632 336054
rect 292580 335990 292632 335996
rect 292488 334416 292540 334422
rect 292488 334358 292540 334364
rect 292500 3602 292528 334358
rect 292684 326398 292712 337742
rect 292948 336184 293000 336190
rect 292948 336126 293000 336132
rect 292764 335708 292816 335714
rect 292764 335650 292816 335656
rect 292776 334286 292804 335650
rect 292960 335458 292988 336126
rect 293052 335918 293080 337742
rect 293040 335912 293092 335918
rect 293040 335854 293092 335860
rect 292868 335430 292988 335458
rect 292868 334422 292896 335430
rect 293144 334762 293172 337878
rect 293132 334756 293184 334762
rect 293132 334698 293184 334704
rect 293236 334642 293264 338014
rect 293374 337770 293402 338028
rect 293512 338014 293572 338042
rect 293374 337742 293448 337770
rect 293420 336734 293448 337742
rect 293408 336728 293460 336734
rect 293408 336670 293460 336676
rect 293408 335640 293460 335646
rect 293408 335582 293460 335588
rect 292960 334614 293264 334642
rect 292856 334416 292908 334422
rect 292856 334358 292908 334364
rect 292764 334280 292816 334286
rect 292764 334222 292816 334228
rect 292672 326392 292724 326398
rect 292672 326334 292724 326340
rect 292960 325694 292988 334614
rect 293224 334416 293276 334422
rect 293420 334370 293448 335582
rect 293224 334358 293276 334364
rect 293132 333260 293184 333266
rect 293132 333202 293184 333208
rect 292960 325666 293080 325694
rect 293052 304298 293080 325666
rect 293040 304292 293092 304298
rect 293040 304234 293092 304240
rect 293144 302938 293172 333202
rect 293132 302932 293184 302938
rect 293132 302874 293184 302880
rect 293236 12170 293264 334358
rect 293328 334342 293448 334370
rect 293328 13122 293356 334342
rect 293408 334280 293460 334286
rect 293408 334222 293460 334228
rect 293420 307086 293448 334222
rect 293512 319462 293540 338014
rect 293650 337906 293678 338028
rect 293788 338014 293848 338042
rect 293650 337878 293724 337906
rect 293592 337816 293644 337822
rect 293592 337758 293644 337764
rect 293604 327826 293632 337758
rect 293696 333266 293724 337878
rect 293788 335782 293816 338014
rect 293926 337770 293954 338028
rect 293880 337742 293954 337770
rect 294064 338014 294124 338042
rect 293776 335776 293828 335782
rect 293776 335718 293828 335724
rect 293776 334756 293828 334762
rect 293776 334698 293828 334704
rect 293684 333260 293736 333266
rect 293684 333202 293736 333208
rect 293788 327826 293816 334698
rect 293592 327820 293644 327826
rect 293592 327762 293644 327768
rect 293776 327820 293828 327826
rect 293776 327762 293828 327768
rect 293880 327706 293908 337742
rect 294064 335374 294092 338014
rect 294202 337770 294230 338028
rect 294340 338014 294400 338042
rect 294202 337742 294276 337770
rect 294248 335986 294276 337742
rect 294144 335980 294196 335986
rect 294144 335922 294196 335928
rect 294236 335980 294288 335986
rect 294236 335922 294288 335928
rect 294052 335368 294104 335374
rect 294052 335310 294104 335316
rect 294156 328030 294184 335922
rect 294144 328024 294196 328030
rect 294144 327966 294196 327972
rect 293604 327678 293908 327706
rect 293500 319456 293552 319462
rect 293500 319398 293552 319404
rect 293604 318102 293632 327678
rect 293684 327616 293736 327622
rect 293684 327558 293736 327564
rect 293592 318096 293644 318102
rect 293592 318038 293644 318044
rect 293408 307080 293460 307086
rect 293408 307022 293460 307028
rect 293696 305658 293724 327558
rect 294340 316034 294368 338014
rect 294570 337770 294598 338028
rect 294662 337906 294690 338028
rect 294800 338014 294860 338042
rect 294662 337878 294736 337906
rect 294570 337742 294644 337770
rect 294420 335844 294472 335850
rect 294420 335786 294472 335792
rect 294432 326534 294460 335786
rect 294616 335458 294644 337742
rect 294708 336530 294736 337878
rect 294696 336524 294748 336530
rect 294696 336466 294748 336472
rect 294800 335578 294828 338014
rect 294938 337770 294966 338028
rect 295076 338014 295136 338042
rect 294938 337742 295012 337770
rect 294788 335572 294840 335578
rect 294788 335514 294840 335520
rect 294616 335430 294920 335458
rect 294696 335368 294748 335374
rect 294696 335310 294748 335316
rect 294604 335232 294656 335238
rect 294604 335174 294656 335180
rect 294420 326528 294472 326534
rect 294420 326470 294472 326476
rect 294616 320958 294644 335174
rect 294708 325694 294736 335310
rect 294708 325666 294828 325694
rect 294604 320952 294656 320958
rect 294604 320894 294656 320900
rect 294156 316006 294368 316034
rect 293684 305652 293736 305658
rect 293684 305594 293736 305600
rect 293316 13116 293368 13122
rect 293316 13058 293368 13064
rect 293224 12164 293276 12170
rect 293224 12106 293276 12112
rect 294156 7750 294184 316006
rect 294800 12374 294828 325666
rect 294788 12368 294840 12374
rect 294788 12310 294840 12316
rect 294892 12306 294920 335430
rect 294880 12300 294932 12306
rect 294880 12242 294932 12248
rect 294880 12164 294932 12170
rect 294880 12106 294932 12112
rect 294144 7744 294196 7750
rect 294144 7686 294196 7692
rect 293684 5296 293736 5302
rect 293684 5238 293736 5244
rect 292580 5228 292632 5234
rect 292580 5170 292632 5176
rect 292488 3596 292540 3602
rect 292488 3538 292540 3544
rect 292396 3460 292448 3466
rect 292396 3402 292448 3408
rect 292592 480 292620 5170
rect 293696 480 293724 5238
rect 294892 480 294920 12106
rect 294984 12102 295012 337742
rect 295076 333266 295104 338014
rect 295214 337770 295242 338028
rect 295168 337742 295242 337770
rect 295352 338014 295412 338042
rect 295064 333260 295116 333266
rect 295064 333202 295116 333208
rect 295168 330562 295196 337742
rect 295248 335572 295300 335578
rect 295248 335514 295300 335520
rect 295076 330534 295196 330562
rect 294972 12096 295024 12102
rect 294972 12038 295024 12044
rect 295076 7614 295104 330534
rect 295260 316034 295288 335514
rect 295352 335374 295380 338014
rect 295490 337770 295518 338028
rect 295674 337770 295702 338028
rect 295766 337906 295794 338028
rect 295904 338014 295964 338042
rect 295766 337878 295840 337906
rect 295490 337742 295564 337770
rect 295674 337742 295748 337770
rect 295536 336462 295564 337742
rect 295524 336456 295576 336462
rect 295524 336398 295576 336404
rect 295340 335368 295392 335374
rect 295340 335310 295392 335316
rect 295720 330478 295748 337742
rect 295812 333198 295840 337878
rect 295904 335510 295932 338014
rect 296042 337770 296070 338028
rect 296226 337906 296254 338028
rect 296364 338014 296424 338042
rect 296226 337878 296300 337906
rect 296168 337816 296220 337822
rect 296042 337742 296116 337770
rect 296168 337758 296220 337764
rect 295892 335504 295944 335510
rect 295892 335446 295944 335452
rect 295984 335436 296036 335442
rect 295984 335378 296036 335384
rect 295892 335368 295944 335374
rect 295892 335310 295944 335316
rect 295800 333192 295852 333198
rect 295800 333134 295852 333140
rect 295708 330472 295760 330478
rect 295708 330414 295760 330420
rect 295168 316006 295288 316034
rect 295168 7682 295196 316006
rect 295904 12034 295932 335310
rect 295892 12028 295944 12034
rect 295892 11970 295944 11976
rect 295156 7676 295208 7682
rect 295156 7618 295208 7624
rect 295064 7608 295116 7614
rect 295064 7550 295116 7556
rect 295996 4554 296024 335378
rect 296088 316742 296116 337742
rect 296076 316736 296128 316742
rect 296076 316678 296128 316684
rect 296180 315314 296208 337758
rect 296272 335322 296300 337878
rect 296364 335442 296392 338014
rect 296502 337822 296530 338028
rect 296640 338014 296700 338042
rect 296490 337816 296542 337822
rect 296490 337758 296542 337764
rect 296444 335504 296496 335510
rect 296444 335446 296496 335452
rect 296352 335436 296404 335442
rect 296352 335378 296404 335384
rect 296272 335294 296392 335322
rect 296260 333192 296312 333198
rect 296260 333134 296312 333140
rect 296168 315308 296220 315314
rect 296168 315250 296220 315256
rect 296272 11966 296300 333134
rect 296260 11960 296312 11966
rect 296260 11902 296312 11908
rect 296364 11898 296392 335294
rect 296456 331906 296484 335446
rect 296444 331900 296496 331906
rect 296444 331842 296496 331848
rect 296640 330562 296668 338014
rect 296778 337770 296806 338028
rect 296962 337770 296990 338028
rect 297054 337906 297082 338028
rect 297192 338014 297252 338042
rect 297054 337878 297128 337906
rect 296778 337742 296852 337770
rect 296962 337742 297036 337770
rect 296824 335714 296852 337742
rect 296812 335708 296864 335714
rect 296812 335650 296864 335656
rect 297008 334490 297036 337742
rect 296996 334484 297048 334490
rect 296996 334426 297048 334432
rect 297100 334422 297128 337878
rect 297192 335578 297220 338014
rect 297330 337770 297358 338028
rect 297468 338014 297528 338042
rect 297330 337742 297404 337770
rect 297272 336388 297324 336394
rect 297272 336330 297324 336336
rect 297180 335572 297232 335578
rect 297180 335514 297232 335520
rect 297088 334416 297140 334422
rect 297088 334358 297140 334364
rect 297284 331214 297312 336330
rect 297376 335220 297404 337742
rect 297468 335374 297496 338014
rect 297606 337770 297634 338028
rect 297744 338014 297804 338042
rect 297606 337742 297680 337770
rect 297652 336258 297680 337742
rect 297640 336252 297692 336258
rect 297640 336194 297692 336200
rect 297456 335368 297508 335374
rect 297456 335310 297508 335316
rect 297376 335192 297680 335220
rect 297456 334552 297508 334558
rect 297456 334494 297508 334500
rect 297284 331186 297404 331214
rect 296456 330534 296668 330562
rect 296352 11892 296404 11898
rect 296352 11834 296404 11840
rect 296456 11830 296484 330534
rect 296628 330472 296680 330478
rect 296628 330414 296680 330420
rect 296640 323610 296668 330414
rect 296628 323604 296680 323610
rect 296628 323546 296680 323552
rect 296444 11824 296496 11830
rect 296444 11766 296496 11772
rect 297272 5160 297324 5166
rect 297272 5102 297324 5108
rect 296076 5092 296128 5098
rect 296076 5034 296128 5040
rect 295984 4548 296036 4554
rect 295984 4490 296036 4496
rect 296088 480 296116 5034
rect 297284 480 297312 5102
rect 297376 4214 297404 331186
rect 297468 297430 297496 334494
rect 297548 334484 297600 334490
rect 297548 334426 297600 334432
rect 297560 324970 297588 334426
rect 297548 324964 297600 324970
rect 297548 324906 297600 324912
rect 297652 322250 297680 335192
rect 297640 322244 297692 322250
rect 297640 322186 297692 322192
rect 297744 314022 297772 338014
rect 297882 337770 297910 338028
rect 297836 337742 297910 337770
rect 298020 338014 298080 338042
rect 298204 338014 298264 338042
rect 297836 334558 297864 337742
rect 297916 335368 297968 335374
rect 297916 335310 297968 335316
rect 297824 334552 297876 334558
rect 297824 334494 297876 334500
rect 297824 334416 297876 334422
rect 297824 334358 297876 334364
rect 297732 314016 297784 314022
rect 297732 313958 297784 313964
rect 297836 301510 297864 334358
rect 297824 301504 297876 301510
rect 297824 301446 297876 301452
rect 297928 300150 297956 335310
rect 298020 334558 298048 338014
rect 298204 334694 298232 338014
rect 298342 337770 298370 338028
rect 298480 338014 298540 338042
rect 298342 337742 298416 337770
rect 298192 334688 298244 334694
rect 298192 334630 298244 334636
rect 298008 334552 298060 334558
rect 298008 334494 298060 334500
rect 298388 333130 298416 337742
rect 298480 335510 298508 338014
rect 298618 337770 298646 338028
rect 298572 337742 298646 337770
rect 298802 337770 298830 338028
rect 298894 337872 298922 338028
rect 299032 338014 299092 338042
rect 298894 337844 298968 337872
rect 298802 337742 298876 337770
rect 298468 335504 298520 335510
rect 298468 335446 298520 335452
rect 298376 333124 298428 333130
rect 298376 333066 298428 333072
rect 298572 329118 298600 337742
rect 298744 335436 298796 335442
rect 298744 335378 298796 335384
rect 298652 333192 298704 333198
rect 298652 333134 298704 333140
rect 298560 329112 298612 329118
rect 298560 329054 298612 329060
rect 297916 300144 297968 300150
rect 297916 300086 297968 300092
rect 297456 297424 297508 297430
rect 297456 297366 297508 297372
rect 298664 4486 298692 333134
rect 298756 320890 298784 335378
rect 298848 330562 298876 337742
rect 298940 333198 298968 337844
rect 299032 335442 299060 338014
rect 299170 337770 299198 338028
rect 299124 337742 299198 337770
rect 299308 338014 299368 338042
rect 299020 335436 299072 335442
rect 299020 335378 299072 335384
rect 298928 333192 298980 333198
rect 298928 333134 298980 333140
rect 299020 333124 299072 333130
rect 299020 333066 299072 333072
rect 298848 330534 298968 330562
rect 298836 330472 298888 330478
rect 298836 330414 298888 330420
rect 298744 320884 298796 320890
rect 298744 320826 298796 320832
rect 298848 13530 298876 330414
rect 298940 13598 298968 330534
rect 298928 13592 298980 13598
rect 298928 13534 298980 13540
rect 298836 13524 298888 13530
rect 298836 13466 298888 13472
rect 299032 11762 299060 333066
rect 299124 330954 299152 337742
rect 299204 335368 299256 335374
rect 299204 335310 299256 335316
rect 299112 330948 299164 330954
rect 299112 330890 299164 330896
rect 299216 330698 299244 335310
rect 299124 330670 299244 330698
rect 299020 11756 299072 11762
rect 299020 11698 299072 11704
rect 299124 8906 299152 330670
rect 299308 330562 299336 338014
rect 299446 337770 299474 338028
rect 299400 337742 299474 337770
rect 299584 338014 299644 338042
rect 299400 335374 299428 337742
rect 299584 335510 299612 338014
rect 299814 337770 299842 338028
rect 299906 337906 299934 338028
rect 299906 337878 299980 337906
rect 299814 337742 299888 337770
rect 299480 335504 299532 335510
rect 299480 335446 299532 335452
rect 299572 335504 299624 335510
rect 299572 335446 299624 335452
rect 299388 335368 299440 335374
rect 299388 335310 299440 335316
rect 299492 335220 299520 335446
rect 299216 330534 299336 330562
rect 299400 335192 299520 335220
rect 299112 8900 299164 8906
rect 299112 8842 299164 8848
rect 299216 4690 299244 330534
rect 299400 316034 299428 335192
rect 299860 330410 299888 337742
rect 299952 333198 299980 337878
rect 300090 337770 300118 338028
rect 300182 337906 300210 338028
rect 300182 337878 300256 337906
rect 300090 337742 300164 337770
rect 300032 337680 300084 337686
rect 300032 337622 300084 337628
rect 299940 333192 299992 333198
rect 299940 333134 299992 333140
rect 299848 330404 299900 330410
rect 299848 330346 299900 330352
rect 299308 316006 299428 316034
rect 299204 4684 299256 4690
rect 299204 4626 299256 4632
rect 299308 4622 299336 316006
rect 300044 13326 300072 337622
rect 300136 13394 300164 337742
rect 300228 333130 300256 337878
rect 300366 337770 300394 338028
rect 300458 337890 300486 338028
rect 300446 337884 300498 337890
rect 300446 337826 300498 337832
rect 300642 337770 300670 338028
rect 300734 337890 300762 338028
rect 300872 338014 300932 338042
rect 300722 337884 300774 337890
rect 300722 337826 300774 337832
rect 300366 337742 300532 337770
rect 300642 337742 300716 337770
rect 300308 335504 300360 335510
rect 300308 335446 300360 335452
rect 300216 333124 300268 333130
rect 300216 333066 300268 333072
rect 300320 330562 300348 335446
rect 300400 333192 300452 333198
rect 300400 333134 300452 333140
rect 300228 330534 300348 330562
rect 300228 13462 300256 330534
rect 300308 330268 300360 330274
rect 300308 330210 300360 330216
rect 300216 13456 300268 13462
rect 300216 13398 300268 13404
rect 300124 13388 300176 13394
rect 300124 13330 300176 13336
rect 300032 13320 300084 13326
rect 300032 13262 300084 13268
rect 300320 9518 300348 330210
rect 300412 9654 300440 333134
rect 300400 9648 300452 9654
rect 300400 9590 300452 9596
rect 300504 9586 300532 337742
rect 300584 333124 300636 333130
rect 300584 333066 300636 333072
rect 300492 9580 300544 9586
rect 300492 9522 300544 9528
rect 300308 9512 300360 9518
rect 300308 9454 300360 9460
rect 300596 5438 300624 333066
rect 300688 330562 300716 337742
rect 300872 335374 300900 338014
rect 301010 337906 301038 338028
rect 301148 338014 301208 338042
rect 301010 337878 301084 337906
rect 300860 335368 300912 335374
rect 300860 335310 300912 335316
rect 300688 330534 300808 330562
rect 300676 330404 300728 330410
rect 300676 330346 300728 330352
rect 300688 5506 300716 330346
rect 300676 5500 300728 5506
rect 300676 5442 300728 5448
rect 300584 5432 300636 5438
rect 300584 5374 300636 5380
rect 300780 5370 300808 330534
rect 301056 330478 301084 337878
rect 301148 335510 301176 338014
rect 301286 337906 301314 338028
rect 301424 338014 301484 338042
rect 301286 337878 301360 337906
rect 301136 335504 301188 335510
rect 301136 335446 301188 335452
rect 301332 331158 301360 337878
rect 301424 335578 301452 338014
rect 301654 337770 301682 338028
rect 301746 337890 301774 338028
rect 301884 338014 301944 338042
rect 301734 337884 301786 337890
rect 301734 337826 301786 337832
rect 301654 337742 301728 337770
rect 301596 335844 301648 335850
rect 301596 335786 301648 335792
rect 301412 335572 301464 335578
rect 301412 335514 301464 335520
rect 301412 335368 301464 335374
rect 301412 335310 301464 335316
rect 301320 331152 301372 331158
rect 301320 331094 301372 331100
rect 301044 330472 301096 330478
rect 301044 330414 301096 330420
rect 301320 13796 301372 13802
rect 301320 13738 301372 13744
rect 301332 9382 301360 13738
rect 301424 13258 301452 335310
rect 301608 331214 301636 335786
rect 301516 331186 301636 331214
rect 301412 13252 301464 13258
rect 301412 13194 301464 13200
rect 301516 13122 301544 331186
rect 301596 331152 301648 331158
rect 301596 331094 301648 331100
rect 301608 13190 301636 331094
rect 301700 13802 301728 337742
rect 301780 335504 301832 335510
rect 301780 335446 301832 335452
rect 301688 13796 301740 13802
rect 301688 13738 301740 13744
rect 301688 13660 301740 13666
rect 301688 13602 301740 13608
rect 301596 13184 301648 13190
rect 301596 13126 301648 13132
rect 301504 13116 301556 13122
rect 301504 13058 301556 13064
rect 301320 9376 301372 9382
rect 301320 9318 301372 9324
rect 301700 9314 301728 13602
rect 301792 9450 301820 335446
rect 301884 335374 301912 338014
rect 302022 337770 302050 338028
rect 301976 337742 302050 337770
rect 302160 338014 302220 338042
rect 301872 335368 301924 335374
rect 301872 335310 301924 335316
rect 301976 330562 302004 337742
rect 302160 335850 302188 338014
rect 302298 337822 302326 338028
rect 302436 338014 302496 338042
rect 302286 337816 302338 337822
rect 302286 337758 302338 337764
rect 302148 335844 302200 335850
rect 302148 335786 302200 335792
rect 302056 335572 302108 335578
rect 302056 335514 302108 335520
rect 301884 330534 302004 330562
rect 301884 13666 301912 330534
rect 301964 330472 302016 330478
rect 301964 330414 302016 330420
rect 301872 13660 301924 13666
rect 301872 13602 301924 13608
rect 301872 13048 301924 13054
rect 301872 12990 301924 12996
rect 301780 9444 301832 9450
rect 301780 9386 301832 9392
rect 301688 9308 301740 9314
rect 301688 9250 301740 9256
rect 300768 5364 300820 5370
rect 300768 5306 300820 5312
rect 300768 5024 300820 5030
rect 300768 4966 300820 4972
rect 299664 4956 299716 4962
rect 299664 4898 299716 4904
rect 299296 4616 299348 4622
rect 299296 4558 299348 4564
rect 298652 4480 298704 4486
rect 298652 4422 298704 4428
rect 297364 4208 297416 4214
rect 297364 4150 297416 4156
rect 298468 4208 298520 4214
rect 298468 4150 298520 4156
rect 298480 480 298508 4150
rect 299676 480 299704 4898
rect 300780 480 300808 4966
rect 301884 3482 301912 12990
rect 301976 5302 302004 330414
rect 301964 5296 302016 5302
rect 301964 5238 302016 5244
rect 302068 5234 302096 335514
rect 302436 335442 302464 338014
rect 302574 337770 302602 338028
rect 302528 337742 302602 337770
rect 302758 337770 302786 338028
rect 302850 337906 302878 338028
rect 302988 338014 303048 338042
rect 302850 337878 302924 337906
rect 302758 337742 302832 337770
rect 302424 335436 302476 335442
rect 302424 335378 302476 335384
rect 302148 335368 302200 335374
rect 302148 335310 302200 335316
rect 302056 5228 302108 5234
rect 302056 5170 302108 5176
rect 302160 5166 302188 335310
rect 302528 330546 302556 337742
rect 302700 335640 302752 335646
rect 302700 335582 302752 335588
rect 302516 330540 302568 330546
rect 302516 330482 302568 330488
rect 302148 5160 302200 5166
rect 302148 5102 302200 5108
rect 302712 4758 302740 335582
rect 302804 5030 302832 337742
rect 302896 330478 302924 337878
rect 302988 335510 303016 338014
rect 303126 337770 303154 338028
rect 303264 338014 303324 338042
rect 303448 338014 303508 338042
rect 303126 337742 303200 337770
rect 302976 335504 303028 335510
rect 302976 335446 303028 335452
rect 303068 335436 303120 335442
rect 303068 335378 303120 335384
rect 302976 335368 303028 335374
rect 302976 335310 303028 335316
rect 302884 330472 302936 330478
rect 302884 330414 302936 330420
rect 302884 327140 302936 327146
rect 302884 327082 302936 327088
rect 302896 311166 302924 327082
rect 302884 311160 302936 311166
rect 302884 311102 302936 311108
rect 302988 9110 303016 335310
rect 303080 9246 303108 335378
rect 303172 330562 303200 337742
rect 303264 335374 303292 338014
rect 303344 337816 303396 337822
rect 303344 337758 303396 337764
rect 303252 335368 303304 335374
rect 303252 335310 303304 335316
rect 303172 330534 303292 330562
rect 303160 330472 303212 330478
rect 303160 330414 303212 330420
rect 303068 9240 303120 9246
rect 303068 9182 303120 9188
rect 303172 9178 303200 330414
rect 303160 9172 303212 9178
rect 303160 9114 303212 9120
rect 302976 9104 303028 9110
rect 302976 9046 303028 9052
rect 302792 5024 302844 5030
rect 302792 4966 302844 4972
rect 303264 4962 303292 330534
rect 303356 5098 303384 337758
rect 303448 327146 303476 338014
rect 303586 337770 303614 338028
rect 303540 337742 303614 337770
rect 303770 337770 303798 338028
rect 303862 337958 303890 338028
rect 303850 337952 303902 337958
rect 303850 337894 303902 337900
rect 304046 337770 304074 338028
rect 304138 337906 304166 338028
rect 304276 338014 304336 338042
rect 304138 337878 304212 337906
rect 303770 337742 303844 337770
rect 304046 337742 304120 337770
rect 303540 335646 303568 337742
rect 303528 335640 303580 335646
rect 303528 335582 303580 335588
rect 303528 335504 303580 335510
rect 303528 335446 303580 335452
rect 303540 327758 303568 335446
rect 303816 330478 303844 337742
rect 304092 334558 304120 337742
rect 304184 335374 304212 337878
rect 304172 335368 304224 335374
rect 304172 335310 304224 335316
rect 304080 334552 304132 334558
rect 304080 334494 304132 334500
rect 303804 330472 303856 330478
rect 303804 330414 303856 330420
rect 303528 327752 303580 327758
rect 303528 327694 303580 327700
rect 303436 327140 303488 327146
rect 303436 327082 303488 327088
rect 304276 313954 304304 338014
rect 304414 337822 304442 338028
rect 304552 338014 304612 338042
rect 304402 337816 304454 337822
rect 304402 337758 304454 337764
rect 304552 335442 304580 338014
rect 304690 337770 304718 338028
rect 304644 337742 304718 337770
rect 304828 338014 304888 338042
rect 304540 335436 304592 335442
rect 304540 335378 304592 335384
rect 304356 335368 304408 335374
rect 304356 335310 304408 335316
rect 304264 313948 304316 313954
rect 304264 313890 304316 313896
rect 304368 8974 304396 335310
rect 304448 334552 304500 334558
rect 304448 334494 304500 334500
rect 304460 330562 304488 334494
rect 304460 330534 304580 330562
rect 304448 330472 304500 330478
rect 304448 330414 304500 330420
rect 304460 9042 304488 330414
rect 304448 9036 304500 9042
rect 304448 8978 304500 8984
rect 304356 8968 304408 8974
rect 304356 8910 304408 8916
rect 303344 5092 303396 5098
rect 303344 5034 303396 5040
rect 303252 4956 303304 4962
rect 303252 4898 303304 4904
rect 303160 4888 303212 4894
rect 303160 4830 303212 4836
rect 302700 4752 302752 4758
rect 302700 4694 302752 4700
rect 301884 3454 302004 3482
rect 301976 480 302004 3454
rect 303172 480 303200 4830
rect 304552 4826 304580 330534
rect 304356 4820 304408 4826
rect 304356 4762 304408 4768
rect 304540 4820 304592 4826
rect 304540 4762 304592 4768
rect 304368 480 304396 4762
rect 304644 3505 304672 337742
rect 304828 330698 304856 338014
rect 305828 337952 305880 337958
rect 305828 337894 305880 337900
rect 305000 337816 305052 337822
rect 305000 337758 305052 337764
rect 304908 335436 304960 335442
rect 304908 335378 304960 335384
rect 304736 330670 304856 330698
rect 304630 3496 304686 3505
rect 304630 3431 304686 3440
rect 304736 3369 304764 330670
rect 304920 330562 304948 335378
rect 304828 330534 304948 330562
rect 304828 3641 304856 330534
rect 305012 330460 305040 337758
rect 305736 335912 305788 335918
rect 305736 335854 305788 335860
rect 305092 335844 305144 335850
rect 305092 335786 305144 335792
rect 305104 330614 305132 335786
rect 305184 335708 305236 335714
rect 305184 335650 305236 335656
rect 305092 330608 305144 330614
rect 305092 330550 305144 330556
rect 304920 330432 305040 330460
rect 304920 3777 304948 330432
rect 305196 329186 305224 335650
rect 305644 334756 305696 334762
rect 305644 334698 305696 334704
rect 305000 329180 305052 329186
rect 305000 329122 305052 329128
rect 305184 329180 305236 329186
rect 305184 329122 305236 329128
rect 305012 16574 305040 329122
rect 305012 16546 305592 16574
rect 304906 3768 304962 3777
rect 304906 3703 304962 3712
rect 304814 3632 304870 3641
rect 304814 3567 304870 3576
rect 304722 3360 304778 3369
rect 304722 3295 304778 3304
rect 305564 480 305592 16546
rect 305656 14618 305684 334698
rect 305748 181490 305776 335854
rect 305840 294642 305868 337894
rect 305920 337884 305972 337890
rect 305920 337826 305972 337832
rect 305932 296002 305960 337826
rect 306288 335776 306340 335782
rect 306288 335718 306340 335724
rect 306300 334762 306328 335718
rect 306288 334756 306340 334762
rect 306288 334698 306340 334704
rect 306392 325650 306420 369815
rect 306470 368520 306526 368529
rect 306470 368455 306526 368464
rect 306380 325644 306432 325650
rect 306380 325586 306432 325592
rect 306484 313274 306512 368455
rect 306562 367296 306618 367305
rect 306562 367231 306618 367240
rect 306472 313268 306524 313274
rect 306472 313210 306524 313216
rect 306576 299470 306604 367231
rect 307036 364334 307064 372671
rect 307128 365702 307156 374031
rect 307666 371376 307722 371385
rect 307666 371311 307722 371320
rect 307680 371278 307708 371311
rect 307668 371272 307720 371278
rect 307668 371214 307720 371220
rect 320824 371272 320876 371278
rect 320824 371214 320876 371220
rect 307666 366072 307722 366081
rect 307666 366007 307722 366016
rect 307680 365770 307708 366007
rect 307668 365764 307720 365770
rect 307668 365706 307720 365712
rect 307116 365696 307168 365702
rect 307116 365638 307168 365644
rect 307666 364712 307722 364721
rect 307666 364647 307722 364656
rect 307680 364410 307708 364647
rect 307668 364404 307720 364410
rect 307668 364346 307720 364352
rect 316684 364404 316736 364410
rect 316684 364346 316736 364352
rect 307036 364306 307156 364334
rect 306654 361720 306710 361729
rect 306654 361655 306710 361664
rect 306564 299464 306616 299470
rect 306564 299406 306616 299412
rect 305920 295996 305972 296002
rect 305920 295938 305972 295944
rect 305828 294636 305880 294642
rect 305828 294578 305880 294584
rect 306668 245614 306696 361655
rect 306746 360496 306802 360505
rect 306746 360431 306802 360440
rect 306656 245608 306708 245614
rect 306656 245550 306708 245556
rect 306760 233238 306788 360431
rect 306838 359136 306894 359145
rect 306838 359071 306894 359080
rect 306748 233232 306800 233238
rect 306748 233174 306800 233180
rect 306852 219434 306880 359071
rect 306930 357912 306986 357921
rect 306930 357847 306986 357856
rect 306840 219428 306892 219434
rect 306840 219370 306892 219376
rect 306944 206990 306972 357847
rect 307128 353258 307156 364306
rect 307298 363352 307354 363361
rect 307298 363287 307354 363296
rect 307312 362982 307340 363287
rect 307300 362976 307352 362982
rect 307300 362918 307352 362924
rect 307666 356552 307722 356561
rect 307666 356487 307722 356496
rect 307680 356386 307708 356487
rect 307668 356380 307720 356386
rect 307668 356322 307720 356328
rect 309784 356380 309836 356386
rect 309784 356322 309836 356328
rect 307666 355192 307722 355201
rect 307666 355127 307722 355136
rect 307680 354754 307708 355127
rect 307668 354748 307720 354754
rect 307668 354690 307720 354696
rect 307666 353832 307722 353841
rect 307666 353767 307722 353776
rect 307116 353252 307168 353258
rect 307116 353194 307168 353200
rect 307574 352472 307630 352481
rect 307574 352407 307630 352416
rect 307482 351248 307538 351257
rect 307482 351183 307538 351192
rect 307390 349888 307446 349897
rect 307390 349823 307446 349832
rect 307298 348528 307354 348537
rect 307298 348463 307354 348472
rect 307022 346624 307078 346633
rect 307022 346559 307078 346568
rect 307036 336394 307064 346559
rect 307206 345264 307262 345273
rect 307206 345199 307262 345208
rect 307220 345014 307248 345199
rect 307128 344986 307248 345014
rect 307024 336388 307076 336394
rect 307024 336330 307076 336336
rect 307024 335912 307076 335918
rect 307024 335854 307076 335860
rect 306932 206984 306984 206990
rect 306932 206926 306984 206932
rect 305736 181484 305788 181490
rect 305736 181426 305788 181432
rect 307036 60722 307064 335854
rect 307128 73166 307156 344986
rect 307206 343904 307262 343913
rect 307206 343839 307262 343848
rect 307220 339794 307248 343839
rect 307208 339788 307260 339794
rect 307208 339730 307260 339736
rect 307206 339688 307262 339697
rect 307206 339623 307262 339632
rect 307220 339522 307248 339623
rect 307208 339516 307260 339522
rect 307208 339458 307260 339464
rect 307206 338328 307262 338337
rect 307206 338263 307262 338272
rect 307220 338162 307248 338263
rect 307208 338156 307260 338162
rect 307208 338098 307260 338104
rect 307208 336388 307260 336394
rect 307208 336330 307260 336336
rect 307220 86970 307248 336330
rect 307312 113150 307340 348463
rect 307404 126954 307432 349823
rect 307496 139398 307524 351183
rect 307588 153202 307616 352407
rect 307680 348106 307708 353767
rect 307680 348078 307800 348106
rect 307666 347984 307722 347993
rect 307666 347919 307722 347928
rect 307680 347818 307708 347919
rect 307668 347812 307720 347818
rect 307668 347754 307720 347760
rect 307772 347698 307800 348078
rect 307680 347670 307800 347698
rect 307680 167006 307708 347670
rect 307760 335096 307812 335102
rect 307760 335038 307812 335044
rect 307668 167000 307720 167006
rect 307668 166942 307720 166948
rect 307576 153196 307628 153202
rect 307576 153138 307628 153144
rect 307484 139392 307536 139398
rect 307484 139334 307536 139340
rect 307392 126948 307444 126954
rect 307392 126890 307444 126896
rect 307300 113144 307352 113150
rect 307300 113086 307352 113092
rect 307208 86964 307260 86970
rect 307208 86906 307260 86912
rect 307116 73160 307168 73166
rect 307116 73102 307168 73108
rect 307024 60716 307076 60722
rect 307024 60658 307076 60664
rect 305644 14612 305696 14618
rect 305644 14554 305696 14560
rect 306748 14612 306800 14618
rect 306748 14554 306800 14560
rect 306760 480 306788 14554
rect 307772 4214 307800 335038
rect 309140 335028 309192 335034
rect 309140 334970 309192 334976
rect 309152 16574 309180 334970
rect 309796 193186 309824 356322
rect 312544 336728 312596 336734
rect 312544 336670 312596 336676
rect 311900 325168 311952 325174
rect 311900 325110 311952 325116
rect 309784 193180 309836 193186
rect 309784 193122 309836 193128
rect 309152 16546 310284 16574
rect 307944 8424 307996 8430
rect 307944 8366 307996 8372
rect 307760 4208 307812 4214
rect 307760 4150 307812 4156
rect 307956 480 307984 8366
rect 309048 4208 309100 4214
rect 309048 4150 309100 4156
rect 309060 480 309088 4150
rect 310256 480 310284 16546
rect 311440 8492 311492 8498
rect 311440 8434 311492 8440
rect 311452 480 311480 8434
rect 311912 6914 311940 325110
rect 312556 14482 312584 336670
rect 313924 335980 313976 335986
rect 313924 335922 313976 335928
rect 313280 335164 313332 335170
rect 313280 335106 313332 335112
rect 313292 16574 313320 335106
rect 313292 16546 313872 16574
rect 312544 14476 312596 14482
rect 312544 14418 312596 14424
rect 311912 6886 312676 6914
rect 312648 480 312676 6886
rect 313844 480 313872 16546
rect 313936 15910 313964 335922
rect 316040 333668 316092 333674
rect 316040 333610 316092 333616
rect 313924 15904 313976 15910
rect 313924 15846 313976 15852
rect 315028 8560 315080 8566
rect 315028 8502 315080 8508
rect 315040 480 315068 8502
rect 316052 4214 316080 333610
rect 316132 321156 316184 321162
rect 316132 321098 316184 321104
rect 316144 16574 316172 321098
rect 316696 273222 316724 364346
rect 320836 340202 320864 371214
rect 461584 365764 461636 365770
rect 461584 365706 461636 365712
rect 331864 362976 331916 362982
rect 331864 362918 331916 362924
rect 324964 354748 325016 354754
rect 324964 354690 325016 354696
rect 323584 347812 323636 347818
rect 323584 347754 323636 347760
rect 320824 340196 320876 340202
rect 320824 340138 320876 340144
rect 318064 339516 318116 339522
rect 318064 339458 318116 339464
rect 316684 273216 316736 273222
rect 316684 273158 316736 273164
rect 318076 20670 318104 339458
rect 320824 336524 320876 336530
rect 320824 336466 320876 336472
rect 320180 332240 320232 332246
rect 320180 332182 320232 332188
rect 318800 319660 318852 319666
rect 318800 319602 318852 319608
rect 318064 20664 318116 20670
rect 318064 20606 318116 20612
rect 318812 16574 318840 319602
rect 320192 16574 320220 332182
rect 320836 17270 320864 336466
rect 322204 336456 322256 336462
rect 322204 336398 322256 336404
rect 322216 18630 322244 336398
rect 322940 323876 322992 323882
rect 322940 323818 322992 323824
rect 322204 18624 322256 18630
rect 322204 18566 322256 18572
rect 320824 17264 320876 17270
rect 320824 17206 320876 17212
rect 322952 16574 322980 323818
rect 323596 100706 323624 347754
rect 324320 333532 324372 333538
rect 324320 333474 324372 333480
rect 323584 100700 323636 100706
rect 323584 100642 323636 100648
rect 324332 16574 324360 333474
rect 324976 179382 325004 354690
rect 327724 336320 327776 336326
rect 327724 336262 327776 336268
rect 327080 330880 327132 330886
rect 327080 330822 327132 330828
rect 325700 312656 325752 312662
rect 325700 312598 325752 312604
rect 324964 179376 325016 179382
rect 324964 179318 325016 179324
rect 325712 16574 325740 312598
rect 327092 16574 327120 330822
rect 327736 21418 327764 336262
rect 331220 328024 331272 328030
rect 331220 327966 331272 327972
rect 329840 318300 329892 318306
rect 329840 318242 329892 318248
rect 327724 21412 327776 21418
rect 327724 21354 327776 21360
rect 329852 16574 329880 318242
rect 331232 16574 331260 327966
rect 331876 259418 331904 362918
rect 460204 342304 460256 342310
rect 460204 342246 460256 342252
rect 406384 338156 406436 338162
rect 406384 338098 406436 338104
rect 336004 336184 336056 336190
rect 336004 336126 336056 336132
rect 333980 334960 334032 334966
rect 333980 334902 334032 334908
rect 332600 330812 332652 330818
rect 332600 330754 332652 330760
rect 331864 259412 331916 259418
rect 331864 259354 331916 259360
rect 316144 16546 316264 16574
rect 318812 16546 319760 16574
rect 320192 16546 320956 16574
rect 322952 16546 323348 16574
rect 324332 16546 324452 16574
rect 325712 16546 326844 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 331232 16546 331628 16574
rect 316040 4208 316092 4214
rect 316040 4150 316092 4156
rect 316236 480 316264 16546
rect 318524 8628 318576 8634
rect 318524 8570 318576 8576
rect 317328 4208 317380 4214
rect 317328 4150 317380 4156
rect 317340 480 317368 4150
rect 318536 480 318564 8570
rect 319732 480 319760 16546
rect 320928 480 320956 16546
rect 322112 8696 322164 8702
rect 322112 8638 322164 8644
rect 322124 480 322152 8638
rect 323320 480 323348 16546
rect 324424 480 324452 16546
rect 325608 8764 325660 8770
rect 325608 8706 325660 8712
rect 325620 480 325648 8706
rect 326816 480 326844 16546
rect 328012 480 328040 16546
rect 329196 8832 329248 8838
rect 329196 8774 329248 8780
rect 329208 480 329236 8774
rect 330404 480 330432 16546
rect 331600 480 331628 16546
rect 332612 3482 332640 330754
rect 332692 316872 332744 316878
rect 332692 316814 332744 316820
rect 332704 4214 332732 316814
rect 333992 16574 334020 334902
rect 335360 334892 335412 334898
rect 335360 334834 335412 334840
rect 335372 16574 335400 334834
rect 336016 22778 336044 336126
rect 400864 336116 400916 336122
rect 400864 336058 400916 336064
rect 368480 334824 368532 334830
rect 368480 334766 368532 334772
rect 338120 333600 338172 333606
rect 338120 333542 338172 333548
rect 336740 321088 336792 321094
rect 336740 321030 336792 321036
rect 336004 22772 336056 22778
rect 336004 22714 336056 22720
rect 336752 16574 336780 321030
rect 338132 16574 338160 333542
rect 342260 332172 342312 332178
rect 342260 332114 342312 332120
rect 339500 329384 339552 329390
rect 339500 329326 339552 329332
rect 339512 16574 339540 329326
rect 340880 309868 340932 309874
rect 340880 309810 340932 309816
rect 340892 16574 340920 309810
rect 342272 16574 342300 332114
rect 347780 332104 347832 332110
rect 347780 332046 347832 332052
rect 346400 326664 346452 326670
rect 346400 326606 346452 326612
rect 343640 314084 343692 314090
rect 343640 314026 343692 314032
rect 343652 16574 343680 314026
rect 346412 16574 346440 326606
rect 347792 16574 347820 332046
rect 357440 330744 357492 330750
rect 357440 330686 357492 330692
rect 353300 327956 353352 327962
rect 353300 327898 353352 327904
rect 349160 325100 349212 325106
rect 349160 325042 349212 325048
rect 333992 16546 335124 16574
rect 335372 16546 336320 16574
rect 336752 16546 337516 16574
rect 338132 16546 338712 16574
rect 339512 16546 339908 16574
rect 340892 16546 341012 16574
rect 342272 16546 343404 16574
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 332692 4208 332744 4214
rect 332692 4150 332744 4156
rect 333888 4208 333940 4214
rect 333888 4150 333940 4156
rect 332612 3454 332732 3482
rect 332704 480 332732 3454
rect 333900 480 333928 4150
rect 335096 480 335124 16546
rect 336292 480 336320 16546
rect 337488 480 337516 16546
rect 338684 480 338712 16546
rect 339880 480 339908 16546
rect 340984 480 341012 16546
rect 342168 5704 342220 5710
rect 342168 5646 342220 5652
rect 342180 480 342208 5646
rect 343376 480 343404 16546
rect 344572 480 344600 16546
rect 345756 5772 345808 5778
rect 345756 5714 345808 5720
rect 345768 480 345796 5714
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 4214 349200 325042
rect 350540 293276 350592 293282
rect 350540 293218 350592 293224
rect 350552 16574 350580 293218
rect 353312 16574 353340 327898
rect 354680 312588 354732 312594
rect 354680 312530 354732 312536
rect 354692 16574 354720 312530
rect 350552 16546 351684 16574
rect 353312 16546 354076 16574
rect 354692 16546 355272 16574
rect 349252 5840 349304 5846
rect 349252 5782 349304 5788
rect 349160 4208 349212 4214
rect 349160 4150 349212 4156
rect 349264 480 349292 5782
rect 350448 4208 350500 4214
rect 350448 4150 350500 4156
rect 350460 480 350488 4150
rect 351656 480 351684 16546
rect 352840 5908 352892 5914
rect 352840 5850 352892 5856
rect 352852 480 352880 5850
rect 354048 480 354076 16546
rect 355244 480 355272 16546
rect 356336 5976 356388 5982
rect 356336 5918 356388 5924
rect 356348 480 356376 5918
rect 357452 3482 357480 330686
rect 365720 329316 365772 329322
rect 365720 329258 365772 329264
rect 357532 325032 357584 325038
rect 357532 324974 357584 324980
rect 357544 4214 357572 324974
rect 360200 323808 360252 323814
rect 360200 323750 360252 323756
rect 360212 16574 360240 323750
rect 361580 291848 361632 291854
rect 361580 291790 361632 291796
rect 361592 16574 361620 291790
rect 365732 16574 365760 329258
rect 368492 16574 368520 334766
rect 372620 333464 372672 333470
rect 372620 333406 372672 333412
rect 372632 16574 372660 333406
rect 375380 326596 375432 326602
rect 375380 326538 375432 326544
rect 375392 16574 375420 326538
rect 393320 323740 393372 323746
rect 393320 323682 393372 323688
rect 379520 322448 379572 322454
rect 379520 322390 379572 322396
rect 379532 16574 379560 322390
rect 382280 319592 382332 319598
rect 382280 319534 382332 319540
rect 360212 16546 361160 16574
rect 361592 16546 362356 16574
rect 365732 16546 365852 16574
rect 368492 16546 369440 16574
rect 372632 16546 372936 16574
rect 375392 16546 376524 16574
rect 379532 16546 380020 16574
rect 359924 6044 359976 6050
rect 359924 5986 359976 5992
rect 357532 4208 357584 4214
rect 357532 4150 357584 4156
rect 358728 4208 358780 4214
rect 358728 4150 358780 4156
rect 357452 3454 357572 3482
rect 357544 480 357572 3454
rect 358740 480 358768 4150
rect 359936 480 359964 5986
rect 361132 480 361160 16546
rect 362328 480 362356 16546
rect 364616 9784 364668 9790
rect 364616 9726 364668 9732
rect 363512 6112 363564 6118
rect 363512 6054 363564 6060
rect 363524 480 363552 6054
rect 364628 480 364656 9726
rect 365824 480 365852 16546
rect 368204 9852 368256 9858
rect 368204 9794 368256 9800
rect 367008 6860 367060 6866
rect 367008 6802 367060 6808
rect 367020 480 367048 6802
rect 368216 480 368244 9794
rect 369412 480 369440 16546
rect 371700 9920 371752 9926
rect 371700 9862 371752 9868
rect 370596 6792 370648 6798
rect 370596 6734 370648 6740
rect 370608 480 370636 6734
rect 371712 480 371740 9862
rect 372908 480 372936 16546
rect 374000 9988 374052 9994
rect 374000 9930 374052 9936
rect 374012 4214 374040 9930
rect 374092 6724 374144 6730
rect 374092 6666 374144 6672
rect 374000 4208 374052 4214
rect 374000 4150 374052 4156
rect 374104 480 374132 6666
rect 375288 4208 375340 4214
rect 375288 4150 375340 4156
rect 375300 480 375328 4150
rect 376496 480 376524 16546
rect 378876 10056 378928 10062
rect 378876 9998 378928 10004
rect 377680 6656 377732 6662
rect 377680 6598 377732 6604
rect 377692 480 377720 6598
rect 378888 480 378916 9998
rect 379992 480 380020 16546
rect 381176 6588 381228 6594
rect 381176 6530 381228 6536
rect 381188 480 381216 6530
rect 382292 4214 382320 319534
rect 386420 315444 386472 315450
rect 386420 315386 386472 315392
rect 386432 16574 386460 315386
rect 390560 308508 390612 308514
rect 390560 308450 390612 308456
rect 390572 16574 390600 308450
rect 393332 16574 393360 323682
rect 397460 321020 397512 321026
rect 397460 320962 397512 320968
rect 397472 16574 397500 320962
rect 400220 318232 400272 318238
rect 400220 318174 400272 318180
rect 400232 16574 400260 318174
rect 386432 16546 387196 16574
rect 390572 16546 390692 16574
rect 393332 16546 394280 16574
rect 397472 16546 397776 16574
rect 400232 16546 400812 16574
rect 385960 10192 386012 10198
rect 385960 10134 386012 10140
rect 382372 10124 382424 10130
rect 382372 10066 382424 10072
rect 382280 4208 382332 4214
rect 382280 4150 382332 4156
rect 382384 480 382412 10066
rect 384764 6520 384816 6526
rect 384764 6462 384816 6468
rect 383568 4208 383620 4214
rect 383568 4150 383620 4156
rect 383580 480 383608 4150
rect 384776 480 384804 6462
rect 385972 480 386000 10134
rect 387168 480 387196 16546
rect 389456 10260 389508 10266
rect 389456 10202 389508 10208
rect 388260 6452 388312 6458
rect 388260 6394 388312 6400
rect 388272 480 388300 6394
rect 389468 480 389496 10202
rect 390664 480 390692 16546
rect 393044 11008 393096 11014
rect 393044 10950 393096 10956
rect 391848 6384 391900 6390
rect 391848 6326 391900 6332
rect 391860 480 391888 6326
rect 393056 480 393084 10950
rect 394252 480 394280 16546
rect 396540 10940 396592 10946
rect 396540 10882 396592 10888
rect 395344 6316 395396 6322
rect 395344 6258 395396 6264
rect 395356 480 395384 6258
rect 396552 480 396580 10882
rect 397748 480 397776 16546
rect 398840 10872 398892 10878
rect 398840 10814 398892 10820
rect 398852 4214 398880 10814
rect 398932 6248 398984 6254
rect 398932 6190 398984 6196
rect 398840 4208 398892 4214
rect 398840 4150 398892 4156
rect 398944 480 398972 6190
rect 400128 4208 400180 4214
rect 400128 4150 400180 4156
rect 400140 480 400168 4150
rect 400784 3482 400812 16546
rect 400876 6254 400904 336058
rect 405740 332036 405792 332042
rect 405740 331978 405792 331984
rect 404360 307148 404412 307154
rect 404360 307090 404412 307096
rect 404372 16574 404400 307090
rect 405752 16574 405780 331978
rect 404372 16546 404860 16574
rect 405752 16546 406056 16574
rect 403624 10804 403676 10810
rect 403624 10746 403676 10752
rect 400864 6248 400916 6254
rect 400864 6190 400916 6196
rect 402520 6180 402572 6186
rect 402520 6122 402572 6128
rect 400784 3454 401364 3482
rect 401336 480 401364 3454
rect 402532 480 402560 6122
rect 403636 480 403664 10746
rect 404832 480 404860 16546
rect 406028 480 406056 16546
rect 406396 6866 406424 338098
rect 426440 333396 426492 333402
rect 426440 333338 426492 333344
rect 423680 330676 423732 330682
rect 423680 330618 423732 330624
rect 419540 329248 419592 329254
rect 419540 329190 419592 329196
rect 415492 327888 415544 327894
rect 415492 327830 415544 327836
rect 412640 326528 412692 326534
rect 412640 326470 412692 326476
rect 407120 305720 407172 305726
rect 407120 305662 407172 305668
rect 406384 6860 406436 6866
rect 406384 6802 406436 6808
rect 407132 2854 407160 305662
rect 412652 16574 412680 326470
rect 412652 16546 413140 16574
rect 407212 10736 407264 10742
rect 407212 10678 407264 10684
rect 407120 2848 407172 2854
rect 407120 2790 407172 2796
rect 407224 480 407252 10678
rect 410800 10668 410852 10674
rect 410800 10610 410852 10616
rect 409604 6248 409656 6254
rect 409604 6190 409656 6196
rect 408408 2848 408460 2854
rect 408408 2790 408460 2796
rect 408420 480 408448 2790
rect 409616 480 409644 6190
rect 410812 480 410840 10610
rect 411904 2848 411956 2854
rect 411904 2790 411956 2796
rect 411916 480 411944 2790
rect 413112 480 413140 16546
rect 414296 10600 414348 10606
rect 414296 10542 414348 10548
rect 414308 480 414336 10542
rect 415504 2990 415532 327830
rect 419552 16574 419580 329190
rect 419552 16546 420224 16574
rect 417884 10532 417936 10538
rect 417884 10474 417936 10480
rect 415492 2984 415544 2990
rect 415492 2926 415544 2932
rect 416688 2984 416740 2990
rect 416688 2926 416740 2932
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 415504 480 415532 2790
rect 416700 480 416728 2926
rect 417896 480 417924 10474
rect 418988 2916 419040 2922
rect 418988 2858 419040 2864
rect 419000 480 419028 2858
rect 420196 480 420224 16546
rect 421380 10464 421432 10470
rect 421380 10406 421432 10412
rect 421392 480 421420 10406
rect 423692 3482 423720 330618
rect 426452 16574 426480 333338
rect 434720 333328 434772 333334
rect 434720 333270 434772 333276
rect 430580 323672 430632 323678
rect 430580 323614 430632 323620
rect 430592 16574 430620 323614
rect 433340 322380 433392 322386
rect 433340 322322 433392 322328
rect 432052 311228 432104 311234
rect 432052 311170 432104 311176
rect 426452 16546 427308 16574
rect 430592 16546 430896 16574
rect 423772 10396 423824 10402
rect 423772 10338 423824 10344
rect 423784 4214 423812 10338
rect 423772 4208 423824 4214
rect 423772 4150 423824 4156
rect 424968 4208 425020 4214
rect 424968 4150 425020 4156
rect 423692 3454 423812 3482
rect 422576 3052 422628 3058
rect 422576 2994 422628 3000
rect 422588 480 422616 2994
rect 423784 480 423812 3454
rect 424980 480 425008 4150
rect 426164 3120 426216 3126
rect 426164 3062 426216 3068
rect 426176 480 426204 3062
rect 427280 480 427308 16546
rect 428464 10328 428516 10334
rect 428464 10270 428516 10276
rect 428476 480 428504 10270
rect 429660 3188 429712 3194
rect 429660 3130 429712 3136
rect 429672 480 429700 3130
rect 430868 480 430896 16546
rect 432064 480 432092 311170
rect 433352 16574 433380 322322
rect 434732 16574 434760 333270
rect 441620 326460 441672 326466
rect 441620 326402 441672 326408
rect 438860 319524 438912 319530
rect 438860 319466 438912 319472
rect 438872 16574 438900 319466
rect 441632 16574 441660 326402
rect 458180 320952 458232 320958
rect 458180 320894 458232 320900
rect 448520 318164 448572 318170
rect 448520 318106 448572 318112
rect 445760 309800 445812 309806
rect 445760 309742 445812 309748
rect 445772 16574 445800 309742
rect 433352 16546 434484 16574
rect 434732 16546 435588 16574
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 445772 16546 446260 16574
rect 433248 3256 433300 3262
rect 433248 3198 433300 3204
rect 433260 480 433288 3198
rect 434456 480 434484 16546
rect 435560 480 435588 16546
rect 437940 7540 437992 7546
rect 437940 7482 437992 7488
rect 436744 3324 436796 3330
rect 436744 3266 436796 3272
rect 436756 480 436784 3266
rect 437952 480 437980 7482
rect 439148 480 439176 16546
rect 441528 8288 441580 8294
rect 441528 8230 441580 8236
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 440344 480 440372 3334
rect 441540 480 441568 8230
rect 442644 480 442672 16546
rect 445024 8220 445076 8226
rect 445024 8162 445076 8168
rect 443828 4140 443880 4146
rect 443828 4082 443880 4088
rect 443840 480 443868 4082
rect 445036 480 445064 8162
rect 446232 480 446260 16546
rect 447416 4072 447468 4078
rect 447416 4014 447468 4020
rect 447428 480 447456 4014
rect 448532 3398 448560 318106
rect 452660 316804 452712 316810
rect 452660 316746 452712 316752
rect 452672 16574 452700 316746
rect 456892 308440 456944 308446
rect 456892 308382 456944 308388
rect 452672 16546 453344 16574
rect 448612 8152 448664 8158
rect 448612 8094 448664 8100
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 448624 480 448652 8094
rect 452108 8084 452160 8090
rect 452108 8026 452160 8032
rect 450912 4004 450964 4010
rect 450912 3946 450964 3952
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 450924 480 450952 3946
rect 452120 480 452148 8026
rect 453316 480 453344 16546
rect 455696 8016 455748 8022
rect 455696 7958 455748 7964
rect 454500 3936 454552 3942
rect 454500 3878 454552 3884
rect 454512 480 454540 3878
rect 455708 480 455736 7958
rect 456904 480 456932 308382
rect 458192 16574 458220 320894
rect 459560 307080 459612 307086
rect 459560 307022 459612 307028
rect 459572 16574 459600 307022
rect 460216 46918 460244 342246
rect 461596 285666 461624 365706
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 340196 580224 340202
rect 580172 340138 580224 340144
rect 580184 338609 580212 340138
rect 580170 338600 580226 338609
rect 580170 338535 580226 338544
rect 479524 336048 479576 336054
rect 479524 335990 479576 335996
rect 465172 331968 465224 331974
rect 465172 331910 465224 331916
rect 463700 322312 463752 322318
rect 463700 322254 463752 322260
rect 461584 285660 461636 285666
rect 461584 285602 461636 285608
rect 460204 46912 460256 46918
rect 460204 46854 460256 46860
rect 462320 22772 462372 22778
rect 462320 22714 462372 22720
rect 462332 16574 462360 22714
rect 463712 16574 463740 322254
rect 465184 16574 465212 331910
rect 466460 315376 466512 315382
rect 466460 315318 466512 315324
rect 466472 16574 466500 315318
rect 458192 16546 459232 16574
rect 459572 16546 460428 16574
rect 462332 16546 462820 16574
rect 463712 16546 464016 16574
rect 465184 16546 466316 16574
rect 466472 16546 467512 16574
rect 458088 3868 458140 3874
rect 458088 3810 458140 3816
rect 458100 480 458128 3810
rect 459204 480 459232 16546
rect 460400 480 460428 16546
rect 461584 3800 461636 3806
rect 461584 3742 461636 3748
rect 461596 480 461624 3742
rect 462792 480 462820 16546
rect 463988 480 464016 16546
rect 465172 3732 465224 3738
rect 465172 3674 465224 3680
rect 465184 480 465212 3674
rect 466288 480 466316 16546
rect 467484 480 467512 16546
rect 471060 12436 471112 12442
rect 471060 12378 471112 12384
rect 469864 7948 469916 7954
rect 469864 7890 469916 7896
rect 468668 3664 468720 3670
rect 468668 3606 468720 3612
rect 468680 480 468708 3606
rect 469876 480 469904 7890
rect 471072 480 471100 12378
rect 473360 12368 473412 12374
rect 473360 12310 473412 12316
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 472268 480 472296 3538
rect 473372 3534 473400 12310
rect 478144 12300 478196 12306
rect 478144 12242 478196 12248
rect 473452 7880 473504 7886
rect 473452 7822 473504 7828
rect 473360 3528 473412 3534
rect 473360 3470 473412 3476
rect 473464 480 473492 7822
rect 476948 7812 477000 7818
rect 476948 7754 477000 7760
rect 474556 3528 474608 3534
rect 474556 3470 474608 3476
rect 474568 480 474596 3470
rect 475752 3460 475804 3466
rect 475752 3402 475804 3408
rect 475764 480 475792 3402
rect 476960 480 476988 7754
rect 478156 480 478184 12242
rect 479536 5574 479564 335990
rect 489920 334756 489972 334762
rect 489920 334698 489972 334704
rect 484400 327820 484452 327826
rect 484400 327762 484452 327768
rect 481640 326392 481692 326398
rect 481640 326334 481692 326340
rect 479524 5568 479576 5574
rect 479524 5510 479576 5516
rect 480536 5568 480588 5574
rect 480536 5510 480588 5516
rect 479340 3392 479392 3398
rect 479340 3334 479392 3340
rect 479352 480 479380 3334
rect 480548 480 480576 5510
rect 481652 3482 481680 326334
rect 481732 305652 481784 305658
rect 481732 305594 481784 305600
rect 481744 16574 481772 305594
rect 483020 181484 483072 181490
rect 483020 181426 483072 181432
rect 483032 16574 483060 181426
rect 484412 16574 484440 327762
rect 488540 319456 488592 319462
rect 488540 319398 488592 319404
rect 485780 304292 485832 304298
rect 485780 304234 485832 304240
rect 485792 16574 485820 304234
rect 488552 16574 488580 319398
rect 481744 16546 482876 16574
rect 483032 16546 484072 16574
rect 484412 16546 485268 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 481652 3454 481772 3482
rect 481744 480 481772 3454
rect 482848 480 482876 16546
rect 484044 480 484072 16546
rect 485240 480 485268 16546
rect 486436 480 486464 16546
rect 487620 14476 487672 14482
rect 487620 14418 487672 14424
rect 487632 480 487660 14418
rect 488828 480 488856 16546
rect 489932 3534 489960 334698
rect 525064 334688 525116 334694
rect 525064 334630 525116 334636
rect 500960 333260 501012 333266
rect 500960 333202 501012 333208
rect 491300 318096 491352 318102
rect 491300 318038 491352 318044
rect 490012 302932 490064 302938
rect 490012 302874 490064 302880
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 1442 490052 302874
rect 491312 16574 491340 318038
rect 498200 17264 498252 17270
rect 498200 17206 498252 17212
rect 491312 16546 492352 16574
rect 491116 3528 491168 3534
rect 491116 3470 491168 3476
rect 489932 1414 490052 1442
rect 489932 480 489960 1414
rect 491128 480 491156 3470
rect 492324 480 492352 16546
rect 494704 15904 494756 15910
rect 494704 15846 494756 15852
rect 493508 12232 493560 12238
rect 493508 12174 493560 12180
rect 493520 480 493548 12174
rect 494716 480 494744 15846
rect 497096 12164 497148 12170
rect 497096 12106 497148 12112
rect 495900 7744 495952 7750
rect 495900 7686 495952 7692
rect 495912 480 495940 7686
rect 497108 480 497136 12106
rect 498212 480 498240 17206
rect 500972 16574 501000 333202
rect 507860 331900 507912 331906
rect 507860 331842 507912 331848
rect 506480 323604 506532 323610
rect 506480 323546 506532 323552
rect 505100 18624 505152 18630
rect 505100 18566 505152 18572
rect 505112 16574 505140 18566
rect 500972 16546 501828 16574
rect 505112 16546 505416 16574
rect 500592 12096 500644 12102
rect 500592 12038 500644 12044
rect 499396 7676 499448 7682
rect 499396 7618 499448 7624
rect 499408 480 499436 7618
rect 500604 480 500632 12038
rect 501800 480 501828 16546
rect 504180 12028 504232 12034
rect 504180 11970 504232 11976
rect 502984 7608 503036 7614
rect 502984 7550 503036 7556
rect 502996 480 503024 7550
rect 504192 480 504220 11970
rect 505388 480 505416 16546
rect 506492 480 506520 323546
rect 507872 16574 507900 331842
rect 514760 330608 514812 330614
rect 514760 330550 514812 330556
rect 509240 316736 509292 316742
rect 509240 316678 509292 316684
rect 509252 16574 509280 316678
rect 513380 315308 513432 315314
rect 513380 315250 513432 315256
rect 513392 16574 513420 315250
rect 507872 16546 508912 16574
rect 509252 16546 510108 16574
rect 513392 16546 513604 16574
rect 507676 11960 507728 11966
rect 507676 11902 507728 11908
rect 507688 480 507716 11902
rect 508884 480 508912 16546
rect 510080 480 510108 16546
rect 511264 11892 511316 11898
rect 511264 11834 511316 11840
rect 511276 480 511304 11834
rect 512460 4548 512512 4554
rect 512460 4490 512512 4496
rect 512472 480 512500 4490
rect 513576 480 513604 16546
rect 514772 3466 514800 330550
rect 518900 329180 518952 329186
rect 518900 329122 518952 329128
rect 516140 324964 516192 324970
rect 516140 324906 516192 324912
rect 516152 16574 516180 324906
rect 517520 301504 517572 301510
rect 517520 301446 517572 301452
rect 517532 16574 517560 301446
rect 518912 16574 518940 329122
rect 520280 322244 520332 322250
rect 520280 322186 520332 322192
rect 520292 16574 520320 322186
rect 522304 314016 522356 314022
rect 522304 313958 522356 313964
rect 521660 300144 521712 300150
rect 521660 300086 521712 300092
rect 521672 16574 521700 300086
rect 516152 16546 517192 16574
rect 517532 16546 518388 16574
rect 518912 16546 519584 16574
rect 520292 16546 520780 16574
rect 521672 16546 521884 16574
rect 514852 11824 514904 11830
rect 514852 11766 514904 11772
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514864 1442 514892 11766
rect 515956 3460 516008 3466
rect 515956 3402 516008 3408
rect 514772 1414 514892 1442
rect 514772 480 514800 1414
rect 515968 480 515996 3402
rect 517164 480 517192 16546
rect 518360 480 518388 16546
rect 519556 480 519584 16546
rect 520752 480 520780 16546
rect 521856 480 521884 16546
rect 522316 3534 522344 313958
rect 524420 297424 524472 297430
rect 524420 297366 524472 297372
rect 523132 21412 523184 21418
rect 523132 21354 523184 21360
rect 523144 6914 523172 21354
rect 524432 16574 524460 297366
rect 524432 16546 525012 16574
rect 523052 6886 523172 6914
rect 522304 3528 522356 3534
rect 522304 3470 522356 3476
rect 523052 480 523080 6886
rect 524236 3528 524288 3534
rect 524236 3470 524288 3476
rect 524984 3482 525012 16546
rect 525076 3602 525104 334630
rect 525800 334620 525852 334626
rect 525800 334562 525852 334568
rect 525812 16574 525840 334562
rect 564440 330540 564492 330546
rect 564440 330482 564492 330488
rect 529204 329112 529256 329118
rect 529204 329054 529256 329060
rect 525812 16546 526668 16574
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 524248 480 524276 3470
rect 524984 3454 525472 3482
rect 525444 480 525472 3454
rect 526640 480 526668 16546
rect 529020 11756 529072 11762
rect 529020 11698 529072 11704
rect 527824 3596 527876 3602
rect 527824 3538 527876 3544
rect 527836 480 527864 3538
rect 529032 480 529060 11698
rect 529216 3058 529244 329054
rect 533344 320884 533396 320890
rect 533344 320826 533396 320832
rect 532516 13592 532568 13598
rect 532516 13534 532568 13540
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 529204 3052 529256 3058
rect 529204 2994 529256 3000
rect 530136 480 530164 4558
rect 531320 3052 531372 3058
rect 531320 2994 531372 3000
rect 531332 480 531360 2994
rect 532528 480 532556 13534
rect 533356 3534 533384 320826
rect 556160 295996 556212 296002
rect 556160 295938 556212 295944
rect 536104 13524 536156 13530
rect 536104 13466 536156 13472
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 533344 3528 533396 3534
rect 533344 3470 533396 3476
rect 533724 480 533752 4626
rect 534908 3528 534960 3534
rect 534908 3470 534960 3476
rect 534920 480 534948 3470
rect 536116 480 536144 13466
rect 539600 13456 539652 13462
rect 539600 13398 539652 13404
rect 538404 8900 538456 8906
rect 538404 8842 538456 8848
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 538416 480 538444 8842
rect 539612 480 539640 13398
rect 543188 13388 543240 13394
rect 543188 13330 543240 13336
rect 541992 9648 542044 9654
rect 541992 9590 542044 9596
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 540808 480 540836 5442
rect 542004 480 542032 9590
rect 543200 480 543228 13330
rect 546684 13320 546736 13326
rect 546684 13262 546736 13268
rect 545488 9580 545540 9586
rect 545488 9522 545540 9528
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 544396 480 544424 5374
rect 545500 480 545528 9522
rect 546696 480 546724 13262
rect 550272 13252 550324 13258
rect 550272 13194 550324 13200
rect 549076 9512 549128 9518
rect 549076 9454 549128 9460
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 547892 480 547920 5306
rect 549088 480 549116 9454
rect 550284 480 550312 13194
rect 553768 13184 553820 13190
rect 553768 13126 553820 13132
rect 552664 9444 552716 9450
rect 552664 9386 552716 9392
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 551480 480 551508 5238
rect 552676 480 552704 9386
rect 553780 480 553808 13126
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 554976 480 555004 5170
rect 556172 3534 556200 295938
rect 560852 13116 560904 13122
rect 560852 13058 560904 13064
rect 556252 9376 556304 9382
rect 556252 9318 556304 9324
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 1442 556292 9318
rect 559748 9308 559800 9314
rect 559748 9250 559800 9256
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3528 557408 3534
rect 557356 3470 557408 3476
rect 556172 1414 556292 1442
rect 556172 480 556200 1414
rect 557368 480 557396 3470
rect 558564 480 558592 5102
rect 559760 480 559788 9250
rect 560864 480 560892 13058
rect 563244 9240 563296 9246
rect 563244 9182 563296 9188
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 562060 480 562088 5034
rect 563256 480 563284 9182
rect 564452 480 564480 330482
rect 566464 327752 566516 327758
rect 566464 327694 566516 327700
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 565648 480 565676 4966
rect 566476 4146 566504 327694
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 576124 313948 576176 313954
rect 576124 313890 576176 313896
rect 571340 311160 571392 311166
rect 571340 311102 571392 311108
rect 571352 16574 571380 311102
rect 574100 294636 574152 294642
rect 574100 294578 574152 294584
rect 574112 16574 574140 294578
rect 571352 16546 571564 16574
rect 574112 16546 575152 16574
rect 566832 9172 566884 9178
rect 566832 9114 566884 9120
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 566844 480 566872 9114
rect 570328 9104 570380 9110
rect 570328 9046 570380 9052
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 568040 480 568068 4082
rect 569144 480 569172 4898
rect 570340 480 570368 9046
rect 571536 480 571564 16546
rect 573916 9036 573968 9042
rect 573916 8978 573968 8984
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 572732 480 572760 4830
rect 573928 480 573956 8978
rect 575124 480 575152 16546
rect 576136 3942 576164 313890
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 285660 580224 285666
rect 580172 285602 580224 285608
rect 580184 285433 580212 285602
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576124 3936 576176 3942
rect 576124 3878 576176 3884
rect 576320 480 576348 4762
rect 577424 480 577452 8910
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 578608 3936 578660 3942
rect 578608 3878 578660 3884
rect 578620 480 578648 3878
rect 579802 3768 579858 3777
rect 579802 3703 579858 3712
rect 579816 480 579844 3703
rect 580998 3632 581054 3641
rect 580998 3567 581054 3576
rect 581012 480 581040 3567
rect 582194 3496 582250 3505
rect 582194 3431 582250 3440
rect 582208 480 582236 3431
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3422 671200 3478 671256
rect 3330 645088 3386 645144
rect 2778 619132 2834 619168
rect 2778 619112 2780 619132
rect 2780 619112 2832 619132
rect 2832 619112 2834 619132
rect 2962 593000 3018 593056
rect 2870 540776 2926 540832
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3330 501744 3386 501800
rect 3238 488688 3294 488744
rect 3146 475632 3202 475688
rect 3054 462576 3110 462632
rect 2962 449520 3018 449576
rect 2870 436600 2926 436656
rect 2778 423544 2834 423600
rect 3514 658144 3570 658200
rect 3606 632032 3662 632088
rect 3422 410508 3478 410544
rect 3422 410488 3424 410508
rect 3424 410488 3476 410508
rect 3476 410488 3478 410508
rect 3698 606056 3754 606112
rect 3790 579944 3846 580000
rect 3422 397432 3478 397488
rect 3882 566888 3938 566944
rect 3974 553832 4030 553888
rect 4066 527856 4122 527912
rect 3514 384376 3570 384432
rect 580170 697176 580226 697232
rect 232042 407224 232098 407280
rect 232042 404640 232098 404696
rect 232042 403280 232098 403336
rect 232042 402056 232098 402112
rect 232042 400696 232098 400752
rect 232042 399472 232098 399528
rect 232042 398112 232098 398168
rect 232042 396888 232098 396944
rect 232042 395528 232098 395584
rect 231950 394304 232006 394360
rect 232042 392944 232098 393000
rect 232042 391720 232098 391776
rect 232042 390360 232098 390416
rect 232042 389036 232044 389056
rect 232044 389036 232096 389056
rect 232096 389036 232098 389056
rect 232042 389000 232098 389036
rect 231950 387776 232006 387832
rect 232042 386416 232098 386472
rect 232042 385192 232098 385248
rect 232042 383832 232098 383888
rect 231858 382608 231914 382664
rect 232042 381248 232098 381304
rect 580170 683848 580226 683904
rect 307022 407768 307078 407824
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 307114 406408 307170 406464
rect 580170 670656 580226 670692
rect 580262 657328 580318 657384
rect 580170 644000 580226 644056
rect 307206 405048 307262 405104
rect 306930 386144 306986 386200
rect 306838 384920 306894 384976
rect 306746 380840 306802 380896
rect 232042 380024 232098 380080
rect 306838 380024 306894 380080
rect 307206 403824 307262 403880
rect 579986 630808 580042 630864
rect 307298 402464 307354 402520
rect 307298 401104 307354 401160
rect 307206 399608 307262 399664
rect 307482 398384 307538 398440
rect 307390 397160 307446 397216
rect 307298 395664 307354 395720
rect 307482 394304 307538 394360
rect 307482 392944 307538 393000
rect 307574 391856 307630 391912
rect 580170 590960 580226 591016
rect 579986 577632 580042 577688
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 444760 580226 444816
rect 580078 431568 580134 431624
rect 580078 418240 580134 418296
rect 232042 378664 232098 378720
rect 307022 378664 307078 378720
rect 232042 377440 232098 377496
rect 307666 390496 307722 390552
rect 307666 388864 307722 388920
rect 307666 387504 307722 387560
rect 307666 383596 307668 383616
rect 307668 383596 307720 383616
rect 307720 383596 307722 383616
rect 307666 383560 307722 383596
rect 307666 382220 307722 382256
rect 307666 382200 307668 382220
rect 307668 382200 307720 382220
rect 307720 382200 307722 382220
rect 580078 404912 580134 404968
rect 580078 391720 580134 391776
rect 580354 617480 580410 617536
rect 580446 604152 580502 604208
rect 580538 564304 580594 564360
rect 580630 551112 580686 551168
rect 580722 511264 580778 511320
rect 580814 497936 580870 497992
rect 580906 458088 580962 458144
rect 580170 378392 580226 378448
rect 307114 377304 307170 377360
rect 232042 376080 232098 376136
rect 307666 376080 307722 376136
rect 232042 374856 232098 374912
rect 307114 374040 307170 374096
rect 232042 373496 232098 373552
rect 307022 372680 307078 372736
rect 3514 371320 3570 371376
rect 3054 332288 3110 332344
rect 3054 319232 3110 319288
rect 3146 306176 3202 306232
rect 3146 293156 3148 293176
rect 3148 293156 3200 293176
rect 3200 293156 3202 293176
rect 3146 293120 3202 293156
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3238 227976 3294 228032
rect 3238 214920 3294 214976
rect 232042 372136 232098 372192
rect 233146 370912 233202 370968
rect 233054 369552 233110 369608
rect 232042 368328 232098 368384
rect 232042 366968 232098 367024
rect 232778 365744 232834 365800
rect 3606 358400 3662 358456
rect 3422 345344 3478 345400
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3330 175888 3386 175944
rect 3330 149776 3386 149832
rect 3146 123664 3202 123720
rect 3146 84632 3202 84688
rect 2870 58520 2926 58576
rect 232686 364384 232742 364440
rect 232042 363160 232098 363216
rect 4066 162832 4122 162888
rect 3974 136720 4030 136776
rect 3882 110608 3938 110664
rect 3790 97552 3846 97608
rect 3698 71576 3754 71632
rect 3606 45464 3662 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 6458 3304 6514 3360
rect 15934 3576 15990 3632
rect 14738 3440 14794 3496
rect 20626 3712 20682 3768
rect 232042 361800 232098 361856
rect 232594 360576 232650 360632
rect 232686 359216 232742 359272
rect 232042 357992 232098 358048
rect 232042 356632 232098 356688
rect 232594 355272 232650 355328
rect 232042 354048 232098 354104
rect 232042 352688 232098 352744
rect 232042 351464 232098 351520
rect 232502 350104 232558 350160
rect 232042 348880 232098 348936
rect 232042 347520 232098 347576
rect 232042 346296 232098 346352
rect 231858 344936 231914 344992
rect 232042 343732 232098 343768
rect 232042 343712 232044 343732
rect 232044 343712 232096 343732
rect 232096 343712 232098 343732
rect 232042 342352 232098 342408
rect 232042 341128 232098 341184
rect 232042 339768 232098 339824
rect 232042 338544 232098 338600
rect 306378 369824 306434 369880
rect 306286 342352 306342 342408
rect 235262 3304 235318 3360
rect 236734 3576 236790 3632
rect 236458 3440 236514 3496
rect 238206 3712 238262 3768
rect 240598 326304 240654 326360
rect 240782 326032 240838 326088
rect 304630 3440 304686 3496
rect 304906 3712 304962 3768
rect 304814 3576 304870 3632
rect 304722 3304 304778 3360
rect 306470 368464 306526 368520
rect 306562 367240 306618 367296
rect 307666 371320 307722 371376
rect 307666 366016 307722 366072
rect 307666 364656 307722 364712
rect 306654 361664 306710 361720
rect 306746 360440 306802 360496
rect 306838 359080 306894 359136
rect 306930 357856 306986 357912
rect 307298 363296 307354 363352
rect 307666 356496 307722 356552
rect 307666 355136 307722 355192
rect 307666 353776 307722 353832
rect 307574 352416 307630 352472
rect 307482 351192 307538 351248
rect 307390 349832 307446 349888
rect 307298 348472 307354 348528
rect 307022 346568 307078 346624
rect 307206 345208 307262 345264
rect 307206 343848 307262 343904
rect 307206 339632 307262 339688
rect 307206 338272 307262 338328
rect 307666 347928 307722 347984
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 338544 580226 338600
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 285368 580226 285424
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 579802 3712 579858 3768
rect 580998 3576 581054 3632
rect 582194 3440 582250 3496
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3366 684314 3372 684316
rect -960 684254 3372 684314
rect -960 684164 480 684254
rect 3366 684252 3372 684254
rect 3436 684252 3442 684316
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 580257 657386 580323 657389
rect 583520 657386 584960 657476
rect 580257 657384 584960 657386
rect 580257 657328 580262 657384
rect 580318 657328 584960 657384
rect 580257 657326 584960 657328
rect 580257 657323 580323 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 3325 645146 3391 645149
rect -960 645144 3391 645146
rect -960 645088 3330 645144
rect 3386 645088 3391 645144
rect -960 645086 3391 645088
rect -960 644996 480 645086
rect 3325 645083 3391 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 580349 617538 580415 617541
rect 583520 617538 584960 617628
rect 580349 617536 584960 617538
rect 580349 617480 580354 617536
rect 580410 617480 584960 617536
rect 580349 617478 584960 617480
rect 580349 617475 580415 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3693 606114 3759 606117
rect -960 606112 3759 606114
rect -960 606056 3698 606112
rect 3754 606056 3759 606112
rect -960 606054 3759 606056
rect -960 605964 480 606054
rect 3693 606051 3759 606054
rect 580441 604210 580507 604213
rect 583520 604210 584960 604300
rect 580441 604208 584960 604210
rect 580441 604152 580446 604208
rect 580502 604152 584960 604208
rect 580441 604150 584960 604152
rect 580441 604147 580507 604150
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 2957 593058 3023 593061
rect -960 593056 3023 593058
rect -960 593000 2962 593056
rect 3018 593000 3023 593056
rect -960 592998 3023 593000
rect -960 592908 480 592998
rect 2957 592995 3023 592998
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3785 580002 3851 580005
rect -960 580000 3851 580002
rect -960 579944 3790 580000
rect 3846 579944 3851 580000
rect -960 579942 3851 579944
rect -960 579852 480 579942
rect 3785 579939 3851 579942
rect 579981 577690 580047 577693
rect 583520 577690 584960 577780
rect 579981 577688 584960 577690
rect 579981 577632 579986 577688
rect 580042 577632 584960 577688
rect 579981 577630 584960 577632
rect 579981 577627 580047 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3877 566946 3943 566949
rect -960 566944 3943 566946
rect -960 566888 3882 566944
rect 3938 566888 3943 566944
rect -960 566886 3943 566888
rect -960 566796 480 566886
rect 3877 566883 3943 566886
rect 580533 564362 580599 564365
rect 583520 564362 584960 564452
rect 580533 564360 584960 564362
rect 580533 564304 580538 564360
rect 580594 564304 584960 564360
rect 580533 564302 584960 564304
rect 580533 564299 580599 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3969 553890 4035 553893
rect -960 553888 4035 553890
rect -960 553832 3974 553888
rect 4030 553832 4035 553888
rect -960 553830 4035 553832
rect -960 553740 480 553830
rect 3969 553827 4035 553830
rect 580625 551170 580691 551173
rect 583520 551170 584960 551260
rect 580625 551168 584960 551170
rect 580625 551112 580630 551168
rect 580686 551112 584960 551168
rect 580625 551110 584960 551112
rect 580625 551107 580691 551110
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 2865 540834 2931 540837
rect -960 540832 2931 540834
rect -960 540776 2870 540832
rect 2926 540776 2931 540832
rect -960 540774 2931 540776
rect -960 540684 480 540774
rect 2865 540771 2931 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 4061 527914 4127 527917
rect -960 527912 4127 527914
rect -960 527856 4066 527912
rect 4122 527856 4127 527912
rect -960 527854 4127 527856
rect -960 527764 480 527854
rect 4061 527851 4127 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580717 511322 580783 511325
rect 583520 511322 584960 511412
rect 580717 511320 584960 511322
rect 580717 511264 580722 511320
rect 580778 511264 584960 511320
rect 580717 511262 584960 511264
rect 580717 511259 580783 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 580809 497994 580875 497997
rect 583520 497994 584960 498084
rect 580809 497992 584960 497994
rect 580809 497936 580814 497992
rect 580870 497936 584960 497992
rect 580809 497934 584960 497936
rect 580809 497931 580875 497934
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect 3233 488746 3299 488749
rect -960 488744 3299 488746
rect -960 488688 3238 488744
rect 3294 488688 3299 488744
rect -960 488686 3299 488688
rect -960 488596 480 488686
rect 3233 488683 3299 488686
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3141 475690 3207 475693
rect -960 475688 3207 475690
rect -960 475632 3146 475688
rect 3202 475632 3207 475688
rect -960 475630 3207 475632
rect -960 475540 480 475630
rect 3141 475627 3207 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580901 458146 580967 458149
rect 583520 458146 584960 458236
rect 580901 458144 584960 458146
rect 580901 458088 580906 458144
rect 580962 458088 584960 458144
rect 580901 458086 584960 458088
rect 580901 458083 580967 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2957 449578 3023 449581
rect -960 449576 3023 449578
rect -960 449520 2962 449576
rect 3018 449520 3023 449576
rect -960 449518 3023 449520
rect -960 449428 480 449518
rect 2957 449515 3023 449518
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect -960 436658 480 436748
rect 2865 436658 2931 436661
rect -960 436656 2931 436658
rect -960 436600 2870 436656
rect 2926 436600 2931 436656
rect -960 436598 2931 436600
rect -960 436508 480 436598
rect 2865 436595 2931 436598
rect 580073 431626 580139 431629
rect 583520 431626 584960 431716
rect 580073 431624 584960 431626
rect 580073 431568 580078 431624
rect 580134 431568 584960 431624
rect 580073 431566 584960 431568
rect 580073 431563 580139 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 580073 418298 580139 418301
rect 583520 418298 584960 418388
rect 580073 418296 584960 418298
rect 580073 418240 580078 418296
rect 580134 418240 584960 418296
rect 580073 418238 584960 418240
rect 580073 418235 580139 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 307017 407826 307083 407829
rect 304950 407824 307083 407826
rect 304950 407768 307022 407824
rect 307078 407768 307083 407824
rect 304950 407766 307083 407768
rect 232037 407282 232103 407285
rect 232037 407280 235060 407282
rect 232037 407224 232042 407280
rect 232098 407224 235060 407280
rect 304950 407252 305010 407766
rect 307017 407763 307083 407766
rect 232037 407222 235060 407224
rect 232037 407219 232103 407222
rect 307109 406466 307175 406469
rect 304950 406464 307175 406466
rect 304950 406408 307114 406464
rect 307170 406408 307175 406464
rect 304950 406406 307175 406408
rect 304950 405892 305010 406406
rect 307109 406403 307175 406406
rect 3366 405724 3372 405788
rect 3436 405786 3442 405788
rect 235030 405786 235090 405892
rect 3436 405726 235090 405786
rect 3436 405724 3442 405726
rect 307201 405106 307267 405109
rect 304950 405104 307267 405106
rect 304950 405048 307206 405104
rect 307262 405048 307267 405104
rect 304950 405046 307267 405048
rect 232037 404698 232103 404701
rect 232037 404696 235060 404698
rect 232037 404640 232042 404696
rect 232098 404640 235060 404696
rect 232037 404638 235060 404640
rect 232037 404635 232103 404638
rect 304950 404532 305010 405046
rect 307201 405043 307267 405046
rect 580073 404970 580139 404973
rect 583520 404970 584960 405060
rect 580073 404968 584960 404970
rect 580073 404912 580078 404968
rect 580134 404912 584960 404968
rect 580073 404910 584960 404912
rect 580073 404907 580139 404910
rect 583520 404820 584960 404910
rect 307201 403882 307267 403885
rect 304950 403880 307267 403882
rect 304950 403824 307206 403880
rect 307262 403824 307267 403880
rect 304950 403822 307267 403824
rect 232037 403338 232103 403341
rect 232037 403336 235060 403338
rect 232037 403280 232042 403336
rect 232098 403280 235060 403336
rect 304950 403308 305010 403822
rect 307201 403819 307267 403822
rect 232037 403278 235060 403280
rect 232037 403275 232103 403278
rect 307293 402522 307359 402525
rect 304950 402520 307359 402522
rect 304950 402464 307298 402520
rect 307354 402464 307359 402520
rect 304950 402462 307359 402464
rect 232037 402114 232103 402117
rect 232037 402112 235060 402114
rect 232037 402056 232042 402112
rect 232098 402056 235060 402112
rect 232037 402054 235060 402056
rect 232037 402051 232103 402054
rect 304950 401948 305010 402462
rect 307293 402459 307359 402462
rect 307293 401162 307359 401165
rect 304950 401160 307359 401162
rect 304950 401104 307298 401160
rect 307354 401104 307359 401160
rect 304950 401102 307359 401104
rect 232037 400754 232103 400757
rect 232037 400752 235060 400754
rect 232037 400696 232042 400752
rect 232098 400696 235060 400752
rect 232037 400694 235060 400696
rect 232037 400691 232103 400694
rect 304950 400588 305010 401102
rect 307293 401099 307359 401102
rect 307201 399666 307267 399669
rect 304950 399664 307267 399666
rect 304950 399608 307206 399664
rect 307262 399608 307267 399664
rect 304950 399606 307267 399608
rect 232037 399530 232103 399533
rect 232037 399528 235060 399530
rect 232037 399472 232042 399528
rect 232098 399472 235060 399528
rect 232037 399470 235060 399472
rect 232037 399467 232103 399470
rect 304950 399228 305010 399606
rect 307201 399603 307267 399606
rect 307477 398442 307543 398445
rect 304950 398440 307543 398442
rect 304950 398384 307482 398440
rect 307538 398384 307543 398440
rect 304950 398382 307543 398384
rect 232037 398170 232103 398173
rect 232037 398168 235060 398170
rect 232037 398112 232042 398168
rect 232098 398112 235060 398168
rect 232037 398110 235060 398112
rect 232037 398107 232103 398110
rect 304950 398004 305010 398382
rect 307477 398379 307543 398382
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 307385 397218 307451 397221
rect 304950 397216 307451 397218
rect 304950 397160 307390 397216
rect 307446 397160 307451 397216
rect 304950 397158 307451 397160
rect 232037 396946 232103 396949
rect 232037 396944 235060 396946
rect 232037 396888 232042 396944
rect 232098 396888 235060 396944
rect 232037 396886 235060 396888
rect 232037 396883 232103 396886
rect 304950 396644 305010 397158
rect 307385 397155 307451 397158
rect 307293 395722 307359 395725
rect 304950 395720 307359 395722
rect 304950 395664 307298 395720
rect 307354 395664 307359 395720
rect 304950 395662 307359 395664
rect 232037 395586 232103 395589
rect 232037 395584 235060 395586
rect 232037 395528 232042 395584
rect 232098 395528 235060 395584
rect 232037 395526 235060 395528
rect 232037 395523 232103 395526
rect 304950 395284 305010 395662
rect 307293 395659 307359 395662
rect 231945 394362 232011 394365
rect 307477 394362 307543 394365
rect 231945 394360 235060 394362
rect 231945 394304 231950 394360
rect 232006 394304 235060 394360
rect 231945 394302 235060 394304
rect 304950 394360 307543 394362
rect 304950 394304 307482 394360
rect 307538 394304 307543 394360
rect 304950 394302 307543 394304
rect 231945 394299 232011 394302
rect 304950 394060 305010 394302
rect 307477 394299 307543 394302
rect 232037 393002 232103 393005
rect 307477 393002 307543 393005
rect 232037 393000 235060 393002
rect 232037 392944 232042 393000
rect 232098 392944 235060 393000
rect 232037 392942 235060 392944
rect 304950 393000 307543 393002
rect 304950 392944 307482 393000
rect 307538 392944 307543 393000
rect 304950 392942 307543 392944
rect 232037 392939 232103 392942
rect 304950 392700 305010 392942
rect 307477 392939 307543 392942
rect 307569 391914 307635 391917
rect 304950 391912 307635 391914
rect 304950 391856 307574 391912
rect 307630 391856 307635 391912
rect 304950 391854 307635 391856
rect 232037 391778 232103 391781
rect 232037 391776 235060 391778
rect 232037 391720 232042 391776
rect 232098 391720 235060 391776
rect 232037 391718 235060 391720
rect 232037 391715 232103 391718
rect 304950 391340 305010 391854
rect 307569 391851 307635 391854
rect 580073 391778 580139 391781
rect 583520 391778 584960 391868
rect 580073 391776 584960 391778
rect 580073 391720 580078 391776
rect 580134 391720 584960 391776
rect 580073 391718 584960 391720
rect 580073 391715 580139 391718
rect 583520 391628 584960 391718
rect 307661 390554 307727 390557
rect 304950 390552 307727 390554
rect 304950 390496 307666 390552
rect 307722 390496 307727 390552
rect 304950 390494 307727 390496
rect 232037 390418 232103 390421
rect 232037 390416 235060 390418
rect 232037 390360 232042 390416
rect 232098 390360 235060 390416
rect 232037 390358 235060 390360
rect 232037 390355 232103 390358
rect 304950 389980 305010 390494
rect 307661 390491 307727 390494
rect 232037 389058 232103 389061
rect 232037 389056 235060 389058
rect 232037 389000 232042 389056
rect 232098 389000 235060 389056
rect 232037 388998 235060 389000
rect 232037 388995 232103 388998
rect 307661 388922 307727 388925
rect 304950 388920 307727 388922
rect 304950 388864 307666 388920
rect 307722 388864 307727 388920
rect 304950 388862 307727 388864
rect 304950 388756 305010 388862
rect 307661 388859 307727 388862
rect 231945 387834 232011 387837
rect 231945 387832 235060 387834
rect 231945 387776 231950 387832
rect 232006 387776 235060 387832
rect 231945 387774 235060 387776
rect 231945 387771 232011 387774
rect 307661 387562 307727 387565
rect 304950 387560 307727 387562
rect 304950 387504 307666 387560
rect 307722 387504 307727 387560
rect 304950 387502 307727 387504
rect 304950 387396 305010 387502
rect 307661 387499 307727 387502
rect 232037 386474 232103 386477
rect 232037 386472 235060 386474
rect 232037 386416 232042 386472
rect 232098 386416 235060 386472
rect 232037 386414 235060 386416
rect 232037 386411 232103 386414
rect 306925 386202 306991 386205
rect 304950 386200 306991 386202
rect 304950 386144 306930 386200
rect 306986 386144 306991 386200
rect 304950 386142 306991 386144
rect 304950 386036 305010 386142
rect 306925 386139 306991 386142
rect 232037 385250 232103 385253
rect 232037 385248 235060 385250
rect 232037 385192 232042 385248
rect 232098 385192 235060 385248
rect 232037 385190 235060 385192
rect 232037 385187 232103 385190
rect 306833 384978 306899 384981
rect 304950 384976 306899 384978
rect 304950 384920 306838 384976
rect 306894 384920 306899 384976
rect 304950 384918 306899 384920
rect 304950 384812 305010 384918
rect 306833 384915 306899 384918
rect -960 384434 480 384524
rect 3509 384434 3575 384437
rect -960 384432 3575 384434
rect -960 384376 3514 384432
rect 3570 384376 3575 384432
rect -960 384374 3575 384376
rect -960 384284 480 384374
rect 3509 384371 3575 384374
rect 232037 383890 232103 383893
rect 232037 383888 235060 383890
rect 232037 383832 232042 383888
rect 232098 383832 235060 383888
rect 232037 383830 235060 383832
rect 232037 383827 232103 383830
rect 307661 383618 307727 383621
rect 304950 383616 307727 383618
rect 304950 383560 307666 383616
rect 307722 383560 307727 383616
rect 304950 383558 307727 383560
rect 304950 383452 305010 383558
rect 307661 383555 307727 383558
rect 231853 382666 231919 382669
rect 231853 382664 235060 382666
rect 231853 382608 231858 382664
rect 231914 382608 235060 382664
rect 231853 382606 235060 382608
rect 231853 382603 231919 382606
rect 307661 382258 307727 382261
rect 304950 382256 307727 382258
rect 304950 382200 307666 382256
rect 307722 382200 307727 382256
rect 304950 382198 307727 382200
rect 304950 382092 305010 382198
rect 307661 382195 307727 382198
rect 232037 381306 232103 381309
rect 232037 381304 235060 381306
rect 232037 381248 232042 381304
rect 232098 381248 235060 381304
rect 232037 381246 235060 381248
rect 232037 381243 232103 381246
rect 306741 380898 306807 380901
rect 304950 380896 306807 380898
rect 304950 380840 306746 380896
rect 306802 380840 306807 380896
rect 304950 380838 306807 380840
rect 304950 380732 305010 380838
rect 306741 380835 306807 380838
rect 232037 380082 232103 380085
rect 306833 380082 306899 380085
rect 232037 380080 235060 380082
rect 232037 380024 232042 380080
rect 232098 380024 235060 380080
rect 232037 380022 235060 380024
rect 304950 380080 306899 380082
rect 304950 380024 306838 380080
rect 306894 380024 306899 380080
rect 304950 380022 306899 380024
rect 232037 380019 232103 380022
rect 304950 379508 305010 380022
rect 306833 380019 306899 380022
rect 232037 378722 232103 378725
rect 307017 378722 307083 378725
rect 232037 378720 235060 378722
rect 232037 378664 232042 378720
rect 232098 378664 235060 378720
rect 232037 378662 235060 378664
rect 304950 378720 307083 378722
rect 304950 378664 307022 378720
rect 307078 378664 307083 378720
rect 304950 378662 307083 378664
rect 232037 378659 232103 378662
rect 304950 378148 305010 378662
rect 307017 378659 307083 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 232037 377498 232103 377501
rect 232037 377496 235060 377498
rect 232037 377440 232042 377496
rect 232098 377440 235060 377496
rect 232037 377438 235060 377440
rect 232037 377435 232103 377438
rect 307109 377362 307175 377365
rect 304950 377360 307175 377362
rect 304950 377304 307114 377360
rect 307170 377304 307175 377360
rect 304950 377302 307175 377304
rect 304950 376788 305010 377302
rect 307109 377299 307175 377302
rect 232037 376138 232103 376141
rect 307661 376138 307727 376141
rect 232037 376136 235060 376138
rect 232037 376080 232042 376136
rect 232098 376080 235060 376136
rect 232037 376078 235060 376080
rect 304950 376136 307727 376138
rect 304950 376080 307666 376136
rect 307722 376080 307727 376136
rect 304950 376078 307727 376080
rect 232037 376075 232103 376078
rect 304950 375564 305010 376078
rect 307661 376075 307727 376078
rect 232037 374914 232103 374917
rect 232037 374912 235060 374914
rect 232037 374856 232042 374912
rect 232098 374856 235060 374912
rect 232037 374854 235060 374856
rect 232037 374851 232103 374854
rect 304766 374098 304826 374204
rect 307109 374098 307175 374101
rect 304766 374096 307175 374098
rect 304766 374040 307114 374096
rect 307170 374040 307175 374096
rect 304766 374038 307175 374040
rect 307109 374035 307175 374038
rect 232037 373554 232103 373557
rect 232037 373552 235060 373554
rect 232037 373496 232042 373552
rect 232098 373496 235060 373552
rect 232037 373494 235060 373496
rect 232037 373491 232103 373494
rect 304766 372738 304826 372844
rect 307017 372738 307083 372741
rect 304766 372736 307083 372738
rect 304766 372680 307022 372736
rect 307078 372680 307083 372736
rect 304766 372678 307083 372680
rect 307017 372675 307083 372678
rect 232037 372194 232103 372197
rect 232037 372192 235060 372194
rect 232037 372136 232042 372192
rect 232098 372136 235060 372192
rect 232037 372134 235060 372136
rect 232037 372131 232103 372134
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect 304766 371378 304826 371484
rect 307661 371378 307727 371381
rect 304766 371376 307727 371378
rect 304766 371320 307666 371376
rect 307722 371320 307727 371376
rect 304766 371318 307727 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 307661 371315 307727 371318
rect 233141 370970 233207 370973
rect 233141 370968 235060 370970
rect 233141 370912 233146 370968
rect 233202 370912 235060 370968
rect 233141 370910 235060 370912
rect 233141 370907 233207 370910
rect 304766 369882 304826 370260
rect 306373 369882 306439 369885
rect 304766 369880 306439 369882
rect 304766 369824 306378 369880
rect 306434 369824 306439 369880
rect 304766 369822 306439 369824
rect 306373 369819 306439 369822
rect 233049 369610 233115 369613
rect 233049 369608 235060 369610
rect 233049 369552 233054 369608
rect 233110 369552 235060 369608
rect 233049 369550 235060 369552
rect 233049 369547 233115 369550
rect 304766 368522 304826 368900
rect 306465 368522 306531 368525
rect 304766 368520 306531 368522
rect 304766 368464 306470 368520
rect 306526 368464 306531 368520
rect 304766 368462 306531 368464
rect 306465 368459 306531 368462
rect 232037 368386 232103 368389
rect 232037 368384 235060 368386
rect 232037 368328 232042 368384
rect 232098 368328 235060 368384
rect 232037 368326 235060 368328
rect 232037 368323 232103 368326
rect 304766 367298 304826 367540
rect 306557 367298 306623 367301
rect 304766 367296 306623 367298
rect 304766 367240 306562 367296
rect 306618 367240 306623 367296
rect 304766 367238 306623 367240
rect 306557 367235 306623 367238
rect 232037 367026 232103 367029
rect 232037 367024 235060 367026
rect 232037 366968 232042 367024
rect 232098 366968 235060 367024
rect 232037 366966 235060 366968
rect 232037 366963 232103 366966
rect 304766 366074 304826 366316
rect 307661 366074 307727 366077
rect 304766 366072 307727 366074
rect 304766 366016 307666 366072
rect 307722 366016 307727 366072
rect 304766 366014 307727 366016
rect 307661 366011 307727 366014
rect 232773 365802 232839 365805
rect 232773 365800 235060 365802
rect 232773 365744 232778 365800
rect 232834 365744 235060 365800
rect 232773 365742 235060 365744
rect 232773 365739 232839 365742
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 304766 364714 304826 364956
rect 307661 364714 307727 364717
rect 304766 364712 307727 364714
rect 304766 364656 307666 364712
rect 307722 364656 307727 364712
rect 304766 364654 307727 364656
rect 307661 364651 307727 364654
rect 232681 364442 232747 364445
rect 232681 364440 235060 364442
rect 232681 364384 232686 364440
rect 232742 364384 235060 364440
rect 232681 364382 235060 364384
rect 232681 364379 232747 364382
rect 304766 363354 304826 363596
rect 307293 363354 307359 363357
rect 304766 363352 307359 363354
rect 304766 363296 307298 363352
rect 307354 363296 307359 363352
rect 304766 363294 307359 363296
rect 307293 363291 307359 363294
rect 232037 363218 232103 363221
rect 232037 363216 235060 363218
rect 232037 363160 232042 363216
rect 232098 363160 235060 363216
rect 232037 363158 235060 363160
rect 232037 363155 232103 363158
rect 232037 361858 232103 361861
rect 232037 361856 235060 361858
rect 232037 361800 232042 361856
rect 232098 361800 235060 361856
rect 232037 361798 235060 361800
rect 232037 361795 232103 361798
rect 304766 361722 304826 362236
rect 306649 361722 306715 361725
rect 304766 361720 306715 361722
rect 304766 361664 306654 361720
rect 306710 361664 306715 361720
rect 304766 361662 306715 361664
rect 306649 361659 306715 361662
rect 232589 360634 232655 360637
rect 232589 360632 235060 360634
rect 232589 360576 232594 360632
rect 232650 360576 235060 360632
rect 232589 360574 235060 360576
rect 232589 360571 232655 360574
rect 304766 360498 304826 361012
rect 306741 360498 306807 360501
rect 304766 360496 306807 360498
rect 304766 360440 306746 360496
rect 306802 360440 306807 360496
rect 304766 360438 306807 360440
rect 306741 360435 306807 360438
rect 232681 359274 232747 359277
rect 232681 359272 235060 359274
rect 232681 359216 232686 359272
rect 232742 359216 235060 359272
rect 232681 359214 235060 359216
rect 232681 359211 232747 359214
rect 304766 359138 304826 359652
rect 306833 359138 306899 359141
rect 304766 359136 306899 359138
rect 304766 359080 306838 359136
rect 306894 359080 306899 359136
rect 304766 359078 306899 359080
rect 306833 359075 306899 359078
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 232037 358050 232103 358053
rect 232037 358048 235060 358050
rect 232037 357992 232042 358048
rect 232098 357992 235060 358048
rect 232037 357990 235060 357992
rect 232037 357987 232103 357990
rect 304766 357914 304826 358292
rect 306925 357914 306991 357917
rect 304766 357912 306991 357914
rect 304766 357856 306930 357912
rect 306986 357856 306991 357912
rect 304766 357854 306991 357856
rect 306925 357851 306991 357854
rect 232037 356690 232103 356693
rect 232037 356688 235060 356690
rect 232037 356632 232042 356688
rect 232098 356632 235060 356688
rect 232037 356630 235060 356632
rect 232037 356627 232103 356630
rect 304766 356554 304826 357068
rect 307661 356554 307727 356557
rect 304766 356552 307727 356554
rect 304766 356496 307666 356552
rect 307722 356496 307727 356552
rect 304766 356494 307727 356496
rect 307661 356491 307727 356494
rect 232589 355330 232655 355333
rect 232589 355328 235060 355330
rect 232589 355272 232594 355328
rect 232650 355272 235060 355328
rect 232589 355270 235060 355272
rect 232589 355267 232655 355270
rect 304766 355194 304826 355708
rect 307661 355194 307727 355197
rect 304766 355192 307727 355194
rect 304766 355136 307666 355192
rect 307722 355136 307727 355192
rect 304766 355134 307727 355136
rect 307661 355131 307727 355134
rect 232037 354106 232103 354109
rect 232037 354104 235060 354106
rect 232037 354048 232042 354104
rect 232098 354048 235060 354104
rect 232037 354046 235060 354048
rect 232037 354043 232103 354046
rect 304766 353834 304826 354348
rect 307661 353834 307727 353837
rect 304766 353832 307727 353834
rect 304766 353776 307666 353832
rect 307722 353776 307727 353832
rect 304766 353774 307727 353776
rect 307661 353771 307727 353774
rect 232037 352746 232103 352749
rect 232037 352744 235060 352746
rect 232037 352688 232042 352744
rect 232098 352688 235060 352744
rect 232037 352686 235060 352688
rect 232037 352683 232103 352686
rect 304766 352474 304826 352988
rect 307569 352474 307635 352477
rect 304766 352472 307635 352474
rect 304766 352416 307574 352472
rect 307630 352416 307635 352472
rect 304766 352414 307635 352416
rect 307569 352411 307635 352414
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 232037 351522 232103 351525
rect 232037 351520 235060 351522
rect 232037 351464 232042 351520
rect 232098 351464 235060 351520
rect 232037 351462 235060 351464
rect 232037 351459 232103 351462
rect 304766 351250 304826 351764
rect 307477 351250 307543 351253
rect 304766 351248 307543 351250
rect 304766 351192 307482 351248
rect 307538 351192 307543 351248
rect 304766 351190 307543 351192
rect 307477 351187 307543 351190
rect 232497 350162 232563 350165
rect 232497 350160 235060 350162
rect 232497 350104 232502 350160
rect 232558 350104 235060 350160
rect 232497 350102 235060 350104
rect 232497 350099 232563 350102
rect 304766 349890 304826 350404
rect 307385 349890 307451 349893
rect 304766 349888 307451 349890
rect 304766 349832 307390 349888
rect 307446 349832 307451 349888
rect 304766 349830 307451 349832
rect 307385 349827 307451 349830
rect 232037 348938 232103 348941
rect 232037 348936 235060 348938
rect 232037 348880 232042 348936
rect 232098 348880 235060 348936
rect 232037 348878 235060 348880
rect 232037 348875 232103 348878
rect 304766 348530 304826 349044
rect 307293 348530 307359 348533
rect 304766 348528 307359 348530
rect 304766 348472 307298 348528
rect 307354 348472 307359 348528
rect 304766 348470 307359 348472
rect 307293 348467 307359 348470
rect 307661 347986 307727 347989
rect 304950 347984 307727 347986
rect 304950 347928 307666 347984
rect 307722 347928 307727 347984
rect 304950 347926 307727 347928
rect 304950 347820 305010 347926
rect 307661 347923 307727 347926
rect 232037 347578 232103 347581
rect 232037 347576 235060 347578
rect 232037 347520 232042 347576
rect 232098 347520 235060 347576
rect 232037 347518 235060 347520
rect 232037 347515 232103 347518
rect 307017 346626 307083 346629
rect 304950 346624 307083 346626
rect 304950 346568 307022 346624
rect 307078 346568 307083 346624
rect 304950 346566 307083 346568
rect 304950 346460 305010 346566
rect 307017 346563 307083 346566
rect 232037 346354 232103 346357
rect 232037 346352 235060 346354
rect 232037 346296 232042 346352
rect 232098 346296 235060 346352
rect 232037 346294 235060 346296
rect 232037 346291 232103 346294
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 307201 345266 307267 345269
rect 304950 345264 307267 345266
rect 304950 345208 307206 345264
rect 307262 345208 307267 345264
rect 304950 345206 307267 345208
rect 304950 345100 305010 345206
rect 307201 345203 307267 345206
rect 231853 344994 231919 344997
rect 231853 344992 235060 344994
rect 231853 344936 231858 344992
rect 231914 344936 235060 344992
rect 231853 344934 235060 344936
rect 231853 344931 231919 344934
rect 307201 343906 307267 343909
rect 304950 343904 307267 343906
rect 304950 343848 307206 343904
rect 307262 343848 307267 343904
rect 304950 343846 307267 343848
rect 232037 343770 232103 343773
rect 232037 343768 235060 343770
rect 232037 343712 232042 343768
rect 232098 343712 235060 343768
rect 304950 343740 305010 343846
rect 307201 343843 307267 343846
rect 232037 343710 235060 343712
rect 232037 343707 232103 343710
rect 232037 342410 232103 342413
rect 304766 342410 304826 342516
rect 306281 342410 306347 342413
rect 232037 342408 235060 342410
rect 232037 342352 232042 342408
rect 232098 342352 235060 342408
rect 232037 342350 235060 342352
rect 304766 342408 306347 342410
rect 304766 342352 306286 342408
rect 306342 342352 306347 342408
rect 304766 342350 306347 342352
rect 232037 342347 232103 342350
rect 306281 342347 306347 342350
rect 232037 341186 232103 341189
rect 232037 341184 235060 341186
rect 232037 341128 232042 341184
rect 232098 341128 235060 341184
rect 232037 341126 235060 341128
rect 232037 341123 232103 341126
rect 304766 340914 304826 341156
rect 306966 340914 306972 340916
rect 304766 340854 306972 340914
rect 306966 340852 306972 340854
rect 307036 340852 307042 340916
rect 232037 339826 232103 339829
rect 232037 339824 235060 339826
rect 232037 339768 232042 339824
rect 232098 339768 235060 339824
rect 232037 339766 235060 339768
rect 232037 339763 232103 339766
rect 304766 339690 304826 339796
rect 307201 339690 307267 339693
rect 304766 339688 307267 339690
rect 304766 339632 307206 339688
rect 307262 339632 307267 339688
rect 304766 339630 307267 339632
rect 307201 339627 307267 339630
rect 232037 338602 232103 338605
rect 580165 338602 580231 338605
rect 583520 338602 584960 338692
rect 232037 338600 235060 338602
rect 232037 338544 232042 338600
rect 232098 338544 235060 338600
rect 580165 338600 584960 338602
rect 232037 338542 235060 338544
rect 232037 338539 232103 338542
rect 304766 338330 304826 338572
rect 580165 338544 580170 338600
rect 580226 338544 584960 338600
rect 580165 338542 584960 338544
rect 580165 338539 580231 338542
rect 583520 338452 584960 338542
rect 307201 338330 307267 338333
rect 304766 338328 307267 338330
rect 304766 338272 307206 338328
rect 307262 338272 307267 338328
rect 304766 338270 307267 338272
rect 307201 338267 307267 338270
rect -960 332346 480 332436
rect 3049 332346 3115 332349
rect -960 332344 3115 332346
rect -960 332288 3054 332344
rect 3110 332288 3115 332344
rect -960 332286 3115 332288
rect -960 332196 480 332286
rect 3049 332283 3115 332286
rect 240593 326362 240659 326365
rect 240593 326360 240794 326362
rect 240593 326304 240598 326360
rect 240654 326304 240794 326360
rect 240593 326302 240794 326304
rect 240593 326299 240659 326302
rect 240734 326093 240794 326302
rect 240734 326088 240843 326093
rect 240734 326032 240782 326088
rect 240838 326032 240843 326088
rect 240734 326030 240843 326032
rect 240777 326027 240843 326030
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3049 319290 3115 319293
rect -960 319288 3115 319290
rect -960 319232 3054 319288
rect 3110 319232 3115 319288
rect -960 319230 3115 319232
rect -960 319140 480 319230
rect 3049 319227 3115 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3141 306234 3207 306237
rect -960 306232 3207 306234
rect -960 306176 3146 306232
rect 3202 306176 3207 306232
rect -960 306174 3207 306176
rect -960 306084 480 306174
rect 3141 306171 3207 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3141 293178 3207 293181
rect -960 293176 3207 293178
rect -960 293120 3146 293176
rect 3202 293120 3207 293176
rect -960 293118 3207 293120
rect -960 293028 480 293118
rect 3141 293115 3207 293118
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect -960 280122 480 280212
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3233 228034 3299 228037
rect -960 228032 3299 228034
rect -960 227976 3238 228032
rect 3294 227976 3299 228032
rect -960 227974 3299 227976
rect -960 227884 480 227974
rect 3233 227971 3299 227974
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3233 214978 3299 214981
rect -960 214976 3299 214978
rect -960 214920 3238 214976
rect 3294 214920 3299 214976
rect -960 214918 3299 214920
rect -960 214828 480 214918
rect 3233 214915 3299 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 3325 175946 3391 175949
rect -960 175944 3391 175946
rect -960 175888 3330 175944
rect 3386 175888 3391 175944
rect -960 175886 3391 175888
rect -960 175796 480 175886
rect 3325 175883 3391 175886
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 4061 162890 4127 162893
rect -960 162888 4127 162890
rect -960 162832 4066 162888
rect 4122 162832 4127 162888
rect -960 162830 4127 162832
rect -960 162740 480 162830
rect 4061 162827 4127 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3969 136778 4035 136781
rect -960 136776 4035 136778
rect -960 136720 3974 136776
rect 4030 136720 4035 136776
rect -960 136718 4035 136720
rect -960 136628 480 136718
rect 3969 136715 4035 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3141 123722 3207 123725
rect -960 123720 3207 123722
rect -960 123664 3146 123720
rect 3202 123664 3207 123720
rect -960 123662 3207 123664
rect -960 123572 480 123662
rect 3141 123659 3207 123662
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3877 110666 3943 110669
rect -960 110664 3943 110666
rect -960 110608 3882 110664
rect 3938 110608 3943 110664
rect -960 110606 3943 110608
rect -960 110516 480 110606
rect 3877 110603 3943 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3785 97610 3851 97613
rect -960 97608 3851 97610
rect -960 97552 3790 97608
rect 3846 97552 3851 97608
rect -960 97550 3851 97552
rect -960 97460 480 97550
rect 3785 97547 3851 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3693 71634 3759 71637
rect -960 71632 3759 71634
rect -960 71576 3698 71632
rect 3754 71576 3759 71632
rect -960 71574 3759 71576
rect -960 71484 480 71574
rect 3693 71571 3759 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2865 58578 2931 58581
rect -960 58576 2931 58578
rect -960 58520 2870 58576
rect 2926 58520 2931 58576
rect -960 58518 2931 58520
rect -960 58428 480 58518
rect 2865 58515 2931 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 583520 33146 584960 33236
rect 567150 33086 584960 33146
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 306966 31724 306972 31788
rect 307036 31786 307042 31788
rect 567150 31786 567210 33086
rect 583520 32996 584960 33086
rect 307036 31726 567210 31786
rect 307036 31724 307042 31726
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 20621 3770 20687 3773
rect 238201 3770 238267 3773
rect 20621 3768 238267 3770
rect 20621 3712 20626 3768
rect 20682 3712 238206 3768
rect 238262 3712 238267 3768
rect 20621 3710 238267 3712
rect 20621 3707 20687 3710
rect 238201 3707 238267 3710
rect 304901 3770 304967 3773
rect 579797 3770 579863 3773
rect 304901 3768 579863 3770
rect 304901 3712 304906 3768
rect 304962 3712 579802 3768
rect 579858 3712 579863 3768
rect 304901 3710 579863 3712
rect 304901 3707 304967 3710
rect 579797 3707 579863 3710
rect 15929 3634 15995 3637
rect 236729 3634 236795 3637
rect 15929 3632 236795 3634
rect 15929 3576 15934 3632
rect 15990 3576 236734 3632
rect 236790 3576 236795 3632
rect 15929 3574 236795 3576
rect 15929 3571 15995 3574
rect 236729 3571 236795 3574
rect 304809 3634 304875 3637
rect 580993 3634 581059 3637
rect 304809 3632 581059 3634
rect 304809 3576 304814 3632
rect 304870 3576 580998 3632
rect 581054 3576 581059 3632
rect 304809 3574 581059 3576
rect 304809 3571 304875 3574
rect 580993 3571 581059 3574
rect 14733 3498 14799 3501
rect 236453 3498 236519 3501
rect 14733 3496 236519 3498
rect 14733 3440 14738 3496
rect 14794 3440 236458 3496
rect 236514 3440 236519 3496
rect 14733 3438 236519 3440
rect 14733 3435 14799 3438
rect 236453 3435 236519 3438
rect 304625 3498 304691 3501
rect 582189 3498 582255 3501
rect 304625 3496 582255 3498
rect 304625 3440 304630 3496
rect 304686 3440 582194 3496
rect 582250 3440 582255 3496
rect 304625 3438 582255 3440
rect 304625 3435 304691 3438
rect 582189 3435 582255 3438
rect 6453 3362 6519 3365
rect 235257 3362 235323 3365
rect 6453 3360 235323 3362
rect 6453 3304 6458 3360
rect 6514 3304 235262 3360
rect 235318 3304 235323 3360
rect 6453 3302 235323 3304
rect 6453 3299 6519 3302
rect 235257 3299 235323 3302
rect 304717 3362 304783 3365
rect 583385 3362 583451 3365
rect 304717 3360 583451 3362
rect 304717 3304 304722 3360
rect 304778 3304 583390 3360
rect 583446 3304 583451 3360
rect 304717 3302 583451 3304
rect 304717 3299 304783 3302
rect 583385 3299 583451 3302
<< via3 >>
rect 3372 684252 3436 684316
rect 3372 405724 3436 405788
rect 306972 340852 307036 340916
rect 306972 31724 307036 31788
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 680254 -7976 710862
rect -8576 680018 -8394 680254
rect -8158 680018 -7976 680254
rect -8576 679934 -7976 680018
rect -8576 679698 -8394 679934
rect -8158 679698 -7976 679934
rect -8576 644254 -7976 679698
rect -8576 644018 -8394 644254
rect -8158 644018 -7976 644254
rect -8576 643934 -7976 644018
rect -8576 643698 -8394 643934
rect -8158 643698 -7976 643934
rect -8576 608254 -7976 643698
rect -8576 608018 -8394 608254
rect -8158 608018 -7976 608254
rect -8576 607934 -7976 608018
rect -8576 607698 -8394 607934
rect -8158 607698 -7976 607934
rect -8576 572254 -7976 607698
rect -8576 572018 -8394 572254
rect -8158 572018 -7976 572254
rect -8576 571934 -7976 572018
rect -8576 571698 -8394 571934
rect -8158 571698 -7976 571934
rect -8576 536254 -7976 571698
rect -8576 536018 -8394 536254
rect -8158 536018 -7976 536254
rect -8576 535934 -7976 536018
rect -8576 535698 -8394 535934
rect -8158 535698 -7976 535934
rect -8576 500254 -7976 535698
rect -8576 500018 -8394 500254
rect -8158 500018 -7976 500254
rect -8576 499934 -7976 500018
rect -8576 499698 -8394 499934
rect -8158 499698 -7976 499934
rect -8576 464254 -7976 499698
rect -8576 464018 -8394 464254
rect -8158 464018 -7976 464254
rect -8576 463934 -7976 464018
rect -8576 463698 -8394 463934
rect -8158 463698 -7976 463934
rect -8576 428254 -7976 463698
rect -8576 428018 -8394 428254
rect -8158 428018 -7976 428254
rect -8576 427934 -7976 428018
rect -8576 427698 -8394 427934
rect -8158 427698 -7976 427934
rect -8576 392254 -7976 427698
rect -8576 392018 -8394 392254
rect -8158 392018 -7976 392254
rect -8576 391934 -7976 392018
rect -8576 391698 -8394 391934
rect -8158 391698 -7976 391934
rect -8576 356254 -7976 391698
rect -8576 356018 -8394 356254
rect -8158 356018 -7976 356254
rect -8576 355934 -7976 356018
rect -8576 355698 -8394 355934
rect -8158 355698 -7976 355934
rect -8576 320254 -7976 355698
rect -8576 320018 -8394 320254
rect -8158 320018 -7976 320254
rect -8576 319934 -7976 320018
rect -8576 319698 -8394 319934
rect -8158 319698 -7976 319934
rect -8576 284254 -7976 319698
rect -8576 284018 -8394 284254
rect -8158 284018 -7976 284254
rect -8576 283934 -7976 284018
rect -8576 283698 -8394 283934
rect -8158 283698 -7976 283934
rect -8576 248254 -7976 283698
rect -8576 248018 -8394 248254
rect -8158 248018 -7976 248254
rect -8576 247934 -7976 248018
rect -8576 247698 -8394 247934
rect -8158 247698 -7976 247934
rect -8576 212254 -7976 247698
rect -8576 212018 -8394 212254
rect -8158 212018 -7976 212254
rect -8576 211934 -7976 212018
rect -8576 211698 -8394 211934
rect -8158 211698 -7976 211934
rect -8576 176254 -7976 211698
rect -8576 176018 -8394 176254
rect -8158 176018 -7976 176254
rect -8576 175934 -7976 176018
rect -8576 175698 -8394 175934
rect -8158 175698 -7976 175934
rect -8576 140254 -7976 175698
rect -8576 140018 -8394 140254
rect -8158 140018 -7976 140254
rect -8576 139934 -7976 140018
rect -8576 139698 -8394 139934
rect -8158 139698 -7976 139934
rect -8576 104254 -7976 139698
rect -8576 104018 -8394 104254
rect -8158 104018 -7976 104254
rect -8576 103934 -7976 104018
rect -8576 103698 -8394 103934
rect -8158 103698 -7976 103934
rect -8576 68254 -7976 103698
rect -8576 68018 -8394 68254
rect -8158 68018 -7976 68254
rect -8576 67934 -7976 68018
rect -8576 67698 -8394 67934
rect -8158 67698 -7976 67934
rect -8576 32254 -7976 67698
rect -8576 32018 -8394 32254
rect -8158 32018 -7976 32254
rect -8576 31934 -7976 32018
rect -8576 31698 -8394 31934
rect -8158 31698 -7976 31934
rect -8576 -6926 -7976 31698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 698254 -7036 709922
rect 12604 710478 13204 711440
rect 12604 710242 12786 710478
rect 13022 710242 13204 710478
rect 12604 710158 13204 710242
rect 12604 709922 12786 710158
rect 13022 709922 13204 710158
rect -7636 698018 -7454 698254
rect -7218 698018 -7036 698254
rect -7636 697934 -7036 698018
rect -7636 697698 -7454 697934
rect -7218 697698 -7036 697934
rect -7636 662254 -7036 697698
rect -7636 662018 -7454 662254
rect -7218 662018 -7036 662254
rect -7636 661934 -7036 662018
rect -7636 661698 -7454 661934
rect -7218 661698 -7036 661934
rect -7636 626254 -7036 661698
rect -7636 626018 -7454 626254
rect -7218 626018 -7036 626254
rect -7636 625934 -7036 626018
rect -7636 625698 -7454 625934
rect -7218 625698 -7036 625934
rect -7636 590254 -7036 625698
rect -7636 590018 -7454 590254
rect -7218 590018 -7036 590254
rect -7636 589934 -7036 590018
rect -7636 589698 -7454 589934
rect -7218 589698 -7036 589934
rect -7636 554254 -7036 589698
rect -7636 554018 -7454 554254
rect -7218 554018 -7036 554254
rect -7636 553934 -7036 554018
rect -7636 553698 -7454 553934
rect -7218 553698 -7036 553934
rect -7636 518254 -7036 553698
rect -7636 518018 -7454 518254
rect -7218 518018 -7036 518254
rect -7636 517934 -7036 518018
rect -7636 517698 -7454 517934
rect -7218 517698 -7036 517934
rect -7636 482254 -7036 517698
rect -7636 482018 -7454 482254
rect -7218 482018 -7036 482254
rect -7636 481934 -7036 482018
rect -7636 481698 -7454 481934
rect -7218 481698 -7036 481934
rect -7636 446254 -7036 481698
rect -7636 446018 -7454 446254
rect -7218 446018 -7036 446254
rect -7636 445934 -7036 446018
rect -7636 445698 -7454 445934
rect -7218 445698 -7036 445934
rect -7636 410254 -7036 445698
rect -7636 410018 -7454 410254
rect -7218 410018 -7036 410254
rect -7636 409934 -7036 410018
rect -7636 409698 -7454 409934
rect -7218 409698 -7036 409934
rect -7636 374254 -7036 409698
rect -7636 374018 -7454 374254
rect -7218 374018 -7036 374254
rect -7636 373934 -7036 374018
rect -7636 373698 -7454 373934
rect -7218 373698 -7036 373934
rect -7636 338254 -7036 373698
rect -7636 338018 -7454 338254
rect -7218 338018 -7036 338254
rect -7636 337934 -7036 338018
rect -7636 337698 -7454 337934
rect -7218 337698 -7036 337934
rect -7636 302254 -7036 337698
rect -7636 302018 -7454 302254
rect -7218 302018 -7036 302254
rect -7636 301934 -7036 302018
rect -7636 301698 -7454 301934
rect -7218 301698 -7036 301934
rect -7636 266254 -7036 301698
rect -7636 266018 -7454 266254
rect -7218 266018 -7036 266254
rect -7636 265934 -7036 266018
rect -7636 265698 -7454 265934
rect -7218 265698 -7036 265934
rect -7636 230254 -7036 265698
rect -7636 230018 -7454 230254
rect -7218 230018 -7036 230254
rect -7636 229934 -7036 230018
rect -7636 229698 -7454 229934
rect -7218 229698 -7036 229934
rect -7636 194254 -7036 229698
rect -7636 194018 -7454 194254
rect -7218 194018 -7036 194254
rect -7636 193934 -7036 194018
rect -7636 193698 -7454 193934
rect -7218 193698 -7036 193934
rect -7636 158254 -7036 193698
rect -7636 158018 -7454 158254
rect -7218 158018 -7036 158254
rect -7636 157934 -7036 158018
rect -7636 157698 -7454 157934
rect -7218 157698 -7036 157934
rect -7636 122254 -7036 157698
rect -7636 122018 -7454 122254
rect -7218 122018 -7036 122254
rect -7636 121934 -7036 122018
rect -7636 121698 -7454 121934
rect -7218 121698 -7036 121934
rect -7636 86254 -7036 121698
rect -7636 86018 -7454 86254
rect -7218 86018 -7036 86254
rect -7636 85934 -7036 86018
rect -7636 85698 -7454 85934
rect -7218 85698 -7036 85934
rect -7636 50254 -7036 85698
rect -7636 50018 -7454 50254
rect -7218 50018 -7036 50254
rect -7636 49934 -7036 50018
rect -7636 49698 -7454 49934
rect -7218 49698 -7036 49934
rect -7636 14254 -7036 49698
rect -7636 14018 -7454 14254
rect -7218 14018 -7036 14254
rect -7636 13934 -7036 14018
rect -7636 13698 -7454 13934
rect -7218 13698 -7036 13934
rect -7636 -5986 -7036 13698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 676654 -6096 708982
rect -6696 676418 -6514 676654
rect -6278 676418 -6096 676654
rect -6696 676334 -6096 676418
rect -6696 676098 -6514 676334
rect -6278 676098 -6096 676334
rect -6696 640654 -6096 676098
rect -6696 640418 -6514 640654
rect -6278 640418 -6096 640654
rect -6696 640334 -6096 640418
rect -6696 640098 -6514 640334
rect -6278 640098 -6096 640334
rect -6696 604654 -6096 640098
rect -6696 604418 -6514 604654
rect -6278 604418 -6096 604654
rect -6696 604334 -6096 604418
rect -6696 604098 -6514 604334
rect -6278 604098 -6096 604334
rect -6696 568654 -6096 604098
rect -6696 568418 -6514 568654
rect -6278 568418 -6096 568654
rect -6696 568334 -6096 568418
rect -6696 568098 -6514 568334
rect -6278 568098 -6096 568334
rect -6696 532654 -6096 568098
rect -6696 532418 -6514 532654
rect -6278 532418 -6096 532654
rect -6696 532334 -6096 532418
rect -6696 532098 -6514 532334
rect -6278 532098 -6096 532334
rect -6696 496654 -6096 532098
rect -6696 496418 -6514 496654
rect -6278 496418 -6096 496654
rect -6696 496334 -6096 496418
rect -6696 496098 -6514 496334
rect -6278 496098 -6096 496334
rect -6696 460654 -6096 496098
rect -6696 460418 -6514 460654
rect -6278 460418 -6096 460654
rect -6696 460334 -6096 460418
rect -6696 460098 -6514 460334
rect -6278 460098 -6096 460334
rect -6696 424654 -6096 460098
rect -6696 424418 -6514 424654
rect -6278 424418 -6096 424654
rect -6696 424334 -6096 424418
rect -6696 424098 -6514 424334
rect -6278 424098 -6096 424334
rect -6696 388654 -6096 424098
rect -6696 388418 -6514 388654
rect -6278 388418 -6096 388654
rect -6696 388334 -6096 388418
rect -6696 388098 -6514 388334
rect -6278 388098 -6096 388334
rect -6696 352654 -6096 388098
rect -6696 352418 -6514 352654
rect -6278 352418 -6096 352654
rect -6696 352334 -6096 352418
rect -6696 352098 -6514 352334
rect -6278 352098 -6096 352334
rect -6696 316654 -6096 352098
rect -6696 316418 -6514 316654
rect -6278 316418 -6096 316654
rect -6696 316334 -6096 316418
rect -6696 316098 -6514 316334
rect -6278 316098 -6096 316334
rect -6696 280654 -6096 316098
rect -6696 280418 -6514 280654
rect -6278 280418 -6096 280654
rect -6696 280334 -6096 280418
rect -6696 280098 -6514 280334
rect -6278 280098 -6096 280334
rect -6696 244654 -6096 280098
rect -6696 244418 -6514 244654
rect -6278 244418 -6096 244654
rect -6696 244334 -6096 244418
rect -6696 244098 -6514 244334
rect -6278 244098 -6096 244334
rect -6696 208654 -6096 244098
rect -6696 208418 -6514 208654
rect -6278 208418 -6096 208654
rect -6696 208334 -6096 208418
rect -6696 208098 -6514 208334
rect -6278 208098 -6096 208334
rect -6696 172654 -6096 208098
rect -6696 172418 -6514 172654
rect -6278 172418 -6096 172654
rect -6696 172334 -6096 172418
rect -6696 172098 -6514 172334
rect -6278 172098 -6096 172334
rect -6696 136654 -6096 172098
rect -6696 136418 -6514 136654
rect -6278 136418 -6096 136654
rect -6696 136334 -6096 136418
rect -6696 136098 -6514 136334
rect -6278 136098 -6096 136334
rect -6696 100654 -6096 136098
rect -6696 100418 -6514 100654
rect -6278 100418 -6096 100654
rect -6696 100334 -6096 100418
rect -6696 100098 -6514 100334
rect -6278 100098 -6096 100334
rect -6696 64654 -6096 100098
rect -6696 64418 -6514 64654
rect -6278 64418 -6096 64654
rect -6696 64334 -6096 64418
rect -6696 64098 -6514 64334
rect -6278 64098 -6096 64334
rect -6696 28654 -6096 64098
rect -6696 28418 -6514 28654
rect -6278 28418 -6096 28654
rect -6696 28334 -6096 28418
rect -6696 28098 -6514 28334
rect -6278 28098 -6096 28334
rect -6696 -5046 -6096 28098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 694654 -5156 708042
rect 9004 708598 9604 709560
rect 9004 708362 9186 708598
rect 9422 708362 9604 708598
rect 9004 708278 9604 708362
rect 9004 708042 9186 708278
rect 9422 708042 9604 708278
rect -5756 694418 -5574 694654
rect -5338 694418 -5156 694654
rect -5756 694334 -5156 694418
rect -5756 694098 -5574 694334
rect -5338 694098 -5156 694334
rect -5756 658654 -5156 694098
rect -5756 658418 -5574 658654
rect -5338 658418 -5156 658654
rect -5756 658334 -5156 658418
rect -5756 658098 -5574 658334
rect -5338 658098 -5156 658334
rect -5756 622654 -5156 658098
rect -5756 622418 -5574 622654
rect -5338 622418 -5156 622654
rect -5756 622334 -5156 622418
rect -5756 622098 -5574 622334
rect -5338 622098 -5156 622334
rect -5756 586654 -5156 622098
rect -5756 586418 -5574 586654
rect -5338 586418 -5156 586654
rect -5756 586334 -5156 586418
rect -5756 586098 -5574 586334
rect -5338 586098 -5156 586334
rect -5756 550654 -5156 586098
rect -5756 550418 -5574 550654
rect -5338 550418 -5156 550654
rect -5756 550334 -5156 550418
rect -5756 550098 -5574 550334
rect -5338 550098 -5156 550334
rect -5756 514654 -5156 550098
rect -5756 514418 -5574 514654
rect -5338 514418 -5156 514654
rect -5756 514334 -5156 514418
rect -5756 514098 -5574 514334
rect -5338 514098 -5156 514334
rect -5756 478654 -5156 514098
rect -5756 478418 -5574 478654
rect -5338 478418 -5156 478654
rect -5756 478334 -5156 478418
rect -5756 478098 -5574 478334
rect -5338 478098 -5156 478334
rect -5756 442654 -5156 478098
rect -5756 442418 -5574 442654
rect -5338 442418 -5156 442654
rect -5756 442334 -5156 442418
rect -5756 442098 -5574 442334
rect -5338 442098 -5156 442334
rect -5756 406654 -5156 442098
rect -5756 406418 -5574 406654
rect -5338 406418 -5156 406654
rect -5756 406334 -5156 406418
rect -5756 406098 -5574 406334
rect -5338 406098 -5156 406334
rect -5756 370654 -5156 406098
rect -5756 370418 -5574 370654
rect -5338 370418 -5156 370654
rect -5756 370334 -5156 370418
rect -5756 370098 -5574 370334
rect -5338 370098 -5156 370334
rect -5756 334654 -5156 370098
rect -5756 334418 -5574 334654
rect -5338 334418 -5156 334654
rect -5756 334334 -5156 334418
rect -5756 334098 -5574 334334
rect -5338 334098 -5156 334334
rect -5756 298654 -5156 334098
rect -5756 298418 -5574 298654
rect -5338 298418 -5156 298654
rect -5756 298334 -5156 298418
rect -5756 298098 -5574 298334
rect -5338 298098 -5156 298334
rect -5756 262654 -5156 298098
rect -5756 262418 -5574 262654
rect -5338 262418 -5156 262654
rect -5756 262334 -5156 262418
rect -5756 262098 -5574 262334
rect -5338 262098 -5156 262334
rect -5756 226654 -5156 262098
rect -5756 226418 -5574 226654
rect -5338 226418 -5156 226654
rect -5756 226334 -5156 226418
rect -5756 226098 -5574 226334
rect -5338 226098 -5156 226334
rect -5756 190654 -5156 226098
rect -5756 190418 -5574 190654
rect -5338 190418 -5156 190654
rect -5756 190334 -5156 190418
rect -5756 190098 -5574 190334
rect -5338 190098 -5156 190334
rect -5756 154654 -5156 190098
rect -5756 154418 -5574 154654
rect -5338 154418 -5156 154654
rect -5756 154334 -5156 154418
rect -5756 154098 -5574 154334
rect -5338 154098 -5156 154334
rect -5756 118654 -5156 154098
rect -5756 118418 -5574 118654
rect -5338 118418 -5156 118654
rect -5756 118334 -5156 118418
rect -5756 118098 -5574 118334
rect -5338 118098 -5156 118334
rect -5756 82654 -5156 118098
rect -5756 82418 -5574 82654
rect -5338 82418 -5156 82654
rect -5756 82334 -5156 82418
rect -5756 82098 -5574 82334
rect -5338 82098 -5156 82334
rect -5756 46654 -5156 82098
rect -5756 46418 -5574 46654
rect -5338 46418 -5156 46654
rect -5756 46334 -5156 46418
rect -5756 46098 -5574 46334
rect -5338 46098 -5156 46334
rect -5756 10654 -5156 46098
rect -5756 10418 -5574 10654
rect -5338 10418 -5156 10654
rect -5756 10334 -5156 10418
rect -5756 10098 -5574 10334
rect -5338 10098 -5156 10334
rect -5756 -4106 -5156 10098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 673054 -4216 707102
rect -4816 672818 -4634 673054
rect -4398 672818 -4216 673054
rect -4816 672734 -4216 672818
rect -4816 672498 -4634 672734
rect -4398 672498 -4216 672734
rect -4816 637054 -4216 672498
rect -4816 636818 -4634 637054
rect -4398 636818 -4216 637054
rect -4816 636734 -4216 636818
rect -4816 636498 -4634 636734
rect -4398 636498 -4216 636734
rect -4816 601054 -4216 636498
rect -4816 600818 -4634 601054
rect -4398 600818 -4216 601054
rect -4816 600734 -4216 600818
rect -4816 600498 -4634 600734
rect -4398 600498 -4216 600734
rect -4816 565054 -4216 600498
rect -4816 564818 -4634 565054
rect -4398 564818 -4216 565054
rect -4816 564734 -4216 564818
rect -4816 564498 -4634 564734
rect -4398 564498 -4216 564734
rect -4816 529054 -4216 564498
rect -4816 528818 -4634 529054
rect -4398 528818 -4216 529054
rect -4816 528734 -4216 528818
rect -4816 528498 -4634 528734
rect -4398 528498 -4216 528734
rect -4816 493054 -4216 528498
rect -4816 492818 -4634 493054
rect -4398 492818 -4216 493054
rect -4816 492734 -4216 492818
rect -4816 492498 -4634 492734
rect -4398 492498 -4216 492734
rect -4816 457054 -4216 492498
rect -4816 456818 -4634 457054
rect -4398 456818 -4216 457054
rect -4816 456734 -4216 456818
rect -4816 456498 -4634 456734
rect -4398 456498 -4216 456734
rect -4816 421054 -4216 456498
rect -4816 420818 -4634 421054
rect -4398 420818 -4216 421054
rect -4816 420734 -4216 420818
rect -4816 420498 -4634 420734
rect -4398 420498 -4216 420734
rect -4816 385054 -4216 420498
rect -4816 384818 -4634 385054
rect -4398 384818 -4216 385054
rect -4816 384734 -4216 384818
rect -4816 384498 -4634 384734
rect -4398 384498 -4216 384734
rect -4816 349054 -4216 384498
rect -4816 348818 -4634 349054
rect -4398 348818 -4216 349054
rect -4816 348734 -4216 348818
rect -4816 348498 -4634 348734
rect -4398 348498 -4216 348734
rect -4816 313054 -4216 348498
rect -4816 312818 -4634 313054
rect -4398 312818 -4216 313054
rect -4816 312734 -4216 312818
rect -4816 312498 -4634 312734
rect -4398 312498 -4216 312734
rect -4816 277054 -4216 312498
rect -4816 276818 -4634 277054
rect -4398 276818 -4216 277054
rect -4816 276734 -4216 276818
rect -4816 276498 -4634 276734
rect -4398 276498 -4216 276734
rect -4816 241054 -4216 276498
rect -4816 240818 -4634 241054
rect -4398 240818 -4216 241054
rect -4816 240734 -4216 240818
rect -4816 240498 -4634 240734
rect -4398 240498 -4216 240734
rect -4816 205054 -4216 240498
rect -4816 204818 -4634 205054
rect -4398 204818 -4216 205054
rect -4816 204734 -4216 204818
rect -4816 204498 -4634 204734
rect -4398 204498 -4216 204734
rect -4816 169054 -4216 204498
rect -4816 168818 -4634 169054
rect -4398 168818 -4216 169054
rect -4816 168734 -4216 168818
rect -4816 168498 -4634 168734
rect -4398 168498 -4216 168734
rect -4816 133054 -4216 168498
rect -4816 132818 -4634 133054
rect -4398 132818 -4216 133054
rect -4816 132734 -4216 132818
rect -4816 132498 -4634 132734
rect -4398 132498 -4216 132734
rect -4816 97054 -4216 132498
rect -4816 96818 -4634 97054
rect -4398 96818 -4216 97054
rect -4816 96734 -4216 96818
rect -4816 96498 -4634 96734
rect -4398 96498 -4216 96734
rect -4816 61054 -4216 96498
rect -4816 60818 -4634 61054
rect -4398 60818 -4216 61054
rect -4816 60734 -4216 60818
rect -4816 60498 -4634 60734
rect -4398 60498 -4216 60734
rect -4816 25054 -4216 60498
rect -4816 24818 -4634 25054
rect -4398 24818 -4216 25054
rect -4816 24734 -4216 24818
rect -4816 24498 -4634 24734
rect -4398 24498 -4216 24734
rect -4816 -3166 -4216 24498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 691054 -3276 706162
rect 5404 706718 6004 707680
rect 5404 706482 5586 706718
rect 5822 706482 6004 706718
rect 5404 706398 6004 706482
rect 5404 706162 5586 706398
rect 5822 706162 6004 706398
rect -3876 690818 -3694 691054
rect -3458 690818 -3276 691054
rect -3876 690734 -3276 690818
rect -3876 690498 -3694 690734
rect -3458 690498 -3276 690734
rect -3876 655054 -3276 690498
rect -3876 654818 -3694 655054
rect -3458 654818 -3276 655054
rect -3876 654734 -3276 654818
rect -3876 654498 -3694 654734
rect -3458 654498 -3276 654734
rect -3876 619054 -3276 654498
rect -3876 618818 -3694 619054
rect -3458 618818 -3276 619054
rect -3876 618734 -3276 618818
rect -3876 618498 -3694 618734
rect -3458 618498 -3276 618734
rect -3876 583054 -3276 618498
rect -3876 582818 -3694 583054
rect -3458 582818 -3276 583054
rect -3876 582734 -3276 582818
rect -3876 582498 -3694 582734
rect -3458 582498 -3276 582734
rect -3876 547054 -3276 582498
rect -3876 546818 -3694 547054
rect -3458 546818 -3276 547054
rect -3876 546734 -3276 546818
rect -3876 546498 -3694 546734
rect -3458 546498 -3276 546734
rect -3876 511054 -3276 546498
rect -3876 510818 -3694 511054
rect -3458 510818 -3276 511054
rect -3876 510734 -3276 510818
rect -3876 510498 -3694 510734
rect -3458 510498 -3276 510734
rect -3876 475054 -3276 510498
rect -3876 474818 -3694 475054
rect -3458 474818 -3276 475054
rect -3876 474734 -3276 474818
rect -3876 474498 -3694 474734
rect -3458 474498 -3276 474734
rect -3876 439054 -3276 474498
rect -3876 438818 -3694 439054
rect -3458 438818 -3276 439054
rect -3876 438734 -3276 438818
rect -3876 438498 -3694 438734
rect -3458 438498 -3276 438734
rect -3876 403054 -3276 438498
rect -3876 402818 -3694 403054
rect -3458 402818 -3276 403054
rect -3876 402734 -3276 402818
rect -3876 402498 -3694 402734
rect -3458 402498 -3276 402734
rect -3876 367054 -3276 402498
rect -3876 366818 -3694 367054
rect -3458 366818 -3276 367054
rect -3876 366734 -3276 366818
rect -3876 366498 -3694 366734
rect -3458 366498 -3276 366734
rect -3876 331054 -3276 366498
rect -3876 330818 -3694 331054
rect -3458 330818 -3276 331054
rect -3876 330734 -3276 330818
rect -3876 330498 -3694 330734
rect -3458 330498 -3276 330734
rect -3876 295054 -3276 330498
rect -3876 294818 -3694 295054
rect -3458 294818 -3276 295054
rect -3876 294734 -3276 294818
rect -3876 294498 -3694 294734
rect -3458 294498 -3276 294734
rect -3876 259054 -3276 294498
rect -3876 258818 -3694 259054
rect -3458 258818 -3276 259054
rect -3876 258734 -3276 258818
rect -3876 258498 -3694 258734
rect -3458 258498 -3276 258734
rect -3876 223054 -3276 258498
rect -3876 222818 -3694 223054
rect -3458 222818 -3276 223054
rect -3876 222734 -3276 222818
rect -3876 222498 -3694 222734
rect -3458 222498 -3276 222734
rect -3876 187054 -3276 222498
rect -3876 186818 -3694 187054
rect -3458 186818 -3276 187054
rect -3876 186734 -3276 186818
rect -3876 186498 -3694 186734
rect -3458 186498 -3276 186734
rect -3876 151054 -3276 186498
rect -3876 150818 -3694 151054
rect -3458 150818 -3276 151054
rect -3876 150734 -3276 150818
rect -3876 150498 -3694 150734
rect -3458 150498 -3276 150734
rect -3876 115054 -3276 150498
rect -3876 114818 -3694 115054
rect -3458 114818 -3276 115054
rect -3876 114734 -3276 114818
rect -3876 114498 -3694 114734
rect -3458 114498 -3276 114734
rect -3876 79054 -3276 114498
rect -3876 78818 -3694 79054
rect -3458 78818 -3276 79054
rect -3876 78734 -3276 78818
rect -3876 78498 -3694 78734
rect -3458 78498 -3276 78734
rect -3876 43054 -3276 78498
rect -3876 42818 -3694 43054
rect -3458 42818 -3276 43054
rect -3876 42734 -3276 42818
rect -3876 42498 -3694 42734
rect -3458 42498 -3276 42734
rect -3876 7054 -3276 42498
rect -3876 6818 -3694 7054
rect -3458 6818 -3276 7054
rect -3876 6734 -3276 6818
rect -3876 6498 -3694 6734
rect -3458 6498 -3276 6734
rect -3876 -2226 -3276 6498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 669454 -2336 705222
rect -2936 669218 -2754 669454
rect -2518 669218 -2336 669454
rect -2936 669134 -2336 669218
rect -2936 668898 -2754 669134
rect -2518 668898 -2336 669134
rect -2936 633454 -2336 668898
rect -2936 633218 -2754 633454
rect -2518 633218 -2336 633454
rect -2936 633134 -2336 633218
rect -2936 632898 -2754 633134
rect -2518 632898 -2336 633134
rect -2936 597454 -2336 632898
rect -2936 597218 -2754 597454
rect -2518 597218 -2336 597454
rect -2936 597134 -2336 597218
rect -2936 596898 -2754 597134
rect -2518 596898 -2336 597134
rect -2936 561454 -2336 596898
rect -2936 561218 -2754 561454
rect -2518 561218 -2336 561454
rect -2936 561134 -2336 561218
rect -2936 560898 -2754 561134
rect -2518 560898 -2336 561134
rect -2936 525454 -2336 560898
rect -2936 525218 -2754 525454
rect -2518 525218 -2336 525454
rect -2936 525134 -2336 525218
rect -2936 524898 -2754 525134
rect -2518 524898 -2336 525134
rect -2936 489454 -2336 524898
rect -2936 489218 -2754 489454
rect -2518 489218 -2336 489454
rect -2936 489134 -2336 489218
rect -2936 488898 -2754 489134
rect -2518 488898 -2336 489134
rect -2936 453454 -2336 488898
rect -2936 453218 -2754 453454
rect -2518 453218 -2336 453454
rect -2936 453134 -2336 453218
rect -2936 452898 -2754 453134
rect -2518 452898 -2336 453134
rect -2936 417454 -2336 452898
rect -2936 417218 -2754 417454
rect -2518 417218 -2336 417454
rect -2936 417134 -2336 417218
rect -2936 416898 -2754 417134
rect -2518 416898 -2336 417134
rect -2936 381454 -2336 416898
rect -2936 381218 -2754 381454
rect -2518 381218 -2336 381454
rect -2936 381134 -2336 381218
rect -2936 380898 -2754 381134
rect -2518 380898 -2336 381134
rect -2936 345454 -2336 380898
rect -2936 345218 -2754 345454
rect -2518 345218 -2336 345454
rect -2936 345134 -2336 345218
rect -2936 344898 -2754 345134
rect -2518 344898 -2336 345134
rect -2936 309454 -2336 344898
rect -2936 309218 -2754 309454
rect -2518 309218 -2336 309454
rect -2936 309134 -2336 309218
rect -2936 308898 -2754 309134
rect -2518 308898 -2336 309134
rect -2936 273454 -2336 308898
rect -2936 273218 -2754 273454
rect -2518 273218 -2336 273454
rect -2936 273134 -2336 273218
rect -2936 272898 -2754 273134
rect -2518 272898 -2336 273134
rect -2936 237454 -2336 272898
rect -2936 237218 -2754 237454
rect -2518 237218 -2336 237454
rect -2936 237134 -2336 237218
rect -2936 236898 -2754 237134
rect -2518 236898 -2336 237134
rect -2936 201454 -2336 236898
rect -2936 201218 -2754 201454
rect -2518 201218 -2336 201454
rect -2936 201134 -2336 201218
rect -2936 200898 -2754 201134
rect -2518 200898 -2336 201134
rect -2936 165454 -2336 200898
rect -2936 165218 -2754 165454
rect -2518 165218 -2336 165454
rect -2936 165134 -2336 165218
rect -2936 164898 -2754 165134
rect -2518 164898 -2336 165134
rect -2936 129454 -2336 164898
rect -2936 129218 -2754 129454
rect -2518 129218 -2336 129454
rect -2936 129134 -2336 129218
rect -2936 128898 -2754 129134
rect -2518 128898 -2336 129134
rect -2936 93454 -2336 128898
rect -2936 93218 -2754 93454
rect -2518 93218 -2336 93454
rect -2936 93134 -2336 93218
rect -2936 92898 -2754 93134
rect -2518 92898 -2336 93134
rect -2936 57454 -2336 92898
rect -2936 57218 -2754 57454
rect -2518 57218 -2336 57454
rect -2936 57134 -2336 57218
rect -2936 56898 -2754 57134
rect -2518 56898 -2336 57134
rect -2936 21454 -2336 56898
rect -2936 21218 -2754 21454
rect -2518 21218 -2336 21454
rect -2936 21134 -2336 21218
rect -2936 20898 -2754 21134
rect -2518 20898 -2336 21134
rect -2936 -1286 -2336 20898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 687454 -1396 704282
rect -1996 687218 -1814 687454
rect -1578 687218 -1396 687454
rect -1996 687134 -1396 687218
rect -1996 686898 -1814 687134
rect -1578 686898 -1396 687134
rect -1996 651454 -1396 686898
rect -1996 651218 -1814 651454
rect -1578 651218 -1396 651454
rect -1996 651134 -1396 651218
rect -1996 650898 -1814 651134
rect -1578 650898 -1396 651134
rect -1996 615454 -1396 650898
rect -1996 615218 -1814 615454
rect -1578 615218 -1396 615454
rect -1996 615134 -1396 615218
rect -1996 614898 -1814 615134
rect -1578 614898 -1396 615134
rect -1996 579454 -1396 614898
rect -1996 579218 -1814 579454
rect -1578 579218 -1396 579454
rect -1996 579134 -1396 579218
rect -1996 578898 -1814 579134
rect -1578 578898 -1396 579134
rect -1996 543454 -1396 578898
rect -1996 543218 -1814 543454
rect -1578 543218 -1396 543454
rect -1996 543134 -1396 543218
rect -1996 542898 -1814 543134
rect -1578 542898 -1396 543134
rect -1996 507454 -1396 542898
rect -1996 507218 -1814 507454
rect -1578 507218 -1396 507454
rect -1996 507134 -1396 507218
rect -1996 506898 -1814 507134
rect -1578 506898 -1396 507134
rect -1996 471454 -1396 506898
rect -1996 471218 -1814 471454
rect -1578 471218 -1396 471454
rect -1996 471134 -1396 471218
rect -1996 470898 -1814 471134
rect -1578 470898 -1396 471134
rect -1996 435454 -1396 470898
rect -1996 435218 -1814 435454
rect -1578 435218 -1396 435454
rect -1996 435134 -1396 435218
rect -1996 434898 -1814 435134
rect -1578 434898 -1396 435134
rect -1996 399454 -1396 434898
rect -1996 399218 -1814 399454
rect -1578 399218 -1396 399454
rect -1996 399134 -1396 399218
rect -1996 398898 -1814 399134
rect -1578 398898 -1396 399134
rect -1996 363454 -1396 398898
rect -1996 363218 -1814 363454
rect -1578 363218 -1396 363454
rect -1996 363134 -1396 363218
rect -1996 362898 -1814 363134
rect -1578 362898 -1396 363134
rect -1996 327454 -1396 362898
rect -1996 327218 -1814 327454
rect -1578 327218 -1396 327454
rect -1996 327134 -1396 327218
rect -1996 326898 -1814 327134
rect -1578 326898 -1396 327134
rect -1996 291454 -1396 326898
rect -1996 291218 -1814 291454
rect -1578 291218 -1396 291454
rect -1996 291134 -1396 291218
rect -1996 290898 -1814 291134
rect -1578 290898 -1396 291134
rect -1996 255454 -1396 290898
rect -1996 255218 -1814 255454
rect -1578 255218 -1396 255454
rect -1996 255134 -1396 255218
rect -1996 254898 -1814 255134
rect -1578 254898 -1396 255134
rect -1996 219454 -1396 254898
rect -1996 219218 -1814 219454
rect -1578 219218 -1396 219454
rect -1996 219134 -1396 219218
rect -1996 218898 -1814 219134
rect -1578 218898 -1396 219134
rect -1996 183454 -1396 218898
rect -1996 183218 -1814 183454
rect -1578 183218 -1396 183454
rect -1996 183134 -1396 183218
rect -1996 182898 -1814 183134
rect -1578 182898 -1396 183134
rect -1996 147454 -1396 182898
rect -1996 147218 -1814 147454
rect -1578 147218 -1396 147454
rect -1996 147134 -1396 147218
rect -1996 146898 -1814 147134
rect -1578 146898 -1396 147134
rect -1996 111454 -1396 146898
rect -1996 111218 -1814 111454
rect -1578 111218 -1396 111454
rect -1996 111134 -1396 111218
rect -1996 110898 -1814 111134
rect -1578 110898 -1396 111134
rect -1996 75454 -1396 110898
rect -1996 75218 -1814 75454
rect -1578 75218 -1396 75454
rect -1996 75134 -1396 75218
rect -1996 74898 -1814 75134
rect -1578 74898 -1396 75134
rect -1996 39454 -1396 74898
rect -1996 39218 -1814 39454
rect -1578 39218 -1396 39454
rect -1996 39134 -1396 39218
rect -1996 38898 -1814 39134
rect -1578 38898 -1396 39134
rect -1996 3454 -1396 38898
rect -1996 3218 -1814 3454
rect -1578 3218 -1396 3454
rect -1996 3134 -1396 3218
rect -1996 2898 -1814 3134
rect -1578 2898 -1396 3134
rect -1996 -346 -1396 2898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 1804 704838 2404 705800
rect 1804 704602 1986 704838
rect 2222 704602 2404 704838
rect 1804 704518 2404 704602
rect 1804 704282 1986 704518
rect 2222 704282 2404 704518
rect 1804 687454 2404 704282
rect 1804 687218 1986 687454
rect 2222 687218 2404 687454
rect 1804 687134 2404 687218
rect 1804 686898 1986 687134
rect 2222 686898 2404 687134
rect 1804 651454 2404 686898
rect 5404 691054 6004 706162
rect 5404 690818 5586 691054
rect 5822 690818 6004 691054
rect 5404 690734 6004 690818
rect 5404 690498 5586 690734
rect 5822 690498 6004 690734
rect 3371 684316 3437 684317
rect 3371 684252 3372 684316
rect 3436 684252 3437 684316
rect 3371 684251 3437 684252
rect 1804 651218 1986 651454
rect 2222 651218 2404 651454
rect 1804 651134 2404 651218
rect 1804 650898 1986 651134
rect 2222 650898 2404 651134
rect 1804 615454 2404 650898
rect 1804 615218 1986 615454
rect 2222 615218 2404 615454
rect 1804 615134 2404 615218
rect 1804 614898 1986 615134
rect 2222 614898 2404 615134
rect 1804 579454 2404 614898
rect 1804 579218 1986 579454
rect 2222 579218 2404 579454
rect 1804 579134 2404 579218
rect 1804 578898 1986 579134
rect 2222 578898 2404 579134
rect 1804 543454 2404 578898
rect 1804 543218 1986 543454
rect 2222 543218 2404 543454
rect 1804 543134 2404 543218
rect 1804 542898 1986 543134
rect 2222 542898 2404 543134
rect 1804 507454 2404 542898
rect 1804 507218 1986 507454
rect 2222 507218 2404 507454
rect 1804 507134 2404 507218
rect 1804 506898 1986 507134
rect 2222 506898 2404 507134
rect 1804 471454 2404 506898
rect 1804 471218 1986 471454
rect 2222 471218 2404 471454
rect 1804 471134 2404 471218
rect 1804 470898 1986 471134
rect 2222 470898 2404 471134
rect 1804 435454 2404 470898
rect 1804 435218 1986 435454
rect 2222 435218 2404 435454
rect 1804 435134 2404 435218
rect 1804 434898 1986 435134
rect 2222 434898 2404 435134
rect 1804 399454 2404 434898
rect 3374 405789 3434 684251
rect 5404 655054 6004 690498
rect 5404 654818 5586 655054
rect 5822 654818 6004 655054
rect 5404 654734 6004 654818
rect 5404 654498 5586 654734
rect 5822 654498 6004 654734
rect 5404 619054 6004 654498
rect 5404 618818 5586 619054
rect 5822 618818 6004 619054
rect 5404 618734 6004 618818
rect 5404 618498 5586 618734
rect 5822 618498 6004 618734
rect 5404 583054 6004 618498
rect 5404 582818 5586 583054
rect 5822 582818 6004 583054
rect 5404 582734 6004 582818
rect 5404 582498 5586 582734
rect 5822 582498 6004 582734
rect 5404 547054 6004 582498
rect 5404 546818 5586 547054
rect 5822 546818 6004 547054
rect 5404 546734 6004 546818
rect 5404 546498 5586 546734
rect 5822 546498 6004 546734
rect 5404 511054 6004 546498
rect 5404 510818 5586 511054
rect 5822 510818 6004 511054
rect 5404 510734 6004 510818
rect 5404 510498 5586 510734
rect 5822 510498 6004 510734
rect 5404 475054 6004 510498
rect 5404 474818 5586 475054
rect 5822 474818 6004 475054
rect 5404 474734 6004 474818
rect 5404 474498 5586 474734
rect 5822 474498 6004 474734
rect 5404 439054 6004 474498
rect 5404 438818 5586 439054
rect 5822 438818 6004 439054
rect 5404 438734 6004 438818
rect 5404 438498 5586 438734
rect 5822 438498 6004 438734
rect 3371 405788 3437 405789
rect 3371 405724 3372 405788
rect 3436 405724 3437 405788
rect 3371 405723 3437 405724
rect 1804 399218 1986 399454
rect 2222 399218 2404 399454
rect 1804 399134 2404 399218
rect 1804 398898 1986 399134
rect 2222 398898 2404 399134
rect 1804 363454 2404 398898
rect 1804 363218 1986 363454
rect 2222 363218 2404 363454
rect 1804 363134 2404 363218
rect 1804 362898 1986 363134
rect 2222 362898 2404 363134
rect 1804 327454 2404 362898
rect 1804 327218 1986 327454
rect 2222 327218 2404 327454
rect 1804 327134 2404 327218
rect 1804 326898 1986 327134
rect 2222 326898 2404 327134
rect 1804 291454 2404 326898
rect 1804 291218 1986 291454
rect 2222 291218 2404 291454
rect 1804 291134 2404 291218
rect 1804 290898 1986 291134
rect 2222 290898 2404 291134
rect 1804 255454 2404 290898
rect 1804 255218 1986 255454
rect 2222 255218 2404 255454
rect 1804 255134 2404 255218
rect 1804 254898 1986 255134
rect 2222 254898 2404 255134
rect 1804 219454 2404 254898
rect 1804 219218 1986 219454
rect 2222 219218 2404 219454
rect 1804 219134 2404 219218
rect 1804 218898 1986 219134
rect 2222 218898 2404 219134
rect 1804 183454 2404 218898
rect 1804 183218 1986 183454
rect 2222 183218 2404 183454
rect 1804 183134 2404 183218
rect 1804 182898 1986 183134
rect 2222 182898 2404 183134
rect 1804 147454 2404 182898
rect 1804 147218 1986 147454
rect 2222 147218 2404 147454
rect 1804 147134 2404 147218
rect 1804 146898 1986 147134
rect 2222 146898 2404 147134
rect 1804 111454 2404 146898
rect 1804 111218 1986 111454
rect 2222 111218 2404 111454
rect 1804 111134 2404 111218
rect 1804 110898 1986 111134
rect 2222 110898 2404 111134
rect 1804 75454 2404 110898
rect 1804 75218 1986 75454
rect 2222 75218 2404 75454
rect 1804 75134 2404 75218
rect 1804 74898 1986 75134
rect 2222 74898 2404 75134
rect 1804 39454 2404 74898
rect 1804 39218 1986 39454
rect 2222 39218 2404 39454
rect 1804 39134 2404 39218
rect 1804 38898 1986 39134
rect 2222 38898 2404 39134
rect 1804 3454 2404 38898
rect 1804 3218 1986 3454
rect 2222 3218 2404 3454
rect 1804 3134 2404 3218
rect 1804 2898 1986 3134
rect 2222 2898 2404 3134
rect 1804 -346 2404 2898
rect 1804 -582 1986 -346
rect 2222 -582 2404 -346
rect 1804 -666 2404 -582
rect 1804 -902 1986 -666
rect 2222 -902 2404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 1804 -1864 2404 -902
rect 5404 403054 6004 438498
rect 5404 402818 5586 403054
rect 5822 402818 6004 403054
rect 5404 402734 6004 402818
rect 5404 402498 5586 402734
rect 5822 402498 6004 402734
rect 5404 367054 6004 402498
rect 5404 366818 5586 367054
rect 5822 366818 6004 367054
rect 5404 366734 6004 366818
rect 5404 366498 5586 366734
rect 5822 366498 6004 366734
rect 5404 331054 6004 366498
rect 5404 330818 5586 331054
rect 5822 330818 6004 331054
rect 5404 330734 6004 330818
rect 5404 330498 5586 330734
rect 5822 330498 6004 330734
rect 5404 295054 6004 330498
rect 5404 294818 5586 295054
rect 5822 294818 6004 295054
rect 5404 294734 6004 294818
rect 5404 294498 5586 294734
rect 5822 294498 6004 294734
rect 5404 259054 6004 294498
rect 5404 258818 5586 259054
rect 5822 258818 6004 259054
rect 5404 258734 6004 258818
rect 5404 258498 5586 258734
rect 5822 258498 6004 258734
rect 5404 223054 6004 258498
rect 5404 222818 5586 223054
rect 5822 222818 6004 223054
rect 5404 222734 6004 222818
rect 5404 222498 5586 222734
rect 5822 222498 6004 222734
rect 5404 187054 6004 222498
rect 5404 186818 5586 187054
rect 5822 186818 6004 187054
rect 5404 186734 6004 186818
rect 5404 186498 5586 186734
rect 5822 186498 6004 186734
rect 5404 151054 6004 186498
rect 5404 150818 5586 151054
rect 5822 150818 6004 151054
rect 5404 150734 6004 150818
rect 5404 150498 5586 150734
rect 5822 150498 6004 150734
rect 5404 115054 6004 150498
rect 5404 114818 5586 115054
rect 5822 114818 6004 115054
rect 5404 114734 6004 114818
rect 5404 114498 5586 114734
rect 5822 114498 6004 114734
rect 5404 79054 6004 114498
rect 5404 78818 5586 79054
rect 5822 78818 6004 79054
rect 5404 78734 6004 78818
rect 5404 78498 5586 78734
rect 5822 78498 6004 78734
rect 5404 43054 6004 78498
rect 5404 42818 5586 43054
rect 5822 42818 6004 43054
rect 5404 42734 6004 42818
rect 5404 42498 5586 42734
rect 5822 42498 6004 42734
rect 5404 7054 6004 42498
rect 5404 6818 5586 7054
rect 5822 6818 6004 7054
rect 5404 6734 6004 6818
rect 5404 6498 5586 6734
rect 5822 6498 6004 6734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 5404 -2226 6004 6498
rect 5404 -2462 5586 -2226
rect 5822 -2462 6004 -2226
rect 5404 -2546 6004 -2462
rect 5404 -2782 5586 -2546
rect 5822 -2782 6004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 5404 -3744 6004 -2782
rect 9004 694654 9604 708042
rect 9004 694418 9186 694654
rect 9422 694418 9604 694654
rect 9004 694334 9604 694418
rect 9004 694098 9186 694334
rect 9422 694098 9604 694334
rect 9004 658654 9604 694098
rect 9004 658418 9186 658654
rect 9422 658418 9604 658654
rect 9004 658334 9604 658418
rect 9004 658098 9186 658334
rect 9422 658098 9604 658334
rect 9004 622654 9604 658098
rect 9004 622418 9186 622654
rect 9422 622418 9604 622654
rect 9004 622334 9604 622418
rect 9004 622098 9186 622334
rect 9422 622098 9604 622334
rect 9004 586654 9604 622098
rect 9004 586418 9186 586654
rect 9422 586418 9604 586654
rect 9004 586334 9604 586418
rect 9004 586098 9186 586334
rect 9422 586098 9604 586334
rect 9004 550654 9604 586098
rect 9004 550418 9186 550654
rect 9422 550418 9604 550654
rect 9004 550334 9604 550418
rect 9004 550098 9186 550334
rect 9422 550098 9604 550334
rect 9004 514654 9604 550098
rect 9004 514418 9186 514654
rect 9422 514418 9604 514654
rect 9004 514334 9604 514418
rect 9004 514098 9186 514334
rect 9422 514098 9604 514334
rect 9004 478654 9604 514098
rect 9004 478418 9186 478654
rect 9422 478418 9604 478654
rect 9004 478334 9604 478418
rect 9004 478098 9186 478334
rect 9422 478098 9604 478334
rect 9004 442654 9604 478098
rect 9004 442418 9186 442654
rect 9422 442418 9604 442654
rect 9004 442334 9604 442418
rect 9004 442098 9186 442334
rect 9422 442098 9604 442334
rect 9004 406654 9604 442098
rect 9004 406418 9186 406654
rect 9422 406418 9604 406654
rect 9004 406334 9604 406418
rect 9004 406098 9186 406334
rect 9422 406098 9604 406334
rect 9004 370654 9604 406098
rect 9004 370418 9186 370654
rect 9422 370418 9604 370654
rect 9004 370334 9604 370418
rect 9004 370098 9186 370334
rect 9422 370098 9604 370334
rect 9004 334654 9604 370098
rect 9004 334418 9186 334654
rect 9422 334418 9604 334654
rect 9004 334334 9604 334418
rect 9004 334098 9186 334334
rect 9422 334098 9604 334334
rect 9004 298654 9604 334098
rect 9004 298418 9186 298654
rect 9422 298418 9604 298654
rect 9004 298334 9604 298418
rect 9004 298098 9186 298334
rect 9422 298098 9604 298334
rect 9004 262654 9604 298098
rect 9004 262418 9186 262654
rect 9422 262418 9604 262654
rect 9004 262334 9604 262418
rect 9004 262098 9186 262334
rect 9422 262098 9604 262334
rect 9004 226654 9604 262098
rect 9004 226418 9186 226654
rect 9422 226418 9604 226654
rect 9004 226334 9604 226418
rect 9004 226098 9186 226334
rect 9422 226098 9604 226334
rect 9004 190654 9604 226098
rect 9004 190418 9186 190654
rect 9422 190418 9604 190654
rect 9004 190334 9604 190418
rect 9004 190098 9186 190334
rect 9422 190098 9604 190334
rect 9004 154654 9604 190098
rect 9004 154418 9186 154654
rect 9422 154418 9604 154654
rect 9004 154334 9604 154418
rect 9004 154098 9186 154334
rect 9422 154098 9604 154334
rect 9004 118654 9604 154098
rect 9004 118418 9186 118654
rect 9422 118418 9604 118654
rect 9004 118334 9604 118418
rect 9004 118098 9186 118334
rect 9422 118098 9604 118334
rect 9004 82654 9604 118098
rect 9004 82418 9186 82654
rect 9422 82418 9604 82654
rect 9004 82334 9604 82418
rect 9004 82098 9186 82334
rect 9422 82098 9604 82334
rect 9004 46654 9604 82098
rect 9004 46418 9186 46654
rect 9422 46418 9604 46654
rect 9004 46334 9604 46418
rect 9004 46098 9186 46334
rect 9422 46098 9604 46334
rect 9004 10654 9604 46098
rect 9004 10418 9186 10654
rect 9422 10418 9604 10654
rect 9004 10334 9604 10418
rect 9004 10098 9186 10334
rect 9422 10098 9604 10334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 9004 -4106 9604 10098
rect 9004 -4342 9186 -4106
rect 9422 -4342 9604 -4106
rect 9004 -4426 9604 -4342
rect 9004 -4662 9186 -4426
rect 9422 -4662 9604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 9004 -5624 9604 -4662
rect 12604 698254 13204 709922
rect 30604 711418 31204 711440
rect 30604 711182 30786 711418
rect 31022 711182 31204 711418
rect 30604 711098 31204 711182
rect 30604 710862 30786 711098
rect 31022 710862 31204 711098
rect 27004 709538 27604 709560
rect 27004 709302 27186 709538
rect 27422 709302 27604 709538
rect 27004 709218 27604 709302
rect 27004 708982 27186 709218
rect 27422 708982 27604 709218
rect 23404 707658 24004 707680
rect 23404 707422 23586 707658
rect 23822 707422 24004 707658
rect 23404 707338 24004 707422
rect 23404 707102 23586 707338
rect 23822 707102 24004 707338
rect 12604 698018 12786 698254
rect 13022 698018 13204 698254
rect 12604 697934 13204 698018
rect 12604 697698 12786 697934
rect 13022 697698 13204 697934
rect 12604 662254 13204 697698
rect 12604 662018 12786 662254
rect 13022 662018 13204 662254
rect 12604 661934 13204 662018
rect 12604 661698 12786 661934
rect 13022 661698 13204 661934
rect 12604 626254 13204 661698
rect 12604 626018 12786 626254
rect 13022 626018 13204 626254
rect 12604 625934 13204 626018
rect 12604 625698 12786 625934
rect 13022 625698 13204 625934
rect 12604 590254 13204 625698
rect 12604 590018 12786 590254
rect 13022 590018 13204 590254
rect 12604 589934 13204 590018
rect 12604 589698 12786 589934
rect 13022 589698 13204 589934
rect 12604 554254 13204 589698
rect 12604 554018 12786 554254
rect 13022 554018 13204 554254
rect 12604 553934 13204 554018
rect 12604 553698 12786 553934
rect 13022 553698 13204 553934
rect 12604 518254 13204 553698
rect 12604 518018 12786 518254
rect 13022 518018 13204 518254
rect 12604 517934 13204 518018
rect 12604 517698 12786 517934
rect 13022 517698 13204 517934
rect 12604 482254 13204 517698
rect 12604 482018 12786 482254
rect 13022 482018 13204 482254
rect 12604 481934 13204 482018
rect 12604 481698 12786 481934
rect 13022 481698 13204 481934
rect 12604 446254 13204 481698
rect 12604 446018 12786 446254
rect 13022 446018 13204 446254
rect 12604 445934 13204 446018
rect 12604 445698 12786 445934
rect 13022 445698 13204 445934
rect 12604 410254 13204 445698
rect 12604 410018 12786 410254
rect 13022 410018 13204 410254
rect 12604 409934 13204 410018
rect 12604 409698 12786 409934
rect 13022 409698 13204 409934
rect 12604 374254 13204 409698
rect 12604 374018 12786 374254
rect 13022 374018 13204 374254
rect 12604 373934 13204 374018
rect 12604 373698 12786 373934
rect 13022 373698 13204 373934
rect 12604 338254 13204 373698
rect 12604 338018 12786 338254
rect 13022 338018 13204 338254
rect 12604 337934 13204 338018
rect 12604 337698 12786 337934
rect 13022 337698 13204 337934
rect 12604 302254 13204 337698
rect 12604 302018 12786 302254
rect 13022 302018 13204 302254
rect 12604 301934 13204 302018
rect 12604 301698 12786 301934
rect 13022 301698 13204 301934
rect 12604 266254 13204 301698
rect 12604 266018 12786 266254
rect 13022 266018 13204 266254
rect 12604 265934 13204 266018
rect 12604 265698 12786 265934
rect 13022 265698 13204 265934
rect 12604 230254 13204 265698
rect 12604 230018 12786 230254
rect 13022 230018 13204 230254
rect 12604 229934 13204 230018
rect 12604 229698 12786 229934
rect 13022 229698 13204 229934
rect 12604 194254 13204 229698
rect 12604 194018 12786 194254
rect 13022 194018 13204 194254
rect 12604 193934 13204 194018
rect 12604 193698 12786 193934
rect 13022 193698 13204 193934
rect 12604 158254 13204 193698
rect 12604 158018 12786 158254
rect 13022 158018 13204 158254
rect 12604 157934 13204 158018
rect 12604 157698 12786 157934
rect 13022 157698 13204 157934
rect 12604 122254 13204 157698
rect 12604 122018 12786 122254
rect 13022 122018 13204 122254
rect 12604 121934 13204 122018
rect 12604 121698 12786 121934
rect 13022 121698 13204 121934
rect 12604 86254 13204 121698
rect 12604 86018 12786 86254
rect 13022 86018 13204 86254
rect 12604 85934 13204 86018
rect 12604 85698 12786 85934
rect 13022 85698 13204 85934
rect 12604 50254 13204 85698
rect 12604 50018 12786 50254
rect 13022 50018 13204 50254
rect 12604 49934 13204 50018
rect 12604 49698 12786 49934
rect 13022 49698 13204 49934
rect 12604 14254 13204 49698
rect 12604 14018 12786 14254
rect 13022 14018 13204 14254
rect 12604 13934 13204 14018
rect 12604 13698 12786 13934
rect 13022 13698 13204 13934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 12604 -5986 13204 13698
rect 19804 705778 20404 705800
rect 19804 705542 19986 705778
rect 20222 705542 20404 705778
rect 19804 705458 20404 705542
rect 19804 705222 19986 705458
rect 20222 705222 20404 705458
rect 19804 669454 20404 705222
rect 19804 669218 19986 669454
rect 20222 669218 20404 669454
rect 19804 669134 20404 669218
rect 19804 668898 19986 669134
rect 20222 668898 20404 669134
rect 19804 633454 20404 668898
rect 19804 633218 19986 633454
rect 20222 633218 20404 633454
rect 19804 633134 20404 633218
rect 19804 632898 19986 633134
rect 20222 632898 20404 633134
rect 19804 597454 20404 632898
rect 19804 597218 19986 597454
rect 20222 597218 20404 597454
rect 19804 597134 20404 597218
rect 19804 596898 19986 597134
rect 20222 596898 20404 597134
rect 19804 561454 20404 596898
rect 19804 561218 19986 561454
rect 20222 561218 20404 561454
rect 19804 561134 20404 561218
rect 19804 560898 19986 561134
rect 20222 560898 20404 561134
rect 19804 525454 20404 560898
rect 19804 525218 19986 525454
rect 20222 525218 20404 525454
rect 19804 525134 20404 525218
rect 19804 524898 19986 525134
rect 20222 524898 20404 525134
rect 19804 489454 20404 524898
rect 19804 489218 19986 489454
rect 20222 489218 20404 489454
rect 19804 489134 20404 489218
rect 19804 488898 19986 489134
rect 20222 488898 20404 489134
rect 19804 453454 20404 488898
rect 19804 453218 19986 453454
rect 20222 453218 20404 453454
rect 19804 453134 20404 453218
rect 19804 452898 19986 453134
rect 20222 452898 20404 453134
rect 19804 417454 20404 452898
rect 19804 417218 19986 417454
rect 20222 417218 20404 417454
rect 19804 417134 20404 417218
rect 19804 416898 19986 417134
rect 20222 416898 20404 417134
rect 19804 381454 20404 416898
rect 19804 381218 19986 381454
rect 20222 381218 20404 381454
rect 19804 381134 20404 381218
rect 19804 380898 19986 381134
rect 20222 380898 20404 381134
rect 19804 345454 20404 380898
rect 19804 345218 19986 345454
rect 20222 345218 20404 345454
rect 19804 345134 20404 345218
rect 19804 344898 19986 345134
rect 20222 344898 20404 345134
rect 19804 309454 20404 344898
rect 19804 309218 19986 309454
rect 20222 309218 20404 309454
rect 19804 309134 20404 309218
rect 19804 308898 19986 309134
rect 20222 308898 20404 309134
rect 19804 273454 20404 308898
rect 19804 273218 19986 273454
rect 20222 273218 20404 273454
rect 19804 273134 20404 273218
rect 19804 272898 19986 273134
rect 20222 272898 20404 273134
rect 19804 237454 20404 272898
rect 19804 237218 19986 237454
rect 20222 237218 20404 237454
rect 19804 237134 20404 237218
rect 19804 236898 19986 237134
rect 20222 236898 20404 237134
rect 19804 201454 20404 236898
rect 19804 201218 19986 201454
rect 20222 201218 20404 201454
rect 19804 201134 20404 201218
rect 19804 200898 19986 201134
rect 20222 200898 20404 201134
rect 19804 165454 20404 200898
rect 19804 165218 19986 165454
rect 20222 165218 20404 165454
rect 19804 165134 20404 165218
rect 19804 164898 19986 165134
rect 20222 164898 20404 165134
rect 19804 129454 20404 164898
rect 19804 129218 19986 129454
rect 20222 129218 20404 129454
rect 19804 129134 20404 129218
rect 19804 128898 19986 129134
rect 20222 128898 20404 129134
rect 19804 93454 20404 128898
rect 19804 93218 19986 93454
rect 20222 93218 20404 93454
rect 19804 93134 20404 93218
rect 19804 92898 19986 93134
rect 20222 92898 20404 93134
rect 19804 57454 20404 92898
rect 19804 57218 19986 57454
rect 20222 57218 20404 57454
rect 19804 57134 20404 57218
rect 19804 56898 19986 57134
rect 20222 56898 20404 57134
rect 19804 21454 20404 56898
rect 19804 21218 19986 21454
rect 20222 21218 20404 21454
rect 19804 21134 20404 21218
rect 19804 20898 19986 21134
rect 20222 20898 20404 21134
rect 19804 -1286 20404 20898
rect 19804 -1522 19986 -1286
rect 20222 -1522 20404 -1286
rect 19804 -1606 20404 -1522
rect 19804 -1842 19986 -1606
rect 20222 -1842 20404 -1606
rect 19804 -1864 20404 -1842
rect 23404 673054 24004 707102
rect 23404 672818 23586 673054
rect 23822 672818 24004 673054
rect 23404 672734 24004 672818
rect 23404 672498 23586 672734
rect 23822 672498 24004 672734
rect 23404 637054 24004 672498
rect 23404 636818 23586 637054
rect 23822 636818 24004 637054
rect 23404 636734 24004 636818
rect 23404 636498 23586 636734
rect 23822 636498 24004 636734
rect 23404 601054 24004 636498
rect 23404 600818 23586 601054
rect 23822 600818 24004 601054
rect 23404 600734 24004 600818
rect 23404 600498 23586 600734
rect 23822 600498 24004 600734
rect 23404 565054 24004 600498
rect 23404 564818 23586 565054
rect 23822 564818 24004 565054
rect 23404 564734 24004 564818
rect 23404 564498 23586 564734
rect 23822 564498 24004 564734
rect 23404 529054 24004 564498
rect 23404 528818 23586 529054
rect 23822 528818 24004 529054
rect 23404 528734 24004 528818
rect 23404 528498 23586 528734
rect 23822 528498 24004 528734
rect 23404 493054 24004 528498
rect 23404 492818 23586 493054
rect 23822 492818 24004 493054
rect 23404 492734 24004 492818
rect 23404 492498 23586 492734
rect 23822 492498 24004 492734
rect 23404 457054 24004 492498
rect 23404 456818 23586 457054
rect 23822 456818 24004 457054
rect 23404 456734 24004 456818
rect 23404 456498 23586 456734
rect 23822 456498 24004 456734
rect 23404 421054 24004 456498
rect 23404 420818 23586 421054
rect 23822 420818 24004 421054
rect 23404 420734 24004 420818
rect 23404 420498 23586 420734
rect 23822 420498 24004 420734
rect 23404 385054 24004 420498
rect 23404 384818 23586 385054
rect 23822 384818 24004 385054
rect 23404 384734 24004 384818
rect 23404 384498 23586 384734
rect 23822 384498 24004 384734
rect 23404 349054 24004 384498
rect 23404 348818 23586 349054
rect 23822 348818 24004 349054
rect 23404 348734 24004 348818
rect 23404 348498 23586 348734
rect 23822 348498 24004 348734
rect 23404 313054 24004 348498
rect 23404 312818 23586 313054
rect 23822 312818 24004 313054
rect 23404 312734 24004 312818
rect 23404 312498 23586 312734
rect 23822 312498 24004 312734
rect 23404 277054 24004 312498
rect 23404 276818 23586 277054
rect 23822 276818 24004 277054
rect 23404 276734 24004 276818
rect 23404 276498 23586 276734
rect 23822 276498 24004 276734
rect 23404 241054 24004 276498
rect 23404 240818 23586 241054
rect 23822 240818 24004 241054
rect 23404 240734 24004 240818
rect 23404 240498 23586 240734
rect 23822 240498 24004 240734
rect 23404 205054 24004 240498
rect 23404 204818 23586 205054
rect 23822 204818 24004 205054
rect 23404 204734 24004 204818
rect 23404 204498 23586 204734
rect 23822 204498 24004 204734
rect 23404 169054 24004 204498
rect 23404 168818 23586 169054
rect 23822 168818 24004 169054
rect 23404 168734 24004 168818
rect 23404 168498 23586 168734
rect 23822 168498 24004 168734
rect 23404 133054 24004 168498
rect 23404 132818 23586 133054
rect 23822 132818 24004 133054
rect 23404 132734 24004 132818
rect 23404 132498 23586 132734
rect 23822 132498 24004 132734
rect 23404 97054 24004 132498
rect 23404 96818 23586 97054
rect 23822 96818 24004 97054
rect 23404 96734 24004 96818
rect 23404 96498 23586 96734
rect 23822 96498 24004 96734
rect 23404 61054 24004 96498
rect 23404 60818 23586 61054
rect 23822 60818 24004 61054
rect 23404 60734 24004 60818
rect 23404 60498 23586 60734
rect 23822 60498 24004 60734
rect 23404 25054 24004 60498
rect 23404 24818 23586 25054
rect 23822 24818 24004 25054
rect 23404 24734 24004 24818
rect 23404 24498 23586 24734
rect 23822 24498 24004 24734
rect 23404 -3166 24004 24498
rect 23404 -3402 23586 -3166
rect 23822 -3402 24004 -3166
rect 23404 -3486 24004 -3402
rect 23404 -3722 23586 -3486
rect 23822 -3722 24004 -3486
rect 23404 -3744 24004 -3722
rect 27004 676654 27604 708982
rect 27004 676418 27186 676654
rect 27422 676418 27604 676654
rect 27004 676334 27604 676418
rect 27004 676098 27186 676334
rect 27422 676098 27604 676334
rect 27004 640654 27604 676098
rect 27004 640418 27186 640654
rect 27422 640418 27604 640654
rect 27004 640334 27604 640418
rect 27004 640098 27186 640334
rect 27422 640098 27604 640334
rect 27004 604654 27604 640098
rect 27004 604418 27186 604654
rect 27422 604418 27604 604654
rect 27004 604334 27604 604418
rect 27004 604098 27186 604334
rect 27422 604098 27604 604334
rect 27004 568654 27604 604098
rect 27004 568418 27186 568654
rect 27422 568418 27604 568654
rect 27004 568334 27604 568418
rect 27004 568098 27186 568334
rect 27422 568098 27604 568334
rect 27004 532654 27604 568098
rect 27004 532418 27186 532654
rect 27422 532418 27604 532654
rect 27004 532334 27604 532418
rect 27004 532098 27186 532334
rect 27422 532098 27604 532334
rect 27004 496654 27604 532098
rect 27004 496418 27186 496654
rect 27422 496418 27604 496654
rect 27004 496334 27604 496418
rect 27004 496098 27186 496334
rect 27422 496098 27604 496334
rect 27004 460654 27604 496098
rect 27004 460418 27186 460654
rect 27422 460418 27604 460654
rect 27004 460334 27604 460418
rect 27004 460098 27186 460334
rect 27422 460098 27604 460334
rect 27004 424654 27604 460098
rect 27004 424418 27186 424654
rect 27422 424418 27604 424654
rect 27004 424334 27604 424418
rect 27004 424098 27186 424334
rect 27422 424098 27604 424334
rect 27004 388654 27604 424098
rect 27004 388418 27186 388654
rect 27422 388418 27604 388654
rect 27004 388334 27604 388418
rect 27004 388098 27186 388334
rect 27422 388098 27604 388334
rect 27004 352654 27604 388098
rect 27004 352418 27186 352654
rect 27422 352418 27604 352654
rect 27004 352334 27604 352418
rect 27004 352098 27186 352334
rect 27422 352098 27604 352334
rect 27004 316654 27604 352098
rect 27004 316418 27186 316654
rect 27422 316418 27604 316654
rect 27004 316334 27604 316418
rect 27004 316098 27186 316334
rect 27422 316098 27604 316334
rect 27004 280654 27604 316098
rect 27004 280418 27186 280654
rect 27422 280418 27604 280654
rect 27004 280334 27604 280418
rect 27004 280098 27186 280334
rect 27422 280098 27604 280334
rect 27004 244654 27604 280098
rect 27004 244418 27186 244654
rect 27422 244418 27604 244654
rect 27004 244334 27604 244418
rect 27004 244098 27186 244334
rect 27422 244098 27604 244334
rect 27004 208654 27604 244098
rect 27004 208418 27186 208654
rect 27422 208418 27604 208654
rect 27004 208334 27604 208418
rect 27004 208098 27186 208334
rect 27422 208098 27604 208334
rect 27004 172654 27604 208098
rect 27004 172418 27186 172654
rect 27422 172418 27604 172654
rect 27004 172334 27604 172418
rect 27004 172098 27186 172334
rect 27422 172098 27604 172334
rect 27004 136654 27604 172098
rect 27004 136418 27186 136654
rect 27422 136418 27604 136654
rect 27004 136334 27604 136418
rect 27004 136098 27186 136334
rect 27422 136098 27604 136334
rect 27004 100654 27604 136098
rect 27004 100418 27186 100654
rect 27422 100418 27604 100654
rect 27004 100334 27604 100418
rect 27004 100098 27186 100334
rect 27422 100098 27604 100334
rect 27004 64654 27604 100098
rect 27004 64418 27186 64654
rect 27422 64418 27604 64654
rect 27004 64334 27604 64418
rect 27004 64098 27186 64334
rect 27422 64098 27604 64334
rect 27004 28654 27604 64098
rect 27004 28418 27186 28654
rect 27422 28418 27604 28654
rect 27004 28334 27604 28418
rect 27004 28098 27186 28334
rect 27422 28098 27604 28334
rect 27004 -5046 27604 28098
rect 27004 -5282 27186 -5046
rect 27422 -5282 27604 -5046
rect 27004 -5366 27604 -5282
rect 27004 -5602 27186 -5366
rect 27422 -5602 27604 -5366
rect 27004 -5624 27604 -5602
rect 30604 680254 31204 710862
rect 48604 710478 49204 711440
rect 48604 710242 48786 710478
rect 49022 710242 49204 710478
rect 48604 710158 49204 710242
rect 48604 709922 48786 710158
rect 49022 709922 49204 710158
rect 45004 708598 45604 709560
rect 45004 708362 45186 708598
rect 45422 708362 45604 708598
rect 45004 708278 45604 708362
rect 45004 708042 45186 708278
rect 45422 708042 45604 708278
rect 41404 706718 42004 707680
rect 41404 706482 41586 706718
rect 41822 706482 42004 706718
rect 41404 706398 42004 706482
rect 41404 706162 41586 706398
rect 41822 706162 42004 706398
rect 30604 680018 30786 680254
rect 31022 680018 31204 680254
rect 30604 679934 31204 680018
rect 30604 679698 30786 679934
rect 31022 679698 31204 679934
rect 30604 644254 31204 679698
rect 30604 644018 30786 644254
rect 31022 644018 31204 644254
rect 30604 643934 31204 644018
rect 30604 643698 30786 643934
rect 31022 643698 31204 643934
rect 30604 608254 31204 643698
rect 30604 608018 30786 608254
rect 31022 608018 31204 608254
rect 30604 607934 31204 608018
rect 30604 607698 30786 607934
rect 31022 607698 31204 607934
rect 30604 572254 31204 607698
rect 30604 572018 30786 572254
rect 31022 572018 31204 572254
rect 30604 571934 31204 572018
rect 30604 571698 30786 571934
rect 31022 571698 31204 571934
rect 30604 536254 31204 571698
rect 30604 536018 30786 536254
rect 31022 536018 31204 536254
rect 30604 535934 31204 536018
rect 30604 535698 30786 535934
rect 31022 535698 31204 535934
rect 30604 500254 31204 535698
rect 30604 500018 30786 500254
rect 31022 500018 31204 500254
rect 30604 499934 31204 500018
rect 30604 499698 30786 499934
rect 31022 499698 31204 499934
rect 30604 464254 31204 499698
rect 30604 464018 30786 464254
rect 31022 464018 31204 464254
rect 30604 463934 31204 464018
rect 30604 463698 30786 463934
rect 31022 463698 31204 463934
rect 30604 428254 31204 463698
rect 30604 428018 30786 428254
rect 31022 428018 31204 428254
rect 30604 427934 31204 428018
rect 30604 427698 30786 427934
rect 31022 427698 31204 427934
rect 30604 392254 31204 427698
rect 30604 392018 30786 392254
rect 31022 392018 31204 392254
rect 30604 391934 31204 392018
rect 30604 391698 30786 391934
rect 31022 391698 31204 391934
rect 30604 356254 31204 391698
rect 30604 356018 30786 356254
rect 31022 356018 31204 356254
rect 30604 355934 31204 356018
rect 30604 355698 30786 355934
rect 31022 355698 31204 355934
rect 30604 320254 31204 355698
rect 30604 320018 30786 320254
rect 31022 320018 31204 320254
rect 30604 319934 31204 320018
rect 30604 319698 30786 319934
rect 31022 319698 31204 319934
rect 30604 284254 31204 319698
rect 30604 284018 30786 284254
rect 31022 284018 31204 284254
rect 30604 283934 31204 284018
rect 30604 283698 30786 283934
rect 31022 283698 31204 283934
rect 30604 248254 31204 283698
rect 30604 248018 30786 248254
rect 31022 248018 31204 248254
rect 30604 247934 31204 248018
rect 30604 247698 30786 247934
rect 31022 247698 31204 247934
rect 30604 212254 31204 247698
rect 30604 212018 30786 212254
rect 31022 212018 31204 212254
rect 30604 211934 31204 212018
rect 30604 211698 30786 211934
rect 31022 211698 31204 211934
rect 30604 176254 31204 211698
rect 30604 176018 30786 176254
rect 31022 176018 31204 176254
rect 30604 175934 31204 176018
rect 30604 175698 30786 175934
rect 31022 175698 31204 175934
rect 30604 140254 31204 175698
rect 30604 140018 30786 140254
rect 31022 140018 31204 140254
rect 30604 139934 31204 140018
rect 30604 139698 30786 139934
rect 31022 139698 31204 139934
rect 30604 104254 31204 139698
rect 30604 104018 30786 104254
rect 31022 104018 31204 104254
rect 30604 103934 31204 104018
rect 30604 103698 30786 103934
rect 31022 103698 31204 103934
rect 30604 68254 31204 103698
rect 30604 68018 30786 68254
rect 31022 68018 31204 68254
rect 30604 67934 31204 68018
rect 30604 67698 30786 67934
rect 31022 67698 31204 67934
rect 30604 32254 31204 67698
rect 30604 32018 30786 32254
rect 31022 32018 31204 32254
rect 30604 31934 31204 32018
rect 30604 31698 30786 31934
rect 31022 31698 31204 31934
rect 12604 -6222 12786 -5986
rect 13022 -6222 13204 -5986
rect 12604 -6306 13204 -6222
rect 12604 -6542 12786 -6306
rect 13022 -6542 13204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 12604 -7504 13204 -6542
rect 30604 -6926 31204 31698
rect 37804 704838 38404 705800
rect 37804 704602 37986 704838
rect 38222 704602 38404 704838
rect 37804 704518 38404 704602
rect 37804 704282 37986 704518
rect 38222 704282 38404 704518
rect 37804 687454 38404 704282
rect 37804 687218 37986 687454
rect 38222 687218 38404 687454
rect 37804 687134 38404 687218
rect 37804 686898 37986 687134
rect 38222 686898 38404 687134
rect 37804 651454 38404 686898
rect 37804 651218 37986 651454
rect 38222 651218 38404 651454
rect 37804 651134 38404 651218
rect 37804 650898 37986 651134
rect 38222 650898 38404 651134
rect 37804 615454 38404 650898
rect 37804 615218 37986 615454
rect 38222 615218 38404 615454
rect 37804 615134 38404 615218
rect 37804 614898 37986 615134
rect 38222 614898 38404 615134
rect 37804 579454 38404 614898
rect 37804 579218 37986 579454
rect 38222 579218 38404 579454
rect 37804 579134 38404 579218
rect 37804 578898 37986 579134
rect 38222 578898 38404 579134
rect 37804 543454 38404 578898
rect 37804 543218 37986 543454
rect 38222 543218 38404 543454
rect 37804 543134 38404 543218
rect 37804 542898 37986 543134
rect 38222 542898 38404 543134
rect 37804 507454 38404 542898
rect 37804 507218 37986 507454
rect 38222 507218 38404 507454
rect 37804 507134 38404 507218
rect 37804 506898 37986 507134
rect 38222 506898 38404 507134
rect 37804 471454 38404 506898
rect 37804 471218 37986 471454
rect 38222 471218 38404 471454
rect 37804 471134 38404 471218
rect 37804 470898 37986 471134
rect 38222 470898 38404 471134
rect 37804 435454 38404 470898
rect 37804 435218 37986 435454
rect 38222 435218 38404 435454
rect 37804 435134 38404 435218
rect 37804 434898 37986 435134
rect 38222 434898 38404 435134
rect 37804 399454 38404 434898
rect 37804 399218 37986 399454
rect 38222 399218 38404 399454
rect 37804 399134 38404 399218
rect 37804 398898 37986 399134
rect 38222 398898 38404 399134
rect 37804 363454 38404 398898
rect 37804 363218 37986 363454
rect 38222 363218 38404 363454
rect 37804 363134 38404 363218
rect 37804 362898 37986 363134
rect 38222 362898 38404 363134
rect 37804 327454 38404 362898
rect 37804 327218 37986 327454
rect 38222 327218 38404 327454
rect 37804 327134 38404 327218
rect 37804 326898 37986 327134
rect 38222 326898 38404 327134
rect 37804 291454 38404 326898
rect 37804 291218 37986 291454
rect 38222 291218 38404 291454
rect 37804 291134 38404 291218
rect 37804 290898 37986 291134
rect 38222 290898 38404 291134
rect 37804 255454 38404 290898
rect 37804 255218 37986 255454
rect 38222 255218 38404 255454
rect 37804 255134 38404 255218
rect 37804 254898 37986 255134
rect 38222 254898 38404 255134
rect 37804 219454 38404 254898
rect 37804 219218 37986 219454
rect 38222 219218 38404 219454
rect 37804 219134 38404 219218
rect 37804 218898 37986 219134
rect 38222 218898 38404 219134
rect 37804 183454 38404 218898
rect 37804 183218 37986 183454
rect 38222 183218 38404 183454
rect 37804 183134 38404 183218
rect 37804 182898 37986 183134
rect 38222 182898 38404 183134
rect 37804 147454 38404 182898
rect 37804 147218 37986 147454
rect 38222 147218 38404 147454
rect 37804 147134 38404 147218
rect 37804 146898 37986 147134
rect 38222 146898 38404 147134
rect 37804 111454 38404 146898
rect 37804 111218 37986 111454
rect 38222 111218 38404 111454
rect 37804 111134 38404 111218
rect 37804 110898 37986 111134
rect 38222 110898 38404 111134
rect 37804 75454 38404 110898
rect 37804 75218 37986 75454
rect 38222 75218 38404 75454
rect 37804 75134 38404 75218
rect 37804 74898 37986 75134
rect 38222 74898 38404 75134
rect 37804 39454 38404 74898
rect 37804 39218 37986 39454
rect 38222 39218 38404 39454
rect 37804 39134 38404 39218
rect 37804 38898 37986 39134
rect 38222 38898 38404 39134
rect 37804 3454 38404 38898
rect 37804 3218 37986 3454
rect 38222 3218 38404 3454
rect 37804 3134 38404 3218
rect 37804 2898 37986 3134
rect 38222 2898 38404 3134
rect 37804 -346 38404 2898
rect 37804 -582 37986 -346
rect 38222 -582 38404 -346
rect 37804 -666 38404 -582
rect 37804 -902 37986 -666
rect 38222 -902 38404 -666
rect 37804 -1864 38404 -902
rect 41404 691054 42004 706162
rect 41404 690818 41586 691054
rect 41822 690818 42004 691054
rect 41404 690734 42004 690818
rect 41404 690498 41586 690734
rect 41822 690498 42004 690734
rect 41404 655054 42004 690498
rect 41404 654818 41586 655054
rect 41822 654818 42004 655054
rect 41404 654734 42004 654818
rect 41404 654498 41586 654734
rect 41822 654498 42004 654734
rect 41404 619054 42004 654498
rect 41404 618818 41586 619054
rect 41822 618818 42004 619054
rect 41404 618734 42004 618818
rect 41404 618498 41586 618734
rect 41822 618498 42004 618734
rect 41404 583054 42004 618498
rect 41404 582818 41586 583054
rect 41822 582818 42004 583054
rect 41404 582734 42004 582818
rect 41404 582498 41586 582734
rect 41822 582498 42004 582734
rect 41404 547054 42004 582498
rect 41404 546818 41586 547054
rect 41822 546818 42004 547054
rect 41404 546734 42004 546818
rect 41404 546498 41586 546734
rect 41822 546498 42004 546734
rect 41404 511054 42004 546498
rect 41404 510818 41586 511054
rect 41822 510818 42004 511054
rect 41404 510734 42004 510818
rect 41404 510498 41586 510734
rect 41822 510498 42004 510734
rect 41404 475054 42004 510498
rect 41404 474818 41586 475054
rect 41822 474818 42004 475054
rect 41404 474734 42004 474818
rect 41404 474498 41586 474734
rect 41822 474498 42004 474734
rect 41404 439054 42004 474498
rect 41404 438818 41586 439054
rect 41822 438818 42004 439054
rect 41404 438734 42004 438818
rect 41404 438498 41586 438734
rect 41822 438498 42004 438734
rect 41404 403054 42004 438498
rect 41404 402818 41586 403054
rect 41822 402818 42004 403054
rect 41404 402734 42004 402818
rect 41404 402498 41586 402734
rect 41822 402498 42004 402734
rect 41404 367054 42004 402498
rect 41404 366818 41586 367054
rect 41822 366818 42004 367054
rect 41404 366734 42004 366818
rect 41404 366498 41586 366734
rect 41822 366498 42004 366734
rect 41404 331054 42004 366498
rect 41404 330818 41586 331054
rect 41822 330818 42004 331054
rect 41404 330734 42004 330818
rect 41404 330498 41586 330734
rect 41822 330498 42004 330734
rect 41404 295054 42004 330498
rect 41404 294818 41586 295054
rect 41822 294818 42004 295054
rect 41404 294734 42004 294818
rect 41404 294498 41586 294734
rect 41822 294498 42004 294734
rect 41404 259054 42004 294498
rect 41404 258818 41586 259054
rect 41822 258818 42004 259054
rect 41404 258734 42004 258818
rect 41404 258498 41586 258734
rect 41822 258498 42004 258734
rect 41404 223054 42004 258498
rect 41404 222818 41586 223054
rect 41822 222818 42004 223054
rect 41404 222734 42004 222818
rect 41404 222498 41586 222734
rect 41822 222498 42004 222734
rect 41404 187054 42004 222498
rect 41404 186818 41586 187054
rect 41822 186818 42004 187054
rect 41404 186734 42004 186818
rect 41404 186498 41586 186734
rect 41822 186498 42004 186734
rect 41404 151054 42004 186498
rect 41404 150818 41586 151054
rect 41822 150818 42004 151054
rect 41404 150734 42004 150818
rect 41404 150498 41586 150734
rect 41822 150498 42004 150734
rect 41404 115054 42004 150498
rect 41404 114818 41586 115054
rect 41822 114818 42004 115054
rect 41404 114734 42004 114818
rect 41404 114498 41586 114734
rect 41822 114498 42004 114734
rect 41404 79054 42004 114498
rect 41404 78818 41586 79054
rect 41822 78818 42004 79054
rect 41404 78734 42004 78818
rect 41404 78498 41586 78734
rect 41822 78498 42004 78734
rect 41404 43054 42004 78498
rect 41404 42818 41586 43054
rect 41822 42818 42004 43054
rect 41404 42734 42004 42818
rect 41404 42498 41586 42734
rect 41822 42498 42004 42734
rect 41404 7054 42004 42498
rect 41404 6818 41586 7054
rect 41822 6818 42004 7054
rect 41404 6734 42004 6818
rect 41404 6498 41586 6734
rect 41822 6498 42004 6734
rect 41404 -2226 42004 6498
rect 41404 -2462 41586 -2226
rect 41822 -2462 42004 -2226
rect 41404 -2546 42004 -2462
rect 41404 -2782 41586 -2546
rect 41822 -2782 42004 -2546
rect 41404 -3744 42004 -2782
rect 45004 694654 45604 708042
rect 45004 694418 45186 694654
rect 45422 694418 45604 694654
rect 45004 694334 45604 694418
rect 45004 694098 45186 694334
rect 45422 694098 45604 694334
rect 45004 658654 45604 694098
rect 45004 658418 45186 658654
rect 45422 658418 45604 658654
rect 45004 658334 45604 658418
rect 45004 658098 45186 658334
rect 45422 658098 45604 658334
rect 45004 622654 45604 658098
rect 45004 622418 45186 622654
rect 45422 622418 45604 622654
rect 45004 622334 45604 622418
rect 45004 622098 45186 622334
rect 45422 622098 45604 622334
rect 45004 586654 45604 622098
rect 45004 586418 45186 586654
rect 45422 586418 45604 586654
rect 45004 586334 45604 586418
rect 45004 586098 45186 586334
rect 45422 586098 45604 586334
rect 45004 550654 45604 586098
rect 45004 550418 45186 550654
rect 45422 550418 45604 550654
rect 45004 550334 45604 550418
rect 45004 550098 45186 550334
rect 45422 550098 45604 550334
rect 45004 514654 45604 550098
rect 45004 514418 45186 514654
rect 45422 514418 45604 514654
rect 45004 514334 45604 514418
rect 45004 514098 45186 514334
rect 45422 514098 45604 514334
rect 45004 478654 45604 514098
rect 45004 478418 45186 478654
rect 45422 478418 45604 478654
rect 45004 478334 45604 478418
rect 45004 478098 45186 478334
rect 45422 478098 45604 478334
rect 45004 442654 45604 478098
rect 45004 442418 45186 442654
rect 45422 442418 45604 442654
rect 45004 442334 45604 442418
rect 45004 442098 45186 442334
rect 45422 442098 45604 442334
rect 45004 406654 45604 442098
rect 45004 406418 45186 406654
rect 45422 406418 45604 406654
rect 45004 406334 45604 406418
rect 45004 406098 45186 406334
rect 45422 406098 45604 406334
rect 45004 370654 45604 406098
rect 45004 370418 45186 370654
rect 45422 370418 45604 370654
rect 45004 370334 45604 370418
rect 45004 370098 45186 370334
rect 45422 370098 45604 370334
rect 45004 334654 45604 370098
rect 45004 334418 45186 334654
rect 45422 334418 45604 334654
rect 45004 334334 45604 334418
rect 45004 334098 45186 334334
rect 45422 334098 45604 334334
rect 45004 298654 45604 334098
rect 45004 298418 45186 298654
rect 45422 298418 45604 298654
rect 45004 298334 45604 298418
rect 45004 298098 45186 298334
rect 45422 298098 45604 298334
rect 45004 262654 45604 298098
rect 45004 262418 45186 262654
rect 45422 262418 45604 262654
rect 45004 262334 45604 262418
rect 45004 262098 45186 262334
rect 45422 262098 45604 262334
rect 45004 226654 45604 262098
rect 45004 226418 45186 226654
rect 45422 226418 45604 226654
rect 45004 226334 45604 226418
rect 45004 226098 45186 226334
rect 45422 226098 45604 226334
rect 45004 190654 45604 226098
rect 45004 190418 45186 190654
rect 45422 190418 45604 190654
rect 45004 190334 45604 190418
rect 45004 190098 45186 190334
rect 45422 190098 45604 190334
rect 45004 154654 45604 190098
rect 45004 154418 45186 154654
rect 45422 154418 45604 154654
rect 45004 154334 45604 154418
rect 45004 154098 45186 154334
rect 45422 154098 45604 154334
rect 45004 118654 45604 154098
rect 45004 118418 45186 118654
rect 45422 118418 45604 118654
rect 45004 118334 45604 118418
rect 45004 118098 45186 118334
rect 45422 118098 45604 118334
rect 45004 82654 45604 118098
rect 45004 82418 45186 82654
rect 45422 82418 45604 82654
rect 45004 82334 45604 82418
rect 45004 82098 45186 82334
rect 45422 82098 45604 82334
rect 45004 46654 45604 82098
rect 45004 46418 45186 46654
rect 45422 46418 45604 46654
rect 45004 46334 45604 46418
rect 45004 46098 45186 46334
rect 45422 46098 45604 46334
rect 45004 10654 45604 46098
rect 45004 10418 45186 10654
rect 45422 10418 45604 10654
rect 45004 10334 45604 10418
rect 45004 10098 45186 10334
rect 45422 10098 45604 10334
rect 45004 -4106 45604 10098
rect 45004 -4342 45186 -4106
rect 45422 -4342 45604 -4106
rect 45004 -4426 45604 -4342
rect 45004 -4662 45186 -4426
rect 45422 -4662 45604 -4426
rect 45004 -5624 45604 -4662
rect 48604 698254 49204 709922
rect 66604 711418 67204 711440
rect 66604 711182 66786 711418
rect 67022 711182 67204 711418
rect 66604 711098 67204 711182
rect 66604 710862 66786 711098
rect 67022 710862 67204 711098
rect 63004 709538 63604 709560
rect 63004 709302 63186 709538
rect 63422 709302 63604 709538
rect 63004 709218 63604 709302
rect 63004 708982 63186 709218
rect 63422 708982 63604 709218
rect 59404 707658 60004 707680
rect 59404 707422 59586 707658
rect 59822 707422 60004 707658
rect 59404 707338 60004 707422
rect 59404 707102 59586 707338
rect 59822 707102 60004 707338
rect 48604 698018 48786 698254
rect 49022 698018 49204 698254
rect 48604 697934 49204 698018
rect 48604 697698 48786 697934
rect 49022 697698 49204 697934
rect 48604 662254 49204 697698
rect 48604 662018 48786 662254
rect 49022 662018 49204 662254
rect 48604 661934 49204 662018
rect 48604 661698 48786 661934
rect 49022 661698 49204 661934
rect 48604 626254 49204 661698
rect 48604 626018 48786 626254
rect 49022 626018 49204 626254
rect 48604 625934 49204 626018
rect 48604 625698 48786 625934
rect 49022 625698 49204 625934
rect 48604 590254 49204 625698
rect 48604 590018 48786 590254
rect 49022 590018 49204 590254
rect 48604 589934 49204 590018
rect 48604 589698 48786 589934
rect 49022 589698 49204 589934
rect 48604 554254 49204 589698
rect 48604 554018 48786 554254
rect 49022 554018 49204 554254
rect 48604 553934 49204 554018
rect 48604 553698 48786 553934
rect 49022 553698 49204 553934
rect 48604 518254 49204 553698
rect 48604 518018 48786 518254
rect 49022 518018 49204 518254
rect 48604 517934 49204 518018
rect 48604 517698 48786 517934
rect 49022 517698 49204 517934
rect 48604 482254 49204 517698
rect 48604 482018 48786 482254
rect 49022 482018 49204 482254
rect 48604 481934 49204 482018
rect 48604 481698 48786 481934
rect 49022 481698 49204 481934
rect 48604 446254 49204 481698
rect 48604 446018 48786 446254
rect 49022 446018 49204 446254
rect 48604 445934 49204 446018
rect 48604 445698 48786 445934
rect 49022 445698 49204 445934
rect 48604 410254 49204 445698
rect 48604 410018 48786 410254
rect 49022 410018 49204 410254
rect 48604 409934 49204 410018
rect 48604 409698 48786 409934
rect 49022 409698 49204 409934
rect 48604 374254 49204 409698
rect 48604 374018 48786 374254
rect 49022 374018 49204 374254
rect 48604 373934 49204 374018
rect 48604 373698 48786 373934
rect 49022 373698 49204 373934
rect 48604 338254 49204 373698
rect 48604 338018 48786 338254
rect 49022 338018 49204 338254
rect 48604 337934 49204 338018
rect 48604 337698 48786 337934
rect 49022 337698 49204 337934
rect 48604 302254 49204 337698
rect 48604 302018 48786 302254
rect 49022 302018 49204 302254
rect 48604 301934 49204 302018
rect 48604 301698 48786 301934
rect 49022 301698 49204 301934
rect 48604 266254 49204 301698
rect 48604 266018 48786 266254
rect 49022 266018 49204 266254
rect 48604 265934 49204 266018
rect 48604 265698 48786 265934
rect 49022 265698 49204 265934
rect 48604 230254 49204 265698
rect 48604 230018 48786 230254
rect 49022 230018 49204 230254
rect 48604 229934 49204 230018
rect 48604 229698 48786 229934
rect 49022 229698 49204 229934
rect 48604 194254 49204 229698
rect 48604 194018 48786 194254
rect 49022 194018 49204 194254
rect 48604 193934 49204 194018
rect 48604 193698 48786 193934
rect 49022 193698 49204 193934
rect 48604 158254 49204 193698
rect 48604 158018 48786 158254
rect 49022 158018 49204 158254
rect 48604 157934 49204 158018
rect 48604 157698 48786 157934
rect 49022 157698 49204 157934
rect 48604 122254 49204 157698
rect 48604 122018 48786 122254
rect 49022 122018 49204 122254
rect 48604 121934 49204 122018
rect 48604 121698 48786 121934
rect 49022 121698 49204 121934
rect 48604 86254 49204 121698
rect 48604 86018 48786 86254
rect 49022 86018 49204 86254
rect 48604 85934 49204 86018
rect 48604 85698 48786 85934
rect 49022 85698 49204 85934
rect 48604 50254 49204 85698
rect 48604 50018 48786 50254
rect 49022 50018 49204 50254
rect 48604 49934 49204 50018
rect 48604 49698 48786 49934
rect 49022 49698 49204 49934
rect 48604 14254 49204 49698
rect 48604 14018 48786 14254
rect 49022 14018 49204 14254
rect 48604 13934 49204 14018
rect 48604 13698 48786 13934
rect 49022 13698 49204 13934
rect 30604 -7162 30786 -6926
rect 31022 -7162 31204 -6926
rect 30604 -7246 31204 -7162
rect 30604 -7482 30786 -7246
rect 31022 -7482 31204 -7246
rect 30604 -7504 31204 -7482
rect 48604 -5986 49204 13698
rect 55804 705778 56404 705800
rect 55804 705542 55986 705778
rect 56222 705542 56404 705778
rect 55804 705458 56404 705542
rect 55804 705222 55986 705458
rect 56222 705222 56404 705458
rect 55804 669454 56404 705222
rect 55804 669218 55986 669454
rect 56222 669218 56404 669454
rect 55804 669134 56404 669218
rect 55804 668898 55986 669134
rect 56222 668898 56404 669134
rect 55804 633454 56404 668898
rect 55804 633218 55986 633454
rect 56222 633218 56404 633454
rect 55804 633134 56404 633218
rect 55804 632898 55986 633134
rect 56222 632898 56404 633134
rect 55804 597454 56404 632898
rect 55804 597218 55986 597454
rect 56222 597218 56404 597454
rect 55804 597134 56404 597218
rect 55804 596898 55986 597134
rect 56222 596898 56404 597134
rect 55804 561454 56404 596898
rect 55804 561218 55986 561454
rect 56222 561218 56404 561454
rect 55804 561134 56404 561218
rect 55804 560898 55986 561134
rect 56222 560898 56404 561134
rect 55804 525454 56404 560898
rect 55804 525218 55986 525454
rect 56222 525218 56404 525454
rect 55804 525134 56404 525218
rect 55804 524898 55986 525134
rect 56222 524898 56404 525134
rect 55804 489454 56404 524898
rect 55804 489218 55986 489454
rect 56222 489218 56404 489454
rect 55804 489134 56404 489218
rect 55804 488898 55986 489134
rect 56222 488898 56404 489134
rect 55804 453454 56404 488898
rect 55804 453218 55986 453454
rect 56222 453218 56404 453454
rect 55804 453134 56404 453218
rect 55804 452898 55986 453134
rect 56222 452898 56404 453134
rect 55804 417454 56404 452898
rect 55804 417218 55986 417454
rect 56222 417218 56404 417454
rect 55804 417134 56404 417218
rect 55804 416898 55986 417134
rect 56222 416898 56404 417134
rect 55804 381454 56404 416898
rect 55804 381218 55986 381454
rect 56222 381218 56404 381454
rect 55804 381134 56404 381218
rect 55804 380898 55986 381134
rect 56222 380898 56404 381134
rect 55804 345454 56404 380898
rect 55804 345218 55986 345454
rect 56222 345218 56404 345454
rect 55804 345134 56404 345218
rect 55804 344898 55986 345134
rect 56222 344898 56404 345134
rect 55804 309454 56404 344898
rect 55804 309218 55986 309454
rect 56222 309218 56404 309454
rect 55804 309134 56404 309218
rect 55804 308898 55986 309134
rect 56222 308898 56404 309134
rect 55804 273454 56404 308898
rect 55804 273218 55986 273454
rect 56222 273218 56404 273454
rect 55804 273134 56404 273218
rect 55804 272898 55986 273134
rect 56222 272898 56404 273134
rect 55804 237454 56404 272898
rect 55804 237218 55986 237454
rect 56222 237218 56404 237454
rect 55804 237134 56404 237218
rect 55804 236898 55986 237134
rect 56222 236898 56404 237134
rect 55804 201454 56404 236898
rect 55804 201218 55986 201454
rect 56222 201218 56404 201454
rect 55804 201134 56404 201218
rect 55804 200898 55986 201134
rect 56222 200898 56404 201134
rect 55804 165454 56404 200898
rect 55804 165218 55986 165454
rect 56222 165218 56404 165454
rect 55804 165134 56404 165218
rect 55804 164898 55986 165134
rect 56222 164898 56404 165134
rect 55804 129454 56404 164898
rect 55804 129218 55986 129454
rect 56222 129218 56404 129454
rect 55804 129134 56404 129218
rect 55804 128898 55986 129134
rect 56222 128898 56404 129134
rect 55804 93454 56404 128898
rect 55804 93218 55986 93454
rect 56222 93218 56404 93454
rect 55804 93134 56404 93218
rect 55804 92898 55986 93134
rect 56222 92898 56404 93134
rect 55804 57454 56404 92898
rect 55804 57218 55986 57454
rect 56222 57218 56404 57454
rect 55804 57134 56404 57218
rect 55804 56898 55986 57134
rect 56222 56898 56404 57134
rect 55804 21454 56404 56898
rect 55804 21218 55986 21454
rect 56222 21218 56404 21454
rect 55804 21134 56404 21218
rect 55804 20898 55986 21134
rect 56222 20898 56404 21134
rect 55804 -1286 56404 20898
rect 55804 -1522 55986 -1286
rect 56222 -1522 56404 -1286
rect 55804 -1606 56404 -1522
rect 55804 -1842 55986 -1606
rect 56222 -1842 56404 -1606
rect 55804 -1864 56404 -1842
rect 59404 673054 60004 707102
rect 59404 672818 59586 673054
rect 59822 672818 60004 673054
rect 59404 672734 60004 672818
rect 59404 672498 59586 672734
rect 59822 672498 60004 672734
rect 59404 637054 60004 672498
rect 59404 636818 59586 637054
rect 59822 636818 60004 637054
rect 59404 636734 60004 636818
rect 59404 636498 59586 636734
rect 59822 636498 60004 636734
rect 59404 601054 60004 636498
rect 59404 600818 59586 601054
rect 59822 600818 60004 601054
rect 59404 600734 60004 600818
rect 59404 600498 59586 600734
rect 59822 600498 60004 600734
rect 59404 565054 60004 600498
rect 59404 564818 59586 565054
rect 59822 564818 60004 565054
rect 59404 564734 60004 564818
rect 59404 564498 59586 564734
rect 59822 564498 60004 564734
rect 59404 529054 60004 564498
rect 59404 528818 59586 529054
rect 59822 528818 60004 529054
rect 59404 528734 60004 528818
rect 59404 528498 59586 528734
rect 59822 528498 60004 528734
rect 59404 493054 60004 528498
rect 59404 492818 59586 493054
rect 59822 492818 60004 493054
rect 59404 492734 60004 492818
rect 59404 492498 59586 492734
rect 59822 492498 60004 492734
rect 59404 457054 60004 492498
rect 59404 456818 59586 457054
rect 59822 456818 60004 457054
rect 59404 456734 60004 456818
rect 59404 456498 59586 456734
rect 59822 456498 60004 456734
rect 59404 421054 60004 456498
rect 59404 420818 59586 421054
rect 59822 420818 60004 421054
rect 59404 420734 60004 420818
rect 59404 420498 59586 420734
rect 59822 420498 60004 420734
rect 59404 385054 60004 420498
rect 59404 384818 59586 385054
rect 59822 384818 60004 385054
rect 59404 384734 60004 384818
rect 59404 384498 59586 384734
rect 59822 384498 60004 384734
rect 59404 349054 60004 384498
rect 59404 348818 59586 349054
rect 59822 348818 60004 349054
rect 59404 348734 60004 348818
rect 59404 348498 59586 348734
rect 59822 348498 60004 348734
rect 59404 313054 60004 348498
rect 59404 312818 59586 313054
rect 59822 312818 60004 313054
rect 59404 312734 60004 312818
rect 59404 312498 59586 312734
rect 59822 312498 60004 312734
rect 59404 277054 60004 312498
rect 59404 276818 59586 277054
rect 59822 276818 60004 277054
rect 59404 276734 60004 276818
rect 59404 276498 59586 276734
rect 59822 276498 60004 276734
rect 59404 241054 60004 276498
rect 59404 240818 59586 241054
rect 59822 240818 60004 241054
rect 59404 240734 60004 240818
rect 59404 240498 59586 240734
rect 59822 240498 60004 240734
rect 59404 205054 60004 240498
rect 59404 204818 59586 205054
rect 59822 204818 60004 205054
rect 59404 204734 60004 204818
rect 59404 204498 59586 204734
rect 59822 204498 60004 204734
rect 59404 169054 60004 204498
rect 59404 168818 59586 169054
rect 59822 168818 60004 169054
rect 59404 168734 60004 168818
rect 59404 168498 59586 168734
rect 59822 168498 60004 168734
rect 59404 133054 60004 168498
rect 59404 132818 59586 133054
rect 59822 132818 60004 133054
rect 59404 132734 60004 132818
rect 59404 132498 59586 132734
rect 59822 132498 60004 132734
rect 59404 97054 60004 132498
rect 59404 96818 59586 97054
rect 59822 96818 60004 97054
rect 59404 96734 60004 96818
rect 59404 96498 59586 96734
rect 59822 96498 60004 96734
rect 59404 61054 60004 96498
rect 59404 60818 59586 61054
rect 59822 60818 60004 61054
rect 59404 60734 60004 60818
rect 59404 60498 59586 60734
rect 59822 60498 60004 60734
rect 59404 25054 60004 60498
rect 59404 24818 59586 25054
rect 59822 24818 60004 25054
rect 59404 24734 60004 24818
rect 59404 24498 59586 24734
rect 59822 24498 60004 24734
rect 59404 -3166 60004 24498
rect 59404 -3402 59586 -3166
rect 59822 -3402 60004 -3166
rect 59404 -3486 60004 -3402
rect 59404 -3722 59586 -3486
rect 59822 -3722 60004 -3486
rect 59404 -3744 60004 -3722
rect 63004 676654 63604 708982
rect 63004 676418 63186 676654
rect 63422 676418 63604 676654
rect 63004 676334 63604 676418
rect 63004 676098 63186 676334
rect 63422 676098 63604 676334
rect 63004 640654 63604 676098
rect 63004 640418 63186 640654
rect 63422 640418 63604 640654
rect 63004 640334 63604 640418
rect 63004 640098 63186 640334
rect 63422 640098 63604 640334
rect 63004 604654 63604 640098
rect 63004 604418 63186 604654
rect 63422 604418 63604 604654
rect 63004 604334 63604 604418
rect 63004 604098 63186 604334
rect 63422 604098 63604 604334
rect 63004 568654 63604 604098
rect 63004 568418 63186 568654
rect 63422 568418 63604 568654
rect 63004 568334 63604 568418
rect 63004 568098 63186 568334
rect 63422 568098 63604 568334
rect 63004 532654 63604 568098
rect 63004 532418 63186 532654
rect 63422 532418 63604 532654
rect 63004 532334 63604 532418
rect 63004 532098 63186 532334
rect 63422 532098 63604 532334
rect 63004 496654 63604 532098
rect 63004 496418 63186 496654
rect 63422 496418 63604 496654
rect 63004 496334 63604 496418
rect 63004 496098 63186 496334
rect 63422 496098 63604 496334
rect 63004 460654 63604 496098
rect 63004 460418 63186 460654
rect 63422 460418 63604 460654
rect 63004 460334 63604 460418
rect 63004 460098 63186 460334
rect 63422 460098 63604 460334
rect 63004 424654 63604 460098
rect 63004 424418 63186 424654
rect 63422 424418 63604 424654
rect 63004 424334 63604 424418
rect 63004 424098 63186 424334
rect 63422 424098 63604 424334
rect 63004 388654 63604 424098
rect 63004 388418 63186 388654
rect 63422 388418 63604 388654
rect 63004 388334 63604 388418
rect 63004 388098 63186 388334
rect 63422 388098 63604 388334
rect 63004 352654 63604 388098
rect 63004 352418 63186 352654
rect 63422 352418 63604 352654
rect 63004 352334 63604 352418
rect 63004 352098 63186 352334
rect 63422 352098 63604 352334
rect 63004 316654 63604 352098
rect 63004 316418 63186 316654
rect 63422 316418 63604 316654
rect 63004 316334 63604 316418
rect 63004 316098 63186 316334
rect 63422 316098 63604 316334
rect 63004 280654 63604 316098
rect 63004 280418 63186 280654
rect 63422 280418 63604 280654
rect 63004 280334 63604 280418
rect 63004 280098 63186 280334
rect 63422 280098 63604 280334
rect 63004 244654 63604 280098
rect 63004 244418 63186 244654
rect 63422 244418 63604 244654
rect 63004 244334 63604 244418
rect 63004 244098 63186 244334
rect 63422 244098 63604 244334
rect 63004 208654 63604 244098
rect 63004 208418 63186 208654
rect 63422 208418 63604 208654
rect 63004 208334 63604 208418
rect 63004 208098 63186 208334
rect 63422 208098 63604 208334
rect 63004 172654 63604 208098
rect 63004 172418 63186 172654
rect 63422 172418 63604 172654
rect 63004 172334 63604 172418
rect 63004 172098 63186 172334
rect 63422 172098 63604 172334
rect 63004 136654 63604 172098
rect 63004 136418 63186 136654
rect 63422 136418 63604 136654
rect 63004 136334 63604 136418
rect 63004 136098 63186 136334
rect 63422 136098 63604 136334
rect 63004 100654 63604 136098
rect 63004 100418 63186 100654
rect 63422 100418 63604 100654
rect 63004 100334 63604 100418
rect 63004 100098 63186 100334
rect 63422 100098 63604 100334
rect 63004 64654 63604 100098
rect 63004 64418 63186 64654
rect 63422 64418 63604 64654
rect 63004 64334 63604 64418
rect 63004 64098 63186 64334
rect 63422 64098 63604 64334
rect 63004 28654 63604 64098
rect 63004 28418 63186 28654
rect 63422 28418 63604 28654
rect 63004 28334 63604 28418
rect 63004 28098 63186 28334
rect 63422 28098 63604 28334
rect 63004 -5046 63604 28098
rect 63004 -5282 63186 -5046
rect 63422 -5282 63604 -5046
rect 63004 -5366 63604 -5282
rect 63004 -5602 63186 -5366
rect 63422 -5602 63604 -5366
rect 63004 -5624 63604 -5602
rect 66604 680254 67204 710862
rect 84604 710478 85204 711440
rect 84604 710242 84786 710478
rect 85022 710242 85204 710478
rect 84604 710158 85204 710242
rect 84604 709922 84786 710158
rect 85022 709922 85204 710158
rect 81004 708598 81604 709560
rect 81004 708362 81186 708598
rect 81422 708362 81604 708598
rect 81004 708278 81604 708362
rect 81004 708042 81186 708278
rect 81422 708042 81604 708278
rect 77404 706718 78004 707680
rect 77404 706482 77586 706718
rect 77822 706482 78004 706718
rect 77404 706398 78004 706482
rect 77404 706162 77586 706398
rect 77822 706162 78004 706398
rect 66604 680018 66786 680254
rect 67022 680018 67204 680254
rect 66604 679934 67204 680018
rect 66604 679698 66786 679934
rect 67022 679698 67204 679934
rect 66604 644254 67204 679698
rect 66604 644018 66786 644254
rect 67022 644018 67204 644254
rect 66604 643934 67204 644018
rect 66604 643698 66786 643934
rect 67022 643698 67204 643934
rect 66604 608254 67204 643698
rect 66604 608018 66786 608254
rect 67022 608018 67204 608254
rect 66604 607934 67204 608018
rect 66604 607698 66786 607934
rect 67022 607698 67204 607934
rect 66604 572254 67204 607698
rect 66604 572018 66786 572254
rect 67022 572018 67204 572254
rect 66604 571934 67204 572018
rect 66604 571698 66786 571934
rect 67022 571698 67204 571934
rect 66604 536254 67204 571698
rect 66604 536018 66786 536254
rect 67022 536018 67204 536254
rect 66604 535934 67204 536018
rect 66604 535698 66786 535934
rect 67022 535698 67204 535934
rect 66604 500254 67204 535698
rect 66604 500018 66786 500254
rect 67022 500018 67204 500254
rect 66604 499934 67204 500018
rect 66604 499698 66786 499934
rect 67022 499698 67204 499934
rect 66604 464254 67204 499698
rect 66604 464018 66786 464254
rect 67022 464018 67204 464254
rect 66604 463934 67204 464018
rect 66604 463698 66786 463934
rect 67022 463698 67204 463934
rect 66604 428254 67204 463698
rect 66604 428018 66786 428254
rect 67022 428018 67204 428254
rect 66604 427934 67204 428018
rect 66604 427698 66786 427934
rect 67022 427698 67204 427934
rect 66604 392254 67204 427698
rect 66604 392018 66786 392254
rect 67022 392018 67204 392254
rect 66604 391934 67204 392018
rect 66604 391698 66786 391934
rect 67022 391698 67204 391934
rect 66604 356254 67204 391698
rect 66604 356018 66786 356254
rect 67022 356018 67204 356254
rect 66604 355934 67204 356018
rect 66604 355698 66786 355934
rect 67022 355698 67204 355934
rect 66604 320254 67204 355698
rect 66604 320018 66786 320254
rect 67022 320018 67204 320254
rect 66604 319934 67204 320018
rect 66604 319698 66786 319934
rect 67022 319698 67204 319934
rect 66604 284254 67204 319698
rect 66604 284018 66786 284254
rect 67022 284018 67204 284254
rect 66604 283934 67204 284018
rect 66604 283698 66786 283934
rect 67022 283698 67204 283934
rect 66604 248254 67204 283698
rect 66604 248018 66786 248254
rect 67022 248018 67204 248254
rect 66604 247934 67204 248018
rect 66604 247698 66786 247934
rect 67022 247698 67204 247934
rect 66604 212254 67204 247698
rect 66604 212018 66786 212254
rect 67022 212018 67204 212254
rect 66604 211934 67204 212018
rect 66604 211698 66786 211934
rect 67022 211698 67204 211934
rect 66604 176254 67204 211698
rect 66604 176018 66786 176254
rect 67022 176018 67204 176254
rect 66604 175934 67204 176018
rect 66604 175698 66786 175934
rect 67022 175698 67204 175934
rect 66604 140254 67204 175698
rect 66604 140018 66786 140254
rect 67022 140018 67204 140254
rect 66604 139934 67204 140018
rect 66604 139698 66786 139934
rect 67022 139698 67204 139934
rect 66604 104254 67204 139698
rect 66604 104018 66786 104254
rect 67022 104018 67204 104254
rect 66604 103934 67204 104018
rect 66604 103698 66786 103934
rect 67022 103698 67204 103934
rect 66604 68254 67204 103698
rect 66604 68018 66786 68254
rect 67022 68018 67204 68254
rect 66604 67934 67204 68018
rect 66604 67698 66786 67934
rect 67022 67698 67204 67934
rect 66604 32254 67204 67698
rect 66604 32018 66786 32254
rect 67022 32018 67204 32254
rect 66604 31934 67204 32018
rect 66604 31698 66786 31934
rect 67022 31698 67204 31934
rect 48604 -6222 48786 -5986
rect 49022 -6222 49204 -5986
rect 48604 -6306 49204 -6222
rect 48604 -6542 48786 -6306
rect 49022 -6542 49204 -6306
rect 48604 -7504 49204 -6542
rect 66604 -6926 67204 31698
rect 73804 704838 74404 705800
rect 73804 704602 73986 704838
rect 74222 704602 74404 704838
rect 73804 704518 74404 704602
rect 73804 704282 73986 704518
rect 74222 704282 74404 704518
rect 73804 687454 74404 704282
rect 73804 687218 73986 687454
rect 74222 687218 74404 687454
rect 73804 687134 74404 687218
rect 73804 686898 73986 687134
rect 74222 686898 74404 687134
rect 73804 651454 74404 686898
rect 73804 651218 73986 651454
rect 74222 651218 74404 651454
rect 73804 651134 74404 651218
rect 73804 650898 73986 651134
rect 74222 650898 74404 651134
rect 73804 615454 74404 650898
rect 73804 615218 73986 615454
rect 74222 615218 74404 615454
rect 73804 615134 74404 615218
rect 73804 614898 73986 615134
rect 74222 614898 74404 615134
rect 73804 579454 74404 614898
rect 73804 579218 73986 579454
rect 74222 579218 74404 579454
rect 73804 579134 74404 579218
rect 73804 578898 73986 579134
rect 74222 578898 74404 579134
rect 73804 543454 74404 578898
rect 73804 543218 73986 543454
rect 74222 543218 74404 543454
rect 73804 543134 74404 543218
rect 73804 542898 73986 543134
rect 74222 542898 74404 543134
rect 73804 507454 74404 542898
rect 73804 507218 73986 507454
rect 74222 507218 74404 507454
rect 73804 507134 74404 507218
rect 73804 506898 73986 507134
rect 74222 506898 74404 507134
rect 73804 471454 74404 506898
rect 73804 471218 73986 471454
rect 74222 471218 74404 471454
rect 73804 471134 74404 471218
rect 73804 470898 73986 471134
rect 74222 470898 74404 471134
rect 73804 435454 74404 470898
rect 73804 435218 73986 435454
rect 74222 435218 74404 435454
rect 73804 435134 74404 435218
rect 73804 434898 73986 435134
rect 74222 434898 74404 435134
rect 73804 399454 74404 434898
rect 73804 399218 73986 399454
rect 74222 399218 74404 399454
rect 73804 399134 74404 399218
rect 73804 398898 73986 399134
rect 74222 398898 74404 399134
rect 73804 363454 74404 398898
rect 73804 363218 73986 363454
rect 74222 363218 74404 363454
rect 73804 363134 74404 363218
rect 73804 362898 73986 363134
rect 74222 362898 74404 363134
rect 73804 327454 74404 362898
rect 73804 327218 73986 327454
rect 74222 327218 74404 327454
rect 73804 327134 74404 327218
rect 73804 326898 73986 327134
rect 74222 326898 74404 327134
rect 73804 291454 74404 326898
rect 73804 291218 73986 291454
rect 74222 291218 74404 291454
rect 73804 291134 74404 291218
rect 73804 290898 73986 291134
rect 74222 290898 74404 291134
rect 73804 255454 74404 290898
rect 73804 255218 73986 255454
rect 74222 255218 74404 255454
rect 73804 255134 74404 255218
rect 73804 254898 73986 255134
rect 74222 254898 74404 255134
rect 73804 219454 74404 254898
rect 73804 219218 73986 219454
rect 74222 219218 74404 219454
rect 73804 219134 74404 219218
rect 73804 218898 73986 219134
rect 74222 218898 74404 219134
rect 73804 183454 74404 218898
rect 73804 183218 73986 183454
rect 74222 183218 74404 183454
rect 73804 183134 74404 183218
rect 73804 182898 73986 183134
rect 74222 182898 74404 183134
rect 73804 147454 74404 182898
rect 73804 147218 73986 147454
rect 74222 147218 74404 147454
rect 73804 147134 74404 147218
rect 73804 146898 73986 147134
rect 74222 146898 74404 147134
rect 73804 111454 74404 146898
rect 73804 111218 73986 111454
rect 74222 111218 74404 111454
rect 73804 111134 74404 111218
rect 73804 110898 73986 111134
rect 74222 110898 74404 111134
rect 73804 75454 74404 110898
rect 73804 75218 73986 75454
rect 74222 75218 74404 75454
rect 73804 75134 74404 75218
rect 73804 74898 73986 75134
rect 74222 74898 74404 75134
rect 73804 39454 74404 74898
rect 73804 39218 73986 39454
rect 74222 39218 74404 39454
rect 73804 39134 74404 39218
rect 73804 38898 73986 39134
rect 74222 38898 74404 39134
rect 73804 3454 74404 38898
rect 73804 3218 73986 3454
rect 74222 3218 74404 3454
rect 73804 3134 74404 3218
rect 73804 2898 73986 3134
rect 74222 2898 74404 3134
rect 73804 -346 74404 2898
rect 73804 -582 73986 -346
rect 74222 -582 74404 -346
rect 73804 -666 74404 -582
rect 73804 -902 73986 -666
rect 74222 -902 74404 -666
rect 73804 -1864 74404 -902
rect 77404 691054 78004 706162
rect 77404 690818 77586 691054
rect 77822 690818 78004 691054
rect 77404 690734 78004 690818
rect 77404 690498 77586 690734
rect 77822 690498 78004 690734
rect 77404 655054 78004 690498
rect 77404 654818 77586 655054
rect 77822 654818 78004 655054
rect 77404 654734 78004 654818
rect 77404 654498 77586 654734
rect 77822 654498 78004 654734
rect 77404 619054 78004 654498
rect 77404 618818 77586 619054
rect 77822 618818 78004 619054
rect 77404 618734 78004 618818
rect 77404 618498 77586 618734
rect 77822 618498 78004 618734
rect 77404 583054 78004 618498
rect 77404 582818 77586 583054
rect 77822 582818 78004 583054
rect 77404 582734 78004 582818
rect 77404 582498 77586 582734
rect 77822 582498 78004 582734
rect 77404 547054 78004 582498
rect 77404 546818 77586 547054
rect 77822 546818 78004 547054
rect 77404 546734 78004 546818
rect 77404 546498 77586 546734
rect 77822 546498 78004 546734
rect 77404 511054 78004 546498
rect 77404 510818 77586 511054
rect 77822 510818 78004 511054
rect 77404 510734 78004 510818
rect 77404 510498 77586 510734
rect 77822 510498 78004 510734
rect 77404 475054 78004 510498
rect 77404 474818 77586 475054
rect 77822 474818 78004 475054
rect 77404 474734 78004 474818
rect 77404 474498 77586 474734
rect 77822 474498 78004 474734
rect 77404 439054 78004 474498
rect 77404 438818 77586 439054
rect 77822 438818 78004 439054
rect 77404 438734 78004 438818
rect 77404 438498 77586 438734
rect 77822 438498 78004 438734
rect 77404 403054 78004 438498
rect 77404 402818 77586 403054
rect 77822 402818 78004 403054
rect 77404 402734 78004 402818
rect 77404 402498 77586 402734
rect 77822 402498 78004 402734
rect 77404 367054 78004 402498
rect 77404 366818 77586 367054
rect 77822 366818 78004 367054
rect 77404 366734 78004 366818
rect 77404 366498 77586 366734
rect 77822 366498 78004 366734
rect 77404 331054 78004 366498
rect 77404 330818 77586 331054
rect 77822 330818 78004 331054
rect 77404 330734 78004 330818
rect 77404 330498 77586 330734
rect 77822 330498 78004 330734
rect 77404 295054 78004 330498
rect 77404 294818 77586 295054
rect 77822 294818 78004 295054
rect 77404 294734 78004 294818
rect 77404 294498 77586 294734
rect 77822 294498 78004 294734
rect 77404 259054 78004 294498
rect 77404 258818 77586 259054
rect 77822 258818 78004 259054
rect 77404 258734 78004 258818
rect 77404 258498 77586 258734
rect 77822 258498 78004 258734
rect 77404 223054 78004 258498
rect 77404 222818 77586 223054
rect 77822 222818 78004 223054
rect 77404 222734 78004 222818
rect 77404 222498 77586 222734
rect 77822 222498 78004 222734
rect 77404 187054 78004 222498
rect 77404 186818 77586 187054
rect 77822 186818 78004 187054
rect 77404 186734 78004 186818
rect 77404 186498 77586 186734
rect 77822 186498 78004 186734
rect 77404 151054 78004 186498
rect 77404 150818 77586 151054
rect 77822 150818 78004 151054
rect 77404 150734 78004 150818
rect 77404 150498 77586 150734
rect 77822 150498 78004 150734
rect 77404 115054 78004 150498
rect 77404 114818 77586 115054
rect 77822 114818 78004 115054
rect 77404 114734 78004 114818
rect 77404 114498 77586 114734
rect 77822 114498 78004 114734
rect 77404 79054 78004 114498
rect 77404 78818 77586 79054
rect 77822 78818 78004 79054
rect 77404 78734 78004 78818
rect 77404 78498 77586 78734
rect 77822 78498 78004 78734
rect 77404 43054 78004 78498
rect 77404 42818 77586 43054
rect 77822 42818 78004 43054
rect 77404 42734 78004 42818
rect 77404 42498 77586 42734
rect 77822 42498 78004 42734
rect 77404 7054 78004 42498
rect 77404 6818 77586 7054
rect 77822 6818 78004 7054
rect 77404 6734 78004 6818
rect 77404 6498 77586 6734
rect 77822 6498 78004 6734
rect 77404 -2226 78004 6498
rect 77404 -2462 77586 -2226
rect 77822 -2462 78004 -2226
rect 77404 -2546 78004 -2462
rect 77404 -2782 77586 -2546
rect 77822 -2782 78004 -2546
rect 77404 -3744 78004 -2782
rect 81004 694654 81604 708042
rect 81004 694418 81186 694654
rect 81422 694418 81604 694654
rect 81004 694334 81604 694418
rect 81004 694098 81186 694334
rect 81422 694098 81604 694334
rect 81004 658654 81604 694098
rect 81004 658418 81186 658654
rect 81422 658418 81604 658654
rect 81004 658334 81604 658418
rect 81004 658098 81186 658334
rect 81422 658098 81604 658334
rect 81004 622654 81604 658098
rect 81004 622418 81186 622654
rect 81422 622418 81604 622654
rect 81004 622334 81604 622418
rect 81004 622098 81186 622334
rect 81422 622098 81604 622334
rect 81004 586654 81604 622098
rect 81004 586418 81186 586654
rect 81422 586418 81604 586654
rect 81004 586334 81604 586418
rect 81004 586098 81186 586334
rect 81422 586098 81604 586334
rect 81004 550654 81604 586098
rect 81004 550418 81186 550654
rect 81422 550418 81604 550654
rect 81004 550334 81604 550418
rect 81004 550098 81186 550334
rect 81422 550098 81604 550334
rect 81004 514654 81604 550098
rect 81004 514418 81186 514654
rect 81422 514418 81604 514654
rect 81004 514334 81604 514418
rect 81004 514098 81186 514334
rect 81422 514098 81604 514334
rect 81004 478654 81604 514098
rect 81004 478418 81186 478654
rect 81422 478418 81604 478654
rect 81004 478334 81604 478418
rect 81004 478098 81186 478334
rect 81422 478098 81604 478334
rect 81004 442654 81604 478098
rect 81004 442418 81186 442654
rect 81422 442418 81604 442654
rect 81004 442334 81604 442418
rect 81004 442098 81186 442334
rect 81422 442098 81604 442334
rect 81004 406654 81604 442098
rect 81004 406418 81186 406654
rect 81422 406418 81604 406654
rect 81004 406334 81604 406418
rect 81004 406098 81186 406334
rect 81422 406098 81604 406334
rect 81004 370654 81604 406098
rect 81004 370418 81186 370654
rect 81422 370418 81604 370654
rect 81004 370334 81604 370418
rect 81004 370098 81186 370334
rect 81422 370098 81604 370334
rect 81004 334654 81604 370098
rect 81004 334418 81186 334654
rect 81422 334418 81604 334654
rect 81004 334334 81604 334418
rect 81004 334098 81186 334334
rect 81422 334098 81604 334334
rect 81004 298654 81604 334098
rect 81004 298418 81186 298654
rect 81422 298418 81604 298654
rect 81004 298334 81604 298418
rect 81004 298098 81186 298334
rect 81422 298098 81604 298334
rect 81004 262654 81604 298098
rect 81004 262418 81186 262654
rect 81422 262418 81604 262654
rect 81004 262334 81604 262418
rect 81004 262098 81186 262334
rect 81422 262098 81604 262334
rect 81004 226654 81604 262098
rect 81004 226418 81186 226654
rect 81422 226418 81604 226654
rect 81004 226334 81604 226418
rect 81004 226098 81186 226334
rect 81422 226098 81604 226334
rect 81004 190654 81604 226098
rect 81004 190418 81186 190654
rect 81422 190418 81604 190654
rect 81004 190334 81604 190418
rect 81004 190098 81186 190334
rect 81422 190098 81604 190334
rect 81004 154654 81604 190098
rect 81004 154418 81186 154654
rect 81422 154418 81604 154654
rect 81004 154334 81604 154418
rect 81004 154098 81186 154334
rect 81422 154098 81604 154334
rect 81004 118654 81604 154098
rect 81004 118418 81186 118654
rect 81422 118418 81604 118654
rect 81004 118334 81604 118418
rect 81004 118098 81186 118334
rect 81422 118098 81604 118334
rect 81004 82654 81604 118098
rect 81004 82418 81186 82654
rect 81422 82418 81604 82654
rect 81004 82334 81604 82418
rect 81004 82098 81186 82334
rect 81422 82098 81604 82334
rect 81004 46654 81604 82098
rect 81004 46418 81186 46654
rect 81422 46418 81604 46654
rect 81004 46334 81604 46418
rect 81004 46098 81186 46334
rect 81422 46098 81604 46334
rect 81004 10654 81604 46098
rect 81004 10418 81186 10654
rect 81422 10418 81604 10654
rect 81004 10334 81604 10418
rect 81004 10098 81186 10334
rect 81422 10098 81604 10334
rect 81004 -4106 81604 10098
rect 81004 -4342 81186 -4106
rect 81422 -4342 81604 -4106
rect 81004 -4426 81604 -4342
rect 81004 -4662 81186 -4426
rect 81422 -4662 81604 -4426
rect 81004 -5624 81604 -4662
rect 84604 698254 85204 709922
rect 102604 711418 103204 711440
rect 102604 711182 102786 711418
rect 103022 711182 103204 711418
rect 102604 711098 103204 711182
rect 102604 710862 102786 711098
rect 103022 710862 103204 711098
rect 99004 709538 99604 709560
rect 99004 709302 99186 709538
rect 99422 709302 99604 709538
rect 99004 709218 99604 709302
rect 99004 708982 99186 709218
rect 99422 708982 99604 709218
rect 95404 707658 96004 707680
rect 95404 707422 95586 707658
rect 95822 707422 96004 707658
rect 95404 707338 96004 707422
rect 95404 707102 95586 707338
rect 95822 707102 96004 707338
rect 84604 698018 84786 698254
rect 85022 698018 85204 698254
rect 84604 697934 85204 698018
rect 84604 697698 84786 697934
rect 85022 697698 85204 697934
rect 84604 662254 85204 697698
rect 84604 662018 84786 662254
rect 85022 662018 85204 662254
rect 84604 661934 85204 662018
rect 84604 661698 84786 661934
rect 85022 661698 85204 661934
rect 84604 626254 85204 661698
rect 84604 626018 84786 626254
rect 85022 626018 85204 626254
rect 84604 625934 85204 626018
rect 84604 625698 84786 625934
rect 85022 625698 85204 625934
rect 84604 590254 85204 625698
rect 84604 590018 84786 590254
rect 85022 590018 85204 590254
rect 84604 589934 85204 590018
rect 84604 589698 84786 589934
rect 85022 589698 85204 589934
rect 84604 554254 85204 589698
rect 84604 554018 84786 554254
rect 85022 554018 85204 554254
rect 84604 553934 85204 554018
rect 84604 553698 84786 553934
rect 85022 553698 85204 553934
rect 84604 518254 85204 553698
rect 84604 518018 84786 518254
rect 85022 518018 85204 518254
rect 84604 517934 85204 518018
rect 84604 517698 84786 517934
rect 85022 517698 85204 517934
rect 84604 482254 85204 517698
rect 84604 482018 84786 482254
rect 85022 482018 85204 482254
rect 84604 481934 85204 482018
rect 84604 481698 84786 481934
rect 85022 481698 85204 481934
rect 84604 446254 85204 481698
rect 84604 446018 84786 446254
rect 85022 446018 85204 446254
rect 84604 445934 85204 446018
rect 84604 445698 84786 445934
rect 85022 445698 85204 445934
rect 84604 410254 85204 445698
rect 84604 410018 84786 410254
rect 85022 410018 85204 410254
rect 84604 409934 85204 410018
rect 84604 409698 84786 409934
rect 85022 409698 85204 409934
rect 84604 374254 85204 409698
rect 84604 374018 84786 374254
rect 85022 374018 85204 374254
rect 84604 373934 85204 374018
rect 84604 373698 84786 373934
rect 85022 373698 85204 373934
rect 84604 338254 85204 373698
rect 84604 338018 84786 338254
rect 85022 338018 85204 338254
rect 84604 337934 85204 338018
rect 84604 337698 84786 337934
rect 85022 337698 85204 337934
rect 84604 302254 85204 337698
rect 84604 302018 84786 302254
rect 85022 302018 85204 302254
rect 84604 301934 85204 302018
rect 84604 301698 84786 301934
rect 85022 301698 85204 301934
rect 84604 266254 85204 301698
rect 84604 266018 84786 266254
rect 85022 266018 85204 266254
rect 84604 265934 85204 266018
rect 84604 265698 84786 265934
rect 85022 265698 85204 265934
rect 84604 230254 85204 265698
rect 84604 230018 84786 230254
rect 85022 230018 85204 230254
rect 84604 229934 85204 230018
rect 84604 229698 84786 229934
rect 85022 229698 85204 229934
rect 84604 194254 85204 229698
rect 84604 194018 84786 194254
rect 85022 194018 85204 194254
rect 84604 193934 85204 194018
rect 84604 193698 84786 193934
rect 85022 193698 85204 193934
rect 84604 158254 85204 193698
rect 84604 158018 84786 158254
rect 85022 158018 85204 158254
rect 84604 157934 85204 158018
rect 84604 157698 84786 157934
rect 85022 157698 85204 157934
rect 84604 122254 85204 157698
rect 84604 122018 84786 122254
rect 85022 122018 85204 122254
rect 84604 121934 85204 122018
rect 84604 121698 84786 121934
rect 85022 121698 85204 121934
rect 84604 86254 85204 121698
rect 84604 86018 84786 86254
rect 85022 86018 85204 86254
rect 84604 85934 85204 86018
rect 84604 85698 84786 85934
rect 85022 85698 85204 85934
rect 84604 50254 85204 85698
rect 84604 50018 84786 50254
rect 85022 50018 85204 50254
rect 84604 49934 85204 50018
rect 84604 49698 84786 49934
rect 85022 49698 85204 49934
rect 84604 14254 85204 49698
rect 84604 14018 84786 14254
rect 85022 14018 85204 14254
rect 84604 13934 85204 14018
rect 84604 13698 84786 13934
rect 85022 13698 85204 13934
rect 66604 -7162 66786 -6926
rect 67022 -7162 67204 -6926
rect 66604 -7246 67204 -7162
rect 66604 -7482 66786 -7246
rect 67022 -7482 67204 -7246
rect 66604 -7504 67204 -7482
rect 84604 -5986 85204 13698
rect 91804 705778 92404 705800
rect 91804 705542 91986 705778
rect 92222 705542 92404 705778
rect 91804 705458 92404 705542
rect 91804 705222 91986 705458
rect 92222 705222 92404 705458
rect 91804 669454 92404 705222
rect 91804 669218 91986 669454
rect 92222 669218 92404 669454
rect 91804 669134 92404 669218
rect 91804 668898 91986 669134
rect 92222 668898 92404 669134
rect 91804 633454 92404 668898
rect 91804 633218 91986 633454
rect 92222 633218 92404 633454
rect 91804 633134 92404 633218
rect 91804 632898 91986 633134
rect 92222 632898 92404 633134
rect 91804 597454 92404 632898
rect 91804 597218 91986 597454
rect 92222 597218 92404 597454
rect 91804 597134 92404 597218
rect 91804 596898 91986 597134
rect 92222 596898 92404 597134
rect 91804 561454 92404 596898
rect 91804 561218 91986 561454
rect 92222 561218 92404 561454
rect 91804 561134 92404 561218
rect 91804 560898 91986 561134
rect 92222 560898 92404 561134
rect 91804 525454 92404 560898
rect 91804 525218 91986 525454
rect 92222 525218 92404 525454
rect 91804 525134 92404 525218
rect 91804 524898 91986 525134
rect 92222 524898 92404 525134
rect 91804 489454 92404 524898
rect 91804 489218 91986 489454
rect 92222 489218 92404 489454
rect 91804 489134 92404 489218
rect 91804 488898 91986 489134
rect 92222 488898 92404 489134
rect 91804 453454 92404 488898
rect 91804 453218 91986 453454
rect 92222 453218 92404 453454
rect 91804 453134 92404 453218
rect 91804 452898 91986 453134
rect 92222 452898 92404 453134
rect 91804 417454 92404 452898
rect 91804 417218 91986 417454
rect 92222 417218 92404 417454
rect 91804 417134 92404 417218
rect 91804 416898 91986 417134
rect 92222 416898 92404 417134
rect 91804 381454 92404 416898
rect 91804 381218 91986 381454
rect 92222 381218 92404 381454
rect 91804 381134 92404 381218
rect 91804 380898 91986 381134
rect 92222 380898 92404 381134
rect 91804 345454 92404 380898
rect 91804 345218 91986 345454
rect 92222 345218 92404 345454
rect 91804 345134 92404 345218
rect 91804 344898 91986 345134
rect 92222 344898 92404 345134
rect 91804 309454 92404 344898
rect 91804 309218 91986 309454
rect 92222 309218 92404 309454
rect 91804 309134 92404 309218
rect 91804 308898 91986 309134
rect 92222 308898 92404 309134
rect 91804 273454 92404 308898
rect 91804 273218 91986 273454
rect 92222 273218 92404 273454
rect 91804 273134 92404 273218
rect 91804 272898 91986 273134
rect 92222 272898 92404 273134
rect 91804 237454 92404 272898
rect 91804 237218 91986 237454
rect 92222 237218 92404 237454
rect 91804 237134 92404 237218
rect 91804 236898 91986 237134
rect 92222 236898 92404 237134
rect 91804 201454 92404 236898
rect 91804 201218 91986 201454
rect 92222 201218 92404 201454
rect 91804 201134 92404 201218
rect 91804 200898 91986 201134
rect 92222 200898 92404 201134
rect 91804 165454 92404 200898
rect 91804 165218 91986 165454
rect 92222 165218 92404 165454
rect 91804 165134 92404 165218
rect 91804 164898 91986 165134
rect 92222 164898 92404 165134
rect 91804 129454 92404 164898
rect 91804 129218 91986 129454
rect 92222 129218 92404 129454
rect 91804 129134 92404 129218
rect 91804 128898 91986 129134
rect 92222 128898 92404 129134
rect 91804 93454 92404 128898
rect 91804 93218 91986 93454
rect 92222 93218 92404 93454
rect 91804 93134 92404 93218
rect 91804 92898 91986 93134
rect 92222 92898 92404 93134
rect 91804 57454 92404 92898
rect 91804 57218 91986 57454
rect 92222 57218 92404 57454
rect 91804 57134 92404 57218
rect 91804 56898 91986 57134
rect 92222 56898 92404 57134
rect 91804 21454 92404 56898
rect 91804 21218 91986 21454
rect 92222 21218 92404 21454
rect 91804 21134 92404 21218
rect 91804 20898 91986 21134
rect 92222 20898 92404 21134
rect 91804 -1286 92404 20898
rect 91804 -1522 91986 -1286
rect 92222 -1522 92404 -1286
rect 91804 -1606 92404 -1522
rect 91804 -1842 91986 -1606
rect 92222 -1842 92404 -1606
rect 91804 -1864 92404 -1842
rect 95404 673054 96004 707102
rect 95404 672818 95586 673054
rect 95822 672818 96004 673054
rect 95404 672734 96004 672818
rect 95404 672498 95586 672734
rect 95822 672498 96004 672734
rect 95404 637054 96004 672498
rect 95404 636818 95586 637054
rect 95822 636818 96004 637054
rect 95404 636734 96004 636818
rect 95404 636498 95586 636734
rect 95822 636498 96004 636734
rect 95404 601054 96004 636498
rect 95404 600818 95586 601054
rect 95822 600818 96004 601054
rect 95404 600734 96004 600818
rect 95404 600498 95586 600734
rect 95822 600498 96004 600734
rect 95404 565054 96004 600498
rect 95404 564818 95586 565054
rect 95822 564818 96004 565054
rect 95404 564734 96004 564818
rect 95404 564498 95586 564734
rect 95822 564498 96004 564734
rect 95404 529054 96004 564498
rect 95404 528818 95586 529054
rect 95822 528818 96004 529054
rect 95404 528734 96004 528818
rect 95404 528498 95586 528734
rect 95822 528498 96004 528734
rect 95404 493054 96004 528498
rect 95404 492818 95586 493054
rect 95822 492818 96004 493054
rect 95404 492734 96004 492818
rect 95404 492498 95586 492734
rect 95822 492498 96004 492734
rect 95404 457054 96004 492498
rect 95404 456818 95586 457054
rect 95822 456818 96004 457054
rect 95404 456734 96004 456818
rect 95404 456498 95586 456734
rect 95822 456498 96004 456734
rect 95404 421054 96004 456498
rect 95404 420818 95586 421054
rect 95822 420818 96004 421054
rect 95404 420734 96004 420818
rect 95404 420498 95586 420734
rect 95822 420498 96004 420734
rect 95404 385054 96004 420498
rect 95404 384818 95586 385054
rect 95822 384818 96004 385054
rect 95404 384734 96004 384818
rect 95404 384498 95586 384734
rect 95822 384498 96004 384734
rect 95404 349054 96004 384498
rect 95404 348818 95586 349054
rect 95822 348818 96004 349054
rect 95404 348734 96004 348818
rect 95404 348498 95586 348734
rect 95822 348498 96004 348734
rect 95404 313054 96004 348498
rect 95404 312818 95586 313054
rect 95822 312818 96004 313054
rect 95404 312734 96004 312818
rect 95404 312498 95586 312734
rect 95822 312498 96004 312734
rect 95404 277054 96004 312498
rect 95404 276818 95586 277054
rect 95822 276818 96004 277054
rect 95404 276734 96004 276818
rect 95404 276498 95586 276734
rect 95822 276498 96004 276734
rect 95404 241054 96004 276498
rect 95404 240818 95586 241054
rect 95822 240818 96004 241054
rect 95404 240734 96004 240818
rect 95404 240498 95586 240734
rect 95822 240498 96004 240734
rect 95404 205054 96004 240498
rect 95404 204818 95586 205054
rect 95822 204818 96004 205054
rect 95404 204734 96004 204818
rect 95404 204498 95586 204734
rect 95822 204498 96004 204734
rect 95404 169054 96004 204498
rect 95404 168818 95586 169054
rect 95822 168818 96004 169054
rect 95404 168734 96004 168818
rect 95404 168498 95586 168734
rect 95822 168498 96004 168734
rect 95404 133054 96004 168498
rect 95404 132818 95586 133054
rect 95822 132818 96004 133054
rect 95404 132734 96004 132818
rect 95404 132498 95586 132734
rect 95822 132498 96004 132734
rect 95404 97054 96004 132498
rect 95404 96818 95586 97054
rect 95822 96818 96004 97054
rect 95404 96734 96004 96818
rect 95404 96498 95586 96734
rect 95822 96498 96004 96734
rect 95404 61054 96004 96498
rect 95404 60818 95586 61054
rect 95822 60818 96004 61054
rect 95404 60734 96004 60818
rect 95404 60498 95586 60734
rect 95822 60498 96004 60734
rect 95404 25054 96004 60498
rect 95404 24818 95586 25054
rect 95822 24818 96004 25054
rect 95404 24734 96004 24818
rect 95404 24498 95586 24734
rect 95822 24498 96004 24734
rect 95404 -3166 96004 24498
rect 95404 -3402 95586 -3166
rect 95822 -3402 96004 -3166
rect 95404 -3486 96004 -3402
rect 95404 -3722 95586 -3486
rect 95822 -3722 96004 -3486
rect 95404 -3744 96004 -3722
rect 99004 676654 99604 708982
rect 99004 676418 99186 676654
rect 99422 676418 99604 676654
rect 99004 676334 99604 676418
rect 99004 676098 99186 676334
rect 99422 676098 99604 676334
rect 99004 640654 99604 676098
rect 99004 640418 99186 640654
rect 99422 640418 99604 640654
rect 99004 640334 99604 640418
rect 99004 640098 99186 640334
rect 99422 640098 99604 640334
rect 99004 604654 99604 640098
rect 99004 604418 99186 604654
rect 99422 604418 99604 604654
rect 99004 604334 99604 604418
rect 99004 604098 99186 604334
rect 99422 604098 99604 604334
rect 99004 568654 99604 604098
rect 99004 568418 99186 568654
rect 99422 568418 99604 568654
rect 99004 568334 99604 568418
rect 99004 568098 99186 568334
rect 99422 568098 99604 568334
rect 99004 532654 99604 568098
rect 99004 532418 99186 532654
rect 99422 532418 99604 532654
rect 99004 532334 99604 532418
rect 99004 532098 99186 532334
rect 99422 532098 99604 532334
rect 99004 496654 99604 532098
rect 99004 496418 99186 496654
rect 99422 496418 99604 496654
rect 99004 496334 99604 496418
rect 99004 496098 99186 496334
rect 99422 496098 99604 496334
rect 99004 460654 99604 496098
rect 99004 460418 99186 460654
rect 99422 460418 99604 460654
rect 99004 460334 99604 460418
rect 99004 460098 99186 460334
rect 99422 460098 99604 460334
rect 99004 424654 99604 460098
rect 99004 424418 99186 424654
rect 99422 424418 99604 424654
rect 99004 424334 99604 424418
rect 99004 424098 99186 424334
rect 99422 424098 99604 424334
rect 99004 388654 99604 424098
rect 99004 388418 99186 388654
rect 99422 388418 99604 388654
rect 99004 388334 99604 388418
rect 99004 388098 99186 388334
rect 99422 388098 99604 388334
rect 99004 352654 99604 388098
rect 99004 352418 99186 352654
rect 99422 352418 99604 352654
rect 99004 352334 99604 352418
rect 99004 352098 99186 352334
rect 99422 352098 99604 352334
rect 99004 316654 99604 352098
rect 99004 316418 99186 316654
rect 99422 316418 99604 316654
rect 99004 316334 99604 316418
rect 99004 316098 99186 316334
rect 99422 316098 99604 316334
rect 99004 280654 99604 316098
rect 99004 280418 99186 280654
rect 99422 280418 99604 280654
rect 99004 280334 99604 280418
rect 99004 280098 99186 280334
rect 99422 280098 99604 280334
rect 99004 244654 99604 280098
rect 99004 244418 99186 244654
rect 99422 244418 99604 244654
rect 99004 244334 99604 244418
rect 99004 244098 99186 244334
rect 99422 244098 99604 244334
rect 99004 208654 99604 244098
rect 99004 208418 99186 208654
rect 99422 208418 99604 208654
rect 99004 208334 99604 208418
rect 99004 208098 99186 208334
rect 99422 208098 99604 208334
rect 99004 172654 99604 208098
rect 99004 172418 99186 172654
rect 99422 172418 99604 172654
rect 99004 172334 99604 172418
rect 99004 172098 99186 172334
rect 99422 172098 99604 172334
rect 99004 136654 99604 172098
rect 99004 136418 99186 136654
rect 99422 136418 99604 136654
rect 99004 136334 99604 136418
rect 99004 136098 99186 136334
rect 99422 136098 99604 136334
rect 99004 100654 99604 136098
rect 99004 100418 99186 100654
rect 99422 100418 99604 100654
rect 99004 100334 99604 100418
rect 99004 100098 99186 100334
rect 99422 100098 99604 100334
rect 99004 64654 99604 100098
rect 99004 64418 99186 64654
rect 99422 64418 99604 64654
rect 99004 64334 99604 64418
rect 99004 64098 99186 64334
rect 99422 64098 99604 64334
rect 99004 28654 99604 64098
rect 99004 28418 99186 28654
rect 99422 28418 99604 28654
rect 99004 28334 99604 28418
rect 99004 28098 99186 28334
rect 99422 28098 99604 28334
rect 99004 -5046 99604 28098
rect 99004 -5282 99186 -5046
rect 99422 -5282 99604 -5046
rect 99004 -5366 99604 -5282
rect 99004 -5602 99186 -5366
rect 99422 -5602 99604 -5366
rect 99004 -5624 99604 -5602
rect 102604 680254 103204 710862
rect 120604 710478 121204 711440
rect 120604 710242 120786 710478
rect 121022 710242 121204 710478
rect 120604 710158 121204 710242
rect 120604 709922 120786 710158
rect 121022 709922 121204 710158
rect 117004 708598 117604 709560
rect 117004 708362 117186 708598
rect 117422 708362 117604 708598
rect 117004 708278 117604 708362
rect 117004 708042 117186 708278
rect 117422 708042 117604 708278
rect 113404 706718 114004 707680
rect 113404 706482 113586 706718
rect 113822 706482 114004 706718
rect 113404 706398 114004 706482
rect 113404 706162 113586 706398
rect 113822 706162 114004 706398
rect 102604 680018 102786 680254
rect 103022 680018 103204 680254
rect 102604 679934 103204 680018
rect 102604 679698 102786 679934
rect 103022 679698 103204 679934
rect 102604 644254 103204 679698
rect 102604 644018 102786 644254
rect 103022 644018 103204 644254
rect 102604 643934 103204 644018
rect 102604 643698 102786 643934
rect 103022 643698 103204 643934
rect 102604 608254 103204 643698
rect 102604 608018 102786 608254
rect 103022 608018 103204 608254
rect 102604 607934 103204 608018
rect 102604 607698 102786 607934
rect 103022 607698 103204 607934
rect 102604 572254 103204 607698
rect 102604 572018 102786 572254
rect 103022 572018 103204 572254
rect 102604 571934 103204 572018
rect 102604 571698 102786 571934
rect 103022 571698 103204 571934
rect 102604 536254 103204 571698
rect 102604 536018 102786 536254
rect 103022 536018 103204 536254
rect 102604 535934 103204 536018
rect 102604 535698 102786 535934
rect 103022 535698 103204 535934
rect 102604 500254 103204 535698
rect 102604 500018 102786 500254
rect 103022 500018 103204 500254
rect 102604 499934 103204 500018
rect 102604 499698 102786 499934
rect 103022 499698 103204 499934
rect 102604 464254 103204 499698
rect 102604 464018 102786 464254
rect 103022 464018 103204 464254
rect 102604 463934 103204 464018
rect 102604 463698 102786 463934
rect 103022 463698 103204 463934
rect 102604 428254 103204 463698
rect 102604 428018 102786 428254
rect 103022 428018 103204 428254
rect 102604 427934 103204 428018
rect 102604 427698 102786 427934
rect 103022 427698 103204 427934
rect 102604 392254 103204 427698
rect 102604 392018 102786 392254
rect 103022 392018 103204 392254
rect 102604 391934 103204 392018
rect 102604 391698 102786 391934
rect 103022 391698 103204 391934
rect 102604 356254 103204 391698
rect 102604 356018 102786 356254
rect 103022 356018 103204 356254
rect 102604 355934 103204 356018
rect 102604 355698 102786 355934
rect 103022 355698 103204 355934
rect 102604 320254 103204 355698
rect 102604 320018 102786 320254
rect 103022 320018 103204 320254
rect 102604 319934 103204 320018
rect 102604 319698 102786 319934
rect 103022 319698 103204 319934
rect 102604 284254 103204 319698
rect 102604 284018 102786 284254
rect 103022 284018 103204 284254
rect 102604 283934 103204 284018
rect 102604 283698 102786 283934
rect 103022 283698 103204 283934
rect 102604 248254 103204 283698
rect 102604 248018 102786 248254
rect 103022 248018 103204 248254
rect 102604 247934 103204 248018
rect 102604 247698 102786 247934
rect 103022 247698 103204 247934
rect 102604 212254 103204 247698
rect 102604 212018 102786 212254
rect 103022 212018 103204 212254
rect 102604 211934 103204 212018
rect 102604 211698 102786 211934
rect 103022 211698 103204 211934
rect 102604 176254 103204 211698
rect 102604 176018 102786 176254
rect 103022 176018 103204 176254
rect 102604 175934 103204 176018
rect 102604 175698 102786 175934
rect 103022 175698 103204 175934
rect 102604 140254 103204 175698
rect 102604 140018 102786 140254
rect 103022 140018 103204 140254
rect 102604 139934 103204 140018
rect 102604 139698 102786 139934
rect 103022 139698 103204 139934
rect 102604 104254 103204 139698
rect 102604 104018 102786 104254
rect 103022 104018 103204 104254
rect 102604 103934 103204 104018
rect 102604 103698 102786 103934
rect 103022 103698 103204 103934
rect 102604 68254 103204 103698
rect 102604 68018 102786 68254
rect 103022 68018 103204 68254
rect 102604 67934 103204 68018
rect 102604 67698 102786 67934
rect 103022 67698 103204 67934
rect 102604 32254 103204 67698
rect 102604 32018 102786 32254
rect 103022 32018 103204 32254
rect 102604 31934 103204 32018
rect 102604 31698 102786 31934
rect 103022 31698 103204 31934
rect 84604 -6222 84786 -5986
rect 85022 -6222 85204 -5986
rect 84604 -6306 85204 -6222
rect 84604 -6542 84786 -6306
rect 85022 -6542 85204 -6306
rect 84604 -7504 85204 -6542
rect 102604 -6926 103204 31698
rect 109804 704838 110404 705800
rect 109804 704602 109986 704838
rect 110222 704602 110404 704838
rect 109804 704518 110404 704602
rect 109804 704282 109986 704518
rect 110222 704282 110404 704518
rect 109804 687454 110404 704282
rect 109804 687218 109986 687454
rect 110222 687218 110404 687454
rect 109804 687134 110404 687218
rect 109804 686898 109986 687134
rect 110222 686898 110404 687134
rect 109804 651454 110404 686898
rect 109804 651218 109986 651454
rect 110222 651218 110404 651454
rect 109804 651134 110404 651218
rect 109804 650898 109986 651134
rect 110222 650898 110404 651134
rect 109804 615454 110404 650898
rect 109804 615218 109986 615454
rect 110222 615218 110404 615454
rect 109804 615134 110404 615218
rect 109804 614898 109986 615134
rect 110222 614898 110404 615134
rect 109804 579454 110404 614898
rect 109804 579218 109986 579454
rect 110222 579218 110404 579454
rect 109804 579134 110404 579218
rect 109804 578898 109986 579134
rect 110222 578898 110404 579134
rect 109804 543454 110404 578898
rect 109804 543218 109986 543454
rect 110222 543218 110404 543454
rect 109804 543134 110404 543218
rect 109804 542898 109986 543134
rect 110222 542898 110404 543134
rect 109804 507454 110404 542898
rect 109804 507218 109986 507454
rect 110222 507218 110404 507454
rect 109804 507134 110404 507218
rect 109804 506898 109986 507134
rect 110222 506898 110404 507134
rect 109804 471454 110404 506898
rect 109804 471218 109986 471454
rect 110222 471218 110404 471454
rect 109804 471134 110404 471218
rect 109804 470898 109986 471134
rect 110222 470898 110404 471134
rect 109804 435454 110404 470898
rect 109804 435218 109986 435454
rect 110222 435218 110404 435454
rect 109804 435134 110404 435218
rect 109804 434898 109986 435134
rect 110222 434898 110404 435134
rect 109804 399454 110404 434898
rect 109804 399218 109986 399454
rect 110222 399218 110404 399454
rect 109804 399134 110404 399218
rect 109804 398898 109986 399134
rect 110222 398898 110404 399134
rect 109804 363454 110404 398898
rect 109804 363218 109986 363454
rect 110222 363218 110404 363454
rect 109804 363134 110404 363218
rect 109804 362898 109986 363134
rect 110222 362898 110404 363134
rect 109804 327454 110404 362898
rect 109804 327218 109986 327454
rect 110222 327218 110404 327454
rect 109804 327134 110404 327218
rect 109804 326898 109986 327134
rect 110222 326898 110404 327134
rect 109804 291454 110404 326898
rect 109804 291218 109986 291454
rect 110222 291218 110404 291454
rect 109804 291134 110404 291218
rect 109804 290898 109986 291134
rect 110222 290898 110404 291134
rect 109804 255454 110404 290898
rect 109804 255218 109986 255454
rect 110222 255218 110404 255454
rect 109804 255134 110404 255218
rect 109804 254898 109986 255134
rect 110222 254898 110404 255134
rect 109804 219454 110404 254898
rect 109804 219218 109986 219454
rect 110222 219218 110404 219454
rect 109804 219134 110404 219218
rect 109804 218898 109986 219134
rect 110222 218898 110404 219134
rect 109804 183454 110404 218898
rect 109804 183218 109986 183454
rect 110222 183218 110404 183454
rect 109804 183134 110404 183218
rect 109804 182898 109986 183134
rect 110222 182898 110404 183134
rect 109804 147454 110404 182898
rect 109804 147218 109986 147454
rect 110222 147218 110404 147454
rect 109804 147134 110404 147218
rect 109804 146898 109986 147134
rect 110222 146898 110404 147134
rect 109804 111454 110404 146898
rect 109804 111218 109986 111454
rect 110222 111218 110404 111454
rect 109804 111134 110404 111218
rect 109804 110898 109986 111134
rect 110222 110898 110404 111134
rect 109804 75454 110404 110898
rect 109804 75218 109986 75454
rect 110222 75218 110404 75454
rect 109804 75134 110404 75218
rect 109804 74898 109986 75134
rect 110222 74898 110404 75134
rect 109804 39454 110404 74898
rect 109804 39218 109986 39454
rect 110222 39218 110404 39454
rect 109804 39134 110404 39218
rect 109804 38898 109986 39134
rect 110222 38898 110404 39134
rect 109804 3454 110404 38898
rect 109804 3218 109986 3454
rect 110222 3218 110404 3454
rect 109804 3134 110404 3218
rect 109804 2898 109986 3134
rect 110222 2898 110404 3134
rect 109804 -346 110404 2898
rect 109804 -582 109986 -346
rect 110222 -582 110404 -346
rect 109804 -666 110404 -582
rect 109804 -902 109986 -666
rect 110222 -902 110404 -666
rect 109804 -1864 110404 -902
rect 113404 691054 114004 706162
rect 113404 690818 113586 691054
rect 113822 690818 114004 691054
rect 113404 690734 114004 690818
rect 113404 690498 113586 690734
rect 113822 690498 114004 690734
rect 113404 655054 114004 690498
rect 113404 654818 113586 655054
rect 113822 654818 114004 655054
rect 113404 654734 114004 654818
rect 113404 654498 113586 654734
rect 113822 654498 114004 654734
rect 113404 619054 114004 654498
rect 113404 618818 113586 619054
rect 113822 618818 114004 619054
rect 113404 618734 114004 618818
rect 113404 618498 113586 618734
rect 113822 618498 114004 618734
rect 113404 583054 114004 618498
rect 113404 582818 113586 583054
rect 113822 582818 114004 583054
rect 113404 582734 114004 582818
rect 113404 582498 113586 582734
rect 113822 582498 114004 582734
rect 113404 547054 114004 582498
rect 113404 546818 113586 547054
rect 113822 546818 114004 547054
rect 113404 546734 114004 546818
rect 113404 546498 113586 546734
rect 113822 546498 114004 546734
rect 113404 511054 114004 546498
rect 113404 510818 113586 511054
rect 113822 510818 114004 511054
rect 113404 510734 114004 510818
rect 113404 510498 113586 510734
rect 113822 510498 114004 510734
rect 113404 475054 114004 510498
rect 113404 474818 113586 475054
rect 113822 474818 114004 475054
rect 113404 474734 114004 474818
rect 113404 474498 113586 474734
rect 113822 474498 114004 474734
rect 113404 439054 114004 474498
rect 113404 438818 113586 439054
rect 113822 438818 114004 439054
rect 113404 438734 114004 438818
rect 113404 438498 113586 438734
rect 113822 438498 114004 438734
rect 113404 403054 114004 438498
rect 113404 402818 113586 403054
rect 113822 402818 114004 403054
rect 113404 402734 114004 402818
rect 113404 402498 113586 402734
rect 113822 402498 114004 402734
rect 113404 367054 114004 402498
rect 113404 366818 113586 367054
rect 113822 366818 114004 367054
rect 113404 366734 114004 366818
rect 113404 366498 113586 366734
rect 113822 366498 114004 366734
rect 113404 331054 114004 366498
rect 113404 330818 113586 331054
rect 113822 330818 114004 331054
rect 113404 330734 114004 330818
rect 113404 330498 113586 330734
rect 113822 330498 114004 330734
rect 113404 295054 114004 330498
rect 113404 294818 113586 295054
rect 113822 294818 114004 295054
rect 113404 294734 114004 294818
rect 113404 294498 113586 294734
rect 113822 294498 114004 294734
rect 113404 259054 114004 294498
rect 113404 258818 113586 259054
rect 113822 258818 114004 259054
rect 113404 258734 114004 258818
rect 113404 258498 113586 258734
rect 113822 258498 114004 258734
rect 113404 223054 114004 258498
rect 113404 222818 113586 223054
rect 113822 222818 114004 223054
rect 113404 222734 114004 222818
rect 113404 222498 113586 222734
rect 113822 222498 114004 222734
rect 113404 187054 114004 222498
rect 113404 186818 113586 187054
rect 113822 186818 114004 187054
rect 113404 186734 114004 186818
rect 113404 186498 113586 186734
rect 113822 186498 114004 186734
rect 113404 151054 114004 186498
rect 113404 150818 113586 151054
rect 113822 150818 114004 151054
rect 113404 150734 114004 150818
rect 113404 150498 113586 150734
rect 113822 150498 114004 150734
rect 113404 115054 114004 150498
rect 113404 114818 113586 115054
rect 113822 114818 114004 115054
rect 113404 114734 114004 114818
rect 113404 114498 113586 114734
rect 113822 114498 114004 114734
rect 113404 79054 114004 114498
rect 113404 78818 113586 79054
rect 113822 78818 114004 79054
rect 113404 78734 114004 78818
rect 113404 78498 113586 78734
rect 113822 78498 114004 78734
rect 113404 43054 114004 78498
rect 113404 42818 113586 43054
rect 113822 42818 114004 43054
rect 113404 42734 114004 42818
rect 113404 42498 113586 42734
rect 113822 42498 114004 42734
rect 113404 7054 114004 42498
rect 113404 6818 113586 7054
rect 113822 6818 114004 7054
rect 113404 6734 114004 6818
rect 113404 6498 113586 6734
rect 113822 6498 114004 6734
rect 113404 -2226 114004 6498
rect 113404 -2462 113586 -2226
rect 113822 -2462 114004 -2226
rect 113404 -2546 114004 -2462
rect 113404 -2782 113586 -2546
rect 113822 -2782 114004 -2546
rect 113404 -3744 114004 -2782
rect 117004 694654 117604 708042
rect 117004 694418 117186 694654
rect 117422 694418 117604 694654
rect 117004 694334 117604 694418
rect 117004 694098 117186 694334
rect 117422 694098 117604 694334
rect 117004 658654 117604 694098
rect 117004 658418 117186 658654
rect 117422 658418 117604 658654
rect 117004 658334 117604 658418
rect 117004 658098 117186 658334
rect 117422 658098 117604 658334
rect 117004 622654 117604 658098
rect 117004 622418 117186 622654
rect 117422 622418 117604 622654
rect 117004 622334 117604 622418
rect 117004 622098 117186 622334
rect 117422 622098 117604 622334
rect 117004 586654 117604 622098
rect 117004 586418 117186 586654
rect 117422 586418 117604 586654
rect 117004 586334 117604 586418
rect 117004 586098 117186 586334
rect 117422 586098 117604 586334
rect 117004 550654 117604 586098
rect 117004 550418 117186 550654
rect 117422 550418 117604 550654
rect 117004 550334 117604 550418
rect 117004 550098 117186 550334
rect 117422 550098 117604 550334
rect 117004 514654 117604 550098
rect 117004 514418 117186 514654
rect 117422 514418 117604 514654
rect 117004 514334 117604 514418
rect 117004 514098 117186 514334
rect 117422 514098 117604 514334
rect 117004 478654 117604 514098
rect 117004 478418 117186 478654
rect 117422 478418 117604 478654
rect 117004 478334 117604 478418
rect 117004 478098 117186 478334
rect 117422 478098 117604 478334
rect 117004 442654 117604 478098
rect 117004 442418 117186 442654
rect 117422 442418 117604 442654
rect 117004 442334 117604 442418
rect 117004 442098 117186 442334
rect 117422 442098 117604 442334
rect 117004 406654 117604 442098
rect 117004 406418 117186 406654
rect 117422 406418 117604 406654
rect 117004 406334 117604 406418
rect 117004 406098 117186 406334
rect 117422 406098 117604 406334
rect 117004 370654 117604 406098
rect 117004 370418 117186 370654
rect 117422 370418 117604 370654
rect 117004 370334 117604 370418
rect 117004 370098 117186 370334
rect 117422 370098 117604 370334
rect 117004 334654 117604 370098
rect 117004 334418 117186 334654
rect 117422 334418 117604 334654
rect 117004 334334 117604 334418
rect 117004 334098 117186 334334
rect 117422 334098 117604 334334
rect 117004 298654 117604 334098
rect 117004 298418 117186 298654
rect 117422 298418 117604 298654
rect 117004 298334 117604 298418
rect 117004 298098 117186 298334
rect 117422 298098 117604 298334
rect 117004 262654 117604 298098
rect 117004 262418 117186 262654
rect 117422 262418 117604 262654
rect 117004 262334 117604 262418
rect 117004 262098 117186 262334
rect 117422 262098 117604 262334
rect 117004 226654 117604 262098
rect 117004 226418 117186 226654
rect 117422 226418 117604 226654
rect 117004 226334 117604 226418
rect 117004 226098 117186 226334
rect 117422 226098 117604 226334
rect 117004 190654 117604 226098
rect 117004 190418 117186 190654
rect 117422 190418 117604 190654
rect 117004 190334 117604 190418
rect 117004 190098 117186 190334
rect 117422 190098 117604 190334
rect 117004 154654 117604 190098
rect 117004 154418 117186 154654
rect 117422 154418 117604 154654
rect 117004 154334 117604 154418
rect 117004 154098 117186 154334
rect 117422 154098 117604 154334
rect 117004 118654 117604 154098
rect 117004 118418 117186 118654
rect 117422 118418 117604 118654
rect 117004 118334 117604 118418
rect 117004 118098 117186 118334
rect 117422 118098 117604 118334
rect 117004 82654 117604 118098
rect 117004 82418 117186 82654
rect 117422 82418 117604 82654
rect 117004 82334 117604 82418
rect 117004 82098 117186 82334
rect 117422 82098 117604 82334
rect 117004 46654 117604 82098
rect 117004 46418 117186 46654
rect 117422 46418 117604 46654
rect 117004 46334 117604 46418
rect 117004 46098 117186 46334
rect 117422 46098 117604 46334
rect 117004 10654 117604 46098
rect 117004 10418 117186 10654
rect 117422 10418 117604 10654
rect 117004 10334 117604 10418
rect 117004 10098 117186 10334
rect 117422 10098 117604 10334
rect 117004 -4106 117604 10098
rect 117004 -4342 117186 -4106
rect 117422 -4342 117604 -4106
rect 117004 -4426 117604 -4342
rect 117004 -4662 117186 -4426
rect 117422 -4662 117604 -4426
rect 117004 -5624 117604 -4662
rect 120604 698254 121204 709922
rect 138604 711418 139204 711440
rect 138604 711182 138786 711418
rect 139022 711182 139204 711418
rect 138604 711098 139204 711182
rect 138604 710862 138786 711098
rect 139022 710862 139204 711098
rect 135004 709538 135604 709560
rect 135004 709302 135186 709538
rect 135422 709302 135604 709538
rect 135004 709218 135604 709302
rect 135004 708982 135186 709218
rect 135422 708982 135604 709218
rect 131404 707658 132004 707680
rect 131404 707422 131586 707658
rect 131822 707422 132004 707658
rect 131404 707338 132004 707422
rect 131404 707102 131586 707338
rect 131822 707102 132004 707338
rect 120604 698018 120786 698254
rect 121022 698018 121204 698254
rect 120604 697934 121204 698018
rect 120604 697698 120786 697934
rect 121022 697698 121204 697934
rect 120604 662254 121204 697698
rect 120604 662018 120786 662254
rect 121022 662018 121204 662254
rect 120604 661934 121204 662018
rect 120604 661698 120786 661934
rect 121022 661698 121204 661934
rect 120604 626254 121204 661698
rect 120604 626018 120786 626254
rect 121022 626018 121204 626254
rect 120604 625934 121204 626018
rect 120604 625698 120786 625934
rect 121022 625698 121204 625934
rect 120604 590254 121204 625698
rect 120604 590018 120786 590254
rect 121022 590018 121204 590254
rect 120604 589934 121204 590018
rect 120604 589698 120786 589934
rect 121022 589698 121204 589934
rect 120604 554254 121204 589698
rect 120604 554018 120786 554254
rect 121022 554018 121204 554254
rect 120604 553934 121204 554018
rect 120604 553698 120786 553934
rect 121022 553698 121204 553934
rect 120604 518254 121204 553698
rect 120604 518018 120786 518254
rect 121022 518018 121204 518254
rect 120604 517934 121204 518018
rect 120604 517698 120786 517934
rect 121022 517698 121204 517934
rect 120604 482254 121204 517698
rect 120604 482018 120786 482254
rect 121022 482018 121204 482254
rect 120604 481934 121204 482018
rect 120604 481698 120786 481934
rect 121022 481698 121204 481934
rect 120604 446254 121204 481698
rect 120604 446018 120786 446254
rect 121022 446018 121204 446254
rect 120604 445934 121204 446018
rect 120604 445698 120786 445934
rect 121022 445698 121204 445934
rect 120604 410254 121204 445698
rect 120604 410018 120786 410254
rect 121022 410018 121204 410254
rect 120604 409934 121204 410018
rect 120604 409698 120786 409934
rect 121022 409698 121204 409934
rect 120604 374254 121204 409698
rect 120604 374018 120786 374254
rect 121022 374018 121204 374254
rect 120604 373934 121204 374018
rect 120604 373698 120786 373934
rect 121022 373698 121204 373934
rect 120604 338254 121204 373698
rect 120604 338018 120786 338254
rect 121022 338018 121204 338254
rect 120604 337934 121204 338018
rect 120604 337698 120786 337934
rect 121022 337698 121204 337934
rect 120604 302254 121204 337698
rect 120604 302018 120786 302254
rect 121022 302018 121204 302254
rect 120604 301934 121204 302018
rect 120604 301698 120786 301934
rect 121022 301698 121204 301934
rect 120604 266254 121204 301698
rect 120604 266018 120786 266254
rect 121022 266018 121204 266254
rect 120604 265934 121204 266018
rect 120604 265698 120786 265934
rect 121022 265698 121204 265934
rect 120604 230254 121204 265698
rect 120604 230018 120786 230254
rect 121022 230018 121204 230254
rect 120604 229934 121204 230018
rect 120604 229698 120786 229934
rect 121022 229698 121204 229934
rect 120604 194254 121204 229698
rect 120604 194018 120786 194254
rect 121022 194018 121204 194254
rect 120604 193934 121204 194018
rect 120604 193698 120786 193934
rect 121022 193698 121204 193934
rect 120604 158254 121204 193698
rect 120604 158018 120786 158254
rect 121022 158018 121204 158254
rect 120604 157934 121204 158018
rect 120604 157698 120786 157934
rect 121022 157698 121204 157934
rect 120604 122254 121204 157698
rect 120604 122018 120786 122254
rect 121022 122018 121204 122254
rect 120604 121934 121204 122018
rect 120604 121698 120786 121934
rect 121022 121698 121204 121934
rect 120604 86254 121204 121698
rect 120604 86018 120786 86254
rect 121022 86018 121204 86254
rect 120604 85934 121204 86018
rect 120604 85698 120786 85934
rect 121022 85698 121204 85934
rect 120604 50254 121204 85698
rect 120604 50018 120786 50254
rect 121022 50018 121204 50254
rect 120604 49934 121204 50018
rect 120604 49698 120786 49934
rect 121022 49698 121204 49934
rect 120604 14254 121204 49698
rect 120604 14018 120786 14254
rect 121022 14018 121204 14254
rect 120604 13934 121204 14018
rect 120604 13698 120786 13934
rect 121022 13698 121204 13934
rect 102604 -7162 102786 -6926
rect 103022 -7162 103204 -6926
rect 102604 -7246 103204 -7162
rect 102604 -7482 102786 -7246
rect 103022 -7482 103204 -7246
rect 102604 -7504 103204 -7482
rect 120604 -5986 121204 13698
rect 127804 705778 128404 705800
rect 127804 705542 127986 705778
rect 128222 705542 128404 705778
rect 127804 705458 128404 705542
rect 127804 705222 127986 705458
rect 128222 705222 128404 705458
rect 127804 669454 128404 705222
rect 127804 669218 127986 669454
rect 128222 669218 128404 669454
rect 127804 669134 128404 669218
rect 127804 668898 127986 669134
rect 128222 668898 128404 669134
rect 127804 633454 128404 668898
rect 127804 633218 127986 633454
rect 128222 633218 128404 633454
rect 127804 633134 128404 633218
rect 127804 632898 127986 633134
rect 128222 632898 128404 633134
rect 127804 597454 128404 632898
rect 127804 597218 127986 597454
rect 128222 597218 128404 597454
rect 127804 597134 128404 597218
rect 127804 596898 127986 597134
rect 128222 596898 128404 597134
rect 127804 561454 128404 596898
rect 127804 561218 127986 561454
rect 128222 561218 128404 561454
rect 127804 561134 128404 561218
rect 127804 560898 127986 561134
rect 128222 560898 128404 561134
rect 127804 525454 128404 560898
rect 127804 525218 127986 525454
rect 128222 525218 128404 525454
rect 127804 525134 128404 525218
rect 127804 524898 127986 525134
rect 128222 524898 128404 525134
rect 127804 489454 128404 524898
rect 127804 489218 127986 489454
rect 128222 489218 128404 489454
rect 127804 489134 128404 489218
rect 127804 488898 127986 489134
rect 128222 488898 128404 489134
rect 127804 453454 128404 488898
rect 127804 453218 127986 453454
rect 128222 453218 128404 453454
rect 127804 453134 128404 453218
rect 127804 452898 127986 453134
rect 128222 452898 128404 453134
rect 127804 417454 128404 452898
rect 127804 417218 127986 417454
rect 128222 417218 128404 417454
rect 127804 417134 128404 417218
rect 127804 416898 127986 417134
rect 128222 416898 128404 417134
rect 127804 381454 128404 416898
rect 127804 381218 127986 381454
rect 128222 381218 128404 381454
rect 127804 381134 128404 381218
rect 127804 380898 127986 381134
rect 128222 380898 128404 381134
rect 127804 345454 128404 380898
rect 127804 345218 127986 345454
rect 128222 345218 128404 345454
rect 127804 345134 128404 345218
rect 127804 344898 127986 345134
rect 128222 344898 128404 345134
rect 127804 309454 128404 344898
rect 127804 309218 127986 309454
rect 128222 309218 128404 309454
rect 127804 309134 128404 309218
rect 127804 308898 127986 309134
rect 128222 308898 128404 309134
rect 127804 273454 128404 308898
rect 127804 273218 127986 273454
rect 128222 273218 128404 273454
rect 127804 273134 128404 273218
rect 127804 272898 127986 273134
rect 128222 272898 128404 273134
rect 127804 237454 128404 272898
rect 127804 237218 127986 237454
rect 128222 237218 128404 237454
rect 127804 237134 128404 237218
rect 127804 236898 127986 237134
rect 128222 236898 128404 237134
rect 127804 201454 128404 236898
rect 127804 201218 127986 201454
rect 128222 201218 128404 201454
rect 127804 201134 128404 201218
rect 127804 200898 127986 201134
rect 128222 200898 128404 201134
rect 127804 165454 128404 200898
rect 127804 165218 127986 165454
rect 128222 165218 128404 165454
rect 127804 165134 128404 165218
rect 127804 164898 127986 165134
rect 128222 164898 128404 165134
rect 127804 129454 128404 164898
rect 127804 129218 127986 129454
rect 128222 129218 128404 129454
rect 127804 129134 128404 129218
rect 127804 128898 127986 129134
rect 128222 128898 128404 129134
rect 127804 93454 128404 128898
rect 127804 93218 127986 93454
rect 128222 93218 128404 93454
rect 127804 93134 128404 93218
rect 127804 92898 127986 93134
rect 128222 92898 128404 93134
rect 127804 57454 128404 92898
rect 127804 57218 127986 57454
rect 128222 57218 128404 57454
rect 127804 57134 128404 57218
rect 127804 56898 127986 57134
rect 128222 56898 128404 57134
rect 127804 21454 128404 56898
rect 127804 21218 127986 21454
rect 128222 21218 128404 21454
rect 127804 21134 128404 21218
rect 127804 20898 127986 21134
rect 128222 20898 128404 21134
rect 127804 -1286 128404 20898
rect 127804 -1522 127986 -1286
rect 128222 -1522 128404 -1286
rect 127804 -1606 128404 -1522
rect 127804 -1842 127986 -1606
rect 128222 -1842 128404 -1606
rect 127804 -1864 128404 -1842
rect 131404 673054 132004 707102
rect 131404 672818 131586 673054
rect 131822 672818 132004 673054
rect 131404 672734 132004 672818
rect 131404 672498 131586 672734
rect 131822 672498 132004 672734
rect 131404 637054 132004 672498
rect 131404 636818 131586 637054
rect 131822 636818 132004 637054
rect 131404 636734 132004 636818
rect 131404 636498 131586 636734
rect 131822 636498 132004 636734
rect 131404 601054 132004 636498
rect 131404 600818 131586 601054
rect 131822 600818 132004 601054
rect 131404 600734 132004 600818
rect 131404 600498 131586 600734
rect 131822 600498 132004 600734
rect 131404 565054 132004 600498
rect 131404 564818 131586 565054
rect 131822 564818 132004 565054
rect 131404 564734 132004 564818
rect 131404 564498 131586 564734
rect 131822 564498 132004 564734
rect 131404 529054 132004 564498
rect 131404 528818 131586 529054
rect 131822 528818 132004 529054
rect 131404 528734 132004 528818
rect 131404 528498 131586 528734
rect 131822 528498 132004 528734
rect 131404 493054 132004 528498
rect 131404 492818 131586 493054
rect 131822 492818 132004 493054
rect 131404 492734 132004 492818
rect 131404 492498 131586 492734
rect 131822 492498 132004 492734
rect 131404 457054 132004 492498
rect 131404 456818 131586 457054
rect 131822 456818 132004 457054
rect 131404 456734 132004 456818
rect 131404 456498 131586 456734
rect 131822 456498 132004 456734
rect 131404 421054 132004 456498
rect 131404 420818 131586 421054
rect 131822 420818 132004 421054
rect 131404 420734 132004 420818
rect 131404 420498 131586 420734
rect 131822 420498 132004 420734
rect 131404 385054 132004 420498
rect 131404 384818 131586 385054
rect 131822 384818 132004 385054
rect 131404 384734 132004 384818
rect 131404 384498 131586 384734
rect 131822 384498 132004 384734
rect 131404 349054 132004 384498
rect 131404 348818 131586 349054
rect 131822 348818 132004 349054
rect 131404 348734 132004 348818
rect 131404 348498 131586 348734
rect 131822 348498 132004 348734
rect 131404 313054 132004 348498
rect 131404 312818 131586 313054
rect 131822 312818 132004 313054
rect 131404 312734 132004 312818
rect 131404 312498 131586 312734
rect 131822 312498 132004 312734
rect 131404 277054 132004 312498
rect 131404 276818 131586 277054
rect 131822 276818 132004 277054
rect 131404 276734 132004 276818
rect 131404 276498 131586 276734
rect 131822 276498 132004 276734
rect 131404 241054 132004 276498
rect 131404 240818 131586 241054
rect 131822 240818 132004 241054
rect 131404 240734 132004 240818
rect 131404 240498 131586 240734
rect 131822 240498 132004 240734
rect 131404 205054 132004 240498
rect 131404 204818 131586 205054
rect 131822 204818 132004 205054
rect 131404 204734 132004 204818
rect 131404 204498 131586 204734
rect 131822 204498 132004 204734
rect 131404 169054 132004 204498
rect 131404 168818 131586 169054
rect 131822 168818 132004 169054
rect 131404 168734 132004 168818
rect 131404 168498 131586 168734
rect 131822 168498 132004 168734
rect 131404 133054 132004 168498
rect 131404 132818 131586 133054
rect 131822 132818 132004 133054
rect 131404 132734 132004 132818
rect 131404 132498 131586 132734
rect 131822 132498 132004 132734
rect 131404 97054 132004 132498
rect 131404 96818 131586 97054
rect 131822 96818 132004 97054
rect 131404 96734 132004 96818
rect 131404 96498 131586 96734
rect 131822 96498 132004 96734
rect 131404 61054 132004 96498
rect 131404 60818 131586 61054
rect 131822 60818 132004 61054
rect 131404 60734 132004 60818
rect 131404 60498 131586 60734
rect 131822 60498 132004 60734
rect 131404 25054 132004 60498
rect 131404 24818 131586 25054
rect 131822 24818 132004 25054
rect 131404 24734 132004 24818
rect 131404 24498 131586 24734
rect 131822 24498 132004 24734
rect 131404 -3166 132004 24498
rect 131404 -3402 131586 -3166
rect 131822 -3402 132004 -3166
rect 131404 -3486 132004 -3402
rect 131404 -3722 131586 -3486
rect 131822 -3722 132004 -3486
rect 131404 -3744 132004 -3722
rect 135004 676654 135604 708982
rect 135004 676418 135186 676654
rect 135422 676418 135604 676654
rect 135004 676334 135604 676418
rect 135004 676098 135186 676334
rect 135422 676098 135604 676334
rect 135004 640654 135604 676098
rect 135004 640418 135186 640654
rect 135422 640418 135604 640654
rect 135004 640334 135604 640418
rect 135004 640098 135186 640334
rect 135422 640098 135604 640334
rect 135004 604654 135604 640098
rect 135004 604418 135186 604654
rect 135422 604418 135604 604654
rect 135004 604334 135604 604418
rect 135004 604098 135186 604334
rect 135422 604098 135604 604334
rect 135004 568654 135604 604098
rect 135004 568418 135186 568654
rect 135422 568418 135604 568654
rect 135004 568334 135604 568418
rect 135004 568098 135186 568334
rect 135422 568098 135604 568334
rect 135004 532654 135604 568098
rect 135004 532418 135186 532654
rect 135422 532418 135604 532654
rect 135004 532334 135604 532418
rect 135004 532098 135186 532334
rect 135422 532098 135604 532334
rect 135004 496654 135604 532098
rect 135004 496418 135186 496654
rect 135422 496418 135604 496654
rect 135004 496334 135604 496418
rect 135004 496098 135186 496334
rect 135422 496098 135604 496334
rect 135004 460654 135604 496098
rect 135004 460418 135186 460654
rect 135422 460418 135604 460654
rect 135004 460334 135604 460418
rect 135004 460098 135186 460334
rect 135422 460098 135604 460334
rect 135004 424654 135604 460098
rect 135004 424418 135186 424654
rect 135422 424418 135604 424654
rect 135004 424334 135604 424418
rect 135004 424098 135186 424334
rect 135422 424098 135604 424334
rect 135004 388654 135604 424098
rect 135004 388418 135186 388654
rect 135422 388418 135604 388654
rect 135004 388334 135604 388418
rect 135004 388098 135186 388334
rect 135422 388098 135604 388334
rect 135004 352654 135604 388098
rect 135004 352418 135186 352654
rect 135422 352418 135604 352654
rect 135004 352334 135604 352418
rect 135004 352098 135186 352334
rect 135422 352098 135604 352334
rect 135004 316654 135604 352098
rect 135004 316418 135186 316654
rect 135422 316418 135604 316654
rect 135004 316334 135604 316418
rect 135004 316098 135186 316334
rect 135422 316098 135604 316334
rect 135004 280654 135604 316098
rect 135004 280418 135186 280654
rect 135422 280418 135604 280654
rect 135004 280334 135604 280418
rect 135004 280098 135186 280334
rect 135422 280098 135604 280334
rect 135004 244654 135604 280098
rect 135004 244418 135186 244654
rect 135422 244418 135604 244654
rect 135004 244334 135604 244418
rect 135004 244098 135186 244334
rect 135422 244098 135604 244334
rect 135004 208654 135604 244098
rect 135004 208418 135186 208654
rect 135422 208418 135604 208654
rect 135004 208334 135604 208418
rect 135004 208098 135186 208334
rect 135422 208098 135604 208334
rect 135004 172654 135604 208098
rect 135004 172418 135186 172654
rect 135422 172418 135604 172654
rect 135004 172334 135604 172418
rect 135004 172098 135186 172334
rect 135422 172098 135604 172334
rect 135004 136654 135604 172098
rect 135004 136418 135186 136654
rect 135422 136418 135604 136654
rect 135004 136334 135604 136418
rect 135004 136098 135186 136334
rect 135422 136098 135604 136334
rect 135004 100654 135604 136098
rect 135004 100418 135186 100654
rect 135422 100418 135604 100654
rect 135004 100334 135604 100418
rect 135004 100098 135186 100334
rect 135422 100098 135604 100334
rect 135004 64654 135604 100098
rect 135004 64418 135186 64654
rect 135422 64418 135604 64654
rect 135004 64334 135604 64418
rect 135004 64098 135186 64334
rect 135422 64098 135604 64334
rect 135004 28654 135604 64098
rect 135004 28418 135186 28654
rect 135422 28418 135604 28654
rect 135004 28334 135604 28418
rect 135004 28098 135186 28334
rect 135422 28098 135604 28334
rect 135004 -5046 135604 28098
rect 135004 -5282 135186 -5046
rect 135422 -5282 135604 -5046
rect 135004 -5366 135604 -5282
rect 135004 -5602 135186 -5366
rect 135422 -5602 135604 -5366
rect 135004 -5624 135604 -5602
rect 138604 680254 139204 710862
rect 156604 710478 157204 711440
rect 156604 710242 156786 710478
rect 157022 710242 157204 710478
rect 156604 710158 157204 710242
rect 156604 709922 156786 710158
rect 157022 709922 157204 710158
rect 153004 708598 153604 709560
rect 153004 708362 153186 708598
rect 153422 708362 153604 708598
rect 153004 708278 153604 708362
rect 153004 708042 153186 708278
rect 153422 708042 153604 708278
rect 149404 706718 150004 707680
rect 149404 706482 149586 706718
rect 149822 706482 150004 706718
rect 149404 706398 150004 706482
rect 149404 706162 149586 706398
rect 149822 706162 150004 706398
rect 138604 680018 138786 680254
rect 139022 680018 139204 680254
rect 138604 679934 139204 680018
rect 138604 679698 138786 679934
rect 139022 679698 139204 679934
rect 138604 644254 139204 679698
rect 138604 644018 138786 644254
rect 139022 644018 139204 644254
rect 138604 643934 139204 644018
rect 138604 643698 138786 643934
rect 139022 643698 139204 643934
rect 138604 608254 139204 643698
rect 138604 608018 138786 608254
rect 139022 608018 139204 608254
rect 138604 607934 139204 608018
rect 138604 607698 138786 607934
rect 139022 607698 139204 607934
rect 138604 572254 139204 607698
rect 138604 572018 138786 572254
rect 139022 572018 139204 572254
rect 138604 571934 139204 572018
rect 138604 571698 138786 571934
rect 139022 571698 139204 571934
rect 138604 536254 139204 571698
rect 138604 536018 138786 536254
rect 139022 536018 139204 536254
rect 138604 535934 139204 536018
rect 138604 535698 138786 535934
rect 139022 535698 139204 535934
rect 138604 500254 139204 535698
rect 138604 500018 138786 500254
rect 139022 500018 139204 500254
rect 138604 499934 139204 500018
rect 138604 499698 138786 499934
rect 139022 499698 139204 499934
rect 138604 464254 139204 499698
rect 138604 464018 138786 464254
rect 139022 464018 139204 464254
rect 138604 463934 139204 464018
rect 138604 463698 138786 463934
rect 139022 463698 139204 463934
rect 138604 428254 139204 463698
rect 138604 428018 138786 428254
rect 139022 428018 139204 428254
rect 138604 427934 139204 428018
rect 138604 427698 138786 427934
rect 139022 427698 139204 427934
rect 138604 392254 139204 427698
rect 138604 392018 138786 392254
rect 139022 392018 139204 392254
rect 138604 391934 139204 392018
rect 138604 391698 138786 391934
rect 139022 391698 139204 391934
rect 138604 356254 139204 391698
rect 138604 356018 138786 356254
rect 139022 356018 139204 356254
rect 138604 355934 139204 356018
rect 138604 355698 138786 355934
rect 139022 355698 139204 355934
rect 138604 320254 139204 355698
rect 138604 320018 138786 320254
rect 139022 320018 139204 320254
rect 138604 319934 139204 320018
rect 138604 319698 138786 319934
rect 139022 319698 139204 319934
rect 138604 284254 139204 319698
rect 138604 284018 138786 284254
rect 139022 284018 139204 284254
rect 138604 283934 139204 284018
rect 138604 283698 138786 283934
rect 139022 283698 139204 283934
rect 138604 248254 139204 283698
rect 138604 248018 138786 248254
rect 139022 248018 139204 248254
rect 138604 247934 139204 248018
rect 138604 247698 138786 247934
rect 139022 247698 139204 247934
rect 138604 212254 139204 247698
rect 138604 212018 138786 212254
rect 139022 212018 139204 212254
rect 138604 211934 139204 212018
rect 138604 211698 138786 211934
rect 139022 211698 139204 211934
rect 138604 176254 139204 211698
rect 138604 176018 138786 176254
rect 139022 176018 139204 176254
rect 138604 175934 139204 176018
rect 138604 175698 138786 175934
rect 139022 175698 139204 175934
rect 138604 140254 139204 175698
rect 138604 140018 138786 140254
rect 139022 140018 139204 140254
rect 138604 139934 139204 140018
rect 138604 139698 138786 139934
rect 139022 139698 139204 139934
rect 138604 104254 139204 139698
rect 138604 104018 138786 104254
rect 139022 104018 139204 104254
rect 138604 103934 139204 104018
rect 138604 103698 138786 103934
rect 139022 103698 139204 103934
rect 138604 68254 139204 103698
rect 138604 68018 138786 68254
rect 139022 68018 139204 68254
rect 138604 67934 139204 68018
rect 138604 67698 138786 67934
rect 139022 67698 139204 67934
rect 138604 32254 139204 67698
rect 138604 32018 138786 32254
rect 139022 32018 139204 32254
rect 138604 31934 139204 32018
rect 138604 31698 138786 31934
rect 139022 31698 139204 31934
rect 120604 -6222 120786 -5986
rect 121022 -6222 121204 -5986
rect 120604 -6306 121204 -6222
rect 120604 -6542 120786 -6306
rect 121022 -6542 121204 -6306
rect 120604 -7504 121204 -6542
rect 138604 -6926 139204 31698
rect 145804 704838 146404 705800
rect 145804 704602 145986 704838
rect 146222 704602 146404 704838
rect 145804 704518 146404 704602
rect 145804 704282 145986 704518
rect 146222 704282 146404 704518
rect 145804 687454 146404 704282
rect 145804 687218 145986 687454
rect 146222 687218 146404 687454
rect 145804 687134 146404 687218
rect 145804 686898 145986 687134
rect 146222 686898 146404 687134
rect 145804 651454 146404 686898
rect 145804 651218 145986 651454
rect 146222 651218 146404 651454
rect 145804 651134 146404 651218
rect 145804 650898 145986 651134
rect 146222 650898 146404 651134
rect 145804 615454 146404 650898
rect 145804 615218 145986 615454
rect 146222 615218 146404 615454
rect 145804 615134 146404 615218
rect 145804 614898 145986 615134
rect 146222 614898 146404 615134
rect 145804 579454 146404 614898
rect 145804 579218 145986 579454
rect 146222 579218 146404 579454
rect 145804 579134 146404 579218
rect 145804 578898 145986 579134
rect 146222 578898 146404 579134
rect 145804 543454 146404 578898
rect 145804 543218 145986 543454
rect 146222 543218 146404 543454
rect 145804 543134 146404 543218
rect 145804 542898 145986 543134
rect 146222 542898 146404 543134
rect 145804 507454 146404 542898
rect 145804 507218 145986 507454
rect 146222 507218 146404 507454
rect 145804 507134 146404 507218
rect 145804 506898 145986 507134
rect 146222 506898 146404 507134
rect 145804 471454 146404 506898
rect 145804 471218 145986 471454
rect 146222 471218 146404 471454
rect 145804 471134 146404 471218
rect 145804 470898 145986 471134
rect 146222 470898 146404 471134
rect 145804 435454 146404 470898
rect 145804 435218 145986 435454
rect 146222 435218 146404 435454
rect 145804 435134 146404 435218
rect 145804 434898 145986 435134
rect 146222 434898 146404 435134
rect 145804 399454 146404 434898
rect 145804 399218 145986 399454
rect 146222 399218 146404 399454
rect 145804 399134 146404 399218
rect 145804 398898 145986 399134
rect 146222 398898 146404 399134
rect 145804 363454 146404 398898
rect 145804 363218 145986 363454
rect 146222 363218 146404 363454
rect 145804 363134 146404 363218
rect 145804 362898 145986 363134
rect 146222 362898 146404 363134
rect 145804 327454 146404 362898
rect 145804 327218 145986 327454
rect 146222 327218 146404 327454
rect 145804 327134 146404 327218
rect 145804 326898 145986 327134
rect 146222 326898 146404 327134
rect 145804 291454 146404 326898
rect 145804 291218 145986 291454
rect 146222 291218 146404 291454
rect 145804 291134 146404 291218
rect 145804 290898 145986 291134
rect 146222 290898 146404 291134
rect 145804 255454 146404 290898
rect 145804 255218 145986 255454
rect 146222 255218 146404 255454
rect 145804 255134 146404 255218
rect 145804 254898 145986 255134
rect 146222 254898 146404 255134
rect 145804 219454 146404 254898
rect 145804 219218 145986 219454
rect 146222 219218 146404 219454
rect 145804 219134 146404 219218
rect 145804 218898 145986 219134
rect 146222 218898 146404 219134
rect 145804 183454 146404 218898
rect 145804 183218 145986 183454
rect 146222 183218 146404 183454
rect 145804 183134 146404 183218
rect 145804 182898 145986 183134
rect 146222 182898 146404 183134
rect 145804 147454 146404 182898
rect 145804 147218 145986 147454
rect 146222 147218 146404 147454
rect 145804 147134 146404 147218
rect 145804 146898 145986 147134
rect 146222 146898 146404 147134
rect 145804 111454 146404 146898
rect 145804 111218 145986 111454
rect 146222 111218 146404 111454
rect 145804 111134 146404 111218
rect 145804 110898 145986 111134
rect 146222 110898 146404 111134
rect 145804 75454 146404 110898
rect 145804 75218 145986 75454
rect 146222 75218 146404 75454
rect 145804 75134 146404 75218
rect 145804 74898 145986 75134
rect 146222 74898 146404 75134
rect 145804 39454 146404 74898
rect 145804 39218 145986 39454
rect 146222 39218 146404 39454
rect 145804 39134 146404 39218
rect 145804 38898 145986 39134
rect 146222 38898 146404 39134
rect 145804 3454 146404 38898
rect 145804 3218 145986 3454
rect 146222 3218 146404 3454
rect 145804 3134 146404 3218
rect 145804 2898 145986 3134
rect 146222 2898 146404 3134
rect 145804 -346 146404 2898
rect 145804 -582 145986 -346
rect 146222 -582 146404 -346
rect 145804 -666 146404 -582
rect 145804 -902 145986 -666
rect 146222 -902 146404 -666
rect 145804 -1864 146404 -902
rect 149404 691054 150004 706162
rect 149404 690818 149586 691054
rect 149822 690818 150004 691054
rect 149404 690734 150004 690818
rect 149404 690498 149586 690734
rect 149822 690498 150004 690734
rect 149404 655054 150004 690498
rect 149404 654818 149586 655054
rect 149822 654818 150004 655054
rect 149404 654734 150004 654818
rect 149404 654498 149586 654734
rect 149822 654498 150004 654734
rect 149404 619054 150004 654498
rect 149404 618818 149586 619054
rect 149822 618818 150004 619054
rect 149404 618734 150004 618818
rect 149404 618498 149586 618734
rect 149822 618498 150004 618734
rect 149404 583054 150004 618498
rect 149404 582818 149586 583054
rect 149822 582818 150004 583054
rect 149404 582734 150004 582818
rect 149404 582498 149586 582734
rect 149822 582498 150004 582734
rect 149404 547054 150004 582498
rect 149404 546818 149586 547054
rect 149822 546818 150004 547054
rect 149404 546734 150004 546818
rect 149404 546498 149586 546734
rect 149822 546498 150004 546734
rect 149404 511054 150004 546498
rect 149404 510818 149586 511054
rect 149822 510818 150004 511054
rect 149404 510734 150004 510818
rect 149404 510498 149586 510734
rect 149822 510498 150004 510734
rect 149404 475054 150004 510498
rect 149404 474818 149586 475054
rect 149822 474818 150004 475054
rect 149404 474734 150004 474818
rect 149404 474498 149586 474734
rect 149822 474498 150004 474734
rect 149404 439054 150004 474498
rect 149404 438818 149586 439054
rect 149822 438818 150004 439054
rect 149404 438734 150004 438818
rect 149404 438498 149586 438734
rect 149822 438498 150004 438734
rect 149404 403054 150004 438498
rect 149404 402818 149586 403054
rect 149822 402818 150004 403054
rect 149404 402734 150004 402818
rect 149404 402498 149586 402734
rect 149822 402498 150004 402734
rect 149404 367054 150004 402498
rect 149404 366818 149586 367054
rect 149822 366818 150004 367054
rect 149404 366734 150004 366818
rect 149404 366498 149586 366734
rect 149822 366498 150004 366734
rect 149404 331054 150004 366498
rect 149404 330818 149586 331054
rect 149822 330818 150004 331054
rect 149404 330734 150004 330818
rect 149404 330498 149586 330734
rect 149822 330498 150004 330734
rect 149404 295054 150004 330498
rect 149404 294818 149586 295054
rect 149822 294818 150004 295054
rect 149404 294734 150004 294818
rect 149404 294498 149586 294734
rect 149822 294498 150004 294734
rect 149404 259054 150004 294498
rect 149404 258818 149586 259054
rect 149822 258818 150004 259054
rect 149404 258734 150004 258818
rect 149404 258498 149586 258734
rect 149822 258498 150004 258734
rect 149404 223054 150004 258498
rect 149404 222818 149586 223054
rect 149822 222818 150004 223054
rect 149404 222734 150004 222818
rect 149404 222498 149586 222734
rect 149822 222498 150004 222734
rect 149404 187054 150004 222498
rect 149404 186818 149586 187054
rect 149822 186818 150004 187054
rect 149404 186734 150004 186818
rect 149404 186498 149586 186734
rect 149822 186498 150004 186734
rect 149404 151054 150004 186498
rect 149404 150818 149586 151054
rect 149822 150818 150004 151054
rect 149404 150734 150004 150818
rect 149404 150498 149586 150734
rect 149822 150498 150004 150734
rect 149404 115054 150004 150498
rect 149404 114818 149586 115054
rect 149822 114818 150004 115054
rect 149404 114734 150004 114818
rect 149404 114498 149586 114734
rect 149822 114498 150004 114734
rect 149404 79054 150004 114498
rect 149404 78818 149586 79054
rect 149822 78818 150004 79054
rect 149404 78734 150004 78818
rect 149404 78498 149586 78734
rect 149822 78498 150004 78734
rect 149404 43054 150004 78498
rect 149404 42818 149586 43054
rect 149822 42818 150004 43054
rect 149404 42734 150004 42818
rect 149404 42498 149586 42734
rect 149822 42498 150004 42734
rect 149404 7054 150004 42498
rect 149404 6818 149586 7054
rect 149822 6818 150004 7054
rect 149404 6734 150004 6818
rect 149404 6498 149586 6734
rect 149822 6498 150004 6734
rect 149404 -2226 150004 6498
rect 149404 -2462 149586 -2226
rect 149822 -2462 150004 -2226
rect 149404 -2546 150004 -2462
rect 149404 -2782 149586 -2546
rect 149822 -2782 150004 -2546
rect 149404 -3744 150004 -2782
rect 153004 694654 153604 708042
rect 153004 694418 153186 694654
rect 153422 694418 153604 694654
rect 153004 694334 153604 694418
rect 153004 694098 153186 694334
rect 153422 694098 153604 694334
rect 153004 658654 153604 694098
rect 153004 658418 153186 658654
rect 153422 658418 153604 658654
rect 153004 658334 153604 658418
rect 153004 658098 153186 658334
rect 153422 658098 153604 658334
rect 153004 622654 153604 658098
rect 153004 622418 153186 622654
rect 153422 622418 153604 622654
rect 153004 622334 153604 622418
rect 153004 622098 153186 622334
rect 153422 622098 153604 622334
rect 153004 586654 153604 622098
rect 153004 586418 153186 586654
rect 153422 586418 153604 586654
rect 153004 586334 153604 586418
rect 153004 586098 153186 586334
rect 153422 586098 153604 586334
rect 153004 550654 153604 586098
rect 153004 550418 153186 550654
rect 153422 550418 153604 550654
rect 153004 550334 153604 550418
rect 153004 550098 153186 550334
rect 153422 550098 153604 550334
rect 153004 514654 153604 550098
rect 153004 514418 153186 514654
rect 153422 514418 153604 514654
rect 153004 514334 153604 514418
rect 153004 514098 153186 514334
rect 153422 514098 153604 514334
rect 153004 478654 153604 514098
rect 153004 478418 153186 478654
rect 153422 478418 153604 478654
rect 153004 478334 153604 478418
rect 153004 478098 153186 478334
rect 153422 478098 153604 478334
rect 153004 442654 153604 478098
rect 153004 442418 153186 442654
rect 153422 442418 153604 442654
rect 153004 442334 153604 442418
rect 153004 442098 153186 442334
rect 153422 442098 153604 442334
rect 153004 406654 153604 442098
rect 153004 406418 153186 406654
rect 153422 406418 153604 406654
rect 153004 406334 153604 406418
rect 153004 406098 153186 406334
rect 153422 406098 153604 406334
rect 153004 370654 153604 406098
rect 153004 370418 153186 370654
rect 153422 370418 153604 370654
rect 153004 370334 153604 370418
rect 153004 370098 153186 370334
rect 153422 370098 153604 370334
rect 153004 334654 153604 370098
rect 153004 334418 153186 334654
rect 153422 334418 153604 334654
rect 153004 334334 153604 334418
rect 153004 334098 153186 334334
rect 153422 334098 153604 334334
rect 153004 298654 153604 334098
rect 153004 298418 153186 298654
rect 153422 298418 153604 298654
rect 153004 298334 153604 298418
rect 153004 298098 153186 298334
rect 153422 298098 153604 298334
rect 153004 262654 153604 298098
rect 153004 262418 153186 262654
rect 153422 262418 153604 262654
rect 153004 262334 153604 262418
rect 153004 262098 153186 262334
rect 153422 262098 153604 262334
rect 153004 226654 153604 262098
rect 153004 226418 153186 226654
rect 153422 226418 153604 226654
rect 153004 226334 153604 226418
rect 153004 226098 153186 226334
rect 153422 226098 153604 226334
rect 153004 190654 153604 226098
rect 153004 190418 153186 190654
rect 153422 190418 153604 190654
rect 153004 190334 153604 190418
rect 153004 190098 153186 190334
rect 153422 190098 153604 190334
rect 153004 154654 153604 190098
rect 153004 154418 153186 154654
rect 153422 154418 153604 154654
rect 153004 154334 153604 154418
rect 153004 154098 153186 154334
rect 153422 154098 153604 154334
rect 153004 118654 153604 154098
rect 153004 118418 153186 118654
rect 153422 118418 153604 118654
rect 153004 118334 153604 118418
rect 153004 118098 153186 118334
rect 153422 118098 153604 118334
rect 153004 82654 153604 118098
rect 153004 82418 153186 82654
rect 153422 82418 153604 82654
rect 153004 82334 153604 82418
rect 153004 82098 153186 82334
rect 153422 82098 153604 82334
rect 153004 46654 153604 82098
rect 153004 46418 153186 46654
rect 153422 46418 153604 46654
rect 153004 46334 153604 46418
rect 153004 46098 153186 46334
rect 153422 46098 153604 46334
rect 153004 10654 153604 46098
rect 153004 10418 153186 10654
rect 153422 10418 153604 10654
rect 153004 10334 153604 10418
rect 153004 10098 153186 10334
rect 153422 10098 153604 10334
rect 153004 -4106 153604 10098
rect 153004 -4342 153186 -4106
rect 153422 -4342 153604 -4106
rect 153004 -4426 153604 -4342
rect 153004 -4662 153186 -4426
rect 153422 -4662 153604 -4426
rect 153004 -5624 153604 -4662
rect 156604 698254 157204 709922
rect 174604 711418 175204 711440
rect 174604 711182 174786 711418
rect 175022 711182 175204 711418
rect 174604 711098 175204 711182
rect 174604 710862 174786 711098
rect 175022 710862 175204 711098
rect 171004 709538 171604 709560
rect 171004 709302 171186 709538
rect 171422 709302 171604 709538
rect 171004 709218 171604 709302
rect 171004 708982 171186 709218
rect 171422 708982 171604 709218
rect 167404 707658 168004 707680
rect 167404 707422 167586 707658
rect 167822 707422 168004 707658
rect 167404 707338 168004 707422
rect 167404 707102 167586 707338
rect 167822 707102 168004 707338
rect 156604 698018 156786 698254
rect 157022 698018 157204 698254
rect 156604 697934 157204 698018
rect 156604 697698 156786 697934
rect 157022 697698 157204 697934
rect 156604 662254 157204 697698
rect 156604 662018 156786 662254
rect 157022 662018 157204 662254
rect 156604 661934 157204 662018
rect 156604 661698 156786 661934
rect 157022 661698 157204 661934
rect 156604 626254 157204 661698
rect 156604 626018 156786 626254
rect 157022 626018 157204 626254
rect 156604 625934 157204 626018
rect 156604 625698 156786 625934
rect 157022 625698 157204 625934
rect 156604 590254 157204 625698
rect 156604 590018 156786 590254
rect 157022 590018 157204 590254
rect 156604 589934 157204 590018
rect 156604 589698 156786 589934
rect 157022 589698 157204 589934
rect 156604 554254 157204 589698
rect 156604 554018 156786 554254
rect 157022 554018 157204 554254
rect 156604 553934 157204 554018
rect 156604 553698 156786 553934
rect 157022 553698 157204 553934
rect 156604 518254 157204 553698
rect 156604 518018 156786 518254
rect 157022 518018 157204 518254
rect 156604 517934 157204 518018
rect 156604 517698 156786 517934
rect 157022 517698 157204 517934
rect 156604 482254 157204 517698
rect 156604 482018 156786 482254
rect 157022 482018 157204 482254
rect 156604 481934 157204 482018
rect 156604 481698 156786 481934
rect 157022 481698 157204 481934
rect 156604 446254 157204 481698
rect 156604 446018 156786 446254
rect 157022 446018 157204 446254
rect 156604 445934 157204 446018
rect 156604 445698 156786 445934
rect 157022 445698 157204 445934
rect 156604 410254 157204 445698
rect 156604 410018 156786 410254
rect 157022 410018 157204 410254
rect 156604 409934 157204 410018
rect 156604 409698 156786 409934
rect 157022 409698 157204 409934
rect 156604 374254 157204 409698
rect 156604 374018 156786 374254
rect 157022 374018 157204 374254
rect 156604 373934 157204 374018
rect 156604 373698 156786 373934
rect 157022 373698 157204 373934
rect 156604 338254 157204 373698
rect 156604 338018 156786 338254
rect 157022 338018 157204 338254
rect 156604 337934 157204 338018
rect 156604 337698 156786 337934
rect 157022 337698 157204 337934
rect 156604 302254 157204 337698
rect 156604 302018 156786 302254
rect 157022 302018 157204 302254
rect 156604 301934 157204 302018
rect 156604 301698 156786 301934
rect 157022 301698 157204 301934
rect 156604 266254 157204 301698
rect 156604 266018 156786 266254
rect 157022 266018 157204 266254
rect 156604 265934 157204 266018
rect 156604 265698 156786 265934
rect 157022 265698 157204 265934
rect 156604 230254 157204 265698
rect 156604 230018 156786 230254
rect 157022 230018 157204 230254
rect 156604 229934 157204 230018
rect 156604 229698 156786 229934
rect 157022 229698 157204 229934
rect 156604 194254 157204 229698
rect 156604 194018 156786 194254
rect 157022 194018 157204 194254
rect 156604 193934 157204 194018
rect 156604 193698 156786 193934
rect 157022 193698 157204 193934
rect 156604 158254 157204 193698
rect 156604 158018 156786 158254
rect 157022 158018 157204 158254
rect 156604 157934 157204 158018
rect 156604 157698 156786 157934
rect 157022 157698 157204 157934
rect 156604 122254 157204 157698
rect 156604 122018 156786 122254
rect 157022 122018 157204 122254
rect 156604 121934 157204 122018
rect 156604 121698 156786 121934
rect 157022 121698 157204 121934
rect 156604 86254 157204 121698
rect 156604 86018 156786 86254
rect 157022 86018 157204 86254
rect 156604 85934 157204 86018
rect 156604 85698 156786 85934
rect 157022 85698 157204 85934
rect 156604 50254 157204 85698
rect 156604 50018 156786 50254
rect 157022 50018 157204 50254
rect 156604 49934 157204 50018
rect 156604 49698 156786 49934
rect 157022 49698 157204 49934
rect 156604 14254 157204 49698
rect 156604 14018 156786 14254
rect 157022 14018 157204 14254
rect 156604 13934 157204 14018
rect 156604 13698 156786 13934
rect 157022 13698 157204 13934
rect 138604 -7162 138786 -6926
rect 139022 -7162 139204 -6926
rect 138604 -7246 139204 -7162
rect 138604 -7482 138786 -7246
rect 139022 -7482 139204 -7246
rect 138604 -7504 139204 -7482
rect 156604 -5986 157204 13698
rect 163804 705778 164404 705800
rect 163804 705542 163986 705778
rect 164222 705542 164404 705778
rect 163804 705458 164404 705542
rect 163804 705222 163986 705458
rect 164222 705222 164404 705458
rect 163804 669454 164404 705222
rect 163804 669218 163986 669454
rect 164222 669218 164404 669454
rect 163804 669134 164404 669218
rect 163804 668898 163986 669134
rect 164222 668898 164404 669134
rect 163804 633454 164404 668898
rect 163804 633218 163986 633454
rect 164222 633218 164404 633454
rect 163804 633134 164404 633218
rect 163804 632898 163986 633134
rect 164222 632898 164404 633134
rect 163804 597454 164404 632898
rect 163804 597218 163986 597454
rect 164222 597218 164404 597454
rect 163804 597134 164404 597218
rect 163804 596898 163986 597134
rect 164222 596898 164404 597134
rect 163804 561454 164404 596898
rect 163804 561218 163986 561454
rect 164222 561218 164404 561454
rect 163804 561134 164404 561218
rect 163804 560898 163986 561134
rect 164222 560898 164404 561134
rect 163804 525454 164404 560898
rect 163804 525218 163986 525454
rect 164222 525218 164404 525454
rect 163804 525134 164404 525218
rect 163804 524898 163986 525134
rect 164222 524898 164404 525134
rect 163804 489454 164404 524898
rect 163804 489218 163986 489454
rect 164222 489218 164404 489454
rect 163804 489134 164404 489218
rect 163804 488898 163986 489134
rect 164222 488898 164404 489134
rect 163804 453454 164404 488898
rect 163804 453218 163986 453454
rect 164222 453218 164404 453454
rect 163804 453134 164404 453218
rect 163804 452898 163986 453134
rect 164222 452898 164404 453134
rect 163804 417454 164404 452898
rect 163804 417218 163986 417454
rect 164222 417218 164404 417454
rect 163804 417134 164404 417218
rect 163804 416898 163986 417134
rect 164222 416898 164404 417134
rect 163804 381454 164404 416898
rect 163804 381218 163986 381454
rect 164222 381218 164404 381454
rect 163804 381134 164404 381218
rect 163804 380898 163986 381134
rect 164222 380898 164404 381134
rect 163804 345454 164404 380898
rect 163804 345218 163986 345454
rect 164222 345218 164404 345454
rect 163804 345134 164404 345218
rect 163804 344898 163986 345134
rect 164222 344898 164404 345134
rect 163804 309454 164404 344898
rect 163804 309218 163986 309454
rect 164222 309218 164404 309454
rect 163804 309134 164404 309218
rect 163804 308898 163986 309134
rect 164222 308898 164404 309134
rect 163804 273454 164404 308898
rect 163804 273218 163986 273454
rect 164222 273218 164404 273454
rect 163804 273134 164404 273218
rect 163804 272898 163986 273134
rect 164222 272898 164404 273134
rect 163804 237454 164404 272898
rect 163804 237218 163986 237454
rect 164222 237218 164404 237454
rect 163804 237134 164404 237218
rect 163804 236898 163986 237134
rect 164222 236898 164404 237134
rect 163804 201454 164404 236898
rect 163804 201218 163986 201454
rect 164222 201218 164404 201454
rect 163804 201134 164404 201218
rect 163804 200898 163986 201134
rect 164222 200898 164404 201134
rect 163804 165454 164404 200898
rect 163804 165218 163986 165454
rect 164222 165218 164404 165454
rect 163804 165134 164404 165218
rect 163804 164898 163986 165134
rect 164222 164898 164404 165134
rect 163804 129454 164404 164898
rect 163804 129218 163986 129454
rect 164222 129218 164404 129454
rect 163804 129134 164404 129218
rect 163804 128898 163986 129134
rect 164222 128898 164404 129134
rect 163804 93454 164404 128898
rect 163804 93218 163986 93454
rect 164222 93218 164404 93454
rect 163804 93134 164404 93218
rect 163804 92898 163986 93134
rect 164222 92898 164404 93134
rect 163804 57454 164404 92898
rect 163804 57218 163986 57454
rect 164222 57218 164404 57454
rect 163804 57134 164404 57218
rect 163804 56898 163986 57134
rect 164222 56898 164404 57134
rect 163804 21454 164404 56898
rect 163804 21218 163986 21454
rect 164222 21218 164404 21454
rect 163804 21134 164404 21218
rect 163804 20898 163986 21134
rect 164222 20898 164404 21134
rect 163804 -1286 164404 20898
rect 163804 -1522 163986 -1286
rect 164222 -1522 164404 -1286
rect 163804 -1606 164404 -1522
rect 163804 -1842 163986 -1606
rect 164222 -1842 164404 -1606
rect 163804 -1864 164404 -1842
rect 167404 673054 168004 707102
rect 167404 672818 167586 673054
rect 167822 672818 168004 673054
rect 167404 672734 168004 672818
rect 167404 672498 167586 672734
rect 167822 672498 168004 672734
rect 167404 637054 168004 672498
rect 167404 636818 167586 637054
rect 167822 636818 168004 637054
rect 167404 636734 168004 636818
rect 167404 636498 167586 636734
rect 167822 636498 168004 636734
rect 167404 601054 168004 636498
rect 167404 600818 167586 601054
rect 167822 600818 168004 601054
rect 167404 600734 168004 600818
rect 167404 600498 167586 600734
rect 167822 600498 168004 600734
rect 167404 565054 168004 600498
rect 167404 564818 167586 565054
rect 167822 564818 168004 565054
rect 167404 564734 168004 564818
rect 167404 564498 167586 564734
rect 167822 564498 168004 564734
rect 167404 529054 168004 564498
rect 167404 528818 167586 529054
rect 167822 528818 168004 529054
rect 167404 528734 168004 528818
rect 167404 528498 167586 528734
rect 167822 528498 168004 528734
rect 167404 493054 168004 528498
rect 167404 492818 167586 493054
rect 167822 492818 168004 493054
rect 167404 492734 168004 492818
rect 167404 492498 167586 492734
rect 167822 492498 168004 492734
rect 167404 457054 168004 492498
rect 167404 456818 167586 457054
rect 167822 456818 168004 457054
rect 167404 456734 168004 456818
rect 167404 456498 167586 456734
rect 167822 456498 168004 456734
rect 167404 421054 168004 456498
rect 167404 420818 167586 421054
rect 167822 420818 168004 421054
rect 167404 420734 168004 420818
rect 167404 420498 167586 420734
rect 167822 420498 168004 420734
rect 167404 385054 168004 420498
rect 167404 384818 167586 385054
rect 167822 384818 168004 385054
rect 167404 384734 168004 384818
rect 167404 384498 167586 384734
rect 167822 384498 168004 384734
rect 167404 349054 168004 384498
rect 167404 348818 167586 349054
rect 167822 348818 168004 349054
rect 167404 348734 168004 348818
rect 167404 348498 167586 348734
rect 167822 348498 168004 348734
rect 167404 313054 168004 348498
rect 167404 312818 167586 313054
rect 167822 312818 168004 313054
rect 167404 312734 168004 312818
rect 167404 312498 167586 312734
rect 167822 312498 168004 312734
rect 167404 277054 168004 312498
rect 167404 276818 167586 277054
rect 167822 276818 168004 277054
rect 167404 276734 168004 276818
rect 167404 276498 167586 276734
rect 167822 276498 168004 276734
rect 167404 241054 168004 276498
rect 167404 240818 167586 241054
rect 167822 240818 168004 241054
rect 167404 240734 168004 240818
rect 167404 240498 167586 240734
rect 167822 240498 168004 240734
rect 167404 205054 168004 240498
rect 167404 204818 167586 205054
rect 167822 204818 168004 205054
rect 167404 204734 168004 204818
rect 167404 204498 167586 204734
rect 167822 204498 168004 204734
rect 167404 169054 168004 204498
rect 167404 168818 167586 169054
rect 167822 168818 168004 169054
rect 167404 168734 168004 168818
rect 167404 168498 167586 168734
rect 167822 168498 168004 168734
rect 167404 133054 168004 168498
rect 167404 132818 167586 133054
rect 167822 132818 168004 133054
rect 167404 132734 168004 132818
rect 167404 132498 167586 132734
rect 167822 132498 168004 132734
rect 167404 97054 168004 132498
rect 167404 96818 167586 97054
rect 167822 96818 168004 97054
rect 167404 96734 168004 96818
rect 167404 96498 167586 96734
rect 167822 96498 168004 96734
rect 167404 61054 168004 96498
rect 167404 60818 167586 61054
rect 167822 60818 168004 61054
rect 167404 60734 168004 60818
rect 167404 60498 167586 60734
rect 167822 60498 168004 60734
rect 167404 25054 168004 60498
rect 167404 24818 167586 25054
rect 167822 24818 168004 25054
rect 167404 24734 168004 24818
rect 167404 24498 167586 24734
rect 167822 24498 168004 24734
rect 167404 -3166 168004 24498
rect 167404 -3402 167586 -3166
rect 167822 -3402 168004 -3166
rect 167404 -3486 168004 -3402
rect 167404 -3722 167586 -3486
rect 167822 -3722 168004 -3486
rect 167404 -3744 168004 -3722
rect 171004 676654 171604 708982
rect 171004 676418 171186 676654
rect 171422 676418 171604 676654
rect 171004 676334 171604 676418
rect 171004 676098 171186 676334
rect 171422 676098 171604 676334
rect 171004 640654 171604 676098
rect 171004 640418 171186 640654
rect 171422 640418 171604 640654
rect 171004 640334 171604 640418
rect 171004 640098 171186 640334
rect 171422 640098 171604 640334
rect 171004 604654 171604 640098
rect 171004 604418 171186 604654
rect 171422 604418 171604 604654
rect 171004 604334 171604 604418
rect 171004 604098 171186 604334
rect 171422 604098 171604 604334
rect 171004 568654 171604 604098
rect 171004 568418 171186 568654
rect 171422 568418 171604 568654
rect 171004 568334 171604 568418
rect 171004 568098 171186 568334
rect 171422 568098 171604 568334
rect 171004 532654 171604 568098
rect 171004 532418 171186 532654
rect 171422 532418 171604 532654
rect 171004 532334 171604 532418
rect 171004 532098 171186 532334
rect 171422 532098 171604 532334
rect 171004 496654 171604 532098
rect 171004 496418 171186 496654
rect 171422 496418 171604 496654
rect 171004 496334 171604 496418
rect 171004 496098 171186 496334
rect 171422 496098 171604 496334
rect 171004 460654 171604 496098
rect 171004 460418 171186 460654
rect 171422 460418 171604 460654
rect 171004 460334 171604 460418
rect 171004 460098 171186 460334
rect 171422 460098 171604 460334
rect 171004 424654 171604 460098
rect 171004 424418 171186 424654
rect 171422 424418 171604 424654
rect 171004 424334 171604 424418
rect 171004 424098 171186 424334
rect 171422 424098 171604 424334
rect 171004 388654 171604 424098
rect 171004 388418 171186 388654
rect 171422 388418 171604 388654
rect 171004 388334 171604 388418
rect 171004 388098 171186 388334
rect 171422 388098 171604 388334
rect 171004 352654 171604 388098
rect 171004 352418 171186 352654
rect 171422 352418 171604 352654
rect 171004 352334 171604 352418
rect 171004 352098 171186 352334
rect 171422 352098 171604 352334
rect 171004 316654 171604 352098
rect 171004 316418 171186 316654
rect 171422 316418 171604 316654
rect 171004 316334 171604 316418
rect 171004 316098 171186 316334
rect 171422 316098 171604 316334
rect 171004 280654 171604 316098
rect 171004 280418 171186 280654
rect 171422 280418 171604 280654
rect 171004 280334 171604 280418
rect 171004 280098 171186 280334
rect 171422 280098 171604 280334
rect 171004 244654 171604 280098
rect 171004 244418 171186 244654
rect 171422 244418 171604 244654
rect 171004 244334 171604 244418
rect 171004 244098 171186 244334
rect 171422 244098 171604 244334
rect 171004 208654 171604 244098
rect 171004 208418 171186 208654
rect 171422 208418 171604 208654
rect 171004 208334 171604 208418
rect 171004 208098 171186 208334
rect 171422 208098 171604 208334
rect 171004 172654 171604 208098
rect 171004 172418 171186 172654
rect 171422 172418 171604 172654
rect 171004 172334 171604 172418
rect 171004 172098 171186 172334
rect 171422 172098 171604 172334
rect 171004 136654 171604 172098
rect 171004 136418 171186 136654
rect 171422 136418 171604 136654
rect 171004 136334 171604 136418
rect 171004 136098 171186 136334
rect 171422 136098 171604 136334
rect 171004 100654 171604 136098
rect 171004 100418 171186 100654
rect 171422 100418 171604 100654
rect 171004 100334 171604 100418
rect 171004 100098 171186 100334
rect 171422 100098 171604 100334
rect 171004 64654 171604 100098
rect 171004 64418 171186 64654
rect 171422 64418 171604 64654
rect 171004 64334 171604 64418
rect 171004 64098 171186 64334
rect 171422 64098 171604 64334
rect 171004 28654 171604 64098
rect 171004 28418 171186 28654
rect 171422 28418 171604 28654
rect 171004 28334 171604 28418
rect 171004 28098 171186 28334
rect 171422 28098 171604 28334
rect 171004 -5046 171604 28098
rect 171004 -5282 171186 -5046
rect 171422 -5282 171604 -5046
rect 171004 -5366 171604 -5282
rect 171004 -5602 171186 -5366
rect 171422 -5602 171604 -5366
rect 171004 -5624 171604 -5602
rect 174604 680254 175204 710862
rect 192604 710478 193204 711440
rect 192604 710242 192786 710478
rect 193022 710242 193204 710478
rect 192604 710158 193204 710242
rect 192604 709922 192786 710158
rect 193022 709922 193204 710158
rect 189004 708598 189604 709560
rect 189004 708362 189186 708598
rect 189422 708362 189604 708598
rect 189004 708278 189604 708362
rect 189004 708042 189186 708278
rect 189422 708042 189604 708278
rect 185404 706718 186004 707680
rect 185404 706482 185586 706718
rect 185822 706482 186004 706718
rect 185404 706398 186004 706482
rect 185404 706162 185586 706398
rect 185822 706162 186004 706398
rect 174604 680018 174786 680254
rect 175022 680018 175204 680254
rect 174604 679934 175204 680018
rect 174604 679698 174786 679934
rect 175022 679698 175204 679934
rect 174604 644254 175204 679698
rect 174604 644018 174786 644254
rect 175022 644018 175204 644254
rect 174604 643934 175204 644018
rect 174604 643698 174786 643934
rect 175022 643698 175204 643934
rect 174604 608254 175204 643698
rect 174604 608018 174786 608254
rect 175022 608018 175204 608254
rect 174604 607934 175204 608018
rect 174604 607698 174786 607934
rect 175022 607698 175204 607934
rect 174604 572254 175204 607698
rect 174604 572018 174786 572254
rect 175022 572018 175204 572254
rect 174604 571934 175204 572018
rect 174604 571698 174786 571934
rect 175022 571698 175204 571934
rect 174604 536254 175204 571698
rect 174604 536018 174786 536254
rect 175022 536018 175204 536254
rect 174604 535934 175204 536018
rect 174604 535698 174786 535934
rect 175022 535698 175204 535934
rect 174604 500254 175204 535698
rect 174604 500018 174786 500254
rect 175022 500018 175204 500254
rect 174604 499934 175204 500018
rect 174604 499698 174786 499934
rect 175022 499698 175204 499934
rect 174604 464254 175204 499698
rect 174604 464018 174786 464254
rect 175022 464018 175204 464254
rect 174604 463934 175204 464018
rect 174604 463698 174786 463934
rect 175022 463698 175204 463934
rect 174604 428254 175204 463698
rect 174604 428018 174786 428254
rect 175022 428018 175204 428254
rect 174604 427934 175204 428018
rect 174604 427698 174786 427934
rect 175022 427698 175204 427934
rect 174604 392254 175204 427698
rect 174604 392018 174786 392254
rect 175022 392018 175204 392254
rect 174604 391934 175204 392018
rect 174604 391698 174786 391934
rect 175022 391698 175204 391934
rect 174604 356254 175204 391698
rect 174604 356018 174786 356254
rect 175022 356018 175204 356254
rect 174604 355934 175204 356018
rect 174604 355698 174786 355934
rect 175022 355698 175204 355934
rect 174604 320254 175204 355698
rect 174604 320018 174786 320254
rect 175022 320018 175204 320254
rect 174604 319934 175204 320018
rect 174604 319698 174786 319934
rect 175022 319698 175204 319934
rect 174604 284254 175204 319698
rect 174604 284018 174786 284254
rect 175022 284018 175204 284254
rect 174604 283934 175204 284018
rect 174604 283698 174786 283934
rect 175022 283698 175204 283934
rect 174604 248254 175204 283698
rect 174604 248018 174786 248254
rect 175022 248018 175204 248254
rect 174604 247934 175204 248018
rect 174604 247698 174786 247934
rect 175022 247698 175204 247934
rect 174604 212254 175204 247698
rect 174604 212018 174786 212254
rect 175022 212018 175204 212254
rect 174604 211934 175204 212018
rect 174604 211698 174786 211934
rect 175022 211698 175204 211934
rect 174604 176254 175204 211698
rect 174604 176018 174786 176254
rect 175022 176018 175204 176254
rect 174604 175934 175204 176018
rect 174604 175698 174786 175934
rect 175022 175698 175204 175934
rect 174604 140254 175204 175698
rect 174604 140018 174786 140254
rect 175022 140018 175204 140254
rect 174604 139934 175204 140018
rect 174604 139698 174786 139934
rect 175022 139698 175204 139934
rect 174604 104254 175204 139698
rect 174604 104018 174786 104254
rect 175022 104018 175204 104254
rect 174604 103934 175204 104018
rect 174604 103698 174786 103934
rect 175022 103698 175204 103934
rect 174604 68254 175204 103698
rect 174604 68018 174786 68254
rect 175022 68018 175204 68254
rect 174604 67934 175204 68018
rect 174604 67698 174786 67934
rect 175022 67698 175204 67934
rect 174604 32254 175204 67698
rect 174604 32018 174786 32254
rect 175022 32018 175204 32254
rect 174604 31934 175204 32018
rect 174604 31698 174786 31934
rect 175022 31698 175204 31934
rect 156604 -6222 156786 -5986
rect 157022 -6222 157204 -5986
rect 156604 -6306 157204 -6222
rect 156604 -6542 156786 -6306
rect 157022 -6542 157204 -6306
rect 156604 -7504 157204 -6542
rect 174604 -6926 175204 31698
rect 181804 704838 182404 705800
rect 181804 704602 181986 704838
rect 182222 704602 182404 704838
rect 181804 704518 182404 704602
rect 181804 704282 181986 704518
rect 182222 704282 182404 704518
rect 181804 687454 182404 704282
rect 181804 687218 181986 687454
rect 182222 687218 182404 687454
rect 181804 687134 182404 687218
rect 181804 686898 181986 687134
rect 182222 686898 182404 687134
rect 181804 651454 182404 686898
rect 181804 651218 181986 651454
rect 182222 651218 182404 651454
rect 181804 651134 182404 651218
rect 181804 650898 181986 651134
rect 182222 650898 182404 651134
rect 181804 615454 182404 650898
rect 181804 615218 181986 615454
rect 182222 615218 182404 615454
rect 181804 615134 182404 615218
rect 181804 614898 181986 615134
rect 182222 614898 182404 615134
rect 181804 579454 182404 614898
rect 181804 579218 181986 579454
rect 182222 579218 182404 579454
rect 181804 579134 182404 579218
rect 181804 578898 181986 579134
rect 182222 578898 182404 579134
rect 181804 543454 182404 578898
rect 181804 543218 181986 543454
rect 182222 543218 182404 543454
rect 181804 543134 182404 543218
rect 181804 542898 181986 543134
rect 182222 542898 182404 543134
rect 181804 507454 182404 542898
rect 181804 507218 181986 507454
rect 182222 507218 182404 507454
rect 181804 507134 182404 507218
rect 181804 506898 181986 507134
rect 182222 506898 182404 507134
rect 181804 471454 182404 506898
rect 181804 471218 181986 471454
rect 182222 471218 182404 471454
rect 181804 471134 182404 471218
rect 181804 470898 181986 471134
rect 182222 470898 182404 471134
rect 181804 435454 182404 470898
rect 181804 435218 181986 435454
rect 182222 435218 182404 435454
rect 181804 435134 182404 435218
rect 181804 434898 181986 435134
rect 182222 434898 182404 435134
rect 181804 399454 182404 434898
rect 181804 399218 181986 399454
rect 182222 399218 182404 399454
rect 181804 399134 182404 399218
rect 181804 398898 181986 399134
rect 182222 398898 182404 399134
rect 181804 363454 182404 398898
rect 181804 363218 181986 363454
rect 182222 363218 182404 363454
rect 181804 363134 182404 363218
rect 181804 362898 181986 363134
rect 182222 362898 182404 363134
rect 181804 327454 182404 362898
rect 181804 327218 181986 327454
rect 182222 327218 182404 327454
rect 181804 327134 182404 327218
rect 181804 326898 181986 327134
rect 182222 326898 182404 327134
rect 181804 291454 182404 326898
rect 181804 291218 181986 291454
rect 182222 291218 182404 291454
rect 181804 291134 182404 291218
rect 181804 290898 181986 291134
rect 182222 290898 182404 291134
rect 181804 255454 182404 290898
rect 181804 255218 181986 255454
rect 182222 255218 182404 255454
rect 181804 255134 182404 255218
rect 181804 254898 181986 255134
rect 182222 254898 182404 255134
rect 181804 219454 182404 254898
rect 181804 219218 181986 219454
rect 182222 219218 182404 219454
rect 181804 219134 182404 219218
rect 181804 218898 181986 219134
rect 182222 218898 182404 219134
rect 181804 183454 182404 218898
rect 181804 183218 181986 183454
rect 182222 183218 182404 183454
rect 181804 183134 182404 183218
rect 181804 182898 181986 183134
rect 182222 182898 182404 183134
rect 181804 147454 182404 182898
rect 181804 147218 181986 147454
rect 182222 147218 182404 147454
rect 181804 147134 182404 147218
rect 181804 146898 181986 147134
rect 182222 146898 182404 147134
rect 181804 111454 182404 146898
rect 181804 111218 181986 111454
rect 182222 111218 182404 111454
rect 181804 111134 182404 111218
rect 181804 110898 181986 111134
rect 182222 110898 182404 111134
rect 181804 75454 182404 110898
rect 181804 75218 181986 75454
rect 182222 75218 182404 75454
rect 181804 75134 182404 75218
rect 181804 74898 181986 75134
rect 182222 74898 182404 75134
rect 181804 39454 182404 74898
rect 181804 39218 181986 39454
rect 182222 39218 182404 39454
rect 181804 39134 182404 39218
rect 181804 38898 181986 39134
rect 182222 38898 182404 39134
rect 181804 3454 182404 38898
rect 181804 3218 181986 3454
rect 182222 3218 182404 3454
rect 181804 3134 182404 3218
rect 181804 2898 181986 3134
rect 182222 2898 182404 3134
rect 181804 -346 182404 2898
rect 181804 -582 181986 -346
rect 182222 -582 182404 -346
rect 181804 -666 182404 -582
rect 181804 -902 181986 -666
rect 182222 -902 182404 -666
rect 181804 -1864 182404 -902
rect 185404 691054 186004 706162
rect 185404 690818 185586 691054
rect 185822 690818 186004 691054
rect 185404 690734 186004 690818
rect 185404 690498 185586 690734
rect 185822 690498 186004 690734
rect 185404 655054 186004 690498
rect 185404 654818 185586 655054
rect 185822 654818 186004 655054
rect 185404 654734 186004 654818
rect 185404 654498 185586 654734
rect 185822 654498 186004 654734
rect 185404 619054 186004 654498
rect 185404 618818 185586 619054
rect 185822 618818 186004 619054
rect 185404 618734 186004 618818
rect 185404 618498 185586 618734
rect 185822 618498 186004 618734
rect 185404 583054 186004 618498
rect 185404 582818 185586 583054
rect 185822 582818 186004 583054
rect 185404 582734 186004 582818
rect 185404 582498 185586 582734
rect 185822 582498 186004 582734
rect 185404 547054 186004 582498
rect 185404 546818 185586 547054
rect 185822 546818 186004 547054
rect 185404 546734 186004 546818
rect 185404 546498 185586 546734
rect 185822 546498 186004 546734
rect 185404 511054 186004 546498
rect 185404 510818 185586 511054
rect 185822 510818 186004 511054
rect 185404 510734 186004 510818
rect 185404 510498 185586 510734
rect 185822 510498 186004 510734
rect 185404 475054 186004 510498
rect 185404 474818 185586 475054
rect 185822 474818 186004 475054
rect 185404 474734 186004 474818
rect 185404 474498 185586 474734
rect 185822 474498 186004 474734
rect 185404 439054 186004 474498
rect 185404 438818 185586 439054
rect 185822 438818 186004 439054
rect 185404 438734 186004 438818
rect 185404 438498 185586 438734
rect 185822 438498 186004 438734
rect 185404 403054 186004 438498
rect 185404 402818 185586 403054
rect 185822 402818 186004 403054
rect 185404 402734 186004 402818
rect 185404 402498 185586 402734
rect 185822 402498 186004 402734
rect 185404 367054 186004 402498
rect 185404 366818 185586 367054
rect 185822 366818 186004 367054
rect 185404 366734 186004 366818
rect 185404 366498 185586 366734
rect 185822 366498 186004 366734
rect 185404 331054 186004 366498
rect 185404 330818 185586 331054
rect 185822 330818 186004 331054
rect 185404 330734 186004 330818
rect 185404 330498 185586 330734
rect 185822 330498 186004 330734
rect 185404 295054 186004 330498
rect 185404 294818 185586 295054
rect 185822 294818 186004 295054
rect 185404 294734 186004 294818
rect 185404 294498 185586 294734
rect 185822 294498 186004 294734
rect 185404 259054 186004 294498
rect 185404 258818 185586 259054
rect 185822 258818 186004 259054
rect 185404 258734 186004 258818
rect 185404 258498 185586 258734
rect 185822 258498 186004 258734
rect 185404 223054 186004 258498
rect 185404 222818 185586 223054
rect 185822 222818 186004 223054
rect 185404 222734 186004 222818
rect 185404 222498 185586 222734
rect 185822 222498 186004 222734
rect 185404 187054 186004 222498
rect 185404 186818 185586 187054
rect 185822 186818 186004 187054
rect 185404 186734 186004 186818
rect 185404 186498 185586 186734
rect 185822 186498 186004 186734
rect 185404 151054 186004 186498
rect 185404 150818 185586 151054
rect 185822 150818 186004 151054
rect 185404 150734 186004 150818
rect 185404 150498 185586 150734
rect 185822 150498 186004 150734
rect 185404 115054 186004 150498
rect 185404 114818 185586 115054
rect 185822 114818 186004 115054
rect 185404 114734 186004 114818
rect 185404 114498 185586 114734
rect 185822 114498 186004 114734
rect 185404 79054 186004 114498
rect 185404 78818 185586 79054
rect 185822 78818 186004 79054
rect 185404 78734 186004 78818
rect 185404 78498 185586 78734
rect 185822 78498 186004 78734
rect 185404 43054 186004 78498
rect 185404 42818 185586 43054
rect 185822 42818 186004 43054
rect 185404 42734 186004 42818
rect 185404 42498 185586 42734
rect 185822 42498 186004 42734
rect 185404 7054 186004 42498
rect 185404 6818 185586 7054
rect 185822 6818 186004 7054
rect 185404 6734 186004 6818
rect 185404 6498 185586 6734
rect 185822 6498 186004 6734
rect 185404 -2226 186004 6498
rect 185404 -2462 185586 -2226
rect 185822 -2462 186004 -2226
rect 185404 -2546 186004 -2462
rect 185404 -2782 185586 -2546
rect 185822 -2782 186004 -2546
rect 185404 -3744 186004 -2782
rect 189004 694654 189604 708042
rect 189004 694418 189186 694654
rect 189422 694418 189604 694654
rect 189004 694334 189604 694418
rect 189004 694098 189186 694334
rect 189422 694098 189604 694334
rect 189004 658654 189604 694098
rect 189004 658418 189186 658654
rect 189422 658418 189604 658654
rect 189004 658334 189604 658418
rect 189004 658098 189186 658334
rect 189422 658098 189604 658334
rect 189004 622654 189604 658098
rect 189004 622418 189186 622654
rect 189422 622418 189604 622654
rect 189004 622334 189604 622418
rect 189004 622098 189186 622334
rect 189422 622098 189604 622334
rect 189004 586654 189604 622098
rect 189004 586418 189186 586654
rect 189422 586418 189604 586654
rect 189004 586334 189604 586418
rect 189004 586098 189186 586334
rect 189422 586098 189604 586334
rect 189004 550654 189604 586098
rect 189004 550418 189186 550654
rect 189422 550418 189604 550654
rect 189004 550334 189604 550418
rect 189004 550098 189186 550334
rect 189422 550098 189604 550334
rect 189004 514654 189604 550098
rect 189004 514418 189186 514654
rect 189422 514418 189604 514654
rect 189004 514334 189604 514418
rect 189004 514098 189186 514334
rect 189422 514098 189604 514334
rect 189004 478654 189604 514098
rect 189004 478418 189186 478654
rect 189422 478418 189604 478654
rect 189004 478334 189604 478418
rect 189004 478098 189186 478334
rect 189422 478098 189604 478334
rect 189004 442654 189604 478098
rect 189004 442418 189186 442654
rect 189422 442418 189604 442654
rect 189004 442334 189604 442418
rect 189004 442098 189186 442334
rect 189422 442098 189604 442334
rect 189004 406654 189604 442098
rect 189004 406418 189186 406654
rect 189422 406418 189604 406654
rect 189004 406334 189604 406418
rect 189004 406098 189186 406334
rect 189422 406098 189604 406334
rect 189004 370654 189604 406098
rect 189004 370418 189186 370654
rect 189422 370418 189604 370654
rect 189004 370334 189604 370418
rect 189004 370098 189186 370334
rect 189422 370098 189604 370334
rect 189004 334654 189604 370098
rect 189004 334418 189186 334654
rect 189422 334418 189604 334654
rect 189004 334334 189604 334418
rect 189004 334098 189186 334334
rect 189422 334098 189604 334334
rect 189004 298654 189604 334098
rect 189004 298418 189186 298654
rect 189422 298418 189604 298654
rect 189004 298334 189604 298418
rect 189004 298098 189186 298334
rect 189422 298098 189604 298334
rect 189004 262654 189604 298098
rect 189004 262418 189186 262654
rect 189422 262418 189604 262654
rect 189004 262334 189604 262418
rect 189004 262098 189186 262334
rect 189422 262098 189604 262334
rect 189004 226654 189604 262098
rect 189004 226418 189186 226654
rect 189422 226418 189604 226654
rect 189004 226334 189604 226418
rect 189004 226098 189186 226334
rect 189422 226098 189604 226334
rect 189004 190654 189604 226098
rect 189004 190418 189186 190654
rect 189422 190418 189604 190654
rect 189004 190334 189604 190418
rect 189004 190098 189186 190334
rect 189422 190098 189604 190334
rect 189004 154654 189604 190098
rect 189004 154418 189186 154654
rect 189422 154418 189604 154654
rect 189004 154334 189604 154418
rect 189004 154098 189186 154334
rect 189422 154098 189604 154334
rect 189004 118654 189604 154098
rect 189004 118418 189186 118654
rect 189422 118418 189604 118654
rect 189004 118334 189604 118418
rect 189004 118098 189186 118334
rect 189422 118098 189604 118334
rect 189004 82654 189604 118098
rect 189004 82418 189186 82654
rect 189422 82418 189604 82654
rect 189004 82334 189604 82418
rect 189004 82098 189186 82334
rect 189422 82098 189604 82334
rect 189004 46654 189604 82098
rect 189004 46418 189186 46654
rect 189422 46418 189604 46654
rect 189004 46334 189604 46418
rect 189004 46098 189186 46334
rect 189422 46098 189604 46334
rect 189004 10654 189604 46098
rect 189004 10418 189186 10654
rect 189422 10418 189604 10654
rect 189004 10334 189604 10418
rect 189004 10098 189186 10334
rect 189422 10098 189604 10334
rect 189004 -4106 189604 10098
rect 189004 -4342 189186 -4106
rect 189422 -4342 189604 -4106
rect 189004 -4426 189604 -4342
rect 189004 -4662 189186 -4426
rect 189422 -4662 189604 -4426
rect 189004 -5624 189604 -4662
rect 192604 698254 193204 709922
rect 210604 711418 211204 711440
rect 210604 711182 210786 711418
rect 211022 711182 211204 711418
rect 210604 711098 211204 711182
rect 210604 710862 210786 711098
rect 211022 710862 211204 711098
rect 207004 709538 207604 709560
rect 207004 709302 207186 709538
rect 207422 709302 207604 709538
rect 207004 709218 207604 709302
rect 207004 708982 207186 709218
rect 207422 708982 207604 709218
rect 203404 707658 204004 707680
rect 203404 707422 203586 707658
rect 203822 707422 204004 707658
rect 203404 707338 204004 707422
rect 203404 707102 203586 707338
rect 203822 707102 204004 707338
rect 192604 698018 192786 698254
rect 193022 698018 193204 698254
rect 192604 697934 193204 698018
rect 192604 697698 192786 697934
rect 193022 697698 193204 697934
rect 192604 662254 193204 697698
rect 192604 662018 192786 662254
rect 193022 662018 193204 662254
rect 192604 661934 193204 662018
rect 192604 661698 192786 661934
rect 193022 661698 193204 661934
rect 192604 626254 193204 661698
rect 192604 626018 192786 626254
rect 193022 626018 193204 626254
rect 192604 625934 193204 626018
rect 192604 625698 192786 625934
rect 193022 625698 193204 625934
rect 192604 590254 193204 625698
rect 192604 590018 192786 590254
rect 193022 590018 193204 590254
rect 192604 589934 193204 590018
rect 192604 589698 192786 589934
rect 193022 589698 193204 589934
rect 192604 554254 193204 589698
rect 192604 554018 192786 554254
rect 193022 554018 193204 554254
rect 192604 553934 193204 554018
rect 192604 553698 192786 553934
rect 193022 553698 193204 553934
rect 192604 518254 193204 553698
rect 192604 518018 192786 518254
rect 193022 518018 193204 518254
rect 192604 517934 193204 518018
rect 192604 517698 192786 517934
rect 193022 517698 193204 517934
rect 192604 482254 193204 517698
rect 192604 482018 192786 482254
rect 193022 482018 193204 482254
rect 192604 481934 193204 482018
rect 192604 481698 192786 481934
rect 193022 481698 193204 481934
rect 192604 446254 193204 481698
rect 192604 446018 192786 446254
rect 193022 446018 193204 446254
rect 192604 445934 193204 446018
rect 192604 445698 192786 445934
rect 193022 445698 193204 445934
rect 192604 410254 193204 445698
rect 192604 410018 192786 410254
rect 193022 410018 193204 410254
rect 192604 409934 193204 410018
rect 192604 409698 192786 409934
rect 193022 409698 193204 409934
rect 192604 374254 193204 409698
rect 192604 374018 192786 374254
rect 193022 374018 193204 374254
rect 192604 373934 193204 374018
rect 192604 373698 192786 373934
rect 193022 373698 193204 373934
rect 192604 338254 193204 373698
rect 192604 338018 192786 338254
rect 193022 338018 193204 338254
rect 192604 337934 193204 338018
rect 192604 337698 192786 337934
rect 193022 337698 193204 337934
rect 192604 302254 193204 337698
rect 192604 302018 192786 302254
rect 193022 302018 193204 302254
rect 192604 301934 193204 302018
rect 192604 301698 192786 301934
rect 193022 301698 193204 301934
rect 192604 266254 193204 301698
rect 192604 266018 192786 266254
rect 193022 266018 193204 266254
rect 192604 265934 193204 266018
rect 192604 265698 192786 265934
rect 193022 265698 193204 265934
rect 192604 230254 193204 265698
rect 192604 230018 192786 230254
rect 193022 230018 193204 230254
rect 192604 229934 193204 230018
rect 192604 229698 192786 229934
rect 193022 229698 193204 229934
rect 192604 194254 193204 229698
rect 192604 194018 192786 194254
rect 193022 194018 193204 194254
rect 192604 193934 193204 194018
rect 192604 193698 192786 193934
rect 193022 193698 193204 193934
rect 192604 158254 193204 193698
rect 192604 158018 192786 158254
rect 193022 158018 193204 158254
rect 192604 157934 193204 158018
rect 192604 157698 192786 157934
rect 193022 157698 193204 157934
rect 192604 122254 193204 157698
rect 192604 122018 192786 122254
rect 193022 122018 193204 122254
rect 192604 121934 193204 122018
rect 192604 121698 192786 121934
rect 193022 121698 193204 121934
rect 192604 86254 193204 121698
rect 192604 86018 192786 86254
rect 193022 86018 193204 86254
rect 192604 85934 193204 86018
rect 192604 85698 192786 85934
rect 193022 85698 193204 85934
rect 192604 50254 193204 85698
rect 192604 50018 192786 50254
rect 193022 50018 193204 50254
rect 192604 49934 193204 50018
rect 192604 49698 192786 49934
rect 193022 49698 193204 49934
rect 192604 14254 193204 49698
rect 192604 14018 192786 14254
rect 193022 14018 193204 14254
rect 192604 13934 193204 14018
rect 192604 13698 192786 13934
rect 193022 13698 193204 13934
rect 174604 -7162 174786 -6926
rect 175022 -7162 175204 -6926
rect 174604 -7246 175204 -7162
rect 174604 -7482 174786 -7246
rect 175022 -7482 175204 -7246
rect 174604 -7504 175204 -7482
rect 192604 -5986 193204 13698
rect 199804 705778 200404 705800
rect 199804 705542 199986 705778
rect 200222 705542 200404 705778
rect 199804 705458 200404 705542
rect 199804 705222 199986 705458
rect 200222 705222 200404 705458
rect 199804 669454 200404 705222
rect 199804 669218 199986 669454
rect 200222 669218 200404 669454
rect 199804 669134 200404 669218
rect 199804 668898 199986 669134
rect 200222 668898 200404 669134
rect 199804 633454 200404 668898
rect 199804 633218 199986 633454
rect 200222 633218 200404 633454
rect 199804 633134 200404 633218
rect 199804 632898 199986 633134
rect 200222 632898 200404 633134
rect 199804 597454 200404 632898
rect 199804 597218 199986 597454
rect 200222 597218 200404 597454
rect 199804 597134 200404 597218
rect 199804 596898 199986 597134
rect 200222 596898 200404 597134
rect 199804 561454 200404 596898
rect 199804 561218 199986 561454
rect 200222 561218 200404 561454
rect 199804 561134 200404 561218
rect 199804 560898 199986 561134
rect 200222 560898 200404 561134
rect 199804 525454 200404 560898
rect 199804 525218 199986 525454
rect 200222 525218 200404 525454
rect 199804 525134 200404 525218
rect 199804 524898 199986 525134
rect 200222 524898 200404 525134
rect 199804 489454 200404 524898
rect 199804 489218 199986 489454
rect 200222 489218 200404 489454
rect 199804 489134 200404 489218
rect 199804 488898 199986 489134
rect 200222 488898 200404 489134
rect 199804 453454 200404 488898
rect 199804 453218 199986 453454
rect 200222 453218 200404 453454
rect 199804 453134 200404 453218
rect 199804 452898 199986 453134
rect 200222 452898 200404 453134
rect 199804 417454 200404 452898
rect 199804 417218 199986 417454
rect 200222 417218 200404 417454
rect 199804 417134 200404 417218
rect 199804 416898 199986 417134
rect 200222 416898 200404 417134
rect 199804 381454 200404 416898
rect 199804 381218 199986 381454
rect 200222 381218 200404 381454
rect 199804 381134 200404 381218
rect 199804 380898 199986 381134
rect 200222 380898 200404 381134
rect 199804 345454 200404 380898
rect 199804 345218 199986 345454
rect 200222 345218 200404 345454
rect 199804 345134 200404 345218
rect 199804 344898 199986 345134
rect 200222 344898 200404 345134
rect 199804 309454 200404 344898
rect 199804 309218 199986 309454
rect 200222 309218 200404 309454
rect 199804 309134 200404 309218
rect 199804 308898 199986 309134
rect 200222 308898 200404 309134
rect 199804 273454 200404 308898
rect 199804 273218 199986 273454
rect 200222 273218 200404 273454
rect 199804 273134 200404 273218
rect 199804 272898 199986 273134
rect 200222 272898 200404 273134
rect 199804 237454 200404 272898
rect 199804 237218 199986 237454
rect 200222 237218 200404 237454
rect 199804 237134 200404 237218
rect 199804 236898 199986 237134
rect 200222 236898 200404 237134
rect 199804 201454 200404 236898
rect 199804 201218 199986 201454
rect 200222 201218 200404 201454
rect 199804 201134 200404 201218
rect 199804 200898 199986 201134
rect 200222 200898 200404 201134
rect 199804 165454 200404 200898
rect 199804 165218 199986 165454
rect 200222 165218 200404 165454
rect 199804 165134 200404 165218
rect 199804 164898 199986 165134
rect 200222 164898 200404 165134
rect 199804 129454 200404 164898
rect 199804 129218 199986 129454
rect 200222 129218 200404 129454
rect 199804 129134 200404 129218
rect 199804 128898 199986 129134
rect 200222 128898 200404 129134
rect 199804 93454 200404 128898
rect 199804 93218 199986 93454
rect 200222 93218 200404 93454
rect 199804 93134 200404 93218
rect 199804 92898 199986 93134
rect 200222 92898 200404 93134
rect 199804 57454 200404 92898
rect 199804 57218 199986 57454
rect 200222 57218 200404 57454
rect 199804 57134 200404 57218
rect 199804 56898 199986 57134
rect 200222 56898 200404 57134
rect 199804 21454 200404 56898
rect 199804 21218 199986 21454
rect 200222 21218 200404 21454
rect 199804 21134 200404 21218
rect 199804 20898 199986 21134
rect 200222 20898 200404 21134
rect 199804 -1286 200404 20898
rect 199804 -1522 199986 -1286
rect 200222 -1522 200404 -1286
rect 199804 -1606 200404 -1522
rect 199804 -1842 199986 -1606
rect 200222 -1842 200404 -1606
rect 199804 -1864 200404 -1842
rect 203404 673054 204004 707102
rect 203404 672818 203586 673054
rect 203822 672818 204004 673054
rect 203404 672734 204004 672818
rect 203404 672498 203586 672734
rect 203822 672498 204004 672734
rect 203404 637054 204004 672498
rect 203404 636818 203586 637054
rect 203822 636818 204004 637054
rect 203404 636734 204004 636818
rect 203404 636498 203586 636734
rect 203822 636498 204004 636734
rect 203404 601054 204004 636498
rect 203404 600818 203586 601054
rect 203822 600818 204004 601054
rect 203404 600734 204004 600818
rect 203404 600498 203586 600734
rect 203822 600498 204004 600734
rect 203404 565054 204004 600498
rect 203404 564818 203586 565054
rect 203822 564818 204004 565054
rect 203404 564734 204004 564818
rect 203404 564498 203586 564734
rect 203822 564498 204004 564734
rect 203404 529054 204004 564498
rect 203404 528818 203586 529054
rect 203822 528818 204004 529054
rect 203404 528734 204004 528818
rect 203404 528498 203586 528734
rect 203822 528498 204004 528734
rect 203404 493054 204004 528498
rect 203404 492818 203586 493054
rect 203822 492818 204004 493054
rect 203404 492734 204004 492818
rect 203404 492498 203586 492734
rect 203822 492498 204004 492734
rect 203404 457054 204004 492498
rect 203404 456818 203586 457054
rect 203822 456818 204004 457054
rect 203404 456734 204004 456818
rect 203404 456498 203586 456734
rect 203822 456498 204004 456734
rect 203404 421054 204004 456498
rect 203404 420818 203586 421054
rect 203822 420818 204004 421054
rect 203404 420734 204004 420818
rect 203404 420498 203586 420734
rect 203822 420498 204004 420734
rect 203404 385054 204004 420498
rect 203404 384818 203586 385054
rect 203822 384818 204004 385054
rect 203404 384734 204004 384818
rect 203404 384498 203586 384734
rect 203822 384498 204004 384734
rect 203404 349054 204004 384498
rect 203404 348818 203586 349054
rect 203822 348818 204004 349054
rect 203404 348734 204004 348818
rect 203404 348498 203586 348734
rect 203822 348498 204004 348734
rect 203404 313054 204004 348498
rect 203404 312818 203586 313054
rect 203822 312818 204004 313054
rect 203404 312734 204004 312818
rect 203404 312498 203586 312734
rect 203822 312498 204004 312734
rect 203404 277054 204004 312498
rect 203404 276818 203586 277054
rect 203822 276818 204004 277054
rect 203404 276734 204004 276818
rect 203404 276498 203586 276734
rect 203822 276498 204004 276734
rect 203404 241054 204004 276498
rect 203404 240818 203586 241054
rect 203822 240818 204004 241054
rect 203404 240734 204004 240818
rect 203404 240498 203586 240734
rect 203822 240498 204004 240734
rect 203404 205054 204004 240498
rect 203404 204818 203586 205054
rect 203822 204818 204004 205054
rect 203404 204734 204004 204818
rect 203404 204498 203586 204734
rect 203822 204498 204004 204734
rect 203404 169054 204004 204498
rect 203404 168818 203586 169054
rect 203822 168818 204004 169054
rect 203404 168734 204004 168818
rect 203404 168498 203586 168734
rect 203822 168498 204004 168734
rect 203404 133054 204004 168498
rect 203404 132818 203586 133054
rect 203822 132818 204004 133054
rect 203404 132734 204004 132818
rect 203404 132498 203586 132734
rect 203822 132498 204004 132734
rect 203404 97054 204004 132498
rect 203404 96818 203586 97054
rect 203822 96818 204004 97054
rect 203404 96734 204004 96818
rect 203404 96498 203586 96734
rect 203822 96498 204004 96734
rect 203404 61054 204004 96498
rect 203404 60818 203586 61054
rect 203822 60818 204004 61054
rect 203404 60734 204004 60818
rect 203404 60498 203586 60734
rect 203822 60498 204004 60734
rect 203404 25054 204004 60498
rect 203404 24818 203586 25054
rect 203822 24818 204004 25054
rect 203404 24734 204004 24818
rect 203404 24498 203586 24734
rect 203822 24498 204004 24734
rect 203404 -3166 204004 24498
rect 203404 -3402 203586 -3166
rect 203822 -3402 204004 -3166
rect 203404 -3486 204004 -3402
rect 203404 -3722 203586 -3486
rect 203822 -3722 204004 -3486
rect 203404 -3744 204004 -3722
rect 207004 676654 207604 708982
rect 207004 676418 207186 676654
rect 207422 676418 207604 676654
rect 207004 676334 207604 676418
rect 207004 676098 207186 676334
rect 207422 676098 207604 676334
rect 207004 640654 207604 676098
rect 207004 640418 207186 640654
rect 207422 640418 207604 640654
rect 207004 640334 207604 640418
rect 207004 640098 207186 640334
rect 207422 640098 207604 640334
rect 207004 604654 207604 640098
rect 207004 604418 207186 604654
rect 207422 604418 207604 604654
rect 207004 604334 207604 604418
rect 207004 604098 207186 604334
rect 207422 604098 207604 604334
rect 207004 568654 207604 604098
rect 207004 568418 207186 568654
rect 207422 568418 207604 568654
rect 207004 568334 207604 568418
rect 207004 568098 207186 568334
rect 207422 568098 207604 568334
rect 207004 532654 207604 568098
rect 207004 532418 207186 532654
rect 207422 532418 207604 532654
rect 207004 532334 207604 532418
rect 207004 532098 207186 532334
rect 207422 532098 207604 532334
rect 207004 496654 207604 532098
rect 207004 496418 207186 496654
rect 207422 496418 207604 496654
rect 207004 496334 207604 496418
rect 207004 496098 207186 496334
rect 207422 496098 207604 496334
rect 207004 460654 207604 496098
rect 207004 460418 207186 460654
rect 207422 460418 207604 460654
rect 207004 460334 207604 460418
rect 207004 460098 207186 460334
rect 207422 460098 207604 460334
rect 207004 424654 207604 460098
rect 207004 424418 207186 424654
rect 207422 424418 207604 424654
rect 207004 424334 207604 424418
rect 207004 424098 207186 424334
rect 207422 424098 207604 424334
rect 207004 388654 207604 424098
rect 207004 388418 207186 388654
rect 207422 388418 207604 388654
rect 207004 388334 207604 388418
rect 207004 388098 207186 388334
rect 207422 388098 207604 388334
rect 207004 352654 207604 388098
rect 207004 352418 207186 352654
rect 207422 352418 207604 352654
rect 207004 352334 207604 352418
rect 207004 352098 207186 352334
rect 207422 352098 207604 352334
rect 207004 316654 207604 352098
rect 207004 316418 207186 316654
rect 207422 316418 207604 316654
rect 207004 316334 207604 316418
rect 207004 316098 207186 316334
rect 207422 316098 207604 316334
rect 207004 280654 207604 316098
rect 207004 280418 207186 280654
rect 207422 280418 207604 280654
rect 207004 280334 207604 280418
rect 207004 280098 207186 280334
rect 207422 280098 207604 280334
rect 207004 244654 207604 280098
rect 207004 244418 207186 244654
rect 207422 244418 207604 244654
rect 207004 244334 207604 244418
rect 207004 244098 207186 244334
rect 207422 244098 207604 244334
rect 207004 208654 207604 244098
rect 207004 208418 207186 208654
rect 207422 208418 207604 208654
rect 207004 208334 207604 208418
rect 207004 208098 207186 208334
rect 207422 208098 207604 208334
rect 207004 172654 207604 208098
rect 207004 172418 207186 172654
rect 207422 172418 207604 172654
rect 207004 172334 207604 172418
rect 207004 172098 207186 172334
rect 207422 172098 207604 172334
rect 207004 136654 207604 172098
rect 207004 136418 207186 136654
rect 207422 136418 207604 136654
rect 207004 136334 207604 136418
rect 207004 136098 207186 136334
rect 207422 136098 207604 136334
rect 207004 100654 207604 136098
rect 207004 100418 207186 100654
rect 207422 100418 207604 100654
rect 207004 100334 207604 100418
rect 207004 100098 207186 100334
rect 207422 100098 207604 100334
rect 207004 64654 207604 100098
rect 207004 64418 207186 64654
rect 207422 64418 207604 64654
rect 207004 64334 207604 64418
rect 207004 64098 207186 64334
rect 207422 64098 207604 64334
rect 207004 28654 207604 64098
rect 207004 28418 207186 28654
rect 207422 28418 207604 28654
rect 207004 28334 207604 28418
rect 207004 28098 207186 28334
rect 207422 28098 207604 28334
rect 207004 -5046 207604 28098
rect 207004 -5282 207186 -5046
rect 207422 -5282 207604 -5046
rect 207004 -5366 207604 -5282
rect 207004 -5602 207186 -5366
rect 207422 -5602 207604 -5366
rect 207004 -5624 207604 -5602
rect 210604 680254 211204 710862
rect 228604 710478 229204 711440
rect 228604 710242 228786 710478
rect 229022 710242 229204 710478
rect 228604 710158 229204 710242
rect 228604 709922 228786 710158
rect 229022 709922 229204 710158
rect 225004 708598 225604 709560
rect 225004 708362 225186 708598
rect 225422 708362 225604 708598
rect 225004 708278 225604 708362
rect 225004 708042 225186 708278
rect 225422 708042 225604 708278
rect 221404 706718 222004 707680
rect 221404 706482 221586 706718
rect 221822 706482 222004 706718
rect 221404 706398 222004 706482
rect 221404 706162 221586 706398
rect 221822 706162 222004 706398
rect 210604 680018 210786 680254
rect 211022 680018 211204 680254
rect 210604 679934 211204 680018
rect 210604 679698 210786 679934
rect 211022 679698 211204 679934
rect 210604 644254 211204 679698
rect 210604 644018 210786 644254
rect 211022 644018 211204 644254
rect 210604 643934 211204 644018
rect 210604 643698 210786 643934
rect 211022 643698 211204 643934
rect 210604 608254 211204 643698
rect 210604 608018 210786 608254
rect 211022 608018 211204 608254
rect 210604 607934 211204 608018
rect 210604 607698 210786 607934
rect 211022 607698 211204 607934
rect 210604 572254 211204 607698
rect 210604 572018 210786 572254
rect 211022 572018 211204 572254
rect 210604 571934 211204 572018
rect 210604 571698 210786 571934
rect 211022 571698 211204 571934
rect 210604 536254 211204 571698
rect 210604 536018 210786 536254
rect 211022 536018 211204 536254
rect 210604 535934 211204 536018
rect 210604 535698 210786 535934
rect 211022 535698 211204 535934
rect 210604 500254 211204 535698
rect 210604 500018 210786 500254
rect 211022 500018 211204 500254
rect 210604 499934 211204 500018
rect 210604 499698 210786 499934
rect 211022 499698 211204 499934
rect 210604 464254 211204 499698
rect 210604 464018 210786 464254
rect 211022 464018 211204 464254
rect 210604 463934 211204 464018
rect 210604 463698 210786 463934
rect 211022 463698 211204 463934
rect 210604 428254 211204 463698
rect 210604 428018 210786 428254
rect 211022 428018 211204 428254
rect 210604 427934 211204 428018
rect 210604 427698 210786 427934
rect 211022 427698 211204 427934
rect 210604 392254 211204 427698
rect 210604 392018 210786 392254
rect 211022 392018 211204 392254
rect 210604 391934 211204 392018
rect 210604 391698 210786 391934
rect 211022 391698 211204 391934
rect 210604 356254 211204 391698
rect 210604 356018 210786 356254
rect 211022 356018 211204 356254
rect 210604 355934 211204 356018
rect 210604 355698 210786 355934
rect 211022 355698 211204 355934
rect 210604 320254 211204 355698
rect 210604 320018 210786 320254
rect 211022 320018 211204 320254
rect 210604 319934 211204 320018
rect 210604 319698 210786 319934
rect 211022 319698 211204 319934
rect 210604 284254 211204 319698
rect 210604 284018 210786 284254
rect 211022 284018 211204 284254
rect 210604 283934 211204 284018
rect 210604 283698 210786 283934
rect 211022 283698 211204 283934
rect 210604 248254 211204 283698
rect 210604 248018 210786 248254
rect 211022 248018 211204 248254
rect 210604 247934 211204 248018
rect 210604 247698 210786 247934
rect 211022 247698 211204 247934
rect 210604 212254 211204 247698
rect 210604 212018 210786 212254
rect 211022 212018 211204 212254
rect 210604 211934 211204 212018
rect 210604 211698 210786 211934
rect 211022 211698 211204 211934
rect 210604 176254 211204 211698
rect 210604 176018 210786 176254
rect 211022 176018 211204 176254
rect 210604 175934 211204 176018
rect 210604 175698 210786 175934
rect 211022 175698 211204 175934
rect 210604 140254 211204 175698
rect 210604 140018 210786 140254
rect 211022 140018 211204 140254
rect 210604 139934 211204 140018
rect 210604 139698 210786 139934
rect 211022 139698 211204 139934
rect 210604 104254 211204 139698
rect 210604 104018 210786 104254
rect 211022 104018 211204 104254
rect 210604 103934 211204 104018
rect 210604 103698 210786 103934
rect 211022 103698 211204 103934
rect 210604 68254 211204 103698
rect 210604 68018 210786 68254
rect 211022 68018 211204 68254
rect 210604 67934 211204 68018
rect 210604 67698 210786 67934
rect 211022 67698 211204 67934
rect 210604 32254 211204 67698
rect 210604 32018 210786 32254
rect 211022 32018 211204 32254
rect 210604 31934 211204 32018
rect 210604 31698 210786 31934
rect 211022 31698 211204 31934
rect 192604 -6222 192786 -5986
rect 193022 -6222 193204 -5986
rect 192604 -6306 193204 -6222
rect 192604 -6542 192786 -6306
rect 193022 -6542 193204 -6306
rect 192604 -7504 193204 -6542
rect 210604 -6926 211204 31698
rect 217804 704838 218404 705800
rect 217804 704602 217986 704838
rect 218222 704602 218404 704838
rect 217804 704518 218404 704602
rect 217804 704282 217986 704518
rect 218222 704282 218404 704518
rect 217804 687454 218404 704282
rect 217804 687218 217986 687454
rect 218222 687218 218404 687454
rect 217804 687134 218404 687218
rect 217804 686898 217986 687134
rect 218222 686898 218404 687134
rect 217804 651454 218404 686898
rect 217804 651218 217986 651454
rect 218222 651218 218404 651454
rect 217804 651134 218404 651218
rect 217804 650898 217986 651134
rect 218222 650898 218404 651134
rect 217804 615454 218404 650898
rect 217804 615218 217986 615454
rect 218222 615218 218404 615454
rect 217804 615134 218404 615218
rect 217804 614898 217986 615134
rect 218222 614898 218404 615134
rect 217804 579454 218404 614898
rect 217804 579218 217986 579454
rect 218222 579218 218404 579454
rect 217804 579134 218404 579218
rect 217804 578898 217986 579134
rect 218222 578898 218404 579134
rect 217804 543454 218404 578898
rect 217804 543218 217986 543454
rect 218222 543218 218404 543454
rect 217804 543134 218404 543218
rect 217804 542898 217986 543134
rect 218222 542898 218404 543134
rect 217804 507454 218404 542898
rect 217804 507218 217986 507454
rect 218222 507218 218404 507454
rect 217804 507134 218404 507218
rect 217804 506898 217986 507134
rect 218222 506898 218404 507134
rect 217804 471454 218404 506898
rect 217804 471218 217986 471454
rect 218222 471218 218404 471454
rect 217804 471134 218404 471218
rect 217804 470898 217986 471134
rect 218222 470898 218404 471134
rect 217804 435454 218404 470898
rect 217804 435218 217986 435454
rect 218222 435218 218404 435454
rect 217804 435134 218404 435218
rect 217804 434898 217986 435134
rect 218222 434898 218404 435134
rect 217804 399454 218404 434898
rect 217804 399218 217986 399454
rect 218222 399218 218404 399454
rect 217804 399134 218404 399218
rect 217804 398898 217986 399134
rect 218222 398898 218404 399134
rect 217804 363454 218404 398898
rect 217804 363218 217986 363454
rect 218222 363218 218404 363454
rect 217804 363134 218404 363218
rect 217804 362898 217986 363134
rect 218222 362898 218404 363134
rect 217804 327454 218404 362898
rect 217804 327218 217986 327454
rect 218222 327218 218404 327454
rect 217804 327134 218404 327218
rect 217804 326898 217986 327134
rect 218222 326898 218404 327134
rect 217804 291454 218404 326898
rect 217804 291218 217986 291454
rect 218222 291218 218404 291454
rect 217804 291134 218404 291218
rect 217804 290898 217986 291134
rect 218222 290898 218404 291134
rect 217804 255454 218404 290898
rect 217804 255218 217986 255454
rect 218222 255218 218404 255454
rect 217804 255134 218404 255218
rect 217804 254898 217986 255134
rect 218222 254898 218404 255134
rect 217804 219454 218404 254898
rect 217804 219218 217986 219454
rect 218222 219218 218404 219454
rect 217804 219134 218404 219218
rect 217804 218898 217986 219134
rect 218222 218898 218404 219134
rect 217804 183454 218404 218898
rect 217804 183218 217986 183454
rect 218222 183218 218404 183454
rect 217804 183134 218404 183218
rect 217804 182898 217986 183134
rect 218222 182898 218404 183134
rect 217804 147454 218404 182898
rect 217804 147218 217986 147454
rect 218222 147218 218404 147454
rect 217804 147134 218404 147218
rect 217804 146898 217986 147134
rect 218222 146898 218404 147134
rect 217804 111454 218404 146898
rect 217804 111218 217986 111454
rect 218222 111218 218404 111454
rect 217804 111134 218404 111218
rect 217804 110898 217986 111134
rect 218222 110898 218404 111134
rect 217804 75454 218404 110898
rect 217804 75218 217986 75454
rect 218222 75218 218404 75454
rect 217804 75134 218404 75218
rect 217804 74898 217986 75134
rect 218222 74898 218404 75134
rect 217804 39454 218404 74898
rect 217804 39218 217986 39454
rect 218222 39218 218404 39454
rect 217804 39134 218404 39218
rect 217804 38898 217986 39134
rect 218222 38898 218404 39134
rect 217804 3454 218404 38898
rect 217804 3218 217986 3454
rect 218222 3218 218404 3454
rect 217804 3134 218404 3218
rect 217804 2898 217986 3134
rect 218222 2898 218404 3134
rect 217804 -346 218404 2898
rect 217804 -582 217986 -346
rect 218222 -582 218404 -346
rect 217804 -666 218404 -582
rect 217804 -902 217986 -666
rect 218222 -902 218404 -666
rect 217804 -1864 218404 -902
rect 221404 691054 222004 706162
rect 221404 690818 221586 691054
rect 221822 690818 222004 691054
rect 221404 690734 222004 690818
rect 221404 690498 221586 690734
rect 221822 690498 222004 690734
rect 221404 655054 222004 690498
rect 221404 654818 221586 655054
rect 221822 654818 222004 655054
rect 221404 654734 222004 654818
rect 221404 654498 221586 654734
rect 221822 654498 222004 654734
rect 221404 619054 222004 654498
rect 221404 618818 221586 619054
rect 221822 618818 222004 619054
rect 221404 618734 222004 618818
rect 221404 618498 221586 618734
rect 221822 618498 222004 618734
rect 221404 583054 222004 618498
rect 221404 582818 221586 583054
rect 221822 582818 222004 583054
rect 221404 582734 222004 582818
rect 221404 582498 221586 582734
rect 221822 582498 222004 582734
rect 221404 547054 222004 582498
rect 221404 546818 221586 547054
rect 221822 546818 222004 547054
rect 221404 546734 222004 546818
rect 221404 546498 221586 546734
rect 221822 546498 222004 546734
rect 221404 511054 222004 546498
rect 221404 510818 221586 511054
rect 221822 510818 222004 511054
rect 221404 510734 222004 510818
rect 221404 510498 221586 510734
rect 221822 510498 222004 510734
rect 221404 475054 222004 510498
rect 221404 474818 221586 475054
rect 221822 474818 222004 475054
rect 221404 474734 222004 474818
rect 221404 474498 221586 474734
rect 221822 474498 222004 474734
rect 221404 439054 222004 474498
rect 221404 438818 221586 439054
rect 221822 438818 222004 439054
rect 221404 438734 222004 438818
rect 221404 438498 221586 438734
rect 221822 438498 222004 438734
rect 221404 403054 222004 438498
rect 221404 402818 221586 403054
rect 221822 402818 222004 403054
rect 221404 402734 222004 402818
rect 221404 402498 221586 402734
rect 221822 402498 222004 402734
rect 221404 367054 222004 402498
rect 221404 366818 221586 367054
rect 221822 366818 222004 367054
rect 221404 366734 222004 366818
rect 221404 366498 221586 366734
rect 221822 366498 222004 366734
rect 221404 331054 222004 366498
rect 221404 330818 221586 331054
rect 221822 330818 222004 331054
rect 221404 330734 222004 330818
rect 221404 330498 221586 330734
rect 221822 330498 222004 330734
rect 221404 295054 222004 330498
rect 221404 294818 221586 295054
rect 221822 294818 222004 295054
rect 221404 294734 222004 294818
rect 221404 294498 221586 294734
rect 221822 294498 222004 294734
rect 221404 259054 222004 294498
rect 221404 258818 221586 259054
rect 221822 258818 222004 259054
rect 221404 258734 222004 258818
rect 221404 258498 221586 258734
rect 221822 258498 222004 258734
rect 221404 223054 222004 258498
rect 221404 222818 221586 223054
rect 221822 222818 222004 223054
rect 221404 222734 222004 222818
rect 221404 222498 221586 222734
rect 221822 222498 222004 222734
rect 221404 187054 222004 222498
rect 221404 186818 221586 187054
rect 221822 186818 222004 187054
rect 221404 186734 222004 186818
rect 221404 186498 221586 186734
rect 221822 186498 222004 186734
rect 221404 151054 222004 186498
rect 221404 150818 221586 151054
rect 221822 150818 222004 151054
rect 221404 150734 222004 150818
rect 221404 150498 221586 150734
rect 221822 150498 222004 150734
rect 221404 115054 222004 150498
rect 221404 114818 221586 115054
rect 221822 114818 222004 115054
rect 221404 114734 222004 114818
rect 221404 114498 221586 114734
rect 221822 114498 222004 114734
rect 221404 79054 222004 114498
rect 221404 78818 221586 79054
rect 221822 78818 222004 79054
rect 221404 78734 222004 78818
rect 221404 78498 221586 78734
rect 221822 78498 222004 78734
rect 221404 43054 222004 78498
rect 221404 42818 221586 43054
rect 221822 42818 222004 43054
rect 221404 42734 222004 42818
rect 221404 42498 221586 42734
rect 221822 42498 222004 42734
rect 221404 7054 222004 42498
rect 221404 6818 221586 7054
rect 221822 6818 222004 7054
rect 221404 6734 222004 6818
rect 221404 6498 221586 6734
rect 221822 6498 222004 6734
rect 221404 -2226 222004 6498
rect 221404 -2462 221586 -2226
rect 221822 -2462 222004 -2226
rect 221404 -2546 222004 -2462
rect 221404 -2782 221586 -2546
rect 221822 -2782 222004 -2546
rect 221404 -3744 222004 -2782
rect 225004 694654 225604 708042
rect 225004 694418 225186 694654
rect 225422 694418 225604 694654
rect 225004 694334 225604 694418
rect 225004 694098 225186 694334
rect 225422 694098 225604 694334
rect 225004 658654 225604 694098
rect 225004 658418 225186 658654
rect 225422 658418 225604 658654
rect 225004 658334 225604 658418
rect 225004 658098 225186 658334
rect 225422 658098 225604 658334
rect 225004 622654 225604 658098
rect 225004 622418 225186 622654
rect 225422 622418 225604 622654
rect 225004 622334 225604 622418
rect 225004 622098 225186 622334
rect 225422 622098 225604 622334
rect 225004 586654 225604 622098
rect 225004 586418 225186 586654
rect 225422 586418 225604 586654
rect 225004 586334 225604 586418
rect 225004 586098 225186 586334
rect 225422 586098 225604 586334
rect 225004 550654 225604 586098
rect 225004 550418 225186 550654
rect 225422 550418 225604 550654
rect 225004 550334 225604 550418
rect 225004 550098 225186 550334
rect 225422 550098 225604 550334
rect 225004 514654 225604 550098
rect 225004 514418 225186 514654
rect 225422 514418 225604 514654
rect 225004 514334 225604 514418
rect 225004 514098 225186 514334
rect 225422 514098 225604 514334
rect 225004 478654 225604 514098
rect 225004 478418 225186 478654
rect 225422 478418 225604 478654
rect 225004 478334 225604 478418
rect 225004 478098 225186 478334
rect 225422 478098 225604 478334
rect 225004 442654 225604 478098
rect 225004 442418 225186 442654
rect 225422 442418 225604 442654
rect 225004 442334 225604 442418
rect 225004 442098 225186 442334
rect 225422 442098 225604 442334
rect 225004 406654 225604 442098
rect 225004 406418 225186 406654
rect 225422 406418 225604 406654
rect 225004 406334 225604 406418
rect 225004 406098 225186 406334
rect 225422 406098 225604 406334
rect 225004 370654 225604 406098
rect 225004 370418 225186 370654
rect 225422 370418 225604 370654
rect 225004 370334 225604 370418
rect 225004 370098 225186 370334
rect 225422 370098 225604 370334
rect 225004 334654 225604 370098
rect 225004 334418 225186 334654
rect 225422 334418 225604 334654
rect 225004 334334 225604 334418
rect 225004 334098 225186 334334
rect 225422 334098 225604 334334
rect 225004 298654 225604 334098
rect 225004 298418 225186 298654
rect 225422 298418 225604 298654
rect 225004 298334 225604 298418
rect 225004 298098 225186 298334
rect 225422 298098 225604 298334
rect 225004 262654 225604 298098
rect 225004 262418 225186 262654
rect 225422 262418 225604 262654
rect 225004 262334 225604 262418
rect 225004 262098 225186 262334
rect 225422 262098 225604 262334
rect 225004 226654 225604 262098
rect 225004 226418 225186 226654
rect 225422 226418 225604 226654
rect 225004 226334 225604 226418
rect 225004 226098 225186 226334
rect 225422 226098 225604 226334
rect 225004 190654 225604 226098
rect 225004 190418 225186 190654
rect 225422 190418 225604 190654
rect 225004 190334 225604 190418
rect 225004 190098 225186 190334
rect 225422 190098 225604 190334
rect 225004 154654 225604 190098
rect 225004 154418 225186 154654
rect 225422 154418 225604 154654
rect 225004 154334 225604 154418
rect 225004 154098 225186 154334
rect 225422 154098 225604 154334
rect 225004 118654 225604 154098
rect 225004 118418 225186 118654
rect 225422 118418 225604 118654
rect 225004 118334 225604 118418
rect 225004 118098 225186 118334
rect 225422 118098 225604 118334
rect 225004 82654 225604 118098
rect 225004 82418 225186 82654
rect 225422 82418 225604 82654
rect 225004 82334 225604 82418
rect 225004 82098 225186 82334
rect 225422 82098 225604 82334
rect 225004 46654 225604 82098
rect 225004 46418 225186 46654
rect 225422 46418 225604 46654
rect 225004 46334 225604 46418
rect 225004 46098 225186 46334
rect 225422 46098 225604 46334
rect 225004 10654 225604 46098
rect 225004 10418 225186 10654
rect 225422 10418 225604 10654
rect 225004 10334 225604 10418
rect 225004 10098 225186 10334
rect 225422 10098 225604 10334
rect 225004 -4106 225604 10098
rect 225004 -4342 225186 -4106
rect 225422 -4342 225604 -4106
rect 225004 -4426 225604 -4342
rect 225004 -4662 225186 -4426
rect 225422 -4662 225604 -4426
rect 225004 -5624 225604 -4662
rect 228604 698254 229204 709922
rect 246604 711418 247204 711440
rect 246604 711182 246786 711418
rect 247022 711182 247204 711418
rect 246604 711098 247204 711182
rect 246604 710862 246786 711098
rect 247022 710862 247204 711098
rect 243004 709538 243604 709560
rect 243004 709302 243186 709538
rect 243422 709302 243604 709538
rect 243004 709218 243604 709302
rect 243004 708982 243186 709218
rect 243422 708982 243604 709218
rect 239404 707658 240004 707680
rect 239404 707422 239586 707658
rect 239822 707422 240004 707658
rect 239404 707338 240004 707422
rect 239404 707102 239586 707338
rect 239822 707102 240004 707338
rect 228604 698018 228786 698254
rect 229022 698018 229204 698254
rect 228604 697934 229204 698018
rect 228604 697698 228786 697934
rect 229022 697698 229204 697934
rect 228604 662254 229204 697698
rect 228604 662018 228786 662254
rect 229022 662018 229204 662254
rect 228604 661934 229204 662018
rect 228604 661698 228786 661934
rect 229022 661698 229204 661934
rect 228604 626254 229204 661698
rect 228604 626018 228786 626254
rect 229022 626018 229204 626254
rect 228604 625934 229204 626018
rect 228604 625698 228786 625934
rect 229022 625698 229204 625934
rect 228604 590254 229204 625698
rect 228604 590018 228786 590254
rect 229022 590018 229204 590254
rect 228604 589934 229204 590018
rect 228604 589698 228786 589934
rect 229022 589698 229204 589934
rect 228604 554254 229204 589698
rect 228604 554018 228786 554254
rect 229022 554018 229204 554254
rect 228604 553934 229204 554018
rect 228604 553698 228786 553934
rect 229022 553698 229204 553934
rect 228604 518254 229204 553698
rect 228604 518018 228786 518254
rect 229022 518018 229204 518254
rect 228604 517934 229204 518018
rect 228604 517698 228786 517934
rect 229022 517698 229204 517934
rect 228604 482254 229204 517698
rect 228604 482018 228786 482254
rect 229022 482018 229204 482254
rect 228604 481934 229204 482018
rect 228604 481698 228786 481934
rect 229022 481698 229204 481934
rect 228604 446254 229204 481698
rect 228604 446018 228786 446254
rect 229022 446018 229204 446254
rect 228604 445934 229204 446018
rect 228604 445698 228786 445934
rect 229022 445698 229204 445934
rect 228604 410254 229204 445698
rect 228604 410018 228786 410254
rect 229022 410018 229204 410254
rect 228604 409934 229204 410018
rect 235804 705778 236404 705800
rect 235804 705542 235986 705778
rect 236222 705542 236404 705778
rect 235804 705458 236404 705542
rect 235804 705222 235986 705458
rect 236222 705222 236404 705458
rect 235804 669454 236404 705222
rect 235804 669218 235986 669454
rect 236222 669218 236404 669454
rect 235804 669134 236404 669218
rect 235804 668898 235986 669134
rect 236222 668898 236404 669134
rect 235804 633454 236404 668898
rect 235804 633218 235986 633454
rect 236222 633218 236404 633454
rect 235804 633134 236404 633218
rect 235804 632898 235986 633134
rect 236222 632898 236404 633134
rect 235804 597454 236404 632898
rect 235804 597218 235986 597454
rect 236222 597218 236404 597454
rect 235804 597134 236404 597218
rect 235804 596898 235986 597134
rect 236222 596898 236404 597134
rect 235804 561454 236404 596898
rect 235804 561218 235986 561454
rect 236222 561218 236404 561454
rect 235804 561134 236404 561218
rect 235804 560898 235986 561134
rect 236222 560898 236404 561134
rect 235804 525454 236404 560898
rect 235804 525218 235986 525454
rect 236222 525218 236404 525454
rect 235804 525134 236404 525218
rect 235804 524898 235986 525134
rect 236222 524898 236404 525134
rect 235804 489454 236404 524898
rect 235804 489218 235986 489454
rect 236222 489218 236404 489454
rect 235804 489134 236404 489218
rect 235804 488898 235986 489134
rect 236222 488898 236404 489134
rect 235804 453454 236404 488898
rect 235804 453218 235986 453454
rect 236222 453218 236404 453454
rect 235804 453134 236404 453218
rect 235804 452898 235986 453134
rect 236222 452898 236404 453134
rect 235804 417454 236404 452898
rect 235804 417218 235986 417454
rect 236222 417218 236404 417454
rect 235804 417134 236404 417218
rect 235804 416898 235986 417134
rect 236222 416898 236404 417134
rect 235804 410000 236404 416898
rect 239404 673054 240004 707102
rect 239404 672818 239586 673054
rect 239822 672818 240004 673054
rect 239404 672734 240004 672818
rect 239404 672498 239586 672734
rect 239822 672498 240004 672734
rect 239404 637054 240004 672498
rect 239404 636818 239586 637054
rect 239822 636818 240004 637054
rect 239404 636734 240004 636818
rect 239404 636498 239586 636734
rect 239822 636498 240004 636734
rect 239404 601054 240004 636498
rect 239404 600818 239586 601054
rect 239822 600818 240004 601054
rect 239404 600734 240004 600818
rect 239404 600498 239586 600734
rect 239822 600498 240004 600734
rect 239404 565054 240004 600498
rect 239404 564818 239586 565054
rect 239822 564818 240004 565054
rect 239404 564734 240004 564818
rect 239404 564498 239586 564734
rect 239822 564498 240004 564734
rect 239404 529054 240004 564498
rect 239404 528818 239586 529054
rect 239822 528818 240004 529054
rect 239404 528734 240004 528818
rect 239404 528498 239586 528734
rect 239822 528498 240004 528734
rect 239404 493054 240004 528498
rect 239404 492818 239586 493054
rect 239822 492818 240004 493054
rect 239404 492734 240004 492818
rect 239404 492498 239586 492734
rect 239822 492498 240004 492734
rect 239404 457054 240004 492498
rect 239404 456818 239586 457054
rect 239822 456818 240004 457054
rect 239404 456734 240004 456818
rect 239404 456498 239586 456734
rect 239822 456498 240004 456734
rect 239404 421054 240004 456498
rect 239404 420818 239586 421054
rect 239822 420818 240004 421054
rect 239404 420734 240004 420818
rect 239404 420498 239586 420734
rect 239822 420498 240004 420734
rect 239404 410000 240004 420498
rect 243004 676654 243604 708982
rect 243004 676418 243186 676654
rect 243422 676418 243604 676654
rect 243004 676334 243604 676418
rect 243004 676098 243186 676334
rect 243422 676098 243604 676334
rect 243004 640654 243604 676098
rect 243004 640418 243186 640654
rect 243422 640418 243604 640654
rect 243004 640334 243604 640418
rect 243004 640098 243186 640334
rect 243422 640098 243604 640334
rect 243004 604654 243604 640098
rect 243004 604418 243186 604654
rect 243422 604418 243604 604654
rect 243004 604334 243604 604418
rect 243004 604098 243186 604334
rect 243422 604098 243604 604334
rect 243004 568654 243604 604098
rect 243004 568418 243186 568654
rect 243422 568418 243604 568654
rect 243004 568334 243604 568418
rect 243004 568098 243186 568334
rect 243422 568098 243604 568334
rect 243004 532654 243604 568098
rect 243004 532418 243186 532654
rect 243422 532418 243604 532654
rect 243004 532334 243604 532418
rect 243004 532098 243186 532334
rect 243422 532098 243604 532334
rect 243004 496654 243604 532098
rect 243004 496418 243186 496654
rect 243422 496418 243604 496654
rect 243004 496334 243604 496418
rect 243004 496098 243186 496334
rect 243422 496098 243604 496334
rect 243004 460654 243604 496098
rect 243004 460418 243186 460654
rect 243422 460418 243604 460654
rect 243004 460334 243604 460418
rect 243004 460098 243186 460334
rect 243422 460098 243604 460334
rect 243004 424654 243604 460098
rect 243004 424418 243186 424654
rect 243422 424418 243604 424654
rect 243004 424334 243604 424418
rect 243004 424098 243186 424334
rect 243422 424098 243604 424334
rect 243004 410000 243604 424098
rect 246604 680254 247204 710862
rect 264604 710478 265204 711440
rect 264604 710242 264786 710478
rect 265022 710242 265204 710478
rect 264604 710158 265204 710242
rect 264604 709922 264786 710158
rect 265022 709922 265204 710158
rect 261004 708598 261604 709560
rect 261004 708362 261186 708598
rect 261422 708362 261604 708598
rect 261004 708278 261604 708362
rect 261004 708042 261186 708278
rect 261422 708042 261604 708278
rect 257404 706718 258004 707680
rect 257404 706482 257586 706718
rect 257822 706482 258004 706718
rect 257404 706398 258004 706482
rect 257404 706162 257586 706398
rect 257822 706162 258004 706398
rect 246604 680018 246786 680254
rect 247022 680018 247204 680254
rect 246604 679934 247204 680018
rect 246604 679698 246786 679934
rect 247022 679698 247204 679934
rect 246604 644254 247204 679698
rect 246604 644018 246786 644254
rect 247022 644018 247204 644254
rect 246604 643934 247204 644018
rect 246604 643698 246786 643934
rect 247022 643698 247204 643934
rect 246604 608254 247204 643698
rect 246604 608018 246786 608254
rect 247022 608018 247204 608254
rect 246604 607934 247204 608018
rect 246604 607698 246786 607934
rect 247022 607698 247204 607934
rect 246604 572254 247204 607698
rect 246604 572018 246786 572254
rect 247022 572018 247204 572254
rect 246604 571934 247204 572018
rect 246604 571698 246786 571934
rect 247022 571698 247204 571934
rect 246604 536254 247204 571698
rect 246604 536018 246786 536254
rect 247022 536018 247204 536254
rect 246604 535934 247204 536018
rect 246604 535698 246786 535934
rect 247022 535698 247204 535934
rect 246604 500254 247204 535698
rect 246604 500018 246786 500254
rect 247022 500018 247204 500254
rect 246604 499934 247204 500018
rect 246604 499698 246786 499934
rect 247022 499698 247204 499934
rect 246604 464254 247204 499698
rect 246604 464018 246786 464254
rect 247022 464018 247204 464254
rect 246604 463934 247204 464018
rect 246604 463698 246786 463934
rect 247022 463698 247204 463934
rect 246604 428254 247204 463698
rect 246604 428018 246786 428254
rect 247022 428018 247204 428254
rect 246604 427934 247204 428018
rect 246604 427698 246786 427934
rect 247022 427698 247204 427934
rect 246604 410000 247204 427698
rect 253804 704838 254404 705800
rect 253804 704602 253986 704838
rect 254222 704602 254404 704838
rect 253804 704518 254404 704602
rect 253804 704282 253986 704518
rect 254222 704282 254404 704518
rect 253804 687454 254404 704282
rect 253804 687218 253986 687454
rect 254222 687218 254404 687454
rect 253804 687134 254404 687218
rect 253804 686898 253986 687134
rect 254222 686898 254404 687134
rect 253804 651454 254404 686898
rect 253804 651218 253986 651454
rect 254222 651218 254404 651454
rect 253804 651134 254404 651218
rect 253804 650898 253986 651134
rect 254222 650898 254404 651134
rect 253804 615454 254404 650898
rect 253804 615218 253986 615454
rect 254222 615218 254404 615454
rect 253804 615134 254404 615218
rect 253804 614898 253986 615134
rect 254222 614898 254404 615134
rect 253804 579454 254404 614898
rect 253804 579218 253986 579454
rect 254222 579218 254404 579454
rect 253804 579134 254404 579218
rect 253804 578898 253986 579134
rect 254222 578898 254404 579134
rect 253804 543454 254404 578898
rect 253804 543218 253986 543454
rect 254222 543218 254404 543454
rect 253804 543134 254404 543218
rect 253804 542898 253986 543134
rect 254222 542898 254404 543134
rect 253804 507454 254404 542898
rect 253804 507218 253986 507454
rect 254222 507218 254404 507454
rect 253804 507134 254404 507218
rect 253804 506898 253986 507134
rect 254222 506898 254404 507134
rect 253804 471454 254404 506898
rect 253804 471218 253986 471454
rect 254222 471218 254404 471454
rect 253804 471134 254404 471218
rect 253804 470898 253986 471134
rect 254222 470898 254404 471134
rect 253804 435454 254404 470898
rect 253804 435218 253986 435454
rect 254222 435218 254404 435454
rect 253804 435134 254404 435218
rect 253804 434898 253986 435134
rect 254222 434898 254404 435134
rect 253804 410000 254404 434898
rect 257404 691054 258004 706162
rect 257404 690818 257586 691054
rect 257822 690818 258004 691054
rect 257404 690734 258004 690818
rect 257404 690498 257586 690734
rect 257822 690498 258004 690734
rect 257404 655054 258004 690498
rect 257404 654818 257586 655054
rect 257822 654818 258004 655054
rect 257404 654734 258004 654818
rect 257404 654498 257586 654734
rect 257822 654498 258004 654734
rect 257404 619054 258004 654498
rect 257404 618818 257586 619054
rect 257822 618818 258004 619054
rect 257404 618734 258004 618818
rect 257404 618498 257586 618734
rect 257822 618498 258004 618734
rect 257404 583054 258004 618498
rect 257404 582818 257586 583054
rect 257822 582818 258004 583054
rect 257404 582734 258004 582818
rect 257404 582498 257586 582734
rect 257822 582498 258004 582734
rect 257404 547054 258004 582498
rect 257404 546818 257586 547054
rect 257822 546818 258004 547054
rect 257404 546734 258004 546818
rect 257404 546498 257586 546734
rect 257822 546498 258004 546734
rect 257404 511054 258004 546498
rect 257404 510818 257586 511054
rect 257822 510818 258004 511054
rect 257404 510734 258004 510818
rect 257404 510498 257586 510734
rect 257822 510498 258004 510734
rect 257404 475054 258004 510498
rect 257404 474818 257586 475054
rect 257822 474818 258004 475054
rect 257404 474734 258004 474818
rect 257404 474498 257586 474734
rect 257822 474498 258004 474734
rect 257404 439054 258004 474498
rect 257404 438818 257586 439054
rect 257822 438818 258004 439054
rect 257404 438734 258004 438818
rect 257404 438498 257586 438734
rect 257822 438498 258004 438734
rect 257404 410000 258004 438498
rect 261004 694654 261604 708042
rect 261004 694418 261186 694654
rect 261422 694418 261604 694654
rect 261004 694334 261604 694418
rect 261004 694098 261186 694334
rect 261422 694098 261604 694334
rect 261004 658654 261604 694098
rect 261004 658418 261186 658654
rect 261422 658418 261604 658654
rect 261004 658334 261604 658418
rect 261004 658098 261186 658334
rect 261422 658098 261604 658334
rect 261004 622654 261604 658098
rect 261004 622418 261186 622654
rect 261422 622418 261604 622654
rect 261004 622334 261604 622418
rect 261004 622098 261186 622334
rect 261422 622098 261604 622334
rect 261004 586654 261604 622098
rect 261004 586418 261186 586654
rect 261422 586418 261604 586654
rect 261004 586334 261604 586418
rect 261004 586098 261186 586334
rect 261422 586098 261604 586334
rect 261004 550654 261604 586098
rect 261004 550418 261186 550654
rect 261422 550418 261604 550654
rect 261004 550334 261604 550418
rect 261004 550098 261186 550334
rect 261422 550098 261604 550334
rect 261004 514654 261604 550098
rect 261004 514418 261186 514654
rect 261422 514418 261604 514654
rect 261004 514334 261604 514418
rect 261004 514098 261186 514334
rect 261422 514098 261604 514334
rect 261004 478654 261604 514098
rect 261004 478418 261186 478654
rect 261422 478418 261604 478654
rect 261004 478334 261604 478418
rect 261004 478098 261186 478334
rect 261422 478098 261604 478334
rect 261004 442654 261604 478098
rect 261004 442418 261186 442654
rect 261422 442418 261604 442654
rect 261004 442334 261604 442418
rect 261004 442098 261186 442334
rect 261422 442098 261604 442334
rect 261004 410000 261604 442098
rect 264604 698254 265204 709922
rect 282604 711418 283204 711440
rect 282604 711182 282786 711418
rect 283022 711182 283204 711418
rect 282604 711098 283204 711182
rect 282604 710862 282786 711098
rect 283022 710862 283204 711098
rect 279004 709538 279604 709560
rect 279004 709302 279186 709538
rect 279422 709302 279604 709538
rect 279004 709218 279604 709302
rect 279004 708982 279186 709218
rect 279422 708982 279604 709218
rect 275404 707658 276004 707680
rect 275404 707422 275586 707658
rect 275822 707422 276004 707658
rect 275404 707338 276004 707422
rect 275404 707102 275586 707338
rect 275822 707102 276004 707338
rect 264604 698018 264786 698254
rect 265022 698018 265204 698254
rect 264604 697934 265204 698018
rect 264604 697698 264786 697934
rect 265022 697698 265204 697934
rect 264604 662254 265204 697698
rect 264604 662018 264786 662254
rect 265022 662018 265204 662254
rect 264604 661934 265204 662018
rect 264604 661698 264786 661934
rect 265022 661698 265204 661934
rect 264604 626254 265204 661698
rect 264604 626018 264786 626254
rect 265022 626018 265204 626254
rect 264604 625934 265204 626018
rect 264604 625698 264786 625934
rect 265022 625698 265204 625934
rect 264604 590254 265204 625698
rect 264604 590018 264786 590254
rect 265022 590018 265204 590254
rect 264604 589934 265204 590018
rect 264604 589698 264786 589934
rect 265022 589698 265204 589934
rect 264604 554254 265204 589698
rect 264604 554018 264786 554254
rect 265022 554018 265204 554254
rect 264604 553934 265204 554018
rect 264604 553698 264786 553934
rect 265022 553698 265204 553934
rect 264604 518254 265204 553698
rect 264604 518018 264786 518254
rect 265022 518018 265204 518254
rect 264604 517934 265204 518018
rect 264604 517698 264786 517934
rect 265022 517698 265204 517934
rect 264604 482254 265204 517698
rect 264604 482018 264786 482254
rect 265022 482018 265204 482254
rect 264604 481934 265204 482018
rect 264604 481698 264786 481934
rect 265022 481698 265204 481934
rect 264604 446254 265204 481698
rect 264604 446018 264786 446254
rect 265022 446018 265204 446254
rect 264604 445934 265204 446018
rect 264604 445698 264786 445934
rect 265022 445698 265204 445934
rect 264604 410000 265204 445698
rect 271804 705778 272404 705800
rect 271804 705542 271986 705778
rect 272222 705542 272404 705778
rect 271804 705458 272404 705542
rect 271804 705222 271986 705458
rect 272222 705222 272404 705458
rect 271804 669454 272404 705222
rect 271804 669218 271986 669454
rect 272222 669218 272404 669454
rect 271804 669134 272404 669218
rect 271804 668898 271986 669134
rect 272222 668898 272404 669134
rect 271804 633454 272404 668898
rect 271804 633218 271986 633454
rect 272222 633218 272404 633454
rect 271804 633134 272404 633218
rect 271804 632898 271986 633134
rect 272222 632898 272404 633134
rect 271804 597454 272404 632898
rect 271804 597218 271986 597454
rect 272222 597218 272404 597454
rect 271804 597134 272404 597218
rect 271804 596898 271986 597134
rect 272222 596898 272404 597134
rect 271804 561454 272404 596898
rect 271804 561218 271986 561454
rect 272222 561218 272404 561454
rect 271804 561134 272404 561218
rect 271804 560898 271986 561134
rect 272222 560898 272404 561134
rect 271804 525454 272404 560898
rect 271804 525218 271986 525454
rect 272222 525218 272404 525454
rect 271804 525134 272404 525218
rect 271804 524898 271986 525134
rect 272222 524898 272404 525134
rect 271804 489454 272404 524898
rect 271804 489218 271986 489454
rect 272222 489218 272404 489454
rect 271804 489134 272404 489218
rect 271804 488898 271986 489134
rect 272222 488898 272404 489134
rect 271804 453454 272404 488898
rect 271804 453218 271986 453454
rect 272222 453218 272404 453454
rect 271804 453134 272404 453218
rect 271804 452898 271986 453134
rect 272222 452898 272404 453134
rect 271804 417454 272404 452898
rect 271804 417218 271986 417454
rect 272222 417218 272404 417454
rect 271804 417134 272404 417218
rect 271804 416898 271986 417134
rect 272222 416898 272404 417134
rect 271804 410000 272404 416898
rect 275404 673054 276004 707102
rect 275404 672818 275586 673054
rect 275822 672818 276004 673054
rect 275404 672734 276004 672818
rect 275404 672498 275586 672734
rect 275822 672498 276004 672734
rect 275404 637054 276004 672498
rect 275404 636818 275586 637054
rect 275822 636818 276004 637054
rect 275404 636734 276004 636818
rect 275404 636498 275586 636734
rect 275822 636498 276004 636734
rect 275404 601054 276004 636498
rect 275404 600818 275586 601054
rect 275822 600818 276004 601054
rect 275404 600734 276004 600818
rect 275404 600498 275586 600734
rect 275822 600498 276004 600734
rect 275404 565054 276004 600498
rect 275404 564818 275586 565054
rect 275822 564818 276004 565054
rect 275404 564734 276004 564818
rect 275404 564498 275586 564734
rect 275822 564498 276004 564734
rect 275404 529054 276004 564498
rect 275404 528818 275586 529054
rect 275822 528818 276004 529054
rect 275404 528734 276004 528818
rect 275404 528498 275586 528734
rect 275822 528498 276004 528734
rect 275404 493054 276004 528498
rect 275404 492818 275586 493054
rect 275822 492818 276004 493054
rect 275404 492734 276004 492818
rect 275404 492498 275586 492734
rect 275822 492498 276004 492734
rect 275404 457054 276004 492498
rect 275404 456818 275586 457054
rect 275822 456818 276004 457054
rect 275404 456734 276004 456818
rect 275404 456498 275586 456734
rect 275822 456498 276004 456734
rect 275404 421054 276004 456498
rect 275404 420818 275586 421054
rect 275822 420818 276004 421054
rect 275404 420734 276004 420818
rect 275404 420498 275586 420734
rect 275822 420498 276004 420734
rect 275404 410000 276004 420498
rect 279004 676654 279604 708982
rect 279004 676418 279186 676654
rect 279422 676418 279604 676654
rect 279004 676334 279604 676418
rect 279004 676098 279186 676334
rect 279422 676098 279604 676334
rect 279004 640654 279604 676098
rect 279004 640418 279186 640654
rect 279422 640418 279604 640654
rect 279004 640334 279604 640418
rect 279004 640098 279186 640334
rect 279422 640098 279604 640334
rect 279004 604654 279604 640098
rect 279004 604418 279186 604654
rect 279422 604418 279604 604654
rect 279004 604334 279604 604418
rect 279004 604098 279186 604334
rect 279422 604098 279604 604334
rect 279004 568654 279604 604098
rect 279004 568418 279186 568654
rect 279422 568418 279604 568654
rect 279004 568334 279604 568418
rect 279004 568098 279186 568334
rect 279422 568098 279604 568334
rect 279004 532654 279604 568098
rect 279004 532418 279186 532654
rect 279422 532418 279604 532654
rect 279004 532334 279604 532418
rect 279004 532098 279186 532334
rect 279422 532098 279604 532334
rect 279004 496654 279604 532098
rect 279004 496418 279186 496654
rect 279422 496418 279604 496654
rect 279004 496334 279604 496418
rect 279004 496098 279186 496334
rect 279422 496098 279604 496334
rect 279004 460654 279604 496098
rect 279004 460418 279186 460654
rect 279422 460418 279604 460654
rect 279004 460334 279604 460418
rect 279004 460098 279186 460334
rect 279422 460098 279604 460334
rect 279004 424654 279604 460098
rect 279004 424418 279186 424654
rect 279422 424418 279604 424654
rect 279004 424334 279604 424418
rect 279004 424098 279186 424334
rect 279422 424098 279604 424334
rect 279004 410000 279604 424098
rect 282604 680254 283204 710862
rect 300604 710478 301204 711440
rect 300604 710242 300786 710478
rect 301022 710242 301204 710478
rect 300604 710158 301204 710242
rect 300604 709922 300786 710158
rect 301022 709922 301204 710158
rect 297004 708598 297604 709560
rect 297004 708362 297186 708598
rect 297422 708362 297604 708598
rect 297004 708278 297604 708362
rect 297004 708042 297186 708278
rect 297422 708042 297604 708278
rect 293404 706718 294004 707680
rect 293404 706482 293586 706718
rect 293822 706482 294004 706718
rect 293404 706398 294004 706482
rect 293404 706162 293586 706398
rect 293822 706162 294004 706398
rect 282604 680018 282786 680254
rect 283022 680018 283204 680254
rect 282604 679934 283204 680018
rect 282604 679698 282786 679934
rect 283022 679698 283204 679934
rect 282604 644254 283204 679698
rect 282604 644018 282786 644254
rect 283022 644018 283204 644254
rect 282604 643934 283204 644018
rect 282604 643698 282786 643934
rect 283022 643698 283204 643934
rect 282604 608254 283204 643698
rect 282604 608018 282786 608254
rect 283022 608018 283204 608254
rect 282604 607934 283204 608018
rect 282604 607698 282786 607934
rect 283022 607698 283204 607934
rect 282604 572254 283204 607698
rect 282604 572018 282786 572254
rect 283022 572018 283204 572254
rect 282604 571934 283204 572018
rect 282604 571698 282786 571934
rect 283022 571698 283204 571934
rect 282604 536254 283204 571698
rect 282604 536018 282786 536254
rect 283022 536018 283204 536254
rect 282604 535934 283204 536018
rect 282604 535698 282786 535934
rect 283022 535698 283204 535934
rect 282604 500254 283204 535698
rect 282604 500018 282786 500254
rect 283022 500018 283204 500254
rect 282604 499934 283204 500018
rect 282604 499698 282786 499934
rect 283022 499698 283204 499934
rect 282604 464254 283204 499698
rect 282604 464018 282786 464254
rect 283022 464018 283204 464254
rect 282604 463934 283204 464018
rect 282604 463698 282786 463934
rect 283022 463698 283204 463934
rect 282604 428254 283204 463698
rect 282604 428018 282786 428254
rect 283022 428018 283204 428254
rect 282604 427934 283204 428018
rect 282604 427698 282786 427934
rect 283022 427698 283204 427934
rect 282604 410000 283204 427698
rect 289804 704838 290404 705800
rect 289804 704602 289986 704838
rect 290222 704602 290404 704838
rect 289804 704518 290404 704602
rect 289804 704282 289986 704518
rect 290222 704282 290404 704518
rect 289804 687454 290404 704282
rect 289804 687218 289986 687454
rect 290222 687218 290404 687454
rect 289804 687134 290404 687218
rect 289804 686898 289986 687134
rect 290222 686898 290404 687134
rect 289804 651454 290404 686898
rect 289804 651218 289986 651454
rect 290222 651218 290404 651454
rect 289804 651134 290404 651218
rect 289804 650898 289986 651134
rect 290222 650898 290404 651134
rect 289804 615454 290404 650898
rect 289804 615218 289986 615454
rect 290222 615218 290404 615454
rect 289804 615134 290404 615218
rect 289804 614898 289986 615134
rect 290222 614898 290404 615134
rect 289804 579454 290404 614898
rect 289804 579218 289986 579454
rect 290222 579218 290404 579454
rect 289804 579134 290404 579218
rect 289804 578898 289986 579134
rect 290222 578898 290404 579134
rect 289804 543454 290404 578898
rect 289804 543218 289986 543454
rect 290222 543218 290404 543454
rect 289804 543134 290404 543218
rect 289804 542898 289986 543134
rect 290222 542898 290404 543134
rect 289804 507454 290404 542898
rect 289804 507218 289986 507454
rect 290222 507218 290404 507454
rect 289804 507134 290404 507218
rect 289804 506898 289986 507134
rect 290222 506898 290404 507134
rect 289804 471454 290404 506898
rect 289804 471218 289986 471454
rect 290222 471218 290404 471454
rect 289804 471134 290404 471218
rect 289804 470898 289986 471134
rect 290222 470898 290404 471134
rect 289804 435454 290404 470898
rect 289804 435218 289986 435454
rect 290222 435218 290404 435454
rect 289804 435134 290404 435218
rect 289804 434898 289986 435134
rect 290222 434898 290404 435134
rect 289804 410000 290404 434898
rect 293404 691054 294004 706162
rect 293404 690818 293586 691054
rect 293822 690818 294004 691054
rect 293404 690734 294004 690818
rect 293404 690498 293586 690734
rect 293822 690498 294004 690734
rect 293404 655054 294004 690498
rect 293404 654818 293586 655054
rect 293822 654818 294004 655054
rect 293404 654734 294004 654818
rect 293404 654498 293586 654734
rect 293822 654498 294004 654734
rect 293404 619054 294004 654498
rect 293404 618818 293586 619054
rect 293822 618818 294004 619054
rect 293404 618734 294004 618818
rect 293404 618498 293586 618734
rect 293822 618498 294004 618734
rect 293404 583054 294004 618498
rect 293404 582818 293586 583054
rect 293822 582818 294004 583054
rect 293404 582734 294004 582818
rect 293404 582498 293586 582734
rect 293822 582498 294004 582734
rect 293404 547054 294004 582498
rect 293404 546818 293586 547054
rect 293822 546818 294004 547054
rect 293404 546734 294004 546818
rect 293404 546498 293586 546734
rect 293822 546498 294004 546734
rect 293404 511054 294004 546498
rect 293404 510818 293586 511054
rect 293822 510818 294004 511054
rect 293404 510734 294004 510818
rect 293404 510498 293586 510734
rect 293822 510498 294004 510734
rect 293404 475054 294004 510498
rect 293404 474818 293586 475054
rect 293822 474818 294004 475054
rect 293404 474734 294004 474818
rect 293404 474498 293586 474734
rect 293822 474498 294004 474734
rect 293404 439054 294004 474498
rect 293404 438818 293586 439054
rect 293822 438818 294004 439054
rect 293404 438734 294004 438818
rect 293404 438498 293586 438734
rect 293822 438498 294004 438734
rect 293404 410000 294004 438498
rect 297004 694654 297604 708042
rect 297004 694418 297186 694654
rect 297422 694418 297604 694654
rect 297004 694334 297604 694418
rect 297004 694098 297186 694334
rect 297422 694098 297604 694334
rect 297004 658654 297604 694098
rect 297004 658418 297186 658654
rect 297422 658418 297604 658654
rect 297004 658334 297604 658418
rect 297004 658098 297186 658334
rect 297422 658098 297604 658334
rect 297004 622654 297604 658098
rect 297004 622418 297186 622654
rect 297422 622418 297604 622654
rect 297004 622334 297604 622418
rect 297004 622098 297186 622334
rect 297422 622098 297604 622334
rect 297004 586654 297604 622098
rect 297004 586418 297186 586654
rect 297422 586418 297604 586654
rect 297004 586334 297604 586418
rect 297004 586098 297186 586334
rect 297422 586098 297604 586334
rect 297004 550654 297604 586098
rect 297004 550418 297186 550654
rect 297422 550418 297604 550654
rect 297004 550334 297604 550418
rect 297004 550098 297186 550334
rect 297422 550098 297604 550334
rect 297004 514654 297604 550098
rect 297004 514418 297186 514654
rect 297422 514418 297604 514654
rect 297004 514334 297604 514418
rect 297004 514098 297186 514334
rect 297422 514098 297604 514334
rect 297004 478654 297604 514098
rect 297004 478418 297186 478654
rect 297422 478418 297604 478654
rect 297004 478334 297604 478418
rect 297004 478098 297186 478334
rect 297422 478098 297604 478334
rect 297004 442654 297604 478098
rect 297004 442418 297186 442654
rect 297422 442418 297604 442654
rect 297004 442334 297604 442418
rect 297004 442098 297186 442334
rect 297422 442098 297604 442334
rect 297004 410000 297604 442098
rect 300604 698254 301204 709922
rect 318604 711418 319204 711440
rect 318604 711182 318786 711418
rect 319022 711182 319204 711418
rect 318604 711098 319204 711182
rect 318604 710862 318786 711098
rect 319022 710862 319204 711098
rect 315004 709538 315604 709560
rect 315004 709302 315186 709538
rect 315422 709302 315604 709538
rect 315004 709218 315604 709302
rect 315004 708982 315186 709218
rect 315422 708982 315604 709218
rect 311404 707658 312004 707680
rect 311404 707422 311586 707658
rect 311822 707422 312004 707658
rect 311404 707338 312004 707422
rect 311404 707102 311586 707338
rect 311822 707102 312004 707338
rect 300604 698018 300786 698254
rect 301022 698018 301204 698254
rect 300604 697934 301204 698018
rect 300604 697698 300786 697934
rect 301022 697698 301204 697934
rect 300604 662254 301204 697698
rect 300604 662018 300786 662254
rect 301022 662018 301204 662254
rect 300604 661934 301204 662018
rect 300604 661698 300786 661934
rect 301022 661698 301204 661934
rect 300604 626254 301204 661698
rect 300604 626018 300786 626254
rect 301022 626018 301204 626254
rect 300604 625934 301204 626018
rect 300604 625698 300786 625934
rect 301022 625698 301204 625934
rect 300604 590254 301204 625698
rect 300604 590018 300786 590254
rect 301022 590018 301204 590254
rect 300604 589934 301204 590018
rect 300604 589698 300786 589934
rect 301022 589698 301204 589934
rect 300604 554254 301204 589698
rect 300604 554018 300786 554254
rect 301022 554018 301204 554254
rect 300604 553934 301204 554018
rect 300604 553698 300786 553934
rect 301022 553698 301204 553934
rect 300604 518254 301204 553698
rect 300604 518018 300786 518254
rect 301022 518018 301204 518254
rect 300604 517934 301204 518018
rect 300604 517698 300786 517934
rect 301022 517698 301204 517934
rect 300604 482254 301204 517698
rect 300604 482018 300786 482254
rect 301022 482018 301204 482254
rect 300604 481934 301204 482018
rect 300604 481698 300786 481934
rect 301022 481698 301204 481934
rect 300604 446254 301204 481698
rect 300604 446018 300786 446254
rect 301022 446018 301204 446254
rect 300604 445934 301204 446018
rect 300604 445698 300786 445934
rect 301022 445698 301204 445934
rect 300604 410000 301204 445698
rect 307804 705778 308404 705800
rect 307804 705542 307986 705778
rect 308222 705542 308404 705778
rect 307804 705458 308404 705542
rect 307804 705222 307986 705458
rect 308222 705222 308404 705458
rect 307804 669454 308404 705222
rect 307804 669218 307986 669454
rect 308222 669218 308404 669454
rect 307804 669134 308404 669218
rect 307804 668898 307986 669134
rect 308222 668898 308404 669134
rect 307804 633454 308404 668898
rect 307804 633218 307986 633454
rect 308222 633218 308404 633454
rect 307804 633134 308404 633218
rect 307804 632898 307986 633134
rect 308222 632898 308404 633134
rect 307804 597454 308404 632898
rect 307804 597218 307986 597454
rect 308222 597218 308404 597454
rect 307804 597134 308404 597218
rect 307804 596898 307986 597134
rect 308222 596898 308404 597134
rect 307804 561454 308404 596898
rect 307804 561218 307986 561454
rect 308222 561218 308404 561454
rect 307804 561134 308404 561218
rect 307804 560898 307986 561134
rect 308222 560898 308404 561134
rect 307804 525454 308404 560898
rect 307804 525218 307986 525454
rect 308222 525218 308404 525454
rect 307804 525134 308404 525218
rect 307804 524898 307986 525134
rect 308222 524898 308404 525134
rect 307804 489454 308404 524898
rect 307804 489218 307986 489454
rect 308222 489218 308404 489454
rect 307804 489134 308404 489218
rect 307804 488898 307986 489134
rect 308222 488898 308404 489134
rect 307804 453454 308404 488898
rect 307804 453218 307986 453454
rect 308222 453218 308404 453454
rect 307804 453134 308404 453218
rect 307804 452898 307986 453134
rect 308222 452898 308404 453134
rect 307804 417454 308404 452898
rect 307804 417218 307986 417454
rect 308222 417218 308404 417454
rect 307804 417134 308404 417218
rect 307804 416898 307986 417134
rect 308222 416898 308404 417134
rect 228604 409698 228786 409934
rect 229022 409698 229204 409934
rect 228604 374254 229204 409698
rect 228604 374018 228786 374254
rect 229022 374018 229204 374254
rect 228604 373934 229204 374018
rect 228604 373698 228786 373934
rect 229022 373698 229204 373934
rect 228604 338254 229204 373698
rect 307804 381454 308404 416898
rect 307804 381218 307986 381454
rect 308222 381218 308404 381454
rect 307804 381134 308404 381218
rect 307804 380898 307986 381134
rect 308222 380898 308404 381134
rect 307804 345454 308404 380898
rect 307804 345218 307986 345454
rect 308222 345218 308404 345454
rect 307804 345134 308404 345218
rect 307804 344898 307986 345134
rect 308222 344898 308404 345134
rect 306971 340916 307037 340917
rect 306971 340852 306972 340916
rect 307036 340852 307037 340916
rect 306971 340851 307037 340852
rect 228604 338018 228786 338254
rect 229022 338018 229204 338254
rect 228604 337934 229204 338018
rect 228604 337698 228786 337934
rect 229022 337698 229204 337934
rect 228604 302254 229204 337698
rect 228604 302018 228786 302254
rect 229022 302018 229204 302254
rect 228604 301934 229204 302018
rect 228604 301698 228786 301934
rect 229022 301698 229204 301934
rect 228604 266254 229204 301698
rect 228604 266018 228786 266254
rect 229022 266018 229204 266254
rect 228604 265934 229204 266018
rect 228604 265698 228786 265934
rect 229022 265698 229204 265934
rect 228604 230254 229204 265698
rect 228604 230018 228786 230254
rect 229022 230018 229204 230254
rect 228604 229934 229204 230018
rect 228604 229698 228786 229934
rect 229022 229698 229204 229934
rect 228604 194254 229204 229698
rect 228604 194018 228786 194254
rect 229022 194018 229204 194254
rect 228604 193934 229204 194018
rect 228604 193698 228786 193934
rect 229022 193698 229204 193934
rect 228604 158254 229204 193698
rect 228604 158018 228786 158254
rect 229022 158018 229204 158254
rect 228604 157934 229204 158018
rect 228604 157698 228786 157934
rect 229022 157698 229204 157934
rect 228604 122254 229204 157698
rect 228604 122018 228786 122254
rect 229022 122018 229204 122254
rect 228604 121934 229204 122018
rect 228604 121698 228786 121934
rect 229022 121698 229204 121934
rect 228604 86254 229204 121698
rect 228604 86018 228786 86254
rect 229022 86018 229204 86254
rect 228604 85934 229204 86018
rect 228604 85698 228786 85934
rect 229022 85698 229204 85934
rect 228604 50254 229204 85698
rect 228604 50018 228786 50254
rect 229022 50018 229204 50254
rect 228604 49934 229204 50018
rect 228604 49698 228786 49934
rect 229022 49698 229204 49934
rect 228604 14254 229204 49698
rect 228604 14018 228786 14254
rect 229022 14018 229204 14254
rect 228604 13934 229204 14018
rect 228604 13698 228786 13934
rect 229022 13698 229204 13934
rect 210604 -7162 210786 -6926
rect 211022 -7162 211204 -6926
rect 210604 -7246 211204 -7162
rect 210604 -7482 210786 -7246
rect 211022 -7482 211204 -7246
rect 210604 -7504 211204 -7482
rect 228604 -5986 229204 13698
rect 235804 309454 236404 336000
rect 235804 309218 235986 309454
rect 236222 309218 236404 309454
rect 235804 309134 236404 309218
rect 235804 308898 235986 309134
rect 236222 308898 236404 309134
rect 235804 273454 236404 308898
rect 235804 273218 235986 273454
rect 236222 273218 236404 273454
rect 235804 273134 236404 273218
rect 235804 272898 235986 273134
rect 236222 272898 236404 273134
rect 235804 237454 236404 272898
rect 235804 237218 235986 237454
rect 236222 237218 236404 237454
rect 235804 237134 236404 237218
rect 235804 236898 235986 237134
rect 236222 236898 236404 237134
rect 235804 201454 236404 236898
rect 235804 201218 235986 201454
rect 236222 201218 236404 201454
rect 235804 201134 236404 201218
rect 235804 200898 235986 201134
rect 236222 200898 236404 201134
rect 235804 165454 236404 200898
rect 235804 165218 235986 165454
rect 236222 165218 236404 165454
rect 235804 165134 236404 165218
rect 235804 164898 235986 165134
rect 236222 164898 236404 165134
rect 235804 129454 236404 164898
rect 235804 129218 235986 129454
rect 236222 129218 236404 129454
rect 235804 129134 236404 129218
rect 235804 128898 235986 129134
rect 236222 128898 236404 129134
rect 235804 93454 236404 128898
rect 235804 93218 235986 93454
rect 236222 93218 236404 93454
rect 235804 93134 236404 93218
rect 235804 92898 235986 93134
rect 236222 92898 236404 93134
rect 235804 57454 236404 92898
rect 235804 57218 235986 57454
rect 236222 57218 236404 57454
rect 235804 57134 236404 57218
rect 235804 56898 235986 57134
rect 236222 56898 236404 57134
rect 235804 21454 236404 56898
rect 235804 21218 235986 21454
rect 236222 21218 236404 21454
rect 235804 21134 236404 21218
rect 235804 20898 235986 21134
rect 236222 20898 236404 21134
rect 235804 -1286 236404 20898
rect 235804 -1522 235986 -1286
rect 236222 -1522 236404 -1286
rect 235804 -1606 236404 -1522
rect 235804 -1842 235986 -1606
rect 236222 -1842 236404 -1606
rect 235804 -1864 236404 -1842
rect 239404 313054 240004 336000
rect 239404 312818 239586 313054
rect 239822 312818 240004 313054
rect 239404 312734 240004 312818
rect 239404 312498 239586 312734
rect 239822 312498 240004 312734
rect 239404 277054 240004 312498
rect 239404 276818 239586 277054
rect 239822 276818 240004 277054
rect 239404 276734 240004 276818
rect 239404 276498 239586 276734
rect 239822 276498 240004 276734
rect 239404 241054 240004 276498
rect 239404 240818 239586 241054
rect 239822 240818 240004 241054
rect 239404 240734 240004 240818
rect 239404 240498 239586 240734
rect 239822 240498 240004 240734
rect 239404 205054 240004 240498
rect 239404 204818 239586 205054
rect 239822 204818 240004 205054
rect 239404 204734 240004 204818
rect 239404 204498 239586 204734
rect 239822 204498 240004 204734
rect 239404 169054 240004 204498
rect 239404 168818 239586 169054
rect 239822 168818 240004 169054
rect 239404 168734 240004 168818
rect 239404 168498 239586 168734
rect 239822 168498 240004 168734
rect 239404 133054 240004 168498
rect 239404 132818 239586 133054
rect 239822 132818 240004 133054
rect 239404 132734 240004 132818
rect 239404 132498 239586 132734
rect 239822 132498 240004 132734
rect 239404 97054 240004 132498
rect 239404 96818 239586 97054
rect 239822 96818 240004 97054
rect 239404 96734 240004 96818
rect 239404 96498 239586 96734
rect 239822 96498 240004 96734
rect 239404 61054 240004 96498
rect 239404 60818 239586 61054
rect 239822 60818 240004 61054
rect 239404 60734 240004 60818
rect 239404 60498 239586 60734
rect 239822 60498 240004 60734
rect 239404 25054 240004 60498
rect 239404 24818 239586 25054
rect 239822 24818 240004 25054
rect 239404 24734 240004 24818
rect 239404 24498 239586 24734
rect 239822 24498 240004 24734
rect 239404 -3166 240004 24498
rect 239404 -3402 239586 -3166
rect 239822 -3402 240004 -3166
rect 239404 -3486 240004 -3402
rect 239404 -3722 239586 -3486
rect 239822 -3722 240004 -3486
rect 239404 -3744 240004 -3722
rect 243004 316654 243604 336000
rect 243004 316418 243186 316654
rect 243422 316418 243604 316654
rect 243004 316334 243604 316418
rect 243004 316098 243186 316334
rect 243422 316098 243604 316334
rect 243004 280654 243604 316098
rect 243004 280418 243186 280654
rect 243422 280418 243604 280654
rect 243004 280334 243604 280418
rect 243004 280098 243186 280334
rect 243422 280098 243604 280334
rect 243004 244654 243604 280098
rect 243004 244418 243186 244654
rect 243422 244418 243604 244654
rect 243004 244334 243604 244418
rect 243004 244098 243186 244334
rect 243422 244098 243604 244334
rect 243004 208654 243604 244098
rect 243004 208418 243186 208654
rect 243422 208418 243604 208654
rect 243004 208334 243604 208418
rect 243004 208098 243186 208334
rect 243422 208098 243604 208334
rect 243004 172654 243604 208098
rect 243004 172418 243186 172654
rect 243422 172418 243604 172654
rect 243004 172334 243604 172418
rect 243004 172098 243186 172334
rect 243422 172098 243604 172334
rect 243004 136654 243604 172098
rect 243004 136418 243186 136654
rect 243422 136418 243604 136654
rect 243004 136334 243604 136418
rect 243004 136098 243186 136334
rect 243422 136098 243604 136334
rect 243004 100654 243604 136098
rect 243004 100418 243186 100654
rect 243422 100418 243604 100654
rect 243004 100334 243604 100418
rect 243004 100098 243186 100334
rect 243422 100098 243604 100334
rect 243004 64654 243604 100098
rect 243004 64418 243186 64654
rect 243422 64418 243604 64654
rect 243004 64334 243604 64418
rect 243004 64098 243186 64334
rect 243422 64098 243604 64334
rect 243004 28654 243604 64098
rect 243004 28418 243186 28654
rect 243422 28418 243604 28654
rect 243004 28334 243604 28418
rect 243004 28098 243186 28334
rect 243422 28098 243604 28334
rect 243004 -5046 243604 28098
rect 243004 -5282 243186 -5046
rect 243422 -5282 243604 -5046
rect 243004 -5366 243604 -5282
rect 243004 -5602 243186 -5366
rect 243422 -5602 243604 -5366
rect 243004 -5624 243604 -5602
rect 246604 320254 247204 336000
rect 246604 320018 246786 320254
rect 247022 320018 247204 320254
rect 246604 319934 247204 320018
rect 246604 319698 246786 319934
rect 247022 319698 247204 319934
rect 246604 284254 247204 319698
rect 246604 284018 246786 284254
rect 247022 284018 247204 284254
rect 246604 283934 247204 284018
rect 246604 283698 246786 283934
rect 247022 283698 247204 283934
rect 246604 248254 247204 283698
rect 246604 248018 246786 248254
rect 247022 248018 247204 248254
rect 246604 247934 247204 248018
rect 246604 247698 246786 247934
rect 247022 247698 247204 247934
rect 246604 212254 247204 247698
rect 246604 212018 246786 212254
rect 247022 212018 247204 212254
rect 246604 211934 247204 212018
rect 246604 211698 246786 211934
rect 247022 211698 247204 211934
rect 246604 176254 247204 211698
rect 246604 176018 246786 176254
rect 247022 176018 247204 176254
rect 246604 175934 247204 176018
rect 246604 175698 246786 175934
rect 247022 175698 247204 175934
rect 246604 140254 247204 175698
rect 246604 140018 246786 140254
rect 247022 140018 247204 140254
rect 246604 139934 247204 140018
rect 246604 139698 246786 139934
rect 247022 139698 247204 139934
rect 246604 104254 247204 139698
rect 246604 104018 246786 104254
rect 247022 104018 247204 104254
rect 246604 103934 247204 104018
rect 246604 103698 246786 103934
rect 247022 103698 247204 103934
rect 246604 68254 247204 103698
rect 246604 68018 246786 68254
rect 247022 68018 247204 68254
rect 246604 67934 247204 68018
rect 246604 67698 246786 67934
rect 247022 67698 247204 67934
rect 246604 32254 247204 67698
rect 246604 32018 246786 32254
rect 247022 32018 247204 32254
rect 246604 31934 247204 32018
rect 246604 31698 246786 31934
rect 247022 31698 247204 31934
rect 228604 -6222 228786 -5986
rect 229022 -6222 229204 -5986
rect 228604 -6306 229204 -6222
rect 228604 -6542 228786 -6306
rect 229022 -6542 229204 -6306
rect 228604 -7504 229204 -6542
rect 246604 -6926 247204 31698
rect 253804 327454 254404 336000
rect 253804 327218 253986 327454
rect 254222 327218 254404 327454
rect 253804 327134 254404 327218
rect 253804 326898 253986 327134
rect 254222 326898 254404 327134
rect 253804 291454 254404 326898
rect 253804 291218 253986 291454
rect 254222 291218 254404 291454
rect 253804 291134 254404 291218
rect 253804 290898 253986 291134
rect 254222 290898 254404 291134
rect 253804 255454 254404 290898
rect 253804 255218 253986 255454
rect 254222 255218 254404 255454
rect 253804 255134 254404 255218
rect 253804 254898 253986 255134
rect 254222 254898 254404 255134
rect 253804 219454 254404 254898
rect 253804 219218 253986 219454
rect 254222 219218 254404 219454
rect 253804 219134 254404 219218
rect 253804 218898 253986 219134
rect 254222 218898 254404 219134
rect 253804 183454 254404 218898
rect 253804 183218 253986 183454
rect 254222 183218 254404 183454
rect 253804 183134 254404 183218
rect 253804 182898 253986 183134
rect 254222 182898 254404 183134
rect 253804 147454 254404 182898
rect 253804 147218 253986 147454
rect 254222 147218 254404 147454
rect 253804 147134 254404 147218
rect 253804 146898 253986 147134
rect 254222 146898 254404 147134
rect 253804 111454 254404 146898
rect 253804 111218 253986 111454
rect 254222 111218 254404 111454
rect 253804 111134 254404 111218
rect 253804 110898 253986 111134
rect 254222 110898 254404 111134
rect 253804 75454 254404 110898
rect 253804 75218 253986 75454
rect 254222 75218 254404 75454
rect 253804 75134 254404 75218
rect 253804 74898 253986 75134
rect 254222 74898 254404 75134
rect 253804 39454 254404 74898
rect 253804 39218 253986 39454
rect 254222 39218 254404 39454
rect 253804 39134 254404 39218
rect 253804 38898 253986 39134
rect 254222 38898 254404 39134
rect 253804 3454 254404 38898
rect 253804 3218 253986 3454
rect 254222 3218 254404 3454
rect 253804 3134 254404 3218
rect 253804 2898 253986 3134
rect 254222 2898 254404 3134
rect 253804 -346 254404 2898
rect 253804 -582 253986 -346
rect 254222 -582 254404 -346
rect 253804 -666 254404 -582
rect 253804 -902 253986 -666
rect 254222 -902 254404 -666
rect 253804 -1864 254404 -902
rect 257404 331054 258004 336000
rect 257404 330818 257586 331054
rect 257822 330818 258004 331054
rect 257404 330734 258004 330818
rect 257404 330498 257586 330734
rect 257822 330498 258004 330734
rect 257404 295054 258004 330498
rect 257404 294818 257586 295054
rect 257822 294818 258004 295054
rect 257404 294734 258004 294818
rect 257404 294498 257586 294734
rect 257822 294498 258004 294734
rect 257404 259054 258004 294498
rect 257404 258818 257586 259054
rect 257822 258818 258004 259054
rect 257404 258734 258004 258818
rect 257404 258498 257586 258734
rect 257822 258498 258004 258734
rect 257404 223054 258004 258498
rect 257404 222818 257586 223054
rect 257822 222818 258004 223054
rect 257404 222734 258004 222818
rect 257404 222498 257586 222734
rect 257822 222498 258004 222734
rect 257404 187054 258004 222498
rect 257404 186818 257586 187054
rect 257822 186818 258004 187054
rect 257404 186734 258004 186818
rect 257404 186498 257586 186734
rect 257822 186498 258004 186734
rect 257404 151054 258004 186498
rect 257404 150818 257586 151054
rect 257822 150818 258004 151054
rect 257404 150734 258004 150818
rect 257404 150498 257586 150734
rect 257822 150498 258004 150734
rect 257404 115054 258004 150498
rect 257404 114818 257586 115054
rect 257822 114818 258004 115054
rect 257404 114734 258004 114818
rect 257404 114498 257586 114734
rect 257822 114498 258004 114734
rect 257404 79054 258004 114498
rect 257404 78818 257586 79054
rect 257822 78818 258004 79054
rect 257404 78734 258004 78818
rect 257404 78498 257586 78734
rect 257822 78498 258004 78734
rect 257404 43054 258004 78498
rect 257404 42818 257586 43054
rect 257822 42818 258004 43054
rect 257404 42734 258004 42818
rect 257404 42498 257586 42734
rect 257822 42498 258004 42734
rect 257404 7054 258004 42498
rect 257404 6818 257586 7054
rect 257822 6818 258004 7054
rect 257404 6734 258004 6818
rect 257404 6498 257586 6734
rect 257822 6498 258004 6734
rect 257404 -2226 258004 6498
rect 257404 -2462 257586 -2226
rect 257822 -2462 258004 -2226
rect 257404 -2546 258004 -2462
rect 257404 -2782 257586 -2546
rect 257822 -2782 258004 -2546
rect 257404 -3744 258004 -2782
rect 261004 334654 261604 336000
rect 261004 334418 261186 334654
rect 261422 334418 261604 334654
rect 261004 334334 261604 334418
rect 261004 334098 261186 334334
rect 261422 334098 261604 334334
rect 261004 298654 261604 334098
rect 261004 298418 261186 298654
rect 261422 298418 261604 298654
rect 261004 298334 261604 298418
rect 261004 298098 261186 298334
rect 261422 298098 261604 298334
rect 261004 262654 261604 298098
rect 261004 262418 261186 262654
rect 261422 262418 261604 262654
rect 261004 262334 261604 262418
rect 261004 262098 261186 262334
rect 261422 262098 261604 262334
rect 261004 226654 261604 262098
rect 261004 226418 261186 226654
rect 261422 226418 261604 226654
rect 261004 226334 261604 226418
rect 261004 226098 261186 226334
rect 261422 226098 261604 226334
rect 261004 190654 261604 226098
rect 261004 190418 261186 190654
rect 261422 190418 261604 190654
rect 261004 190334 261604 190418
rect 261004 190098 261186 190334
rect 261422 190098 261604 190334
rect 261004 154654 261604 190098
rect 261004 154418 261186 154654
rect 261422 154418 261604 154654
rect 261004 154334 261604 154418
rect 261004 154098 261186 154334
rect 261422 154098 261604 154334
rect 261004 118654 261604 154098
rect 261004 118418 261186 118654
rect 261422 118418 261604 118654
rect 261004 118334 261604 118418
rect 261004 118098 261186 118334
rect 261422 118098 261604 118334
rect 261004 82654 261604 118098
rect 261004 82418 261186 82654
rect 261422 82418 261604 82654
rect 261004 82334 261604 82418
rect 261004 82098 261186 82334
rect 261422 82098 261604 82334
rect 261004 46654 261604 82098
rect 261004 46418 261186 46654
rect 261422 46418 261604 46654
rect 261004 46334 261604 46418
rect 261004 46098 261186 46334
rect 261422 46098 261604 46334
rect 261004 10654 261604 46098
rect 261004 10418 261186 10654
rect 261422 10418 261604 10654
rect 261004 10334 261604 10418
rect 261004 10098 261186 10334
rect 261422 10098 261604 10334
rect 261004 -4106 261604 10098
rect 261004 -4342 261186 -4106
rect 261422 -4342 261604 -4106
rect 261004 -4426 261604 -4342
rect 261004 -4662 261186 -4426
rect 261422 -4662 261604 -4426
rect 261004 -5624 261604 -4662
rect 264604 302254 265204 336000
rect 264604 302018 264786 302254
rect 265022 302018 265204 302254
rect 264604 301934 265204 302018
rect 264604 301698 264786 301934
rect 265022 301698 265204 301934
rect 264604 266254 265204 301698
rect 264604 266018 264786 266254
rect 265022 266018 265204 266254
rect 264604 265934 265204 266018
rect 264604 265698 264786 265934
rect 265022 265698 265204 265934
rect 264604 230254 265204 265698
rect 264604 230018 264786 230254
rect 265022 230018 265204 230254
rect 264604 229934 265204 230018
rect 264604 229698 264786 229934
rect 265022 229698 265204 229934
rect 264604 194254 265204 229698
rect 264604 194018 264786 194254
rect 265022 194018 265204 194254
rect 264604 193934 265204 194018
rect 264604 193698 264786 193934
rect 265022 193698 265204 193934
rect 264604 158254 265204 193698
rect 264604 158018 264786 158254
rect 265022 158018 265204 158254
rect 264604 157934 265204 158018
rect 264604 157698 264786 157934
rect 265022 157698 265204 157934
rect 264604 122254 265204 157698
rect 264604 122018 264786 122254
rect 265022 122018 265204 122254
rect 264604 121934 265204 122018
rect 264604 121698 264786 121934
rect 265022 121698 265204 121934
rect 264604 86254 265204 121698
rect 264604 86018 264786 86254
rect 265022 86018 265204 86254
rect 264604 85934 265204 86018
rect 264604 85698 264786 85934
rect 265022 85698 265204 85934
rect 264604 50254 265204 85698
rect 264604 50018 264786 50254
rect 265022 50018 265204 50254
rect 264604 49934 265204 50018
rect 264604 49698 264786 49934
rect 265022 49698 265204 49934
rect 264604 14254 265204 49698
rect 264604 14018 264786 14254
rect 265022 14018 265204 14254
rect 264604 13934 265204 14018
rect 264604 13698 264786 13934
rect 265022 13698 265204 13934
rect 246604 -7162 246786 -6926
rect 247022 -7162 247204 -6926
rect 246604 -7246 247204 -7162
rect 246604 -7482 246786 -7246
rect 247022 -7482 247204 -7246
rect 246604 -7504 247204 -7482
rect 264604 -5986 265204 13698
rect 271804 309454 272404 336000
rect 271804 309218 271986 309454
rect 272222 309218 272404 309454
rect 271804 309134 272404 309218
rect 271804 308898 271986 309134
rect 272222 308898 272404 309134
rect 271804 273454 272404 308898
rect 271804 273218 271986 273454
rect 272222 273218 272404 273454
rect 271804 273134 272404 273218
rect 271804 272898 271986 273134
rect 272222 272898 272404 273134
rect 271804 237454 272404 272898
rect 271804 237218 271986 237454
rect 272222 237218 272404 237454
rect 271804 237134 272404 237218
rect 271804 236898 271986 237134
rect 272222 236898 272404 237134
rect 271804 201454 272404 236898
rect 271804 201218 271986 201454
rect 272222 201218 272404 201454
rect 271804 201134 272404 201218
rect 271804 200898 271986 201134
rect 272222 200898 272404 201134
rect 271804 165454 272404 200898
rect 271804 165218 271986 165454
rect 272222 165218 272404 165454
rect 271804 165134 272404 165218
rect 271804 164898 271986 165134
rect 272222 164898 272404 165134
rect 271804 129454 272404 164898
rect 271804 129218 271986 129454
rect 272222 129218 272404 129454
rect 271804 129134 272404 129218
rect 271804 128898 271986 129134
rect 272222 128898 272404 129134
rect 271804 93454 272404 128898
rect 271804 93218 271986 93454
rect 272222 93218 272404 93454
rect 271804 93134 272404 93218
rect 271804 92898 271986 93134
rect 272222 92898 272404 93134
rect 271804 57454 272404 92898
rect 271804 57218 271986 57454
rect 272222 57218 272404 57454
rect 271804 57134 272404 57218
rect 271804 56898 271986 57134
rect 272222 56898 272404 57134
rect 271804 21454 272404 56898
rect 271804 21218 271986 21454
rect 272222 21218 272404 21454
rect 271804 21134 272404 21218
rect 271804 20898 271986 21134
rect 272222 20898 272404 21134
rect 271804 -1286 272404 20898
rect 271804 -1522 271986 -1286
rect 272222 -1522 272404 -1286
rect 271804 -1606 272404 -1522
rect 271804 -1842 271986 -1606
rect 272222 -1842 272404 -1606
rect 271804 -1864 272404 -1842
rect 275404 313054 276004 336000
rect 275404 312818 275586 313054
rect 275822 312818 276004 313054
rect 275404 312734 276004 312818
rect 275404 312498 275586 312734
rect 275822 312498 276004 312734
rect 275404 277054 276004 312498
rect 275404 276818 275586 277054
rect 275822 276818 276004 277054
rect 275404 276734 276004 276818
rect 275404 276498 275586 276734
rect 275822 276498 276004 276734
rect 275404 241054 276004 276498
rect 275404 240818 275586 241054
rect 275822 240818 276004 241054
rect 275404 240734 276004 240818
rect 275404 240498 275586 240734
rect 275822 240498 276004 240734
rect 275404 205054 276004 240498
rect 275404 204818 275586 205054
rect 275822 204818 276004 205054
rect 275404 204734 276004 204818
rect 275404 204498 275586 204734
rect 275822 204498 276004 204734
rect 275404 169054 276004 204498
rect 275404 168818 275586 169054
rect 275822 168818 276004 169054
rect 275404 168734 276004 168818
rect 275404 168498 275586 168734
rect 275822 168498 276004 168734
rect 275404 133054 276004 168498
rect 275404 132818 275586 133054
rect 275822 132818 276004 133054
rect 275404 132734 276004 132818
rect 275404 132498 275586 132734
rect 275822 132498 276004 132734
rect 275404 97054 276004 132498
rect 275404 96818 275586 97054
rect 275822 96818 276004 97054
rect 275404 96734 276004 96818
rect 275404 96498 275586 96734
rect 275822 96498 276004 96734
rect 275404 61054 276004 96498
rect 275404 60818 275586 61054
rect 275822 60818 276004 61054
rect 275404 60734 276004 60818
rect 275404 60498 275586 60734
rect 275822 60498 276004 60734
rect 275404 25054 276004 60498
rect 275404 24818 275586 25054
rect 275822 24818 276004 25054
rect 275404 24734 276004 24818
rect 275404 24498 275586 24734
rect 275822 24498 276004 24734
rect 275404 -3166 276004 24498
rect 275404 -3402 275586 -3166
rect 275822 -3402 276004 -3166
rect 275404 -3486 276004 -3402
rect 275404 -3722 275586 -3486
rect 275822 -3722 276004 -3486
rect 275404 -3744 276004 -3722
rect 279004 316654 279604 336000
rect 279004 316418 279186 316654
rect 279422 316418 279604 316654
rect 279004 316334 279604 316418
rect 279004 316098 279186 316334
rect 279422 316098 279604 316334
rect 279004 280654 279604 316098
rect 279004 280418 279186 280654
rect 279422 280418 279604 280654
rect 279004 280334 279604 280418
rect 279004 280098 279186 280334
rect 279422 280098 279604 280334
rect 279004 244654 279604 280098
rect 279004 244418 279186 244654
rect 279422 244418 279604 244654
rect 279004 244334 279604 244418
rect 279004 244098 279186 244334
rect 279422 244098 279604 244334
rect 279004 208654 279604 244098
rect 279004 208418 279186 208654
rect 279422 208418 279604 208654
rect 279004 208334 279604 208418
rect 279004 208098 279186 208334
rect 279422 208098 279604 208334
rect 279004 172654 279604 208098
rect 279004 172418 279186 172654
rect 279422 172418 279604 172654
rect 279004 172334 279604 172418
rect 279004 172098 279186 172334
rect 279422 172098 279604 172334
rect 279004 136654 279604 172098
rect 279004 136418 279186 136654
rect 279422 136418 279604 136654
rect 279004 136334 279604 136418
rect 279004 136098 279186 136334
rect 279422 136098 279604 136334
rect 279004 100654 279604 136098
rect 279004 100418 279186 100654
rect 279422 100418 279604 100654
rect 279004 100334 279604 100418
rect 279004 100098 279186 100334
rect 279422 100098 279604 100334
rect 279004 64654 279604 100098
rect 279004 64418 279186 64654
rect 279422 64418 279604 64654
rect 279004 64334 279604 64418
rect 279004 64098 279186 64334
rect 279422 64098 279604 64334
rect 279004 28654 279604 64098
rect 279004 28418 279186 28654
rect 279422 28418 279604 28654
rect 279004 28334 279604 28418
rect 279004 28098 279186 28334
rect 279422 28098 279604 28334
rect 279004 -5046 279604 28098
rect 279004 -5282 279186 -5046
rect 279422 -5282 279604 -5046
rect 279004 -5366 279604 -5282
rect 279004 -5602 279186 -5366
rect 279422 -5602 279604 -5366
rect 279004 -5624 279604 -5602
rect 282604 320254 283204 336000
rect 282604 320018 282786 320254
rect 283022 320018 283204 320254
rect 282604 319934 283204 320018
rect 282604 319698 282786 319934
rect 283022 319698 283204 319934
rect 282604 284254 283204 319698
rect 282604 284018 282786 284254
rect 283022 284018 283204 284254
rect 282604 283934 283204 284018
rect 282604 283698 282786 283934
rect 283022 283698 283204 283934
rect 282604 248254 283204 283698
rect 282604 248018 282786 248254
rect 283022 248018 283204 248254
rect 282604 247934 283204 248018
rect 282604 247698 282786 247934
rect 283022 247698 283204 247934
rect 282604 212254 283204 247698
rect 282604 212018 282786 212254
rect 283022 212018 283204 212254
rect 282604 211934 283204 212018
rect 282604 211698 282786 211934
rect 283022 211698 283204 211934
rect 282604 176254 283204 211698
rect 282604 176018 282786 176254
rect 283022 176018 283204 176254
rect 282604 175934 283204 176018
rect 282604 175698 282786 175934
rect 283022 175698 283204 175934
rect 282604 140254 283204 175698
rect 282604 140018 282786 140254
rect 283022 140018 283204 140254
rect 282604 139934 283204 140018
rect 282604 139698 282786 139934
rect 283022 139698 283204 139934
rect 282604 104254 283204 139698
rect 282604 104018 282786 104254
rect 283022 104018 283204 104254
rect 282604 103934 283204 104018
rect 282604 103698 282786 103934
rect 283022 103698 283204 103934
rect 282604 68254 283204 103698
rect 282604 68018 282786 68254
rect 283022 68018 283204 68254
rect 282604 67934 283204 68018
rect 282604 67698 282786 67934
rect 283022 67698 283204 67934
rect 282604 32254 283204 67698
rect 282604 32018 282786 32254
rect 283022 32018 283204 32254
rect 282604 31934 283204 32018
rect 282604 31698 282786 31934
rect 283022 31698 283204 31934
rect 264604 -6222 264786 -5986
rect 265022 -6222 265204 -5986
rect 264604 -6306 265204 -6222
rect 264604 -6542 264786 -6306
rect 265022 -6542 265204 -6306
rect 264604 -7504 265204 -6542
rect 282604 -6926 283204 31698
rect 289804 327454 290404 336000
rect 289804 327218 289986 327454
rect 290222 327218 290404 327454
rect 289804 327134 290404 327218
rect 289804 326898 289986 327134
rect 290222 326898 290404 327134
rect 289804 291454 290404 326898
rect 289804 291218 289986 291454
rect 290222 291218 290404 291454
rect 289804 291134 290404 291218
rect 289804 290898 289986 291134
rect 290222 290898 290404 291134
rect 289804 255454 290404 290898
rect 289804 255218 289986 255454
rect 290222 255218 290404 255454
rect 289804 255134 290404 255218
rect 289804 254898 289986 255134
rect 290222 254898 290404 255134
rect 289804 219454 290404 254898
rect 289804 219218 289986 219454
rect 290222 219218 290404 219454
rect 289804 219134 290404 219218
rect 289804 218898 289986 219134
rect 290222 218898 290404 219134
rect 289804 183454 290404 218898
rect 289804 183218 289986 183454
rect 290222 183218 290404 183454
rect 289804 183134 290404 183218
rect 289804 182898 289986 183134
rect 290222 182898 290404 183134
rect 289804 147454 290404 182898
rect 289804 147218 289986 147454
rect 290222 147218 290404 147454
rect 289804 147134 290404 147218
rect 289804 146898 289986 147134
rect 290222 146898 290404 147134
rect 289804 111454 290404 146898
rect 289804 111218 289986 111454
rect 290222 111218 290404 111454
rect 289804 111134 290404 111218
rect 289804 110898 289986 111134
rect 290222 110898 290404 111134
rect 289804 75454 290404 110898
rect 289804 75218 289986 75454
rect 290222 75218 290404 75454
rect 289804 75134 290404 75218
rect 289804 74898 289986 75134
rect 290222 74898 290404 75134
rect 289804 39454 290404 74898
rect 289804 39218 289986 39454
rect 290222 39218 290404 39454
rect 289804 39134 290404 39218
rect 289804 38898 289986 39134
rect 290222 38898 290404 39134
rect 289804 3454 290404 38898
rect 289804 3218 289986 3454
rect 290222 3218 290404 3454
rect 289804 3134 290404 3218
rect 289804 2898 289986 3134
rect 290222 2898 290404 3134
rect 289804 -346 290404 2898
rect 289804 -582 289986 -346
rect 290222 -582 290404 -346
rect 289804 -666 290404 -582
rect 289804 -902 289986 -666
rect 290222 -902 290404 -666
rect 289804 -1864 290404 -902
rect 293404 331054 294004 336000
rect 293404 330818 293586 331054
rect 293822 330818 294004 331054
rect 293404 330734 294004 330818
rect 293404 330498 293586 330734
rect 293822 330498 294004 330734
rect 293404 295054 294004 330498
rect 293404 294818 293586 295054
rect 293822 294818 294004 295054
rect 293404 294734 294004 294818
rect 293404 294498 293586 294734
rect 293822 294498 294004 294734
rect 293404 259054 294004 294498
rect 293404 258818 293586 259054
rect 293822 258818 294004 259054
rect 293404 258734 294004 258818
rect 293404 258498 293586 258734
rect 293822 258498 294004 258734
rect 293404 223054 294004 258498
rect 293404 222818 293586 223054
rect 293822 222818 294004 223054
rect 293404 222734 294004 222818
rect 293404 222498 293586 222734
rect 293822 222498 294004 222734
rect 293404 187054 294004 222498
rect 293404 186818 293586 187054
rect 293822 186818 294004 187054
rect 293404 186734 294004 186818
rect 293404 186498 293586 186734
rect 293822 186498 294004 186734
rect 293404 151054 294004 186498
rect 293404 150818 293586 151054
rect 293822 150818 294004 151054
rect 293404 150734 294004 150818
rect 293404 150498 293586 150734
rect 293822 150498 294004 150734
rect 293404 115054 294004 150498
rect 293404 114818 293586 115054
rect 293822 114818 294004 115054
rect 293404 114734 294004 114818
rect 293404 114498 293586 114734
rect 293822 114498 294004 114734
rect 293404 79054 294004 114498
rect 293404 78818 293586 79054
rect 293822 78818 294004 79054
rect 293404 78734 294004 78818
rect 293404 78498 293586 78734
rect 293822 78498 294004 78734
rect 293404 43054 294004 78498
rect 293404 42818 293586 43054
rect 293822 42818 294004 43054
rect 293404 42734 294004 42818
rect 293404 42498 293586 42734
rect 293822 42498 294004 42734
rect 293404 7054 294004 42498
rect 293404 6818 293586 7054
rect 293822 6818 294004 7054
rect 293404 6734 294004 6818
rect 293404 6498 293586 6734
rect 293822 6498 294004 6734
rect 293404 -2226 294004 6498
rect 293404 -2462 293586 -2226
rect 293822 -2462 294004 -2226
rect 293404 -2546 294004 -2462
rect 293404 -2782 293586 -2546
rect 293822 -2782 294004 -2546
rect 293404 -3744 294004 -2782
rect 297004 334654 297604 336000
rect 297004 334418 297186 334654
rect 297422 334418 297604 334654
rect 297004 334334 297604 334418
rect 297004 334098 297186 334334
rect 297422 334098 297604 334334
rect 297004 298654 297604 334098
rect 297004 298418 297186 298654
rect 297422 298418 297604 298654
rect 297004 298334 297604 298418
rect 297004 298098 297186 298334
rect 297422 298098 297604 298334
rect 297004 262654 297604 298098
rect 297004 262418 297186 262654
rect 297422 262418 297604 262654
rect 297004 262334 297604 262418
rect 297004 262098 297186 262334
rect 297422 262098 297604 262334
rect 297004 226654 297604 262098
rect 297004 226418 297186 226654
rect 297422 226418 297604 226654
rect 297004 226334 297604 226418
rect 297004 226098 297186 226334
rect 297422 226098 297604 226334
rect 297004 190654 297604 226098
rect 297004 190418 297186 190654
rect 297422 190418 297604 190654
rect 297004 190334 297604 190418
rect 297004 190098 297186 190334
rect 297422 190098 297604 190334
rect 297004 154654 297604 190098
rect 297004 154418 297186 154654
rect 297422 154418 297604 154654
rect 297004 154334 297604 154418
rect 297004 154098 297186 154334
rect 297422 154098 297604 154334
rect 297004 118654 297604 154098
rect 297004 118418 297186 118654
rect 297422 118418 297604 118654
rect 297004 118334 297604 118418
rect 297004 118098 297186 118334
rect 297422 118098 297604 118334
rect 297004 82654 297604 118098
rect 297004 82418 297186 82654
rect 297422 82418 297604 82654
rect 297004 82334 297604 82418
rect 297004 82098 297186 82334
rect 297422 82098 297604 82334
rect 297004 46654 297604 82098
rect 297004 46418 297186 46654
rect 297422 46418 297604 46654
rect 297004 46334 297604 46418
rect 297004 46098 297186 46334
rect 297422 46098 297604 46334
rect 297004 10654 297604 46098
rect 297004 10418 297186 10654
rect 297422 10418 297604 10654
rect 297004 10334 297604 10418
rect 297004 10098 297186 10334
rect 297422 10098 297604 10334
rect 297004 -4106 297604 10098
rect 297004 -4342 297186 -4106
rect 297422 -4342 297604 -4106
rect 297004 -4426 297604 -4342
rect 297004 -4662 297186 -4426
rect 297422 -4662 297604 -4426
rect 297004 -5624 297604 -4662
rect 300604 302254 301204 336000
rect 300604 302018 300786 302254
rect 301022 302018 301204 302254
rect 300604 301934 301204 302018
rect 300604 301698 300786 301934
rect 301022 301698 301204 301934
rect 300604 266254 301204 301698
rect 300604 266018 300786 266254
rect 301022 266018 301204 266254
rect 300604 265934 301204 266018
rect 300604 265698 300786 265934
rect 301022 265698 301204 265934
rect 300604 230254 301204 265698
rect 300604 230018 300786 230254
rect 301022 230018 301204 230254
rect 300604 229934 301204 230018
rect 300604 229698 300786 229934
rect 301022 229698 301204 229934
rect 300604 194254 301204 229698
rect 300604 194018 300786 194254
rect 301022 194018 301204 194254
rect 300604 193934 301204 194018
rect 300604 193698 300786 193934
rect 301022 193698 301204 193934
rect 300604 158254 301204 193698
rect 300604 158018 300786 158254
rect 301022 158018 301204 158254
rect 300604 157934 301204 158018
rect 300604 157698 300786 157934
rect 301022 157698 301204 157934
rect 300604 122254 301204 157698
rect 300604 122018 300786 122254
rect 301022 122018 301204 122254
rect 300604 121934 301204 122018
rect 300604 121698 300786 121934
rect 301022 121698 301204 121934
rect 300604 86254 301204 121698
rect 300604 86018 300786 86254
rect 301022 86018 301204 86254
rect 300604 85934 301204 86018
rect 300604 85698 300786 85934
rect 301022 85698 301204 85934
rect 300604 50254 301204 85698
rect 300604 50018 300786 50254
rect 301022 50018 301204 50254
rect 300604 49934 301204 50018
rect 300604 49698 300786 49934
rect 301022 49698 301204 49934
rect 300604 14254 301204 49698
rect 306974 31789 307034 340851
rect 307804 309454 308404 344898
rect 307804 309218 307986 309454
rect 308222 309218 308404 309454
rect 307804 309134 308404 309218
rect 307804 308898 307986 309134
rect 308222 308898 308404 309134
rect 307804 273454 308404 308898
rect 307804 273218 307986 273454
rect 308222 273218 308404 273454
rect 307804 273134 308404 273218
rect 307804 272898 307986 273134
rect 308222 272898 308404 273134
rect 307804 237454 308404 272898
rect 307804 237218 307986 237454
rect 308222 237218 308404 237454
rect 307804 237134 308404 237218
rect 307804 236898 307986 237134
rect 308222 236898 308404 237134
rect 307804 201454 308404 236898
rect 307804 201218 307986 201454
rect 308222 201218 308404 201454
rect 307804 201134 308404 201218
rect 307804 200898 307986 201134
rect 308222 200898 308404 201134
rect 307804 165454 308404 200898
rect 307804 165218 307986 165454
rect 308222 165218 308404 165454
rect 307804 165134 308404 165218
rect 307804 164898 307986 165134
rect 308222 164898 308404 165134
rect 307804 129454 308404 164898
rect 307804 129218 307986 129454
rect 308222 129218 308404 129454
rect 307804 129134 308404 129218
rect 307804 128898 307986 129134
rect 308222 128898 308404 129134
rect 307804 93454 308404 128898
rect 307804 93218 307986 93454
rect 308222 93218 308404 93454
rect 307804 93134 308404 93218
rect 307804 92898 307986 93134
rect 308222 92898 308404 93134
rect 307804 57454 308404 92898
rect 307804 57218 307986 57454
rect 308222 57218 308404 57454
rect 307804 57134 308404 57218
rect 307804 56898 307986 57134
rect 308222 56898 308404 57134
rect 306971 31788 307037 31789
rect 306971 31724 306972 31788
rect 307036 31724 307037 31788
rect 306971 31723 307037 31724
rect 300604 14018 300786 14254
rect 301022 14018 301204 14254
rect 300604 13934 301204 14018
rect 300604 13698 300786 13934
rect 301022 13698 301204 13934
rect 282604 -7162 282786 -6926
rect 283022 -7162 283204 -6926
rect 282604 -7246 283204 -7162
rect 282604 -7482 282786 -7246
rect 283022 -7482 283204 -7246
rect 282604 -7504 283204 -7482
rect 300604 -5986 301204 13698
rect 307804 21454 308404 56898
rect 307804 21218 307986 21454
rect 308222 21218 308404 21454
rect 307804 21134 308404 21218
rect 307804 20898 307986 21134
rect 308222 20898 308404 21134
rect 307804 -1286 308404 20898
rect 307804 -1522 307986 -1286
rect 308222 -1522 308404 -1286
rect 307804 -1606 308404 -1522
rect 307804 -1842 307986 -1606
rect 308222 -1842 308404 -1606
rect 307804 -1864 308404 -1842
rect 311404 673054 312004 707102
rect 311404 672818 311586 673054
rect 311822 672818 312004 673054
rect 311404 672734 312004 672818
rect 311404 672498 311586 672734
rect 311822 672498 312004 672734
rect 311404 637054 312004 672498
rect 311404 636818 311586 637054
rect 311822 636818 312004 637054
rect 311404 636734 312004 636818
rect 311404 636498 311586 636734
rect 311822 636498 312004 636734
rect 311404 601054 312004 636498
rect 311404 600818 311586 601054
rect 311822 600818 312004 601054
rect 311404 600734 312004 600818
rect 311404 600498 311586 600734
rect 311822 600498 312004 600734
rect 311404 565054 312004 600498
rect 311404 564818 311586 565054
rect 311822 564818 312004 565054
rect 311404 564734 312004 564818
rect 311404 564498 311586 564734
rect 311822 564498 312004 564734
rect 311404 529054 312004 564498
rect 311404 528818 311586 529054
rect 311822 528818 312004 529054
rect 311404 528734 312004 528818
rect 311404 528498 311586 528734
rect 311822 528498 312004 528734
rect 311404 493054 312004 528498
rect 311404 492818 311586 493054
rect 311822 492818 312004 493054
rect 311404 492734 312004 492818
rect 311404 492498 311586 492734
rect 311822 492498 312004 492734
rect 311404 457054 312004 492498
rect 311404 456818 311586 457054
rect 311822 456818 312004 457054
rect 311404 456734 312004 456818
rect 311404 456498 311586 456734
rect 311822 456498 312004 456734
rect 311404 421054 312004 456498
rect 311404 420818 311586 421054
rect 311822 420818 312004 421054
rect 311404 420734 312004 420818
rect 311404 420498 311586 420734
rect 311822 420498 312004 420734
rect 311404 385054 312004 420498
rect 311404 384818 311586 385054
rect 311822 384818 312004 385054
rect 311404 384734 312004 384818
rect 311404 384498 311586 384734
rect 311822 384498 312004 384734
rect 311404 349054 312004 384498
rect 311404 348818 311586 349054
rect 311822 348818 312004 349054
rect 311404 348734 312004 348818
rect 311404 348498 311586 348734
rect 311822 348498 312004 348734
rect 311404 313054 312004 348498
rect 311404 312818 311586 313054
rect 311822 312818 312004 313054
rect 311404 312734 312004 312818
rect 311404 312498 311586 312734
rect 311822 312498 312004 312734
rect 311404 277054 312004 312498
rect 311404 276818 311586 277054
rect 311822 276818 312004 277054
rect 311404 276734 312004 276818
rect 311404 276498 311586 276734
rect 311822 276498 312004 276734
rect 311404 241054 312004 276498
rect 311404 240818 311586 241054
rect 311822 240818 312004 241054
rect 311404 240734 312004 240818
rect 311404 240498 311586 240734
rect 311822 240498 312004 240734
rect 311404 205054 312004 240498
rect 311404 204818 311586 205054
rect 311822 204818 312004 205054
rect 311404 204734 312004 204818
rect 311404 204498 311586 204734
rect 311822 204498 312004 204734
rect 311404 169054 312004 204498
rect 311404 168818 311586 169054
rect 311822 168818 312004 169054
rect 311404 168734 312004 168818
rect 311404 168498 311586 168734
rect 311822 168498 312004 168734
rect 311404 133054 312004 168498
rect 311404 132818 311586 133054
rect 311822 132818 312004 133054
rect 311404 132734 312004 132818
rect 311404 132498 311586 132734
rect 311822 132498 312004 132734
rect 311404 97054 312004 132498
rect 311404 96818 311586 97054
rect 311822 96818 312004 97054
rect 311404 96734 312004 96818
rect 311404 96498 311586 96734
rect 311822 96498 312004 96734
rect 311404 61054 312004 96498
rect 311404 60818 311586 61054
rect 311822 60818 312004 61054
rect 311404 60734 312004 60818
rect 311404 60498 311586 60734
rect 311822 60498 312004 60734
rect 311404 25054 312004 60498
rect 311404 24818 311586 25054
rect 311822 24818 312004 25054
rect 311404 24734 312004 24818
rect 311404 24498 311586 24734
rect 311822 24498 312004 24734
rect 311404 -3166 312004 24498
rect 311404 -3402 311586 -3166
rect 311822 -3402 312004 -3166
rect 311404 -3486 312004 -3402
rect 311404 -3722 311586 -3486
rect 311822 -3722 312004 -3486
rect 311404 -3744 312004 -3722
rect 315004 676654 315604 708982
rect 315004 676418 315186 676654
rect 315422 676418 315604 676654
rect 315004 676334 315604 676418
rect 315004 676098 315186 676334
rect 315422 676098 315604 676334
rect 315004 640654 315604 676098
rect 315004 640418 315186 640654
rect 315422 640418 315604 640654
rect 315004 640334 315604 640418
rect 315004 640098 315186 640334
rect 315422 640098 315604 640334
rect 315004 604654 315604 640098
rect 315004 604418 315186 604654
rect 315422 604418 315604 604654
rect 315004 604334 315604 604418
rect 315004 604098 315186 604334
rect 315422 604098 315604 604334
rect 315004 568654 315604 604098
rect 315004 568418 315186 568654
rect 315422 568418 315604 568654
rect 315004 568334 315604 568418
rect 315004 568098 315186 568334
rect 315422 568098 315604 568334
rect 315004 532654 315604 568098
rect 315004 532418 315186 532654
rect 315422 532418 315604 532654
rect 315004 532334 315604 532418
rect 315004 532098 315186 532334
rect 315422 532098 315604 532334
rect 315004 496654 315604 532098
rect 315004 496418 315186 496654
rect 315422 496418 315604 496654
rect 315004 496334 315604 496418
rect 315004 496098 315186 496334
rect 315422 496098 315604 496334
rect 315004 460654 315604 496098
rect 315004 460418 315186 460654
rect 315422 460418 315604 460654
rect 315004 460334 315604 460418
rect 315004 460098 315186 460334
rect 315422 460098 315604 460334
rect 315004 424654 315604 460098
rect 315004 424418 315186 424654
rect 315422 424418 315604 424654
rect 315004 424334 315604 424418
rect 315004 424098 315186 424334
rect 315422 424098 315604 424334
rect 315004 388654 315604 424098
rect 315004 388418 315186 388654
rect 315422 388418 315604 388654
rect 315004 388334 315604 388418
rect 315004 388098 315186 388334
rect 315422 388098 315604 388334
rect 315004 352654 315604 388098
rect 315004 352418 315186 352654
rect 315422 352418 315604 352654
rect 315004 352334 315604 352418
rect 315004 352098 315186 352334
rect 315422 352098 315604 352334
rect 315004 316654 315604 352098
rect 315004 316418 315186 316654
rect 315422 316418 315604 316654
rect 315004 316334 315604 316418
rect 315004 316098 315186 316334
rect 315422 316098 315604 316334
rect 315004 280654 315604 316098
rect 315004 280418 315186 280654
rect 315422 280418 315604 280654
rect 315004 280334 315604 280418
rect 315004 280098 315186 280334
rect 315422 280098 315604 280334
rect 315004 244654 315604 280098
rect 315004 244418 315186 244654
rect 315422 244418 315604 244654
rect 315004 244334 315604 244418
rect 315004 244098 315186 244334
rect 315422 244098 315604 244334
rect 315004 208654 315604 244098
rect 315004 208418 315186 208654
rect 315422 208418 315604 208654
rect 315004 208334 315604 208418
rect 315004 208098 315186 208334
rect 315422 208098 315604 208334
rect 315004 172654 315604 208098
rect 315004 172418 315186 172654
rect 315422 172418 315604 172654
rect 315004 172334 315604 172418
rect 315004 172098 315186 172334
rect 315422 172098 315604 172334
rect 315004 136654 315604 172098
rect 315004 136418 315186 136654
rect 315422 136418 315604 136654
rect 315004 136334 315604 136418
rect 315004 136098 315186 136334
rect 315422 136098 315604 136334
rect 315004 100654 315604 136098
rect 315004 100418 315186 100654
rect 315422 100418 315604 100654
rect 315004 100334 315604 100418
rect 315004 100098 315186 100334
rect 315422 100098 315604 100334
rect 315004 64654 315604 100098
rect 315004 64418 315186 64654
rect 315422 64418 315604 64654
rect 315004 64334 315604 64418
rect 315004 64098 315186 64334
rect 315422 64098 315604 64334
rect 315004 28654 315604 64098
rect 315004 28418 315186 28654
rect 315422 28418 315604 28654
rect 315004 28334 315604 28418
rect 315004 28098 315186 28334
rect 315422 28098 315604 28334
rect 315004 -5046 315604 28098
rect 315004 -5282 315186 -5046
rect 315422 -5282 315604 -5046
rect 315004 -5366 315604 -5282
rect 315004 -5602 315186 -5366
rect 315422 -5602 315604 -5366
rect 315004 -5624 315604 -5602
rect 318604 680254 319204 710862
rect 336604 710478 337204 711440
rect 336604 710242 336786 710478
rect 337022 710242 337204 710478
rect 336604 710158 337204 710242
rect 336604 709922 336786 710158
rect 337022 709922 337204 710158
rect 333004 708598 333604 709560
rect 333004 708362 333186 708598
rect 333422 708362 333604 708598
rect 333004 708278 333604 708362
rect 333004 708042 333186 708278
rect 333422 708042 333604 708278
rect 329404 706718 330004 707680
rect 329404 706482 329586 706718
rect 329822 706482 330004 706718
rect 329404 706398 330004 706482
rect 329404 706162 329586 706398
rect 329822 706162 330004 706398
rect 318604 680018 318786 680254
rect 319022 680018 319204 680254
rect 318604 679934 319204 680018
rect 318604 679698 318786 679934
rect 319022 679698 319204 679934
rect 318604 644254 319204 679698
rect 318604 644018 318786 644254
rect 319022 644018 319204 644254
rect 318604 643934 319204 644018
rect 318604 643698 318786 643934
rect 319022 643698 319204 643934
rect 318604 608254 319204 643698
rect 318604 608018 318786 608254
rect 319022 608018 319204 608254
rect 318604 607934 319204 608018
rect 318604 607698 318786 607934
rect 319022 607698 319204 607934
rect 318604 572254 319204 607698
rect 318604 572018 318786 572254
rect 319022 572018 319204 572254
rect 318604 571934 319204 572018
rect 318604 571698 318786 571934
rect 319022 571698 319204 571934
rect 318604 536254 319204 571698
rect 318604 536018 318786 536254
rect 319022 536018 319204 536254
rect 318604 535934 319204 536018
rect 318604 535698 318786 535934
rect 319022 535698 319204 535934
rect 318604 500254 319204 535698
rect 318604 500018 318786 500254
rect 319022 500018 319204 500254
rect 318604 499934 319204 500018
rect 318604 499698 318786 499934
rect 319022 499698 319204 499934
rect 318604 464254 319204 499698
rect 318604 464018 318786 464254
rect 319022 464018 319204 464254
rect 318604 463934 319204 464018
rect 318604 463698 318786 463934
rect 319022 463698 319204 463934
rect 318604 428254 319204 463698
rect 318604 428018 318786 428254
rect 319022 428018 319204 428254
rect 318604 427934 319204 428018
rect 318604 427698 318786 427934
rect 319022 427698 319204 427934
rect 318604 392254 319204 427698
rect 318604 392018 318786 392254
rect 319022 392018 319204 392254
rect 318604 391934 319204 392018
rect 318604 391698 318786 391934
rect 319022 391698 319204 391934
rect 318604 356254 319204 391698
rect 318604 356018 318786 356254
rect 319022 356018 319204 356254
rect 318604 355934 319204 356018
rect 318604 355698 318786 355934
rect 319022 355698 319204 355934
rect 318604 320254 319204 355698
rect 318604 320018 318786 320254
rect 319022 320018 319204 320254
rect 318604 319934 319204 320018
rect 318604 319698 318786 319934
rect 319022 319698 319204 319934
rect 318604 284254 319204 319698
rect 318604 284018 318786 284254
rect 319022 284018 319204 284254
rect 318604 283934 319204 284018
rect 318604 283698 318786 283934
rect 319022 283698 319204 283934
rect 318604 248254 319204 283698
rect 318604 248018 318786 248254
rect 319022 248018 319204 248254
rect 318604 247934 319204 248018
rect 318604 247698 318786 247934
rect 319022 247698 319204 247934
rect 318604 212254 319204 247698
rect 318604 212018 318786 212254
rect 319022 212018 319204 212254
rect 318604 211934 319204 212018
rect 318604 211698 318786 211934
rect 319022 211698 319204 211934
rect 318604 176254 319204 211698
rect 318604 176018 318786 176254
rect 319022 176018 319204 176254
rect 318604 175934 319204 176018
rect 318604 175698 318786 175934
rect 319022 175698 319204 175934
rect 318604 140254 319204 175698
rect 318604 140018 318786 140254
rect 319022 140018 319204 140254
rect 318604 139934 319204 140018
rect 318604 139698 318786 139934
rect 319022 139698 319204 139934
rect 318604 104254 319204 139698
rect 318604 104018 318786 104254
rect 319022 104018 319204 104254
rect 318604 103934 319204 104018
rect 318604 103698 318786 103934
rect 319022 103698 319204 103934
rect 318604 68254 319204 103698
rect 318604 68018 318786 68254
rect 319022 68018 319204 68254
rect 318604 67934 319204 68018
rect 318604 67698 318786 67934
rect 319022 67698 319204 67934
rect 318604 32254 319204 67698
rect 318604 32018 318786 32254
rect 319022 32018 319204 32254
rect 318604 31934 319204 32018
rect 318604 31698 318786 31934
rect 319022 31698 319204 31934
rect 300604 -6222 300786 -5986
rect 301022 -6222 301204 -5986
rect 300604 -6306 301204 -6222
rect 300604 -6542 300786 -6306
rect 301022 -6542 301204 -6306
rect 300604 -7504 301204 -6542
rect 318604 -6926 319204 31698
rect 325804 704838 326404 705800
rect 325804 704602 325986 704838
rect 326222 704602 326404 704838
rect 325804 704518 326404 704602
rect 325804 704282 325986 704518
rect 326222 704282 326404 704518
rect 325804 687454 326404 704282
rect 325804 687218 325986 687454
rect 326222 687218 326404 687454
rect 325804 687134 326404 687218
rect 325804 686898 325986 687134
rect 326222 686898 326404 687134
rect 325804 651454 326404 686898
rect 325804 651218 325986 651454
rect 326222 651218 326404 651454
rect 325804 651134 326404 651218
rect 325804 650898 325986 651134
rect 326222 650898 326404 651134
rect 325804 615454 326404 650898
rect 325804 615218 325986 615454
rect 326222 615218 326404 615454
rect 325804 615134 326404 615218
rect 325804 614898 325986 615134
rect 326222 614898 326404 615134
rect 325804 579454 326404 614898
rect 325804 579218 325986 579454
rect 326222 579218 326404 579454
rect 325804 579134 326404 579218
rect 325804 578898 325986 579134
rect 326222 578898 326404 579134
rect 325804 543454 326404 578898
rect 325804 543218 325986 543454
rect 326222 543218 326404 543454
rect 325804 543134 326404 543218
rect 325804 542898 325986 543134
rect 326222 542898 326404 543134
rect 325804 507454 326404 542898
rect 325804 507218 325986 507454
rect 326222 507218 326404 507454
rect 325804 507134 326404 507218
rect 325804 506898 325986 507134
rect 326222 506898 326404 507134
rect 325804 471454 326404 506898
rect 325804 471218 325986 471454
rect 326222 471218 326404 471454
rect 325804 471134 326404 471218
rect 325804 470898 325986 471134
rect 326222 470898 326404 471134
rect 325804 435454 326404 470898
rect 325804 435218 325986 435454
rect 326222 435218 326404 435454
rect 325804 435134 326404 435218
rect 325804 434898 325986 435134
rect 326222 434898 326404 435134
rect 325804 399454 326404 434898
rect 325804 399218 325986 399454
rect 326222 399218 326404 399454
rect 325804 399134 326404 399218
rect 325804 398898 325986 399134
rect 326222 398898 326404 399134
rect 325804 363454 326404 398898
rect 325804 363218 325986 363454
rect 326222 363218 326404 363454
rect 325804 363134 326404 363218
rect 325804 362898 325986 363134
rect 326222 362898 326404 363134
rect 325804 327454 326404 362898
rect 325804 327218 325986 327454
rect 326222 327218 326404 327454
rect 325804 327134 326404 327218
rect 325804 326898 325986 327134
rect 326222 326898 326404 327134
rect 325804 291454 326404 326898
rect 325804 291218 325986 291454
rect 326222 291218 326404 291454
rect 325804 291134 326404 291218
rect 325804 290898 325986 291134
rect 326222 290898 326404 291134
rect 325804 255454 326404 290898
rect 325804 255218 325986 255454
rect 326222 255218 326404 255454
rect 325804 255134 326404 255218
rect 325804 254898 325986 255134
rect 326222 254898 326404 255134
rect 325804 219454 326404 254898
rect 325804 219218 325986 219454
rect 326222 219218 326404 219454
rect 325804 219134 326404 219218
rect 325804 218898 325986 219134
rect 326222 218898 326404 219134
rect 325804 183454 326404 218898
rect 325804 183218 325986 183454
rect 326222 183218 326404 183454
rect 325804 183134 326404 183218
rect 325804 182898 325986 183134
rect 326222 182898 326404 183134
rect 325804 147454 326404 182898
rect 325804 147218 325986 147454
rect 326222 147218 326404 147454
rect 325804 147134 326404 147218
rect 325804 146898 325986 147134
rect 326222 146898 326404 147134
rect 325804 111454 326404 146898
rect 325804 111218 325986 111454
rect 326222 111218 326404 111454
rect 325804 111134 326404 111218
rect 325804 110898 325986 111134
rect 326222 110898 326404 111134
rect 325804 75454 326404 110898
rect 325804 75218 325986 75454
rect 326222 75218 326404 75454
rect 325804 75134 326404 75218
rect 325804 74898 325986 75134
rect 326222 74898 326404 75134
rect 325804 39454 326404 74898
rect 325804 39218 325986 39454
rect 326222 39218 326404 39454
rect 325804 39134 326404 39218
rect 325804 38898 325986 39134
rect 326222 38898 326404 39134
rect 325804 3454 326404 38898
rect 325804 3218 325986 3454
rect 326222 3218 326404 3454
rect 325804 3134 326404 3218
rect 325804 2898 325986 3134
rect 326222 2898 326404 3134
rect 325804 -346 326404 2898
rect 325804 -582 325986 -346
rect 326222 -582 326404 -346
rect 325804 -666 326404 -582
rect 325804 -902 325986 -666
rect 326222 -902 326404 -666
rect 325804 -1864 326404 -902
rect 329404 691054 330004 706162
rect 329404 690818 329586 691054
rect 329822 690818 330004 691054
rect 329404 690734 330004 690818
rect 329404 690498 329586 690734
rect 329822 690498 330004 690734
rect 329404 655054 330004 690498
rect 329404 654818 329586 655054
rect 329822 654818 330004 655054
rect 329404 654734 330004 654818
rect 329404 654498 329586 654734
rect 329822 654498 330004 654734
rect 329404 619054 330004 654498
rect 329404 618818 329586 619054
rect 329822 618818 330004 619054
rect 329404 618734 330004 618818
rect 329404 618498 329586 618734
rect 329822 618498 330004 618734
rect 329404 583054 330004 618498
rect 329404 582818 329586 583054
rect 329822 582818 330004 583054
rect 329404 582734 330004 582818
rect 329404 582498 329586 582734
rect 329822 582498 330004 582734
rect 329404 547054 330004 582498
rect 329404 546818 329586 547054
rect 329822 546818 330004 547054
rect 329404 546734 330004 546818
rect 329404 546498 329586 546734
rect 329822 546498 330004 546734
rect 329404 511054 330004 546498
rect 329404 510818 329586 511054
rect 329822 510818 330004 511054
rect 329404 510734 330004 510818
rect 329404 510498 329586 510734
rect 329822 510498 330004 510734
rect 329404 475054 330004 510498
rect 329404 474818 329586 475054
rect 329822 474818 330004 475054
rect 329404 474734 330004 474818
rect 329404 474498 329586 474734
rect 329822 474498 330004 474734
rect 329404 439054 330004 474498
rect 329404 438818 329586 439054
rect 329822 438818 330004 439054
rect 329404 438734 330004 438818
rect 329404 438498 329586 438734
rect 329822 438498 330004 438734
rect 329404 403054 330004 438498
rect 329404 402818 329586 403054
rect 329822 402818 330004 403054
rect 329404 402734 330004 402818
rect 329404 402498 329586 402734
rect 329822 402498 330004 402734
rect 329404 367054 330004 402498
rect 329404 366818 329586 367054
rect 329822 366818 330004 367054
rect 329404 366734 330004 366818
rect 329404 366498 329586 366734
rect 329822 366498 330004 366734
rect 329404 331054 330004 366498
rect 329404 330818 329586 331054
rect 329822 330818 330004 331054
rect 329404 330734 330004 330818
rect 329404 330498 329586 330734
rect 329822 330498 330004 330734
rect 329404 295054 330004 330498
rect 329404 294818 329586 295054
rect 329822 294818 330004 295054
rect 329404 294734 330004 294818
rect 329404 294498 329586 294734
rect 329822 294498 330004 294734
rect 329404 259054 330004 294498
rect 329404 258818 329586 259054
rect 329822 258818 330004 259054
rect 329404 258734 330004 258818
rect 329404 258498 329586 258734
rect 329822 258498 330004 258734
rect 329404 223054 330004 258498
rect 329404 222818 329586 223054
rect 329822 222818 330004 223054
rect 329404 222734 330004 222818
rect 329404 222498 329586 222734
rect 329822 222498 330004 222734
rect 329404 187054 330004 222498
rect 329404 186818 329586 187054
rect 329822 186818 330004 187054
rect 329404 186734 330004 186818
rect 329404 186498 329586 186734
rect 329822 186498 330004 186734
rect 329404 151054 330004 186498
rect 329404 150818 329586 151054
rect 329822 150818 330004 151054
rect 329404 150734 330004 150818
rect 329404 150498 329586 150734
rect 329822 150498 330004 150734
rect 329404 115054 330004 150498
rect 329404 114818 329586 115054
rect 329822 114818 330004 115054
rect 329404 114734 330004 114818
rect 329404 114498 329586 114734
rect 329822 114498 330004 114734
rect 329404 79054 330004 114498
rect 329404 78818 329586 79054
rect 329822 78818 330004 79054
rect 329404 78734 330004 78818
rect 329404 78498 329586 78734
rect 329822 78498 330004 78734
rect 329404 43054 330004 78498
rect 329404 42818 329586 43054
rect 329822 42818 330004 43054
rect 329404 42734 330004 42818
rect 329404 42498 329586 42734
rect 329822 42498 330004 42734
rect 329404 7054 330004 42498
rect 329404 6818 329586 7054
rect 329822 6818 330004 7054
rect 329404 6734 330004 6818
rect 329404 6498 329586 6734
rect 329822 6498 330004 6734
rect 329404 -2226 330004 6498
rect 329404 -2462 329586 -2226
rect 329822 -2462 330004 -2226
rect 329404 -2546 330004 -2462
rect 329404 -2782 329586 -2546
rect 329822 -2782 330004 -2546
rect 329404 -3744 330004 -2782
rect 333004 694654 333604 708042
rect 333004 694418 333186 694654
rect 333422 694418 333604 694654
rect 333004 694334 333604 694418
rect 333004 694098 333186 694334
rect 333422 694098 333604 694334
rect 333004 658654 333604 694098
rect 333004 658418 333186 658654
rect 333422 658418 333604 658654
rect 333004 658334 333604 658418
rect 333004 658098 333186 658334
rect 333422 658098 333604 658334
rect 333004 622654 333604 658098
rect 333004 622418 333186 622654
rect 333422 622418 333604 622654
rect 333004 622334 333604 622418
rect 333004 622098 333186 622334
rect 333422 622098 333604 622334
rect 333004 586654 333604 622098
rect 333004 586418 333186 586654
rect 333422 586418 333604 586654
rect 333004 586334 333604 586418
rect 333004 586098 333186 586334
rect 333422 586098 333604 586334
rect 333004 550654 333604 586098
rect 333004 550418 333186 550654
rect 333422 550418 333604 550654
rect 333004 550334 333604 550418
rect 333004 550098 333186 550334
rect 333422 550098 333604 550334
rect 333004 514654 333604 550098
rect 333004 514418 333186 514654
rect 333422 514418 333604 514654
rect 333004 514334 333604 514418
rect 333004 514098 333186 514334
rect 333422 514098 333604 514334
rect 333004 478654 333604 514098
rect 333004 478418 333186 478654
rect 333422 478418 333604 478654
rect 333004 478334 333604 478418
rect 333004 478098 333186 478334
rect 333422 478098 333604 478334
rect 333004 442654 333604 478098
rect 333004 442418 333186 442654
rect 333422 442418 333604 442654
rect 333004 442334 333604 442418
rect 333004 442098 333186 442334
rect 333422 442098 333604 442334
rect 333004 406654 333604 442098
rect 333004 406418 333186 406654
rect 333422 406418 333604 406654
rect 333004 406334 333604 406418
rect 333004 406098 333186 406334
rect 333422 406098 333604 406334
rect 333004 370654 333604 406098
rect 333004 370418 333186 370654
rect 333422 370418 333604 370654
rect 333004 370334 333604 370418
rect 333004 370098 333186 370334
rect 333422 370098 333604 370334
rect 333004 334654 333604 370098
rect 333004 334418 333186 334654
rect 333422 334418 333604 334654
rect 333004 334334 333604 334418
rect 333004 334098 333186 334334
rect 333422 334098 333604 334334
rect 333004 298654 333604 334098
rect 333004 298418 333186 298654
rect 333422 298418 333604 298654
rect 333004 298334 333604 298418
rect 333004 298098 333186 298334
rect 333422 298098 333604 298334
rect 333004 262654 333604 298098
rect 333004 262418 333186 262654
rect 333422 262418 333604 262654
rect 333004 262334 333604 262418
rect 333004 262098 333186 262334
rect 333422 262098 333604 262334
rect 333004 226654 333604 262098
rect 333004 226418 333186 226654
rect 333422 226418 333604 226654
rect 333004 226334 333604 226418
rect 333004 226098 333186 226334
rect 333422 226098 333604 226334
rect 333004 190654 333604 226098
rect 333004 190418 333186 190654
rect 333422 190418 333604 190654
rect 333004 190334 333604 190418
rect 333004 190098 333186 190334
rect 333422 190098 333604 190334
rect 333004 154654 333604 190098
rect 333004 154418 333186 154654
rect 333422 154418 333604 154654
rect 333004 154334 333604 154418
rect 333004 154098 333186 154334
rect 333422 154098 333604 154334
rect 333004 118654 333604 154098
rect 333004 118418 333186 118654
rect 333422 118418 333604 118654
rect 333004 118334 333604 118418
rect 333004 118098 333186 118334
rect 333422 118098 333604 118334
rect 333004 82654 333604 118098
rect 333004 82418 333186 82654
rect 333422 82418 333604 82654
rect 333004 82334 333604 82418
rect 333004 82098 333186 82334
rect 333422 82098 333604 82334
rect 333004 46654 333604 82098
rect 333004 46418 333186 46654
rect 333422 46418 333604 46654
rect 333004 46334 333604 46418
rect 333004 46098 333186 46334
rect 333422 46098 333604 46334
rect 333004 10654 333604 46098
rect 333004 10418 333186 10654
rect 333422 10418 333604 10654
rect 333004 10334 333604 10418
rect 333004 10098 333186 10334
rect 333422 10098 333604 10334
rect 333004 -4106 333604 10098
rect 333004 -4342 333186 -4106
rect 333422 -4342 333604 -4106
rect 333004 -4426 333604 -4342
rect 333004 -4662 333186 -4426
rect 333422 -4662 333604 -4426
rect 333004 -5624 333604 -4662
rect 336604 698254 337204 709922
rect 354604 711418 355204 711440
rect 354604 711182 354786 711418
rect 355022 711182 355204 711418
rect 354604 711098 355204 711182
rect 354604 710862 354786 711098
rect 355022 710862 355204 711098
rect 351004 709538 351604 709560
rect 351004 709302 351186 709538
rect 351422 709302 351604 709538
rect 351004 709218 351604 709302
rect 351004 708982 351186 709218
rect 351422 708982 351604 709218
rect 347404 707658 348004 707680
rect 347404 707422 347586 707658
rect 347822 707422 348004 707658
rect 347404 707338 348004 707422
rect 347404 707102 347586 707338
rect 347822 707102 348004 707338
rect 336604 698018 336786 698254
rect 337022 698018 337204 698254
rect 336604 697934 337204 698018
rect 336604 697698 336786 697934
rect 337022 697698 337204 697934
rect 336604 662254 337204 697698
rect 336604 662018 336786 662254
rect 337022 662018 337204 662254
rect 336604 661934 337204 662018
rect 336604 661698 336786 661934
rect 337022 661698 337204 661934
rect 336604 626254 337204 661698
rect 336604 626018 336786 626254
rect 337022 626018 337204 626254
rect 336604 625934 337204 626018
rect 336604 625698 336786 625934
rect 337022 625698 337204 625934
rect 336604 590254 337204 625698
rect 336604 590018 336786 590254
rect 337022 590018 337204 590254
rect 336604 589934 337204 590018
rect 336604 589698 336786 589934
rect 337022 589698 337204 589934
rect 336604 554254 337204 589698
rect 336604 554018 336786 554254
rect 337022 554018 337204 554254
rect 336604 553934 337204 554018
rect 336604 553698 336786 553934
rect 337022 553698 337204 553934
rect 336604 518254 337204 553698
rect 336604 518018 336786 518254
rect 337022 518018 337204 518254
rect 336604 517934 337204 518018
rect 336604 517698 336786 517934
rect 337022 517698 337204 517934
rect 336604 482254 337204 517698
rect 336604 482018 336786 482254
rect 337022 482018 337204 482254
rect 336604 481934 337204 482018
rect 336604 481698 336786 481934
rect 337022 481698 337204 481934
rect 336604 446254 337204 481698
rect 336604 446018 336786 446254
rect 337022 446018 337204 446254
rect 336604 445934 337204 446018
rect 336604 445698 336786 445934
rect 337022 445698 337204 445934
rect 336604 410254 337204 445698
rect 336604 410018 336786 410254
rect 337022 410018 337204 410254
rect 336604 409934 337204 410018
rect 336604 409698 336786 409934
rect 337022 409698 337204 409934
rect 336604 374254 337204 409698
rect 336604 374018 336786 374254
rect 337022 374018 337204 374254
rect 336604 373934 337204 374018
rect 336604 373698 336786 373934
rect 337022 373698 337204 373934
rect 336604 338254 337204 373698
rect 336604 338018 336786 338254
rect 337022 338018 337204 338254
rect 336604 337934 337204 338018
rect 336604 337698 336786 337934
rect 337022 337698 337204 337934
rect 336604 302254 337204 337698
rect 336604 302018 336786 302254
rect 337022 302018 337204 302254
rect 336604 301934 337204 302018
rect 336604 301698 336786 301934
rect 337022 301698 337204 301934
rect 336604 266254 337204 301698
rect 336604 266018 336786 266254
rect 337022 266018 337204 266254
rect 336604 265934 337204 266018
rect 336604 265698 336786 265934
rect 337022 265698 337204 265934
rect 336604 230254 337204 265698
rect 336604 230018 336786 230254
rect 337022 230018 337204 230254
rect 336604 229934 337204 230018
rect 336604 229698 336786 229934
rect 337022 229698 337204 229934
rect 336604 194254 337204 229698
rect 336604 194018 336786 194254
rect 337022 194018 337204 194254
rect 336604 193934 337204 194018
rect 336604 193698 336786 193934
rect 337022 193698 337204 193934
rect 336604 158254 337204 193698
rect 336604 158018 336786 158254
rect 337022 158018 337204 158254
rect 336604 157934 337204 158018
rect 336604 157698 336786 157934
rect 337022 157698 337204 157934
rect 336604 122254 337204 157698
rect 336604 122018 336786 122254
rect 337022 122018 337204 122254
rect 336604 121934 337204 122018
rect 336604 121698 336786 121934
rect 337022 121698 337204 121934
rect 336604 86254 337204 121698
rect 336604 86018 336786 86254
rect 337022 86018 337204 86254
rect 336604 85934 337204 86018
rect 336604 85698 336786 85934
rect 337022 85698 337204 85934
rect 336604 50254 337204 85698
rect 336604 50018 336786 50254
rect 337022 50018 337204 50254
rect 336604 49934 337204 50018
rect 336604 49698 336786 49934
rect 337022 49698 337204 49934
rect 336604 14254 337204 49698
rect 336604 14018 336786 14254
rect 337022 14018 337204 14254
rect 336604 13934 337204 14018
rect 336604 13698 336786 13934
rect 337022 13698 337204 13934
rect 318604 -7162 318786 -6926
rect 319022 -7162 319204 -6926
rect 318604 -7246 319204 -7162
rect 318604 -7482 318786 -7246
rect 319022 -7482 319204 -7246
rect 318604 -7504 319204 -7482
rect 336604 -5986 337204 13698
rect 343804 705778 344404 705800
rect 343804 705542 343986 705778
rect 344222 705542 344404 705778
rect 343804 705458 344404 705542
rect 343804 705222 343986 705458
rect 344222 705222 344404 705458
rect 343804 669454 344404 705222
rect 343804 669218 343986 669454
rect 344222 669218 344404 669454
rect 343804 669134 344404 669218
rect 343804 668898 343986 669134
rect 344222 668898 344404 669134
rect 343804 633454 344404 668898
rect 343804 633218 343986 633454
rect 344222 633218 344404 633454
rect 343804 633134 344404 633218
rect 343804 632898 343986 633134
rect 344222 632898 344404 633134
rect 343804 597454 344404 632898
rect 343804 597218 343986 597454
rect 344222 597218 344404 597454
rect 343804 597134 344404 597218
rect 343804 596898 343986 597134
rect 344222 596898 344404 597134
rect 343804 561454 344404 596898
rect 343804 561218 343986 561454
rect 344222 561218 344404 561454
rect 343804 561134 344404 561218
rect 343804 560898 343986 561134
rect 344222 560898 344404 561134
rect 343804 525454 344404 560898
rect 343804 525218 343986 525454
rect 344222 525218 344404 525454
rect 343804 525134 344404 525218
rect 343804 524898 343986 525134
rect 344222 524898 344404 525134
rect 343804 489454 344404 524898
rect 343804 489218 343986 489454
rect 344222 489218 344404 489454
rect 343804 489134 344404 489218
rect 343804 488898 343986 489134
rect 344222 488898 344404 489134
rect 343804 453454 344404 488898
rect 343804 453218 343986 453454
rect 344222 453218 344404 453454
rect 343804 453134 344404 453218
rect 343804 452898 343986 453134
rect 344222 452898 344404 453134
rect 343804 417454 344404 452898
rect 343804 417218 343986 417454
rect 344222 417218 344404 417454
rect 343804 417134 344404 417218
rect 343804 416898 343986 417134
rect 344222 416898 344404 417134
rect 343804 381454 344404 416898
rect 343804 381218 343986 381454
rect 344222 381218 344404 381454
rect 343804 381134 344404 381218
rect 343804 380898 343986 381134
rect 344222 380898 344404 381134
rect 343804 345454 344404 380898
rect 343804 345218 343986 345454
rect 344222 345218 344404 345454
rect 343804 345134 344404 345218
rect 343804 344898 343986 345134
rect 344222 344898 344404 345134
rect 343804 309454 344404 344898
rect 343804 309218 343986 309454
rect 344222 309218 344404 309454
rect 343804 309134 344404 309218
rect 343804 308898 343986 309134
rect 344222 308898 344404 309134
rect 343804 273454 344404 308898
rect 343804 273218 343986 273454
rect 344222 273218 344404 273454
rect 343804 273134 344404 273218
rect 343804 272898 343986 273134
rect 344222 272898 344404 273134
rect 343804 237454 344404 272898
rect 343804 237218 343986 237454
rect 344222 237218 344404 237454
rect 343804 237134 344404 237218
rect 343804 236898 343986 237134
rect 344222 236898 344404 237134
rect 343804 201454 344404 236898
rect 343804 201218 343986 201454
rect 344222 201218 344404 201454
rect 343804 201134 344404 201218
rect 343804 200898 343986 201134
rect 344222 200898 344404 201134
rect 343804 165454 344404 200898
rect 343804 165218 343986 165454
rect 344222 165218 344404 165454
rect 343804 165134 344404 165218
rect 343804 164898 343986 165134
rect 344222 164898 344404 165134
rect 343804 129454 344404 164898
rect 343804 129218 343986 129454
rect 344222 129218 344404 129454
rect 343804 129134 344404 129218
rect 343804 128898 343986 129134
rect 344222 128898 344404 129134
rect 343804 93454 344404 128898
rect 343804 93218 343986 93454
rect 344222 93218 344404 93454
rect 343804 93134 344404 93218
rect 343804 92898 343986 93134
rect 344222 92898 344404 93134
rect 343804 57454 344404 92898
rect 343804 57218 343986 57454
rect 344222 57218 344404 57454
rect 343804 57134 344404 57218
rect 343804 56898 343986 57134
rect 344222 56898 344404 57134
rect 343804 21454 344404 56898
rect 343804 21218 343986 21454
rect 344222 21218 344404 21454
rect 343804 21134 344404 21218
rect 343804 20898 343986 21134
rect 344222 20898 344404 21134
rect 343804 -1286 344404 20898
rect 343804 -1522 343986 -1286
rect 344222 -1522 344404 -1286
rect 343804 -1606 344404 -1522
rect 343804 -1842 343986 -1606
rect 344222 -1842 344404 -1606
rect 343804 -1864 344404 -1842
rect 347404 673054 348004 707102
rect 347404 672818 347586 673054
rect 347822 672818 348004 673054
rect 347404 672734 348004 672818
rect 347404 672498 347586 672734
rect 347822 672498 348004 672734
rect 347404 637054 348004 672498
rect 347404 636818 347586 637054
rect 347822 636818 348004 637054
rect 347404 636734 348004 636818
rect 347404 636498 347586 636734
rect 347822 636498 348004 636734
rect 347404 601054 348004 636498
rect 347404 600818 347586 601054
rect 347822 600818 348004 601054
rect 347404 600734 348004 600818
rect 347404 600498 347586 600734
rect 347822 600498 348004 600734
rect 347404 565054 348004 600498
rect 347404 564818 347586 565054
rect 347822 564818 348004 565054
rect 347404 564734 348004 564818
rect 347404 564498 347586 564734
rect 347822 564498 348004 564734
rect 347404 529054 348004 564498
rect 347404 528818 347586 529054
rect 347822 528818 348004 529054
rect 347404 528734 348004 528818
rect 347404 528498 347586 528734
rect 347822 528498 348004 528734
rect 347404 493054 348004 528498
rect 347404 492818 347586 493054
rect 347822 492818 348004 493054
rect 347404 492734 348004 492818
rect 347404 492498 347586 492734
rect 347822 492498 348004 492734
rect 347404 457054 348004 492498
rect 347404 456818 347586 457054
rect 347822 456818 348004 457054
rect 347404 456734 348004 456818
rect 347404 456498 347586 456734
rect 347822 456498 348004 456734
rect 347404 421054 348004 456498
rect 347404 420818 347586 421054
rect 347822 420818 348004 421054
rect 347404 420734 348004 420818
rect 347404 420498 347586 420734
rect 347822 420498 348004 420734
rect 347404 385054 348004 420498
rect 347404 384818 347586 385054
rect 347822 384818 348004 385054
rect 347404 384734 348004 384818
rect 347404 384498 347586 384734
rect 347822 384498 348004 384734
rect 347404 349054 348004 384498
rect 347404 348818 347586 349054
rect 347822 348818 348004 349054
rect 347404 348734 348004 348818
rect 347404 348498 347586 348734
rect 347822 348498 348004 348734
rect 347404 313054 348004 348498
rect 347404 312818 347586 313054
rect 347822 312818 348004 313054
rect 347404 312734 348004 312818
rect 347404 312498 347586 312734
rect 347822 312498 348004 312734
rect 347404 277054 348004 312498
rect 347404 276818 347586 277054
rect 347822 276818 348004 277054
rect 347404 276734 348004 276818
rect 347404 276498 347586 276734
rect 347822 276498 348004 276734
rect 347404 241054 348004 276498
rect 347404 240818 347586 241054
rect 347822 240818 348004 241054
rect 347404 240734 348004 240818
rect 347404 240498 347586 240734
rect 347822 240498 348004 240734
rect 347404 205054 348004 240498
rect 347404 204818 347586 205054
rect 347822 204818 348004 205054
rect 347404 204734 348004 204818
rect 347404 204498 347586 204734
rect 347822 204498 348004 204734
rect 347404 169054 348004 204498
rect 347404 168818 347586 169054
rect 347822 168818 348004 169054
rect 347404 168734 348004 168818
rect 347404 168498 347586 168734
rect 347822 168498 348004 168734
rect 347404 133054 348004 168498
rect 347404 132818 347586 133054
rect 347822 132818 348004 133054
rect 347404 132734 348004 132818
rect 347404 132498 347586 132734
rect 347822 132498 348004 132734
rect 347404 97054 348004 132498
rect 347404 96818 347586 97054
rect 347822 96818 348004 97054
rect 347404 96734 348004 96818
rect 347404 96498 347586 96734
rect 347822 96498 348004 96734
rect 347404 61054 348004 96498
rect 347404 60818 347586 61054
rect 347822 60818 348004 61054
rect 347404 60734 348004 60818
rect 347404 60498 347586 60734
rect 347822 60498 348004 60734
rect 347404 25054 348004 60498
rect 347404 24818 347586 25054
rect 347822 24818 348004 25054
rect 347404 24734 348004 24818
rect 347404 24498 347586 24734
rect 347822 24498 348004 24734
rect 347404 -3166 348004 24498
rect 347404 -3402 347586 -3166
rect 347822 -3402 348004 -3166
rect 347404 -3486 348004 -3402
rect 347404 -3722 347586 -3486
rect 347822 -3722 348004 -3486
rect 347404 -3744 348004 -3722
rect 351004 676654 351604 708982
rect 351004 676418 351186 676654
rect 351422 676418 351604 676654
rect 351004 676334 351604 676418
rect 351004 676098 351186 676334
rect 351422 676098 351604 676334
rect 351004 640654 351604 676098
rect 351004 640418 351186 640654
rect 351422 640418 351604 640654
rect 351004 640334 351604 640418
rect 351004 640098 351186 640334
rect 351422 640098 351604 640334
rect 351004 604654 351604 640098
rect 351004 604418 351186 604654
rect 351422 604418 351604 604654
rect 351004 604334 351604 604418
rect 351004 604098 351186 604334
rect 351422 604098 351604 604334
rect 351004 568654 351604 604098
rect 351004 568418 351186 568654
rect 351422 568418 351604 568654
rect 351004 568334 351604 568418
rect 351004 568098 351186 568334
rect 351422 568098 351604 568334
rect 351004 532654 351604 568098
rect 351004 532418 351186 532654
rect 351422 532418 351604 532654
rect 351004 532334 351604 532418
rect 351004 532098 351186 532334
rect 351422 532098 351604 532334
rect 351004 496654 351604 532098
rect 351004 496418 351186 496654
rect 351422 496418 351604 496654
rect 351004 496334 351604 496418
rect 351004 496098 351186 496334
rect 351422 496098 351604 496334
rect 351004 460654 351604 496098
rect 351004 460418 351186 460654
rect 351422 460418 351604 460654
rect 351004 460334 351604 460418
rect 351004 460098 351186 460334
rect 351422 460098 351604 460334
rect 351004 424654 351604 460098
rect 351004 424418 351186 424654
rect 351422 424418 351604 424654
rect 351004 424334 351604 424418
rect 351004 424098 351186 424334
rect 351422 424098 351604 424334
rect 351004 388654 351604 424098
rect 351004 388418 351186 388654
rect 351422 388418 351604 388654
rect 351004 388334 351604 388418
rect 351004 388098 351186 388334
rect 351422 388098 351604 388334
rect 351004 352654 351604 388098
rect 351004 352418 351186 352654
rect 351422 352418 351604 352654
rect 351004 352334 351604 352418
rect 351004 352098 351186 352334
rect 351422 352098 351604 352334
rect 351004 316654 351604 352098
rect 351004 316418 351186 316654
rect 351422 316418 351604 316654
rect 351004 316334 351604 316418
rect 351004 316098 351186 316334
rect 351422 316098 351604 316334
rect 351004 280654 351604 316098
rect 351004 280418 351186 280654
rect 351422 280418 351604 280654
rect 351004 280334 351604 280418
rect 351004 280098 351186 280334
rect 351422 280098 351604 280334
rect 351004 244654 351604 280098
rect 351004 244418 351186 244654
rect 351422 244418 351604 244654
rect 351004 244334 351604 244418
rect 351004 244098 351186 244334
rect 351422 244098 351604 244334
rect 351004 208654 351604 244098
rect 351004 208418 351186 208654
rect 351422 208418 351604 208654
rect 351004 208334 351604 208418
rect 351004 208098 351186 208334
rect 351422 208098 351604 208334
rect 351004 172654 351604 208098
rect 351004 172418 351186 172654
rect 351422 172418 351604 172654
rect 351004 172334 351604 172418
rect 351004 172098 351186 172334
rect 351422 172098 351604 172334
rect 351004 136654 351604 172098
rect 351004 136418 351186 136654
rect 351422 136418 351604 136654
rect 351004 136334 351604 136418
rect 351004 136098 351186 136334
rect 351422 136098 351604 136334
rect 351004 100654 351604 136098
rect 351004 100418 351186 100654
rect 351422 100418 351604 100654
rect 351004 100334 351604 100418
rect 351004 100098 351186 100334
rect 351422 100098 351604 100334
rect 351004 64654 351604 100098
rect 351004 64418 351186 64654
rect 351422 64418 351604 64654
rect 351004 64334 351604 64418
rect 351004 64098 351186 64334
rect 351422 64098 351604 64334
rect 351004 28654 351604 64098
rect 351004 28418 351186 28654
rect 351422 28418 351604 28654
rect 351004 28334 351604 28418
rect 351004 28098 351186 28334
rect 351422 28098 351604 28334
rect 351004 -5046 351604 28098
rect 351004 -5282 351186 -5046
rect 351422 -5282 351604 -5046
rect 351004 -5366 351604 -5282
rect 351004 -5602 351186 -5366
rect 351422 -5602 351604 -5366
rect 351004 -5624 351604 -5602
rect 354604 680254 355204 710862
rect 372604 710478 373204 711440
rect 372604 710242 372786 710478
rect 373022 710242 373204 710478
rect 372604 710158 373204 710242
rect 372604 709922 372786 710158
rect 373022 709922 373204 710158
rect 369004 708598 369604 709560
rect 369004 708362 369186 708598
rect 369422 708362 369604 708598
rect 369004 708278 369604 708362
rect 369004 708042 369186 708278
rect 369422 708042 369604 708278
rect 365404 706718 366004 707680
rect 365404 706482 365586 706718
rect 365822 706482 366004 706718
rect 365404 706398 366004 706482
rect 365404 706162 365586 706398
rect 365822 706162 366004 706398
rect 354604 680018 354786 680254
rect 355022 680018 355204 680254
rect 354604 679934 355204 680018
rect 354604 679698 354786 679934
rect 355022 679698 355204 679934
rect 354604 644254 355204 679698
rect 354604 644018 354786 644254
rect 355022 644018 355204 644254
rect 354604 643934 355204 644018
rect 354604 643698 354786 643934
rect 355022 643698 355204 643934
rect 354604 608254 355204 643698
rect 354604 608018 354786 608254
rect 355022 608018 355204 608254
rect 354604 607934 355204 608018
rect 354604 607698 354786 607934
rect 355022 607698 355204 607934
rect 354604 572254 355204 607698
rect 354604 572018 354786 572254
rect 355022 572018 355204 572254
rect 354604 571934 355204 572018
rect 354604 571698 354786 571934
rect 355022 571698 355204 571934
rect 354604 536254 355204 571698
rect 354604 536018 354786 536254
rect 355022 536018 355204 536254
rect 354604 535934 355204 536018
rect 354604 535698 354786 535934
rect 355022 535698 355204 535934
rect 354604 500254 355204 535698
rect 354604 500018 354786 500254
rect 355022 500018 355204 500254
rect 354604 499934 355204 500018
rect 354604 499698 354786 499934
rect 355022 499698 355204 499934
rect 354604 464254 355204 499698
rect 354604 464018 354786 464254
rect 355022 464018 355204 464254
rect 354604 463934 355204 464018
rect 354604 463698 354786 463934
rect 355022 463698 355204 463934
rect 354604 428254 355204 463698
rect 354604 428018 354786 428254
rect 355022 428018 355204 428254
rect 354604 427934 355204 428018
rect 354604 427698 354786 427934
rect 355022 427698 355204 427934
rect 354604 392254 355204 427698
rect 354604 392018 354786 392254
rect 355022 392018 355204 392254
rect 354604 391934 355204 392018
rect 354604 391698 354786 391934
rect 355022 391698 355204 391934
rect 354604 356254 355204 391698
rect 354604 356018 354786 356254
rect 355022 356018 355204 356254
rect 354604 355934 355204 356018
rect 354604 355698 354786 355934
rect 355022 355698 355204 355934
rect 354604 320254 355204 355698
rect 354604 320018 354786 320254
rect 355022 320018 355204 320254
rect 354604 319934 355204 320018
rect 354604 319698 354786 319934
rect 355022 319698 355204 319934
rect 354604 284254 355204 319698
rect 354604 284018 354786 284254
rect 355022 284018 355204 284254
rect 354604 283934 355204 284018
rect 354604 283698 354786 283934
rect 355022 283698 355204 283934
rect 354604 248254 355204 283698
rect 354604 248018 354786 248254
rect 355022 248018 355204 248254
rect 354604 247934 355204 248018
rect 354604 247698 354786 247934
rect 355022 247698 355204 247934
rect 354604 212254 355204 247698
rect 354604 212018 354786 212254
rect 355022 212018 355204 212254
rect 354604 211934 355204 212018
rect 354604 211698 354786 211934
rect 355022 211698 355204 211934
rect 354604 176254 355204 211698
rect 354604 176018 354786 176254
rect 355022 176018 355204 176254
rect 354604 175934 355204 176018
rect 354604 175698 354786 175934
rect 355022 175698 355204 175934
rect 354604 140254 355204 175698
rect 354604 140018 354786 140254
rect 355022 140018 355204 140254
rect 354604 139934 355204 140018
rect 354604 139698 354786 139934
rect 355022 139698 355204 139934
rect 354604 104254 355204 139698
rect 354604 104018 354786 104254
rect 355022 104018 355204 104254
rect 354604 103934 355204 104018
rect 354604 103698 354786 103934
rect 355022 103698 355204 103934
rect 354604 68254 355204 103698
rect 354604 68018 354786 68254
rect 355022 68018 355204 68254
rect 354604 67934 355204 68018
rect 354604 67698 354786 67934
rect 355022 67698 355204 67934
rect 354604 32254 355204 67698
rect 354604 32018 354786 32254
rect 355022 32018 355204 32254
rect 354604 31934 355204 32018
rect 354604 31698 354786 31934
rect 355022 31698 355204 31934
rect 336604 -6222 336786 -5986
rect 337022 -6222 337204 -5986
rect 336604 -6306 337204 -6222
rect 336604 -6542 336786 -6306
rect 337022 -6542 337204 -6306
rect 336604 -7504 337204 -6542
rect 354604 -6926 355204 31698
rect 361804 704838 362404 705800
rect 361804 704602 361986 704838
rect 362222 704602 362404 704838
rect 361804 704518 362404 704602
rect 361804 704282 361986 704518
rect 362222 704282 362404 704518
rect 361804 687454 362404 704282
rect 361804 687218 361986 687454
rect 362222 687218 362404 687454
rect 361804 687134 362404 687218
rect 361804 686898 361986 687134
rect 362222 686898 362404 687134
rect 361804 651454 362404 686898
rect 361804 651218 361986 651454
rect 362222 651218 362404 651454
rect 361804 651134 362404 651218
rect 361804 650898 361986 651134
rect 362222 650898 362404 651134
rect 361804 615454 362404 650898
rect 361804 615218 361986 615454
rect 362222 615218 362404 615454
rect 361804 615134 362404 615218
rect 361804 614898 361986 615134
rect 362222 614898 362404 615134
rect 361804 579454 362404 614898
rect 361804 579218 361986 579454
rect 362222 579218 362404 579454
rect 361804 579134 362404 579218
rect 361804 578898 361986 579134
rect 362222 578898 362404 579134
rect 361804 543454 362404 578898
rect 361804 543218 361986 543454
rect 362222 543218 362404 543454
rect 361804 543134 362404 543218
rect 361804 542898 361986 543134
rect 362222 542898 362404 543134
rect 361804 507454 362404 542898
rect 361804 507218 361986 507454
rect 362222 507218 362404 507454
rect 361804 507134 362404 507218
rect 361804 506898 361986 507134
rect 362222 506898 362404 507134
rect 361804 471454 362404 506898
rect 361804 471218 361986 471454
rect 362222 471218 362404 471454
rect 361804 471134 362404 471218
rect 361804 470898 361986 471134
rect 362222 470898 362404 471134
rect 361804 435454 362404 470898
rect 361804 435218 361986 435454
rect 362222 435218 362404 435454
rect 361804 435134 362404 435218
rect 361804 434898 361986 435134
rect 362222 434898 362404 435134
rect 361804 399454 362404 434898
rect 361804 399218 361986 399454
rect 362222 399218 362404 399454
rect 361804 399134 362404 399218
rect 361804 398898 361986 399134
rect 362222 398898 362404 399134
rect 361804 363454 362404 398898
rect 361804 363218 361986 363454
rect 362222 363218 362404 363454
rect 361804 363134 362404 363218
rect 361804 362898 361986 363134
rect 362222 362898 362404 363134
rect 361804 327454 362404 362898
rect 361804 327218 361986 327454
rect 362222 327218 362404 327454
rect 361804 327134 362404 327218
rect 361804 326898 361986 327134
rect 362222 326898 362404 327134
rect 361804 291454 362404 326898
rect 361804 291218 361986 291454
rect 362222 291218 362404 291454
rect 361804 291134 362404 291218
rect 361804 290898 361986 291134
rect 362222 290898 362404 291134
rect 361804 255454 362404 290898
rect 361804 255218 361986 255454
rect 362222 255218 362404 255454
rect 361804 255134 362404 255218
rect 361804 254898 361986 255134
rect 362222 254898 362404 255134
rect 361804 219454 362404 254898
rect 361804 219218 361986 219454
rect 362222 219218 362404 219454
rect 361804 219134 362404 219218
rect 361804 218898 361986 219134
rect 362222 218898 362404 219134
rect 361804 183454 362404 218898
rect 361804 183218 361986 183454
rect 362222 183218 362404 183454
rect 361804 183134 362404 183218
rect 361804 182898 361986 183134
rect 362222 182898 362404 183134
rect 361804 147454 362404 182898
rect 361804 147218 361986 147454
rect 362222 147218 362404 147454
rect 361804 147134 362404 147218
rect 361804 146898 361986 147134
rect 362222 146898 362404 147134
rect 361804 111454 362404 146898
rect 361804 111218 361986 111454
rect 362222 111218 362404 111454
rect 361804 111134 362404 111218
rect 361804 110898 361986 111134
rect 362222 110898 362404 111134
rect 361804 75454 362404 110898
rect 361804 75218 361986 75454
rect 362222 75218 362404 75454
rect 361804 75134 362404 75218
rect 361804 74898 361986 75134
rect 362222 74898 362404 75134
rect 361804 39454 362404 74898
rect 361804 39218 361986 39454
rect 362222 39218 362404 39454
rect 361804 39134 362404 39218
rect 361804 38898 361986 39134
rect 362222 38898 362404 39134
rect 361804 3454 362404 38898
rect 361804 3218 361986 3454
rect 362222 3218 362404 3454
rect 361804 3134 362404 3218
rect 361804 2898 361986 3134
rect 362222 2898 362404 3134
rect 361804 -346 362404 2898
rect 361804 -582 361986 -346
rect 362222 -582 362404 -346
rect 361804 -666 362404 -582
rect 361804 -902 361986 -666
rect 362222 -902 362404 -666
rect 361804 -1864 362404 -902
rect 365404 691054 366004 706162
rect 365404 690818 365586 691054
rect 365822 690818 366004 691054
rect 365404 690734 366004 690818
rect 365404 690498 365586 690734
rect 365822 690498 366004 690734
rect 365404 655054 366004 690498
rect 365404 654818 365586 655054
rect 365822 654818 366004 655054
rect 365404 654734 366004 654818
rect 365404 654498 365586 654734
rect 365822 654498 366004 654734
rect 365404 619054 366004 654498
rect 365404 618818 365586 619054
rect 365822 618818 366004 619054
rect 365404 618734 366004 618818
rect 365404 618498 365586 618734
rect 365822 618498 366004 618734
rect 365404 583054 366004 618498
rect 365404 582818 365586 583054
rect 365822 582818 366004 583054
rect 365404 582734 366004 582818
rect 365404 582498 365586 582734
rect 365822 582498 366004 582734
rect 365404 547054 366004 582498
rect 365404 546818 365586 547054
rect 365822 546818 366004 547054
rect 365404 546734 366004 546818
rect 365404 546498 365586 546734
rect 365822 546498 366004 546734
rect 365404 511054 366004 546498
rect 365404 510818 365586 511054
rect 365822 510818 366004 511054
rect 365404 510734 366004 510818
rect 365404 510498 365586 510734
rect 365822 510498 366004 510734
rect 365404 475054 366004 510498
rect 365404 474818 365586 475054
rect 365822 474818 366004 475054
rect 365404 474734 366004 474818
rect 365404 474498 365586 474734
rect 365822 474498 366004 474734
rect 365404 439054 366004 474498
rect 365404 438818 365586 439054
rect 365822 438818 366004 439054
rect 365404 438734 366004 438818
rect 365404 438498 365586 438734
rect 365822 438498 366004 438734
rect 365404 403054 366004 438498
rect 365404 402818 365586 403054
rect 365822 402818 366004 403054
rect 365404 402734 366004 402818
rect 365404 402498 365586 402734
rect 365822 402498 366004 402734
rect 365404 367054 366004 402498
rect 365404 366818 365586 367054
rect 365822 366818 366004 367054
rect 365404 366734 366004 366818
rect 365404 366498 365586 366734
rect 365822 366498 366004 366734
rect 365404 331054 366004 366498
rect 365404 330818 365586 331054
rect 365822 330818 366004 331054
rect 365404 330734 366004 330818
rect 365404 330498 365586 330734
rect 365822 330498 366004 330734
rect 365404 295054 366004 330498
rect 365404 294818 365586 295054
rect 365822 294818 366004 295054
rect 365404 294734 366004 294818
rect 365404 294498 365586 294734
rect 365822 294498 366004 294734
rect 365404 259054 366004 294498
rect 365404 258818 365586 259054
rect 365822 258818 366004 259054
rect 365404 258734 366004 258818
rect 365404 258498 365586 258734
rect 365822 258498 366004 258734
rect 365404 223054 366004 258498
rect 365404 222818 365586 223054
rect 365822 222818 366004 223054
rect 365404 222734 366004 222818
rect 365404 222498 365586 222734
rect 365822 222498 366004 222734
rect 365404 187054 366004 222498
rect 365404 186818 365586 187054
rect 365822 186818 366004 187054
rect 365404 186734 366004 186818
rect 365404 186498 365586 186734
rect 365822 186498 366004 186734
rect 365404 151054 366004 186498
rect 365404 150818 365586 151054
rect 365822 150818 366004 151054
rect 365404 150734 366004 150818
rect 365404 150498 365586 150734
rect 365822 150498 366004 150734
rect 365404 115054 366004 150498
rect 365404 114818 365586 115054
rect 365822 114818 366004 115054
rect 365404 114734 366004 114818
rect 365404 114498 365586 114734
rect 365822 114498 366004 114734
rect 365404 79054 366004 114498
rect 365404 78818 365586 79054
rect 365822 78818 366004 79054
rect 365404 78734 366004 78818
rect 365404 78498 365586 78734
rect 365822 78498 366004 78734
rect 365404 43054 366004 78498
rect 365404 42818 365586 43054
rect 365822 42818 366004 43054
rect 365404 42734 366004 42818
rect 365404 42498 365586 42734
rect 365822 42498 366004 42734
rect 365404 7054 366004 42498
rect 365404 6818 365586 7054
rect 365822 6818 366004 7054
rect 365404 6734 366004 6818
rect 365404 6498 365586 6734
rect 365822 6498 366004 6734
rect 365404 -2226 366004 6498
rect 365404 -2462 365586 -2226
rect 365822 -2462 366004 -2226
rect 365404 -2546 366004 -2462
rect 365404 -2782 365586 -2546
rect 365822 -2782 366004 -2546
rect 365404 -3744 366004 -2782
rect 369004 694654 369604 708042
rect 369004 694418 369186 694654
rect 369422 694418 369604 694654
rect 369004 694334 369604 694418
rect 369004 694098 369186 694334
rect 369422 694098 369604 694334
rect 369004 658654 369604 694098
rect 369004 658418 369186 658654
rect 369422 658418 369604 658654
rect 369004 658334 369604 658418
rect 369004 658098 369186 658334
rect 369422 658098 369604 658334
rect 369004 622654 369604 658098
rect 369004 622418 369186 622654
rect 369422 622418 369604 622654
rect 369004 622334 369604 622418
rect 369004 622098 369186 622334
rect 369422 622098 369604 622334
rect 369004 586654 369604 622098
rect 369004 586418 369186 586654
rect 369422 586418 369604 586654
rect 369004 586334 369604 586418
rect 369004 586098 369186 586334
rect 369422 586098 369604 586334
rect 369004 550654 369604 586098
rect 369004 550418 369186 550654
rect 369422 550418 369604 550654
rect 369004 550334 369604 550418
rect 369004 550098 369186 550334
rect 369422 550098 369604 550334
rect 369004 514654 369604 550098
rect 369004 514418 369186 514654
rect 369422 514418 369604 514654
rect 369004 514334 369604 514418
rect 369004 514098 369186 514334
rect 369422 514098 369604 514334
rect 369004 478654 369604 514098
rect 369004 478418 369186 478654
rect 369422 478418 369604 478654
rect 369004 478334 369604 478418
rect 369004 478098 369186 478334
rect 369422 478098 369604 478334
rect 369004 442654 369604 478098
rect 369004 442418 369186 442654
rect 369422 442418 369604 442654
rect 369004 442334 369604 442418
rect 369004 442098 369186 442334
rect 369422 442098 369604 442334
rect 369004 406654 369604 442098
rect 369004 406418 369186 406654
rect 369422 406418 369604 406654
rect 369004 406334 369604 406418
rect 369004 406098 369186 406334
rect 369422 406098 369604 406334
rect 369004 370654 369604 406098
rect 369004 370418 369186 370654
rect 369422 370418 369604 370654
rect 369004 370334 369604 370418
rect 369004 370098 369186 370334
rect 369422 370098 369604 370334
rect 369004 334654 369604 370098
rect 369004 334418 369186 334654
rect 369422 334418 369604 334654
rect 369004 334334 369604 334418
rect 369004 334098 369186 334334
rect 369422 334098 369604 334334
rect 369004 298654 369604 334098
rect 369004 298418 369186 298654
rect 369422 298418 369604 298654
rect 369004 298334 369604 298418
rect 369004 298098 369186 298334
rect 369422 298098 369604 298334
rect 369004 262654 369604 298098
rect 369004 262418 369186 262654
rect 369422 262418 369604 262654
rect 369004 262334 369604 262418
rect 369004 262098 369186 262334
rect 369422 262098 369604 262334
rect 369004 226654 369604 262098
rect 369004 226418 369186 226654
rect 369422 226418 369604 226654
rect 369004 226334 369604 226418
rect 369004 226098 369186 226334
rect 369422 226098 369604 226334
rect 369004 190654 369604 226098
rect 369004 190418 369186 190654
rect 369422 190418 369604 190654
rect 369004 190334 369604 190418
rect 369004 190098 369186 190334
rect 369422 190098 369604 190334
rect 369004 154654 369604 190098
rect 369004 154418 369186 154654
rect 369422 154418 369604 154654
rect 369004 154334 369604 154418
rect 369004 154098 369186 154334
rect 369422 154098 369604 154334
rect 369004 118654 369604 154098
rect 369004 118418 369186 118654
rect 369422 118418 369604 118654
rect 369004 118334 369604 118418
rect 369004 118098 369186 118334
rect 369422 118098 369604 118334
rect 369004 82654 369604 118098
rect 369004 82418 369186 82654
rect 369422 82418 369604 82654
rect 369004 82334 369604 82418
rect 369004 82098 369186 82334
rect 369422 82098 369604 82334
rect 369004 46654 369604 82098
rect 369004 46418 369186 46654
rect 369422 46418 369604 46654
rect 369004 46334 369604 46418
rect 369004 46098 369186 46334
rect 369422 46098 369604 46334
rect 369004 10654 369604 46098
rect 369004 10418 369186 10654
rect 369422 10418 369604 10654
rect 369004 10334 369604 10418
rect 369004 10098 369186 10334
rect 369422 10098 369604 10334
rect 369004 -4106 369604 10098
rect 369004 -4342 369186 -4106
rect 369422 -4342 369604 -4106
rect 369004 -4426 369604 -4342
rect 369004 -4662 369186 -4426
rect 369422 -4662 369604 -4426
rect 369004 -5624 369604 -4662
rect 372604 698254 373204 709922
rect 390604 711418 391204 711440
rect 390604 711182 390786 711418
rect 391022 711182 391204 711418
rect 390604 711098 391204 711182
rect 390604 710862 390786 711098
rect 391022 710862 391204 711098
rect 387004 709538 387604 709560
rect 387004 709302 387186 709538
rect 387422 709302 387604 709538
rect 387004 709218 387604 709302
rect 387004 708982 387186 709218
rect 387422 708982 387604 709218
rect 383404 707658 384004 707680
rect 383404 707422 383586 707658
rect 383822 707422 384004 707658
rect 383404 707338 384004 707422
rect 383404 707102 383586 707338
rect 383822 707102 384004 707338
rect 372604 698018 372786 698254
rect 373022 698018 373204 698254
rect 372604 697934 373204 698018
rect 372604 697698 372786 697934
rect 373022 697698 373204 697934
rect 372604 662254 373204 697698
rect 372604 662018 372786 662254
rect 373022 662018 373204 662254
rect 372604 661934 373204 662018
rect 372604 661698 372786 661934
rect 373022 661698 373204 661934
rect 372604 626254 373204 661698
rect 372604 626018 372786 626254
rect 373022 626018 373204 626254
rect 372604 625934 373204 626018
rect 372604 625698 372786 625934
rect 373022 625698 373204 625934
rect 372604 590254 373204 625698
rect 372604 590018 372786 590254
rect 373022 590018 373204 590254
rect 372604 589934 373204 590018
rect 372604 589698 372786 589934
rect 373022 589698 373204 589934
rect 372604 554254 373204 589698
rect 372604 554018 372786 554254
rect 373022 554018 373204 554254
rect 372604 553934 373204 554018
rect 372604 553698 372786 553934
rect 373022 553698 373204 553934
rect 372604 518254 373204 553698
rect 372604 518018 372786 518254
rect 373022 518018 373204 518254
rect 372604 517934 373204 518018
rect 372604 517698 372786 517934
rect 373022 517698 373204 517934
rect 372604 482254 373204 517698
rect 372604 482018 372786 482254
rect 373022 482018 373204 482254
rect 372604 481934 373204 482018
rect 372604 481698 372786 481934
rect 373022 481698 373204 481934
rect 372604 446254 373204 481698
rect 372604 446018 372786 446254
rect 373022 446018 373204 446254
rect 372604 445934 373204 446018
rect 372604 445698 372786 445934
rect 373022 445698 373204 445934
rect 372604 410254 373204 445698
rect 372604 410018 372786 410254
rect 373022 410018 373204 410254
rect 372604 409934 373204 410018
rect 372604 409698 372786 409934
rect 373022 409698 373204 409934
rect 372604 374254 373204 409698
rect 372604 374018 372786 374254
rect 373022 374018 373204 374254
rect 372604 373934 373204 374018
rect 372604 373698 372786 373934
rect 373022 373698 373204 373934
rect 372604 338254 373204 373698
rect 372604 338018 372786 338254
rect 373022 338018 373204 338254
rect 372604 337934 373204 338018
rect 372604 337698 372786 337934
rect 373022 337698 373204 337934
rect 372604 302254 373204 337698
rect 372604 302018 372786 302254
rect 373022 302018 373204 302254
rect 372604 301934 373204 302018
rect 372604 301698 372786 301934
rect 373022 301698 373204 301934
rect 372604 266254 373204 301698
rect 372604 266018 372786 266254
rect 373022 266018 373204 266254
rect 372604 265934 373204 266018
rect 372604 265698 372786 265934
rect 373022 265698 373204 265934
rect 372604 230254 373204 265698
rect 372604 230018 372786 230254
rect 373022 230018 373204 230254
rect 372604 229934 373204 230018
rect 372604 229698 372786 229934
rect 373022 229698 373204 229934
rect 372604 194254 373204 229698
rect 372604 194018 372786 194254
rect 373022 194018 373204 194254
rect 372604 193934 373204 194018
rect 372604 193698 372786 193934
rect 373022 193698 373204 193934
rect 372604 158254 373204 193698
rect 372604 158018 372786 158254
rect 373022 158018 373204 158254
rect 372604 157934 373204 158018
rect 372604 157698 372786 157934
rect 373022 157698 373204 157934
rect 372604 122254 373204 157698
rect 372604 122018 372786 122254
rect 373022 122018 373204 122254
rect 372604 121934 373204 122018
rect 372604 121698 372786 121934
rect 373022 121698 373204 121934
rect 372604 86254 373204 121698
rect 372604 86018 372786 86254
rect 373022 86018 373204 86254
rect 372604 85934 373204 86018
rect 372604 85698 372786 85934
rect 373022 85698 373204 85934
rect 372604 50254 373204 85698
rect 372604 50018 372786 50254
rect 373022 50018 373204 50254
rect 372604 49934 373204 50018
rect 372604 49698 372786 49934
rect 373022 49698 373204 49934
rect 372604 14254 373204 49698
rect 372604 14018 372786 14254
rect 373022 14018 373204 14254
rect 372604 13934 373204 14018
rect 372604 13698 372786 13934
rect 373022 13698 373204 13934
rect 354604 -7162 354786 -6926
rect 355022 -7162 355204 -6926
rect 354604 -7246 355204 -7162
rect 354604 -7482 354786 -7246
rect 355022 -7482 355204 -7246
rect 354604 -7504 355204 -7482
rect 372604 -5986 373204 13698
rect 379804 705778 380404 705800
rect 379804 705542 379986 705778
rect 380222 705542 380404 705778
rect 379804 705458 380404 705542
rect 379804 705222 379986 705458
rect 380222 705222 380404 705458
rect 379804 669454 380404 705222
rect 379804 669218 379986 669454
rect 380222 669218 380404 669454
rect 379804 669134 380404 669218
rect 379804 668898 379986 669134
rect 380222 668898 380404 669134
rect 379804 633454 380404 668898
rect 379804 633218 379986 633454
rect 380222 633218 380404 633454
rect 379804 633134 380404 633218
rect 379804 632898 379986 633134
rect 380222 632898 380404 633134
rect 379804 597454 380404 632898
rect 379804 597218 379986 597454
rect 380222 597218 380404 597454
rect 379804 597134 380404 597218
rect 379804 596898 379986 597134
rect 380222 596898 380404 597134
rect 379804 561454 380404 596898
rect 379804 561218 379986 561454
rect 380222 561218 380404 561454
rect 379804 561134 380404 561218
rect 379804 560898 379986 561134
rect 380222 560898 380404 561134
rect 379804 525454 380404 560898
rect 379804 525218 379986 525454
rect 380222 525218 380404 525454
rect 379804 525134 380404 525218
rect 379804 524898 379986 525134
rect 380222 524898 380404 525134
rect 379804 489454 380404 524898
rect 379804 489218 379986 489454
rect 380222 489218 380404 489454
rect 379804 489134 380404 489218
rect 379804 488898 379986 489134
rect 380222 488898 380404 489134
rect 379804 453454 380404 488898
rect 379804 453218 379986 453454
rect 380222 453218 380404 453454
rect 379804 453134 380404 453218
rect 379804 452898 379986 453134
rect 380222 452898 380404 453134
rect 379804 417454 380404 452898
rect 379804 417218 379986 417454
rect 380222 417218 380404 417454
rect 379804 417134 380404 417218
rect 379804 416898 379986 417134
rect 380222 416898 380404 417134
rect 379804 381454 380404 416898
rect 379804 381218 379986 381454
rect 380222 381218 380404 381454
rect 379804 381134 380404 381218
rect 379804 380898 379986 381134
rect 380222 380898 380404 381134
rect 379804 345454 380404 380898
rect 379804 345218 379986 345454
rect 380222 345218 380404 345454
rect 379804 345134 380404 345218
rect 379804 344898 379986 345134
rect 380222 344898 380404 345134
rect 379804 309454 380404 344898
rect 379804 309218 379986 309454
rect 380222 309218 380404 309454
rect 379804 309134 380404 309218
rect 379804 308898 379986 309134
rect 380222 308898 380404 309134
rect 379804 273454 380404 308898
rect 379804 273218 379986 273454
rect 380222 273218 380404 273454
rect 379804 273134 380404 273218
rect 379804 272898 379986 273134
rect 380222 272898 380404 273134
rect 379804 237454 380404 272898
rect 379804 237218 379986 237454
rect 380222 237218 380404 237454
rect 379804 237134 380404 237218
rect 379804 236898 379986 237134
rect 380222 236898 380404 237134
rect 379804 201454 380404 236898
rect 379804 201218 379986 201454
rect 380222 201218 380404 201454
rect 379804 201134 380404 201218
rect 379804 200898 379986 201134
rect 380222 200898 380404 201134
rect 379804 165454 380404 200898
rect 379804 165218 379986 165454
rect 380222 165218 380404 165454
rect 379804 165134 380404 165218
rect 379804 164898 379986 165134
rect 380222 164898 380404 165134
rect 379804 129454 380404 164898
rect 379804 129218 379986 129454
rect 380222 129218 380404 129454
rect 379804 129134 380404 129218
rect 379804 128898 379986 129134
rect 380222 128898 380404 129134
rect 379804 93454 380404 128898
rect 379804 93218 379986 93454
rect 380222 93218 380404 93454
rect 379804 93134 380404 93218
rect 379804 92898 379986 93134
rect 380222 92898 380404 93134
rect 379804 57454 380404 92898
rect 379804 57218 379986 57454
rect 380222 57218 380404 57454
rect 379804 57134 380404 57218
rect 379804 56898 379986 57134
rect 380222 56898 380404 57134
rect 379804 21454 380404 56898
rect 379804 21218 379986 21454
rect 380222 21218 380404 21454
rect 379804 21134 380404 21218
rect 379804 20898 379986 21134
rect 380222 20898 380404 21134
rect 379804 -1286 380404 20898
rect 379804 -1522 379986 -1286
rect 380222 -1522 380404 -1286
rect 379804 -1606 380404 -1522
rect 379804 -1842 379986 -1606
rect 380222 -1842 380404 -1606
rect 379804 -1864 380404 -1842
rect 383404 673054 384004 707102
rect 383404 672818 383586 673054
rect 383822 672818 384004 673054
rect 383404 672734 384004 672818
rect 383404 672498 383586 672734
rect 383822 672498 384004 672734
rect 383404 637054 384004 672498
rect 383404 636818 383586 637054
rect 383822 636818 384004 637054
rect 383404 636734 384004 636818
rect 383404 636498 383586 636734
rect 383822 636498 384004 636734
rect 383404 601054 384004 636498
rect 383404 600818 383586 601054
rect 383822 600818 384004 601054
rect 383404 600734 384004 600818
rect 383404 600498 383586 600734
rect 383822 600498 384004 600734
rect 383404 565054 384004 600498
rect 383404 564818 383586 565054
rect 383822 564818 384004 565054
rect 383404 564734 384004 564818
rect 383404 564498 383586 564734
rect 383822 564498 384004 564734
rect 383404 529054 384004 564498
rect 383404 528818 383586 529054
rect 383822 528818 384004 529054
rect 383404 528734 384004 528818
rect 383404 528498 383586 528734
rect 383822 528498 384004 528734
rect 383404 493054 384004 528498
rect 383404 492818 383586 493054
rect 383822 492818 384004 493054
rect 383404 492734 384004 492818
rect 383404 492498 383586 492734
rect 383822 492498 384004 492734
rect 383404 457054 384004 492498
rect 383404 456818 383586 457054
rect 383822 456818 384004 457054
rect 383404 456734 384004 456818
rect 383404 456498 383586 456734
rect 383822 456498 384004 456734
rect 383404 421054 384004 456498
rect 383404 420818 383586 421054
rect 383822 420818 384004 421054
rect 383404 420734 384004 420818
rect 383404 420498 383586 420734
rect 383822 420498 384004 420734
rect 383404 385054 384004 420498
rect 383404 384818 383586 385054
rect 383822 384818 384004 385054
rect 383404 384734 384004 384818
rect 383404 384498 383586 384734
rect 383822 384498 384004 384734
rect 383404 349054 384004 384498
rect 383404 348818 383586 349054
rect 383822 348818 384004 349054
rect 383404 348734 384004 348818
rect 383404 348498 383586 348734
rect 383822 348498 384004 348734
rect 383404 313054 384004 348498
rect 383404 312818 383586 313054
rect 383822 312818 384004 313054
rect 383404 312734 384004 312818
rect 383404 312498 383586 312734
rect 383822 312498 384004 312734
rect 383404 277054 384004 312498
rect 383404 276818 383586 277054
rect 383822 276818 384004 277054
rect 383404 276734 384004 276818
rect 383404 276498 383586 276734
rect 383822 276498 384004 276734
rect 383404 241054 384004 276498
rect 383404 240818 383586 241054
rect 383822 240818 384004 241054
rect 383404 240734 384004 240818
rect 383404 240498 383586 240734
rect 383822 240498 384004 240734
rect 383404 205054 384004 240498
rect 383404 204818 383586 205054
rect 383822 204818 384004 205054
rect 383404 204734 384004 204818
rect 383404 204498 383586 204734
rect 383822 204498 384004 204734
rect 383404 169054 384004 204498
rect 383404 168818 383586 169054
rect 383822 168818 384004 169054
rect 383404 168734 384004 168818
rect 383404 168498 383586 168734
rect 383822 168498 384004 168734
rect 383404 133054 384004 168498
rect 383404 132818 383586 133054
rect 383822 132818 384004 133054
rect 383404 132734 384004 132818
rect 383404 132498 383586 132734
rect 383822 132498 384004 132734
rect 383404 97054 384004 132498
rect 383404 96818 383586 97054
rect 383822 96818 384004 97054
rect 383404 96734 384004 96818
rect 383404 96498 383586 96734
rect 383822 96498 384004 96734
rect 383404 61054 384004 96498
rect 383404 60818 383586 61054
rect 383822 60818 384004 61054
rect 383404 60734 384004 60818
rect 383404 60498 383586 60734
rect 383822 60498 384004 60734
rect 383404 25054 384004 60498
rect 383404 24818 383586 25054
rect 383822 24818 384004 25054
rect 383404 24734 384004 24818
rect 383404 24498 383586 24734
rect 383822 24498 384004 24734
rect 383404 -3166 384004 24498
rect 383404 -3402 383586 -3166
rect 383822 -3402 384004 -3166
rect 383404 -3486 384004 -3402
rect 383404 -3722 383586 -3486
rect 383822 -3722 384004 -3486
rect 383404 -3744 384004 -3722
rect 387004 676654 387604 708982
rect 387004 676418 387186 676654
rect 387422 676418 387604 676654
rect 387004 676334 387604 676418
rect 387004 676098 387186 676334
rect 387422 676098 387604 676334
rect 387004 640654 387604 676098
rect 387004 640418 387186 640654
rect 387422 640418 387604 640654
rect 387004 640334 387604 640418
rect 387004 640098 387186 640334
rect 387422 640098 387604 640334
rect 387004 604654 387604 640098
rect 387004 604418 387186 604654
rect 387422 604418 387604 604654
rect 387004 604334 387604 604418
rect 387004 604098 387186 604334
rect 387422 604098 387604 604334
rect 387004 568654 387604 604098
rect 387004 568418 387186 568654
rect 387422 568418 387604 568654
rect 387004 568334 387604 568418
rect 387004 568098 387186 568334
rect 387422 568098 387604 568334
rect 387004 532654 387604 568098
rect 387004 532418 387186 532654
rect 387422 532418 387604 532654
rect 387004 532334 387604 532418
rect 387004 532098 387186 532334
rect 387422 532098 387604 532334
rect 387004 496654 387604 532098
rect 387004 496418 387186 496654
rect 387422 496418 387604 496654
rect 387004 496334 387604 496418
rect 387004 496098 387186 496334
rect 387422 496098 387604 496334
rect 387004 460654 387604 496098
rect 387004 460418 387186 460654
rect 387422 460418 387604 460654
rect 387004 460334 387604 460418
rect 387004 460098 387186 460334
rect 387422 460098 387604 460334
rect 387004 424654 387604 460098
rect 387004 424418 387186 424654
rect 387422 424418 387604 424654
rect 387004 424334 387604 424418
rect 387004 424098 387186 424334
rect 387422 424098 387604 424334
rect 387004 388654 387604 424098
rect 387004 388418 387186 388654
rect 387422 388418 387604 388654
rect 387004 388334 387604 388418
rect 387004 388098 387186 388334
rect 387422 388098 387604 388334
rect 387004 352654 387604 388098
rect 387004 352418 387186 352654
rect 387422 352418 387604 352654
rect 387004 352334 387604 352418
rect 387004 352098 387186 352334
rect 387422 352098 387604 352334
rect 387004 316654 387604 352098
rect 387004 316418 387186 316654
rect 387422 316418 387604 316654
rect 387004 316334 387604 316418
rect 387004 316098 387186 316334
rect 387422 316098 387604 316334
rect 387004 280654 387604 316098
rect 387004 280418 387186 280654
rect 387422 280418 387604 280654
rect 387004 280334 387604 280418
rect 387004 280098 387186 280334
rect 387422 280098 387604 280334
rect 387004 244654 387604 280098
rect 387004 244418 387186 244654
rect 387422 244418 387604 244654
rect 387004 244334 387604 244418
rect 387004 244098 387186 244334
rect 387422 244098 387604 244334
rect 387004 208654 387604 244098
rect 387004 208418 387186 208654
rect 387422 208418 387604 208654
rect 387004 208334 387604 208418
rect 387004 208098 387186 208334
rect 387422 208098 387604 208334
rect 387004 172654 387604 208098
rect 387004 172418 387186 172654
rect 387422 172418 387604 172654
rect 387004 172334 387604 172418
rect 387004 172098 387186 172334
rect 387422 172098 387604 172334
rect 387004 136654 387604 172098
rect 387004 136418 387186 136654
rect 387422 136418 387604 136654
rect 387004 136334 387604 136418
rect 387004 136098 387186 136334
rect 387422 136098 387604 136334
rect 387004 100654 387604 136098
rect 387004 100418 387186 100654
rect 387422 100418 387604 100654
rect 387004 100334 387604 100418
rect 387004 100098 387186 100334
rect 387422 100098 387604 100334
rect 387004 64654 387604 100098
rect 387004 64418 387186 64654
rect 387422 64418 387604 64654
rect 387004 64334 387604 64418
rect 387004 64098 387186 64334
rect 387422 64098 387604 64334
rect 387004 28654 387604 64098
rect 387004 28418 387186 28654
rect 387422 28418 387604 28654
rect 387004 28334 387604 28418
rect 387004 28098 387186 28334
rect 387422 28098 387604 28334
rect 387004 -5046 387604 28098
rect 387004 -5282 387186 -5046
rect 387422 -5282 387604 -5046
rect 387004 -5366 387604 -5282
rect 387004 -5602 387186 -5366
rect 387422 -5602 387604 -5366
rect 387004 -5624 387604 -5602
rect 390604 680254 391204 710862
rect 408604 710478 409204 711440
rect 408604 710242 408786 710478
rect 409022 710242 409204 710478
rect 408604 710158 409204 710242
rect 408604 709922 408786 710158
rect 409022 709922 409204 710158
rect 405004 708598 405604 709560
rect 405004 708362 405186 708598
rect 405422 708362 405604 708598
rect 405004 708278 405604 708362
rect 405004 708042 405186 708278
rect 405422 708042 405604 708278
rect 401404 706718 402004 707680
rect 401404 706482 401586 706718
rect 401822 706482 402004 706718
rect 401404 706398 402004 706482
rect 401404 706162 401586 706398
rect 401822 706162 402004 706398
rect 390604 680018 390786 680254
rect 391022 680018 391204 680254
rect 390604 679934 391204 680018
rect 390604 679698 390786 679934
rect 391022 679698 391204 679934
rect 390604 644254 391204 679698
rect 390604 644018 390786 644254
rect 391022 644018 391204 644254
rect 390604 643934 391204 644018
rect 390604 643698 390786 643934
rect 391022 643698 391204 643934
rect 390604 608254 391204 643698
rect 390604 608018 390786 608254
rect 391022 608018 391204 608254
rect 390604 607934 391204 608018
rect 390604 607698 390786 607934
rect 391022 607698 391204 607934
rect 390604 572254 391204 607698
rect 390604 572018 390786 572254
rect 391022 572018 391204 572254
rect 390604 571934 391204 572018
rect 390604 571698 390786 571934
rect 391022 571698 391204 571934
rect 390604 536254 391204 571698
rect 390604 536018 390786 536254
rect 391022 536018 391204 536254
rect 390604 535934 391204 536018
rect 390604 535698 390786 535934
rect 391022 535698 391204 535934
rect 390604 500254 391204 535698
rect 390604 500018 390786 500254
rect 391022 500018 391204 500254
rect 390604 499934 391204 500018
rect 390604 499698 390786 499934
rect 391022 499698 391204 499934
rect 390604 464254 391204 499698
rect 390604 464018 390786 464254
rect 391022 464018 391204 464254
rect 390604 463934 391204 464018
rect 390604 463698 390786 463934
rect 391022 463698 391204 463934
rect 390604 428254 391204 463698
rect 390604 428018 390786 428254
rect 391022 428018 391204 428254
rect 390604 427934 391204 428018
rect 390604 427698 390786 427934
rect 391022 427698 391204 427934
rect 390604 392254 391204 427698
rect 390604 392018 390786 392254
rect 391022 392018 391204 392254
rect 390604 391934 391204 392018
rect 390604 391698 390786 391934
rect 391022 391698 391204 391934
rect 390604 356254 391204 391698
rect 390604 356018 390786 356254
rect 391022 356018 391204 356254
rect 390604 355934 391204 356018
rect 390604 355698 390786 355934
rect 391022 355698 391204 355934
rect 390604 320254 391204 355698
rect 390604 320018 390786 320254
rect 391022 320018 391204 320254
rect 390604 319934 391204 320018
rect 390604 319698 390786 319934
rect 391022 319698 391204 319934
rect 390604 284254 391204 319698
rect 390604 284018 390786 284254
rect 391022 284018 391204 284254
rect 390604 283934 391204 284018
rect 390604 283698 390786 283934
rect 391022 283698 391204 283934
rect 390604 248254 391204 283698
rect 390604 248018 390786 248254
rect 391022 248018 391204 248254
rect 390604 247934 391204 248018
rect 390604 247698 390786 247934
rect 391022 247698 391204 247934
rect 390604 212254 391204 247698
rect 390604 212018 390786 212254
rect 391022 212018 391204 212254
rect 390604 211934 391204 212018
rect 390604 211698 390786 211934
rect 391022 211698 391204 211934
rect 390604 176254 391204 211698
rect 390604 176018 390786 176254
rect 391022 176018 391204 176254
rect 390604 175934 391204 176018
rect 390604 175698 390786 175934
rect 391022 175698 391204 175934
rect 390604 140254 391204 175698
rect 390604 140018 390786 140254
rect 391022 140018 391204 140254
rect 390604 139934 391204 140018
rect 390604 139698 390786 139934
rect 391022 139698 391204 139934
rect 390604 104254 391204 139698
rect 390604 104018 390786 104254
rect 391022 104018 391204 104254
rect 390604 103934 391204 104018
rect 390604 103698 390786 103934
rect 391022 103698 391204 103934
rect 390604 68254 391204 103698
rect 390604 68018 390786 68254
rect 391022 68018 391204 68254
rect 390604 67934 391204 68018
rect 390604 67698 390786 67934
rect 391022 67698 391204 67934
rect 390604 32254 391204 67698
rect 390604 32018 390786 32254
rect 391022 32018 391204 32254
rect 390604 31934 391204 32018
rect 390604 31698 390786 31934
rect 391022 31698 391204 31934
rect 372604 -6222 372786 -5986
rect 373022 -6222 373204 -5986
rect 372604 -6306 373204 -6222
rect 372604 -6542 372786 -6306
rect 373022 -6542 373204 -6306
rect 372604 -7504 373204 -6542
rect 390604 -6926 391204 31698
rect 397804 704838 398404 705800
rect 397804 704602 397986 704838
rect 398222 704602 398404 704838
rect 397804 704518 398404 704602
rect 397804 704282 397986 704518
rect 398222 704282 398404 704518
rect 397804 687454 398404 704282
rect 397804 687218 397986 687454
rect 398222 687218 398404 687454
rect 397804 687134 398404 687218
rect 397804 686898 397986 687134
rect 398222 686898 398404 687134
rect 397804 651454 398404 686898
rect 397804 651218 397986 651454
rect 398222 651218 398404 651454
rect 397804 651134 398404 651218
rect 397804 650898 397986 651134
rect 398222 650898 398404 651134
rect 397804 615454 398404 650898
rect 397804 615218 397986 615454
rect 398222 615218 398404 615454
rect 397804 615134 398404 615218
rect 397804 614898 397986 615134
rect 398222 614898 398404 615134
rect 397804 579454 398404 614898
rect 397804 579218 397986 579454
rect 398222 579218 398404 579454
rect 397804 579134 398404 579218
rect 397804 578898 397986 579134
rect 398222 578898 398404 579134
rect 397804 543454 398404 578898
rect 397804 543218 397986 543454
rect 398222 543218 398404 543454
rect 397804 543134 398404 543218
rect 397804 542898 397986 543134
rect 398222 542898 398404 543134
rect 397804 507454 398404 542898
rect 397804 507218 397986 507454
rect 398222 507218 398404 507454
rect 397804 507134 398404 507218
rect 397804 506898 397986 507134
rect 398222 506898 398404 507134
rect 397804 471454 398404 506898
rect 397804 471218 397986 471454
rect 398222 471218 398404 471454
rect 397804 471134 398404 471218
rect 397804 470898 397986 471134
rect 398222 470898 398404 471134
rect 397804 435454 398404 470898
rect 397804 435218 397986 435454
rect 398222 435218 398404 435454
rect 397804 435134 398404 435218
rect 397804 434898 397986 435134
rect 398222 434898 398404 435134
rect 397804 399454 398404 434898
rect 397804 399218 397986 399454
rect 398222 399218 398404 399454
rect 397804 399134 398404 399218
rect 397804 398898 397986 399134
rect 398222 398898 398404 399134
rect 397804 363454 398404 398898
rect 397804 363218 397986 363454
rect 398222 363218 398404 363454
rect 397804 363134 398404 363218
rect 397804 362898 397986 363134
rect 398222 362898 398404 363134
rect 397804 327454 398404 362898
rect 397804 327218 397986 327454
rect 398222 327218 398404 327454
rect 397804 327134 398404 327218
rect 397804 326898 397986 327134
rect 398222 326898 398404 327134
rect 397804 291454 398404 326898
rect 397804 291218 397986 291454
rect 398222 291218 398404 291454
rect 397804 291134 398404 291218
rect 397804 290898 397986 291134
rect 398222 290898 398404 291134
rect 397804 255454 398404 290898
rect 397804 255218 397986 255454
rect 398222 255218 398404 255454
rect 397804 255134 398404 255218
rect 397804 254898 397986 255134
rect 398222 254898 398404 255134
rect 397804 219454 398404 254898
rect 397804 219218 397986 219454
rect 398222 219218 398404 219454
rect 397804 219134 398404 219218
rect 397804 218898 397986 219134
rect 398222 218898 398404 219134
rect 397804 183454 398404 218898
rect 397804 183218 397986 183454
rect 398222 183218 398404 183454
rect 397804 183134 398404 183218
rect 397804 182898 397986 183134
rect 398222 182898 398404 183134
rect 397804 147454 398404 182898
rect 397804 147218 397986 147454
rect 398222 147218 398404 147454
rect 397804 147134 398404 147218
rect 397804 146898 397986 147134
rect 398222 146898 398404 147134
rect 397804 111454 398404 146898
rect 397804 111218 397986 111454
rect 398222 111218 398404 111454
rect 397804 111134 398404 111218
rect 397804 110898 397986 111134
rect 398222 110898 398404 111134
rect 397804 75454 398404 110898
rect 397804 75218 397986 75454
rect 398222 75218 398404 75454
rect 397804 75134 398404 75218
rect 397804 74898 397986 75134
rect 398222 74898 398404 75134
rect 397804 39454 398404 74898
rect 397804 39218 397986 39454
rect 398222 39218 398404 39454
rect 397804 39134 398404 39218
rect 397804 38898 397986 39134
rect 398222 38898 398404 39134
rect 397804 3454 398404 38898
rect 397804 3218 397986 3454
rect 398222 3218 398404 3454
rect 397804 3134 398404 3218
rect 397804 2898 397986 3134
rect 398222 2898 398404 3134
rect 397804 -346 398404 2898
rect 397804 -582 397986 -346
rect 398222 -582 398404 -346
rect 397804 -666 398404 -582
rect 397804 -902 397986 -666
rect 398222 -902 398404 -666
rect 397804 -1864 398404 -902
rect 401404 691054 402004 706162
rect 401404 690818 401586 691054
rect 401822 690818 402004 691054
rect 401404 690734 402004 690818
rect 401404 690498 401586 690734
rect 401822 690498 402004 690734
rect 401404 655054 402004 690498
rect 401404 654818 401586 655054
rect 401822 654818 402004 655054
rect 401404 654734 402004 654818
rect 401404 654498 401586 654734
rect 401822 654498 402004 654734
rect 401404 619054 402004 654498
rect 401404 618818 401586 619054
rect 401822 618818 402004 619054
rect 401404 618734 402004 618818
rect 401404 618498 401586 618734
rect 401822 618498 402004 618734
rect 401404 583054 402004 618498
rect 401404 582818 401586 583054
rect 401822 582818 402004 583054
rect 401404 582734 402004 582818
rect 401404 582498 401586 582734
rect 401822 582498 402004 582734
rect 401404 547054 402004 582498
rect 401404 546818 401586 547054
rect 401822 546818 402004 547054
rect 401404 546734 402004 546818
rect 401404 546498 401586 546734
rect 401822 546498 402004 546734
rect 401404 511054 402004 546498
rect 401404 510818 401586 511054
rect 401822 510818 402004 511054
rect 401404 510734 402004 510818
rect 401404 510498 401586 510734
rect 401822 510498 402004 510734
rect 401404 475054 402004 510498
rect 401404 474818 401586 475054
rect 401822 474818 402004 475054
rect 401404 474734 402004 474818
rect 401404 474498 401586 474734
rect 401822 474498 402004 474734
rect 401404 439054 402004 474498
rect 401404 438818 401586 439054
rect 401822 438818 402004 439054
rect 401404 438734 402004 438818
rect 401404 438498 401586 438734
rect 401822 438498 402004 438734
rect 401404 403054 402004 438498
rect 401404 402818 401586 403054
rect 401822 402818 402004 403054
rect 401404 402734 402004 402818
rect 401404 402498 401586 402734
rect 401822 402498 402004 402734
rect 401404 367054 402004 402498
rect 401404 366818 401586 367054
rect 401822 366818 402004 367054
rect 401404 366734 402004 366818
rect 401404 366498 401586 366734
rect 401822 366498 402004 366734
rect 401404 331054 402004 366498
rect 401404 330818 401586 331054
rect 401822 330818 402004 331054
rect 401404 330734 402004 330818
rect 401404 330498 401586 330734
rect 401822 330498 402004 330734
rect 401404 295054 402004 330498
rect 401404 294818 401586 295054
rect 401822 294818 402004 295054
rect 401404 294734 402004 294818
rect 401404 294498 401586 294734
rect 401822 294498 402004 294734
rect 401404 259054 402004 294498
rect 401404 258818 401586 259054
rect 401822 258818 402004 259054
rect 401404 258734 402004 258818
rect 401404 258498 401586 258734
rect 401822 258498 402004 258734
rect 401404 223054 402004 258498
rect 401404 222818 401586 223054
rect 401822 222818 402004 223054
rect 401404 222734 402004 222818
rect 401404 222498 401586 222734
rect 401822 222498 402004 222734
rect 401404 187054 402004 222498
rect 401404 186818 401586 187054
rect 401822 186818 402004 187054
rect 401404 186734 402004 186818
rect 401404 186498 401586 186734
rect 401822 186498 402004 186734
rect 401404 151054 402004 186498
rect 401404 150818 401586 151054
rect 401822 150818 402004 151054
rect 401404 150734 402004 150818
rect 401404 150498 401586 150734
rect 401822 150498 402004 150734
rect 401404 115054 402004 150498
rect 401404 114818 401586 115054
rect 401822 114818 402004 115054
rect 401404 114734 402004 114818
rect 401404 114498 401586 114734
rect 401822 114498 402004 114734
rect 401404 79054 402004 114498
rect 401404 78818 401586 79054
rect 401822 78818 402004 79054
rect 401404 78734 402004 78818
rect 401404 78498 401586 78734
rect 401822 78498 402004 78734
rect 401404 43054 402004 78498
rect 401404 42818 401586 43054
rect 401822 42818 402004 43054
rect 401404 42734 402004 42818
rect 401404 42498 401586 42734
rect 401822 42498 402004 42734
rect 401404 7054 402004 42498
rect 401404 6818 401586 7054
rect 401822 6818 402004 7054
rect 401404 6734 402004 6818
rect 401404 6498 401586 6734
rect 401822 6498 402004 6734
rect 401404 -2226 402004 6498
rect 401404 -2462 401586 -2226
rect 401822 -2462 402004 -2226
rect 401404 -2546 402004 -2462
rect 401404 -2782 401586 -2546
rect 401822 -2782 402004 -2546
rect 401404 -3744 402004 -2782
rect 405004 694654 405604 708042
rect 405004 694418 405186 694654
rect 405422 694418 405604 694654
rect 405004 694334 405604 694418
rect 405004 694098 405186 694334
rect 405422 694098 405604 694334
rect 405004 658654 405604 694098
rect 405004 658418 405186 658654
rect 405422 658418 405604 658654
rect 405004 658334 405604 658418
rect 405004 658098 405186 658334
rect 405422 658098 405604 658334
rect 405004 622654 405604 658098
rect 405004 622418 405186 622654
rect 405422 622418 405604 622654
rect 405004 622334 405604 622418
rect 405004 622098 405186 622334
rect 405422 622098 405604 622334
rect 405004 586654 405604 622098
rect 405004 586418 405186 586654
rect 405422 586418 405604 586654
rect 405004 586334 405604 586418
rect 405004 586098 405186 586334
rect 405422 586098 405604 586334
rect 405004 550654 405604 586098
rect 405004 550418 405186 550654
rect 405422 550418 405604 550654
rect 405004 550334 405604 550418
rect 405004 550098 405186 550334
rect 405422 550098 405604 550334
rect 405004 514654 405604 550098
rect 405004 514418 405186 514654
rect 405422 514418 405604 514654
rect 405004 514334 405604 514418
rect 405004 514098 405186 514334
rect 405422 514098 405604 514334
rect 405004 478654 405604 514098
rect 405004 478418 405186 478654
rect 405422 478418 405604 478654
rect 405004 478334 405604 478418
rect 405004 478098 405186 478334
rect 405422 478098 405604 478334
rect 405004 442654 405604 478098
rect 405004 442418 405186 442654
rect 405422 442418 405604 442654
rect 405004 442334 405604 442418
rect 405004 442098 405186 442334
rect 405422 442098 405604 442334
rect 405004 406654 405604 442098
rect 405004 406418 405186 406654
rect 405422 406418 405604 406654
rect 405004 406334 405604 406418
rect 405004 406098 405186 406334
rect 405422 406098 405604 406334
rect 405004 370654 405604 406098
rect 405004 370418 405186 370654
rect 405422 370418 405604 370654
rect 405004 370334 405604 370418
rect 405004 370098 405186 370334
rect 405422 370098 405604 370334
rect 405004 334654 405604 370098
rect 405004 334418 405186 334654
rect 405422 334418 405604 334654
rect 405004 334334 405604 334418
rect 405004 334098 405186 334334
rect 405422 334098 405604 334334
rect 405004 298654 405604 334098
rect 405004 298418 405186 298654
rect 405422 298418 405604 298654
rect 405004 298334 405604 298418
rect 405004 298098 405186 298334
rect 405422 298098 405604 298334
rect 405004 262654 405604 298098
rect 405004 262418 405186 262654
rect 405422 262418 405604 262654
rect 405004 262334 405604 262418
rect 405004 262098 405186 262334
rect 405422 262098 405604 262334
rect 405004 226654 405604 262098
rect 405004 226418 405186 226654
rect 405422 226418 405604 226654
rect 405004 226334 405604 226418
rect 405004 226098 405186 226334
rect 405422 226098 405604 226334
rect 405004 190654 405604 226098
rect 405004 190418 405186 190654
rect 405422 190418 405604 190654
rect 405004 190334 405604 190418
rect 405004 190098 405186 190334
rect 405422 190098 405604 190334
rect 405004 154654 405604 190098
rect 405004 154418 405186 154654
rect 405422 154418 405604 154654
rect 405004 154334 405604 154418
rect 405004 154098 405186 154334
rect 405422 154098 405604 154334
rect 405004 118654 405604 154098
rect 405004 118418 405186 118654
rect 405422 118418 405604 118654
rect 405004 118334 405604 118418
rect 405004 118098 405186 118334
rect 405422 118098 405604 118334
rect 405004 82654 405604 118098
rect 405004 82418 405186 82654
rect 405422 82418 405604 82654
rect 405004 82334 405604 82418
rect 405004 82098 405186 82334
rect 405422 82098 405604 82334
rect 405004 46654 405604 82098
rect 405004 46418 405186 46654
rect 405422 46418 405604 46654
rect 405004 46334 405604 46418
rect 405004 46098 405186 46334
rect 405422 46098 405604 46334
rect 405004 10654 405604 46098
rect 405004 10418 405186 10654
rect 405422 10418 405604 10654
rect 405004 10334 405604 10418
rect 405004 10098 405186 10334
rect 405422 10098 405604 10334
rect 405004 -4106 405604 10098
rect 405004 -4342 405186 -4106
rect 405422 -4342 405604 -4106
rect 405004 -4426 405604 -4342
rect 405004 -4662 405186 -4426
rect 405422 -4662 405604 -4426
rect 405004 -5624 405604 -4662
rect 408604 698254 409204 709922
rect 426604 711418 427204 711440
rect 426604 711182 426786 711418
rect 427022 711182 427204 711418
rect 426604 711098 427204 711182
rect 426604 710862 426786 711098
rect 427022 710862 427204 711098
rect 423004 709538 423604 709560
rect 423004 709302 423186 709538
rect 423422 709302 423604 709538
rect 423004 709218 423604 709302
rect 423004 708982 423186 709218
rect 423422 708982 423604 709218
rect 419404 707658 420004 707680
rect 419404 707422 419586 707658
rect 419822 707422 420004 707658
rect 419404 707338 420004 707422
rect 419404 707102 419586 707338
rect 419822 707102 420004 707338
rect 408604 698018 408786 698254
rect 409022 698018 409204 698254
rect 408604 697934 409204 698018
rect 408604 697698 408786 697934
rect 409022 697698 409204 697934
rect 408604 662254 409204 697698
rect 408604 662018 408786 662254
rect 409022 662018 409204 662254
rect 408604 661934 409204 662018
rect 408604 661698 408786 661934
rect 409022 661698 409204 661934
rect 408604 626254 409204 661698
rect 408604 626018 408786 626254
rect 409022 626018 409204 626254
rect 408604 625934 409204 626018
rect 408604 625698 408786 625934
rect 409022 625698 409204 625934
rect 408604 590254 409204 625698
rect 408604 590018 408786 590254
rect 409022 590018 409204 590254
rect 408604 589934 409204 590018
rect 408604 589698 408786 589934
rect 409022 589698 409204 589934
rect 408604 554254 409204 589698
rect 408604 554018 408786 554254
rect 409022 554018 409204 554254
rect 408604 553934 409204 554018
rect 408604 553698 408786 553934
rect 409022 553698 409204 553934
rect 408604 518254 409204 553698
rect 408604 518018 408786 518254
rect 409022 518018 409204 518254
rect 408604 517934 409204 518018
rect 408604 517698 408786 517934
rect 409022 517698 409204 517934
rect 408604 482254 409204 517698
rect 408604 482018 408786 482254
rect 409022 482018 409204 482254
rect 408604 481934 409204 482018
rect 408604 481698 408786 481934
rect 409022 481698 409204 481934
rect 408604 446254 409204 481698
rect 408604 446018 408786 446254
rect 409022 446018 409204 446254
rect 408604 445934 409204 446018
rect 408604 445698 408786 445934
rect 409022 445698 409204 445934
rect 408604 410254 409204 445698
rect 408604 410018 408786 410254
rect 409022 410018 409204 410254
rect 408604 409934 409204 410018
rect 408604 409698 408786 409934
rect 409022 409698 409204 409934
rect 408604 374254 409204 409698
rect 408604 374018 408786 374254
rect 409022 374018 409204 374254
rect 408604 373934 409204 374018
rect 408604 373698 408786 373934
rect 409022 373698 409204 373934
rect 408604 338254 409204 373698
rect 408604 338018 408786 338254
rect 409022 338018 409204 338254
rect 408604 337934 409204 338018
rect 408604 337698 408786 337934
rect 409022 337698 409204 337934
rect 408604 302254 409204 337698
rect 408604 302018 408786 302254
rect 409022 302018 409204 302254
rect 408604 301934 409204 302018
rect 408604 301698 408786 301934
rect 409022 301698 409204 301934
rect 408604 266254 409204 301698
rect 408604 266018 408786 266254
rect 409022 266018 409204 266254
rect 408604 265934 409204 266018
rect 408604 265698 408786 265934
rect 409022 265698 409204 265934
rect 408604 230254 409204 265698
rect 408604 230018 408786 230254
rect 409022 230018 409204 230254
rect 408604 229934 409204 230018
rect 408604 229698 408786 229934
rect 409022 229698 409204 229934
rect 408604 194254 409204 229698
rect 408604 194018 408786 194254
rect 409022 194018 409204 194254
rect 408604 193934 409204 194018
rect 408604 193698 408786 193934
rect 409022 193698 409204 193934
rect 408604 158254 409204 193698
rect 408604 158018 408786 158254
rect 409022 158018 409204 158254
rect 408604 157934 409204 158018
rect 408604 157698 408786 157934
rect 409022 157698 409204 157934
rect 408604 122254 409204 157698
rect 408604 122018 408786 122254
rect 409022 122018 409204 122254
rect 408604 121934 409204 122018
rect 408604 121698 408786 121934
rect 409022 121698 409204 121934
rect 408604 86254 409204 121698
rect 408604 86018 408786 86254
rect 409022 86018 409204 86254
rect 408604 85934 409204 86018
rect 408604 85698 408786 85934
rect 409022 85698 409204 85934
rect 408604 50254 409204 85698
rect 408604 50018 408786 50254
rect 409022 50018 409204 50254
rect 408604 49934 409204 50018
rect 408604 49698 408786 49934
rect 409022 49698 409204 49934
rect 408604 14254 409204 49698
rect 408604 14018 408786 14254
rect 409022 14018 409204 14254
rect 408604 13934 409204 14018
rect 408604 13698 408786 13934
rect 409022 13698 409204 13934
rect 390604 -7162 390786 -6926
rect 391022 -7162 391204 -6926
rect 390604 -7246 391204 -7162
rect 390604 -7482 390786 -7246
rect 391022 -7482 391204 -7246
rect 390604 -7504 391204 -7482
rect 408604 -5986 409204 13698
rect 415804 705778 416404 705800
rect 415804 705542 415986 705778
rect 416222 705542 416404 705778
rect 415804 705458 416404 705542
rect 415804 705222 415986 705458
rect 416222 705222 416404 705458
rect 415804 669454 416404 705222
rect 415804 669218 415986 669454
rect 416222 669218 416404 669454
rect 415804 669134 416404 669218
rect 415804 668898 415986 669134
rect 416222 668898 416404 669134
rect 415804 633454 416404 668898
rect 415804 633218 415986 633454
rect 416222 633218 416404 633454
rect 415804 633134 416404 633218
rect 415804 632898 415986 633134
rect 416222 632898 416404 633134
rect 415804 597454 416404 632898
rect 415804 597218 415986 597454
rect 416222 597218 416404 597454
rect 415804 597134 416404 597218
rect 415804 596898 415986 597134
rect 416222 596898 416404 597134
rect 415804 561454 416404 596898
rect 415804 561218 415986 561454
rect 416222 561218 416404 561454
rect 415804 561134 416404 561218
rect 415804 560898 415986 561134
rect 416222 560898 416404 561134
rect 415804 525454 416404 560898
rect 415804 525218 415986 525454
rect 416222 525218 416404 525454
rect 415804 525134 416404 525218
rect 415804 524898 415986 525134
rect 416222 524898 416404 525134
rect 415804 489454 416404 524898
rect 415804 489218 415986 489454
rect 416222 489218 416404 489454
rect 415804 489134 416404 489218
rect 415804 488898 415986 489134
rect 416222 488898 416404 489134
rect 415804 453454 416404 488898
rect 415804 453218 415986 453454
rect 416222 453218 416404 453454
rect 415804 453134 416404 453218
rect 415804 452898 415986 453134
rect 416222 452898 416404 453134
rect 415804 417454 416404 452898
rect 415804 417218 415986 417454
rect 416222 417218 416404 417454
rect 415804 417134 416404 417218
rect 415804 416898 415986 417134
rect 416222 416898 416404 417134
rect 415804 381454 416404 416898
rect 415804 381218 415986 381454
rect 416222 381218 416404 381454
rect 415804 381134 416404 381218
rect 415804 380898 415986 381134
rect 416222 380898 416404 381134
rect 415804 345454 416404 380898
rect 415804 345218 415986 345454
rect 416222 345218 416404 345454
rect 415804 345134 416404 345218
rect 415804 344898 415986 345134
rect 416222 344898 416404 345134
rect 415804 309454 416404 344898
rect 415804 309218 415986 309454
rect 416222 309218 416404 309454
rect 415804 309134 416404 309218
rect 415804 308898 415986 309134
rect 416222 308898 416404 309134
rect 415804 273454 416404 308898
rect 415804 273218 415986 273454
rect 416222 273218 416404 273454
rect 415804 273134 416404 273218
rect 415804 272898 415986 273134
rect 416222 272898 416404 273134
rect 415804 237454 416404 272898
rect 415804 237218 415986 237454
rect 416222 237218 416404 237454
rect 415804 237134 416404 237218
rect 415804 236898 415986 237134
rect 416222 236898 416404 237134
rect 415804 201454 416404 236898
rect 415804 201218 415986 201454
rect 416222 201218 416404 201454
rect 415804 201134 416404 201218
rect 415804 200898 415986 201134
rect 416222 200898 416404 201134
rect 415804 165454 416404 200898
rect 415804 165218 415986 165454
rect 416222 165218 416404 165454
rect 415804 165134 416404 165218
rect 415804 164898 415986 165134
rect 416222 164898 416404 165134
rect 415804 129454 416404 164898
rect 415804 129218 415986 129454
rect 416222 129218 416404 129454
rect 415804 129134 416404 129218
rect 415804 128898 415986 129134
rect 416222 128898 416404 129134
rect 415804 93454 416404 128898
rect 415804 93218 415986 93454
rect 416222 93218 416404 93454
rect 415804 93134 416404 93218
rect 415804 92898 415986 93134
rect 416222 92898 416404 93134
rect 415804 57454 416404 92898
rect 415804 57218 415986 57454
rect 416222 57218 416404 57454
rect 415804 57134 416404 57218
rect 415804 56898 415986 57134
rect 416222 56898 416404 57134
rect 415804 21454 416404 56898
rect 415804 21218 415986 21454
rect 416222 21218 416404 21454
rect 415804 21134 416404 21218
rect 415804 20898 415986 21134
rect 416222 20898 416404 21134
rect 415804 -1286 416404 20898
rect 415804 -1522 415986 -1286
rect 416222 -1522 416404 -1286
rect 415804 -1606 416404 -1522
rect 415804 -1842 415986 -1606
rect 416222 -1842 416404 -1606
rect 415804 -1864 416404 -1842
rect 419404 673054 420004 707102
rect 419404 672818 419586 673054
rect 419822 672818 420004 673054
rect 419404 672734 420004 672818
rect 419404 672498 419586 672734
rect 419822 672498 420004 672734
rect 419404 637054 420004 672498
rect 419404 636818 419586 637054
rect 419822 636818 420004 637054
rect 419404 636734 420004 636818
rect 419404 636498 419586 636734
rect 419822 636498 420004 636734
rect 419404 601054 420004 636498
rect 419404 600818 419586 601054
rect 419822 600818 420004 601054
rect 419404 600734 420004 600818
rect 419404 600498 419586 600734
rect 419822 600498 420004 600734
rect 419404 565054 420004 600498
rect 419404 564818 419586 565054
rect 419822 564818 420004 565054
rect 419404 564734 420004 564818
rect 419404 564498 419586 564734
rect 419822 564498 420004 564734
rect 419404 529054 420004 564498
rect 419404 528818 419586 529054
rect 419822 528818 420004 529054
rect 419404 528734 420004 528818
rect 419404 528498 419586 528734
rect 419822 528498 420004 528734
rect 419404 493054 420004 528498
rect 419404 492818 419586 493054
rect 419822 492818 420004 493054
rect 419404 492734 420004 492818
rect 419404 492498 419586 492734
rect 419822 492498 420004 492734
rect 419404 457054 420004 492498
rect 419404 456818 419586 457054
rect 419822 456818 420004 457054
rect 419404 456734 420004 456818
rect 419404 456498 419586 456734
rect 419822 456498 420004 456734
rect 419404 421054 420004 456498
rect 419404 420818 419586 421054
rect 419822 420818 420004 421054
rect 419404 420734 420004 420818
rect 419404 420498 419586 420734
rect 419822 420498 420004 420734
rect 419404 385054 420004 420498
rect 419404 384818 419586 385054
rect 419822 384818 420004 385054
rect 419404 384734 420004 384818
rect 419404 384498 419586 384734
rect 419822 384498 420004 384734
rect 419404 349054 420004 384498
rect 419404 348818 419586 349054
rect 419822 348818 420004 349054
rect 419404 348734 420004 348818
rect 419404 348498 419586 348734
rect 419822 348498 420004 348734
rect 419404 313054 420004 348498
rect 419404 312818 419586 313054
rect 419822 312818 420004 313054
rect 419404 312734 420004 312818
rect 419404 312498 419586 312734
rect 419822 312498 420004 312734
rect 419404 277054 420004 312498
rect 419404 276818 419586 277054
rect 419822 276818 420004 277054
rect 419404 276734 420004 276818
rect 419404 276498 419586 276734
rect 419822 276498 420004 276734
rect 419404 241054 420004 276498
rect 419404 240818 419586 241054
rect 419822 240818 420004 241054
rect 419404 240734 420004 240818
rect 419404 240498 419586 240734
rect 419822 240498 420004 240734
rect 419404 205054 420004 240498
rect 419404 204818 419586 205054
rect 419822 204818 420004 205054
rect 419404 204734 420004 204818
rect 419404 204498 419586 204734
rect 419822 204498 420004 204734
rect 419404 169054 420004 204498
rect 419404 168818 419586 169054
rect 419822 168818 420004 169054
rect 419404 168734 420004 168818
rect 419404 168498 419586 168734
rect 419822 168498 420004 168734
rect 419404 133054 420004 168498
rect 419404 132818 419586 133054
rect 419822 132818 420004 133054
rect 419404 132734 420004 132818
rect 419404 132498 419586 132734
rect 419822 132498 420004 132734
rect 419404 97054 420004 132498
rect 419404 96818 419586 97054
rect 419822 96818 420004 97054
rect 419404 96734 420004 96818
rect 419404 96498 419586 96734
rect 419822 96498 420004 96734
rect 419404 61054 420004 96498
rect 419404 60818 419586 61054
rect 419822 60818 420004 61054
rect 419404 60734 420004 60818
rect 419404 60498 419586 60734
rect 419822 60498 420004 60734
rect 419404 25054 420004 60498
rect 419404 24818 419586 25054
rect 419822 24818 420004 25054
rect 419404 24734 420004 24818
rect 419404 24498 419586 24734
rect 419822 24498 420004 24734
rect 419404 -3166 420004 24498
rect 419404 -3402 419586 -3166
rect 419822 -3402 420004 -3166
rect 419404 -3486 420004 -3402
rect 419404 -3722 419586 -3486
rect 419822 -3722 420004 -3486
rect 419404 -3744 420004 -3722
rect 423004 676654 423604 708982
rect 423004 676418 423186 676654
rect 423422 676418 423604 676654
rect 423004 676334 423604 676418
rect 423004 676098 423186 676334
rect 423422 676098 423604 676334
rect 423004 640654 423604 676098
rect 423004 640418 423186 640654
rect 423422 640418 423604 640654
rect 423004 640334 423604 640418
rect 423004 640098 423186 640334
rect 423422 640098 423604 640334
rect 423004 604654 423604 640098
rect 423004 604418 423186 604654
rect 423422 604418 423604 604654
rect 423004 604334 423604 604418
rect 423004 604098 423186 604334
rect 423422 604098 423604 604334
rect 423004 568654 423604 604098
rect 423004 568418 423186 568654
rect 423422 568418 423604 568654
rect 423004 568334 423604 568418
rect 423004 568098 423186 568334
rect 423422 568098 423604 568334
rect 423004 532654 423604 568098
rect 423004 532418 423186 532654
rect 423422 532418 423604 532654
rect 423004 532334 423604 532418
rect 423004 532098 423186 532334
rect 423422 532098 423604 532334
rect 423004 496654 423604 532098
rect 423004 496418 423186 496654
rect 423422 496418 423604 496654
rect 423004 496334 423604 496418
rect 423004 496098 423186 496334
rect 423422 496098 423604 496334
rect 423004 460654 423604 496098
rect 423004 460418 423186 460654
rect 423422 460418 423604 460654
rect 423004 460334 423604 460418
rect 423004 460098 423186 460334
rect 423422 460098 423604 460334
rect 423004 424654 423604 460098
rect 423004 424418 423186 424654
rect 423422 424418 423604 424654
rect 423004 424334 423604 424418
rect 423004 424098 423186 424334
rect 423422 424098 423604 424334
rect 423004 388654 423604 424098
rect 423004 388418 423186 388654
rect 423422 388418 423604 388654
rect 423004 388334 423604 388418
rect 423004 388098 423186 388334
rect 423422 388098 423604 388334
rect 423004 352654 423604 388098
rect 423004 352418 423186 352654
rect 423422 352418 423604 352654
rect 423004 352334 423604 352418
rect 423004 352098 423186 352334
rect 423422 352098 423604 352334
rect 423004 316654 423604 352098
rect 423004 316418 423186 316654
rect 423422 316418 423604 316654
rect 423004 316334 423604 316418
rect 423004 316098 423186 316334
rect 423422 316098 423604 316334
rect 423004 280654 423604 316098
rect 423004 280418 423186 280654
rect 423422 280418 423604 280654
rect 423004 280334 423604 280418
rect 423004 280098 423186 280334
rect 423422 280098 423604 280334
rect 423004 244654 423604 280098
rect 423004 244418 423186 244654
rect 423422 244418 423604 244654
rect 423004 244334 423604 244418
rect 423004 244098 423186 244334
rect 423422 244098 423604 244334
rect 423004 208654 423604 244098
rect 423004 208418 423186 208654
rect 423422 208418 423604 208654
rect 423004 208334 423604 208418
rect 423004 208098 423186 208334
rect 423422 208098 423604 208334
rect 423004 172654 423604 208098
rect 423004 172418 423186 172654
rect 423422 172418 423604 172654
rect 423004 172334 423604 172418
rect 423004 172098 423186 172334
rect 423422 172098 423604 172334
rect 423004 136654 423604 172098
rect 423004 136418 423186 136654
rect 423422 136418 423604 136654
rect 423004 136334 423604 136418
rect 423004 136098 423186 136334
rect 423422 136098 423604 136334
rect 423004 100654 423604 136098
rect 423004 100418 423186 100654
rect 423422 100418 423604 100654
rect 423004 100334 423604 100418
rect 423004 100098 423186 100334
rect 423422 100098 423604 100334
rect 423004 64654 423604 100098
rect 423004 64418 423186 64654
rect 423422 64418 423604 64654
rect 423004 64334 423604 64418
rect 423004 64098 423186 64334
rect 423422 64098 423604 64334
rect 423004 28654 423604 64098
rect 423004 28418 423186 28654
rect 423422 28418 423604 28654
rect 423004 28334 423604 28418
rect 423004 28098 423186 28334
rect 423422 28098 423604 28334
rect 423004 -5046 423604 28098
rect 423004 -5282 423186 -5046
rect 423422 -5282 423604 -5046
rect 423004 -5366 423604 -5282
rect 423004 -5602 423186 -5366
rect 423422 -5602 423604 -5366
rect 423004 -5624 423604 -5602
rect 426604 680254 427204 710862
rect 444604 710478 445204 711440
rect 444604 710242 444786 710478
rect 445022 710242 445204 710478
rect 444604 710158 445204 710242
rect 444604 709922 444786 710158
rect 445022 709922 445204 710158
rect 441004 708598 441604 709560
rect 441004 708362 441186 708598
rect 441422 708362 441604 708598
rect 441004 708278 441604 708362
rect 441004 708042 441186 708278
rect 441422 708042 441604 708278
rect 437404 706718 438004 707680
rect 437404 706482 437586 706718
rect 437822 706482 438004 706718
rect 437404 706398 438004 706482
rect 437404 706162 437586 706398
rect 437822 706162 438004 706398
rect 426604 680018 426786 680254
rect 427022 680018 427204 680254
rect 426604 679934 427204 680018
rect 426604 679698 426786 679934
rect 427022 679698 427204 679934
rect 426604 644254 427204 679698
rect 426604 644018 426786 644254
rect 427022 644018 427204 644254
rect 426604 643934 427204 644018
rect 426604 643698 426786 643934
rect 427022 643698 427204 643934
rect 426604 608254 427204 643698
rect 426604 608018 426786 608254
rect 427022 608018 427204 608254
rect 426604 607934 427204 608018
rect 426604 607698 426786 607934
rect 427022 607698 427204 607934
rect 426604 572254 427204 607698
rect 426604 572018 426786 572254
rect 427022 572018 427204 572254
rect 426604 571934 427204 572018
rect 426604 571698 426786 571934
rect 427022 571698 427204 571934
rect 426604 536254 427204 571698
rect 426604 536018 426786 536254
rect 427022 536018 427204 536254
rect 426604 535934 427204 536018
rect 426604 535698 426786 535934
rect 427022 535698 427204 535934
rect 426604 500254 427204 535698
rect 426604 500018 426786 500254
rect 427022 500018 427204 500254
rect 426604 499934 427204 500018
rect 426604 499698 426786 499934
rect 427022 499698 427204 499934
rect 426604 464254 427204 499698
rect 426604 464018 426786 464254
rect 427022 464018 427204 464254
rect 426604 463934 427204 464018
rect 426604 463698 426786 463934
rect 427022 463698 427204 463934
rect 426604 428254 427204 463698
rect 426604 428018 426786 428254
rect 427022 428018 427204 428254
rect 426604 427934 427204 428018
rect 426604 427698 426786 427934
rect 427022 427698 427204 427934
rect 426604 392254 427204 427698
rect 426604 392018 426786 392254
rect 427022 392018 427204 392254
rect 426604 391934 427204 392018
rect 426604 391698 426786 391934
rect 427022 391698 427204 391934
rect 426604 356254 427204 391698
rect 426604 356018 426786 356254
rect 427022 356018 427204 356254
rect 426604 355934 427204 356018
rect 426604 355698 426786 355934
rect 427022 355698 427204 355934
rect 426604 320254 427204 355698
rect 426604 320018 426786 320254
rect 427022 320018 427204 320254
rect 426604 319934 427204 320018
rect 426604 319698 426786 319934
rect 427022 319698 427204 319934
rect 426604 284254 427204 319698
rect 426604 284018 426786 284254
rect 427022 284018 427204 284254
rect 426604 283934 427204 284018
rect 426604 283698 426786 283934
rect 427022 283698 427204 283934
rect 426604 248254 427204 283698
rect 426604 248018 426786 248254
rect 427022 248018 427204 248254
rect 426604 247934 427204 248018
rect 426604 247698 426786 247934
rect 427022 247698 427204 247934
rect 426604 212254 427204 247698
rect 426604 212018 426786 212254
rect 427022 212018 427204 212254
rect 426604 211934 427204 212018
rect 426604 211698 426786 211934
rect 427022 211698 427204 211934
rect 426604 176254 427204 211698
rect 426604 176018 426786 176254
rect 427022 176018 427204 176254
rect 426604 175934 427204 176018
rect 426604 175698 426786 175934
rect 427022 175698 427204 175934
rect 426604 140254 427204 175698
rect 426604 140018 426786 140254
rect 427022 140018 427204 140254
rect 426604 139934 427204 140018
rect 426604 139698 426786 139934
rect 427022 139698 427204 139934
rect 426604 104254 427204 139698
rect 426604 104018 426786 104254
rect 427022 104018 427204 104254
rect 426604 103934 427204 104018
rect 426604 103698 426786 103934
rect 427022 103698 427204 103934
rect 426604 68254 427204 103698
rect 426604 68018 426786 68254
rect 427022 68018 427204 68254
rect 426604 67934 427204 68018
rect 426604 67698 426786 67934
rect 427022 67698 427204 67934
rect 426604 32254 427204 67698
rect 426604 32018 426786 32254
rect 427022 32018 427204 32254
rect 426604 31934 427204 32018
rect 426604 31698 426786 31934
rect 427022 31698 427204 31934
rect 408604 -6222 408786 -5986
rect 409022 -6222 409204 -5986
rect 408604 -6306 409204 -6222
rect 408604 -6542 408786 -6306
rect 409022 -6542 409204 -6306
rect 408604 -7504 409204 -6542
rect 426604 -6926 427204 31698
rect 433804 704838 434404 705800
rect 433804 704602 433986 704838
rect 434222 704602 434404 704838
rect 433804 704518 434404 704602
rect 433804 704282 433986 704518
rect 434222 704282 434404 704518
rect 433804 687454 434404 704282
rect 433804 687218 433986 687454
rect 434222 687218 434404 687454
rect 433804 687134 434404 687218
rect 433804 686898 433986 687134
rect 434222 686898 434404 687134
rect 433804 651454 434404 686898
rect 433804 651218 433986 651454
rect 434222 651218 434404 651454
rect 433804 651134 434404 651218
rect 433804 650898 433986 651134
rect 434222 650898 434404 651134
rect 433804 615454 434404 650898
rect 433804 615218 433986 615454
rect 434222 615218 434404 615454
rect 433804 615134 434404 615218
rect 433804 614898 433986 615134
rect 434222 614898 434404 615134
rect 433804 579454 434404 614898
rect 433804 579218 433986 579454
rect 434222 579218 434404 579454
rect 433804 579134 434404 579218
rect 433804 578898 433986 579134
rect 434222 578898 434404 579134
rect 433804 543454 434404 578898
rect 433804 543218 433986 543454
rect 434222 543218 434404 543454
rect 433804 543134 434404 543218
rect 433804 542898 433986 543134
rect 434222 542898 434404 543134
rect 433804 507454 434404 542898
rect 433804 507218 433986 507454
rect 434222 507218 434404 507454
rect 433804 507134 434404 507218
rect 433804 506898 433986 507134
rect 434222 506898 434404 507134
rect 433804 471454 434404 506898
rect 433804 471218 433986 471454
rect 434222 471218 434404 471454
rect 433804 471134 434404 471218
rect 433804 470898 433986 471134
rect 434222 470898 434404 471134
rect 433804 435454 434404 470898
rect 433804 435218 433986 435454
rect 434222 435218 434404 435454
rect 433804 435134 434404 435218
rect 433804 434898 433986 435134
rect 434222 434898 434404 435134
rect 433804 399454 434404 434898
rect 433804 399218 433986 399454
rect 434222 399218 434404 399454
rect 433804 399134 434404 399218
rect 433804 398898 433986 399134
rect 434222 398898 434404 399134
rect 433804 363454 434404 398898
rect 433804 363218 433986 363454
rect 434222 363218 434404 363454
rect 433804 363134 434404 363218
rect 433804 362898 433986 363134
rect 434222 362898 434404 363134
rect 433804 327454 434404 362898
rect 433804 327218 433986 327454
rect 434222 327218 434404 327454
rect 433804 327134 434404 327218
rect 433804 326898 433986 327134
rect 434222 326898 434404 327134
rect 433804 291454 434404 326898
rect 433804 291218 433986 291454
rect 434222 291218 434404 291454
rect 433804 291134 434404 291218
rect 433804 290898 433986 291134
rect 434222 290898 434404 291134
rect 433804 255454 434404 290898
rect 433804 255218 433986 255454
rect 434222 255218 434404 255454
rect 433804 255134 434404 255218
rect 433804 254898 433986 255134
rect 434222 254898 434404 255134
rect 433804 219454 434404 254898
rect 433804 219218 433986 219454
rect 434222 219218 434404 219454
rect 433804 219134 434404 219218
rect 433804 218898 433986 219134
rect 434222 218898 434404 219134
rect 433804 183454 434404 218898
rect 433804 183218 433986 183454
rect 434222 183218 434404 183454
rect 433804 183134 434404 183218
rect 433804 182898 433986 183134
rect 434222 182898 434404 183134
rect 433804 147454 434404 182898
rect 433804 147218 433986 147454
rect 434222 147218 434404 147454
rect 433804 147134 434404 147218
rect 433804 146898 433986 147134
rect 434222 146898 434404 147134
rect 433804 111454 434404 146898
rect 433804 111218 433986 111454
rect 434222 111218 434404 111454
rect 433804 111134 434404 111218
rect 433804 110898 433986 111134
rect 434222 110898 434404 111134
rect 433804 75454 434404 110898
rect 433804 75218 433986 75454
rect 434222 75218 434404 75454
rect 433804 75134 434404 75218
rect 433804 74898 433986 75134
rect 434222 74898 434404 75134
rect 433804 39454 434404 74898
rect 433804 39218 433986 39454
rect 434222 39218 434404 39454
rect 433804 39134 434404 39218
rect 433804 38898 433986 39134
rect 434222 38898 434404 39134
rect 433804 3454 434404 38898
rect 433804 3218 433986 3454
rect 434222 3218 434404 3454
rect 433804 3134 434404 3218
rect 433804 2898 433986 3134
rect 434222 2898 434404 3134
rect 433804 -346 434404 2898
rect 433804 -582 433986 -346
rect 434222 -582 434404 -346
rect 433804 -666 434404 -582
rect 433804 -902 433986 -666
rect 434222 -902 434404 -666
rect 433804 -1864 434404 -902
rect 437404 691054 438004 706162
rect 437404 690818 437586 691054
rect 437822 690818 438004 691054
rect 437404 690734 438004 690818
rect 437404 690498 437586 690734
rect 437822 690498 438004 690734
rect 437404 655054 438004 690498
rect 437404 654818 437586 655054
rect 437822 654818 438004 655054
rect 437404 654734 438004 654818
rect 437404 654498 437586 654734
rect 437822 654498 438004 654734
rect 437404 619054 438004 654498
rect 437404 618818 437586 619054
rect 437822 618818 438004 619054
rect 437404 618734 438004 618818
rect 437404 618498 437586 618734
rect 437822 618498 438004 618734
rect 437404 583054 438004 618498
rect 437404 582818 437586 583054
rect 437822 582818 438004 583054
rect 437404 582734 438004 582818
rect 437404 582498 437586 582734
rect 437822 582498 438004 582734
rect 437404 547054 438004 582498
rect 437404 546818 437586 547054
rect 437822 546818 438004 547054
rect 437404 546734 438004 546818
rect 437404 546498 437586 546734
rect 437822 546498 438004 546734
rect 437404 511054 438004 546498
rect 437404 510818 437586 511054
rect 437822 510818 438004 511054
rect 437404 510734 438004 510818
rect 437404 510498 437586 510734
rect 437822 510498 438004 510734
rect 437404 475054 438004 510498
rect 437404 474818 437586 475054
rect 437822 474818 438004 475054
rect 437404 474734 438004 474818
rect 437404 474498 437586 474734
rect 437822 474498 438004 474734
rect 437404 439054 438004 474498
rect 437404 438818 437586 439054
rect 437822 438818 438004 439054
rect 437404 438734 438004 438818
rect 437404 438498 437586 438734
rect 437822 438498 438004 438734
rect 437404 403054 438004 438498
rect 437404 402818 437586 403054
rect 437822 402818 438004 403054
rect 437404 402734 438004 402818
rect 437404 402498 437586 402734
rect 437822 402498 438004 402734
rect 437404 367054 438004 402498
rect 437404 366818 437586 367054
rect 437822 366818 438004 367054
rect 437404 366734 438004 366818
rect 437404 366498 437586 366734
rect 437822 366498 438004 366734
rect 437404 331054 438004 366498
rect 437404 330818 437586 331054
rect 437822 330818 438004 331054
rect 437404 330734 438004 330818
rect 437404 330498 437586 330734
rect 437822 330498 438004 330734
rect 437404 295054 438004 330498
rect 437404 294818 437586 295054
rect 437822 294818 438004 295054
rect 437404 294734 438004 294818
rect 437404 294498 437586 294734
rect 437822 294498 438004 294734
rect 437404 259054 438004 294498
rect 437404 258818 437586 259054
rect 437822 258818 438004 259054
rect 437404 258734 438004 258818
rect 437404 258498 437586 258734
rect 437822 258498 438004 258734
rect 437404 223054 438004 258498
rect 437404 222818 437586 223054
rect 437822 222818 438004 223054
rect 437404 222734 438004 222818
rect 437404 222498 437586 222734
rect 437822 222498 438004 222734
rect 437404 187054 438004 222498
rect 437404 186818 437586 187054
rect 437822 186818 438004 187054
rect 437404 186734 438004 186818
rect 437404 186498 437586 186734
rect 437822 186498 438004 186734
rect 437404 151054 438004 186498
rect 437404 150818 437586 151054
rect 437822 150818 438004 151054
rect 437404 150734 438004 150818
rect 437404 150498 437586 150734
rect 437822 150498 438004 150734
rect 437404 115054 438004 150498
rect 437404 114818 437586 115054
rect 437822 114818 438004 115054
rect 437404 114734 438004 114818
rect 437404 114498 437586 114734
rect 437822 114498 438004 114734
rect 437404 79054 438004 114498
rect 437404 78818 437586 79054
rect 437822 78818 438004 79054
rect 437404 78734 438004 78818
rect 437404 78498 437586 78734
rect 437822 78498 438004 78734
rect 437404 43054 438004 78498
rect 437404 42818 437586 43054
rect 437822 42818 438004 43054
rect 437404 42734 438004 42818
rect 437404 42498 437586 42734
rect 437822 42498 438004 42734
rect 437404 7054 438004 42498
rect 437404 6818 437586 7054
rect 437822 6818 438004 7054
rect 437404 6734 438004 6818
rect 437404 6498 437586 6734
rect 437822 6498 438004 6734
rect 437404 -2226 438004 6498
rect 437404 -2462 437586 -2226
rect 437822 -2462 438004 -2226
rect 437404 -2546 438004 -2462
rect 437404 -2782 437586 -2546
rect 437822 -2782 438004 -2546
rect 437404 -3744 438004 -2782
rect 441004 694654 441604 708042
rect 441004 694418 441186 694654
rect 441422 694418 441604 694654
rect 441004 694334 441604 694418
rect 441004 694098 441186 694334
rect 441422 694098 441604 694334
rect 441004 658654 441604 694098
rect 441004 658418 441186 658654
rect 441422 658418 441604 658654
rect 441004 658334 441604 658418
rect 441004 658098 441186 658334
rect 441422 658098 441604 658334
rect 441004 622654 441604 658098
rect 441004 622418 441186 622654
rect 441422 622418 441604 622654
rect 441004 622334 441604 622418
rect 441004 622098 441186 622334
rect 441422 622098 441604 622334
rect 441004 586654 441604 622098
rect 441004 586418 441186 586654
rect 441422 586418 441604 586654
rect 441004 586334 441604 586418
rect 441004 586098 441186 586334
rect 441422 586098 441604 586334
rect 441004 550654 441604 586098
rect 441004 550418 441186 550654
rect 441422 550418 441604 550654
rect 441004 550334 441604 550418
rect 441004 550098 441186 550334
rect 441422 550098 441604 550334
rect 441004 514654 441604 550098
rect 441004 514418 441186 514654
rect 441422 514418 441604 514654
rect 441004 514334 441604 514418
rect 441004 514098 441186 514334
rect 441422 514098 441604 514334
rect 441004 478654 441604 514098
rect 441004 478418 441186 478654
rect 441422 478418 441604 478654
rect 441004 478334 441604 478418
rect 441004 478098 441186 478334
rect 441422 478098 441604 478334
rect 441004 442654 441604 478098
rect 441004 442418 441186 442654
rect 441422 442418 441604 442654
rect 441004 442334 441604 442418
rect 441004 442098 441186 442334
rect 441422 442098 441604 442334
rect 441004 406654 441604 442098
rect 441004 406418 441186 406654
rect 441422 406418 441604 406654
rect 441004 406334 441604 406418
rect 441004 406098 441186 406334
rect 441422 406098 441604 406334
rect 441004 370654 441604 406098
rect 441004 370418 441186 370654
rect 441422 370418 441604 370654
rect 441004 370334 441604 370418
rect 441004 370098 441186 370334
rect 441422 370098 441604 370334
rect 441004 334654 441604 370098
rect 441004 334418 441186 334654
rect 441422 334418 441604 334654
rect 441004 334334 441604 334418
rect 441004 334098 441186 334334
rect 441422 334098 441604 334334
rect 441004 298654 441604 334098
rect 441004 298418 441186 298654
rect 441422 298418 441604 298654
rect 441004 298334 441604 298418
rect 441004 298098 441186 298334
rect 441422 298098 441604 298334
rect 441004 262654 441604 298098
rect 441004 262418 441186 262654
rect 441422 262418 441604 262654
rect 441004 262334 441604 262418
rect 441004 262098 441186 262334
rect 441422 262098 441604 262334
rect 441004 226654 441604 262098
rect 441004 226418 441186 226654
rect 441422 226418 441604 226654
rect 441004 226334 441604 226418
rect 441004 226098 441186 226334
rect 441422 226098 441604 226334
rect 441004 190654 441604 226098
rect 441004 190418 441186 190654
rect 441422 190418 441604 190654
rect 441004 190334 441604 190418
rect 441004 190098 441186 190334
rect 441422 190098 441604 190334
rect 441004 154654 441604 190098
rect 441004 154418 441186 154654
rect 441422 154418 441604 154654
rect 441004 154334 441604 154418
rect 441004 154098 441186 154334
rect 441422 154098 441604 154334
rect 441004 118654 441604 154098
rect 441004 118418 441186 118654
rect 441422 118418 441604 118654
rect 441004 118334 441604 118418
rect 441004 118098 441186 118334
rect 441422 118098 441604 118334
rect 441004 82654 441604 118098
rect 441004 82418 441186 82654
rect 441422 82418 441604 82654
rect 441004 82334 441604 82418
rect 441004 82098 441186 82334
rect 441422 82098 441604 82334
rect 441004 46654 441604 82098
rect 441004 46418 441186 46654
rect 441422 46418 441604 46654
rect 441004 46334 441604 46418
rect 441004 46098 441186 46334
rect 441422 46098 441604 46334
rect 441004 10654 441604 46098
rect 441004 10418 441186 10654
rect 441422 10418 441604 10654
rect 441004 10334 441604 10418
rect 441004 10098 441186 10334
rect 441422 10098 441604 10334
rect 441004 -4106 441604 10098
rect 441004 -4342 441186 -4106
rect 441422 -4342 441604 -4106
rect 441004 -4426 441604 -4342
rect 441004 -4662 441186 -4426
rect 441422 -4662 441604 -4426
rect 441004 -5624 441604 -4662
rect 444604 698254 445204 709922
rect 462604 711418 463204 711440
rect 462604 711182 462786 711418
rect 463022 711182 463204 711418
rect 462604 711098 463204 711182
rect 462604 710862 462786 711098
rect 463022 710862 463204 711098
rect 459004 709538 459604 709560
rect 459004 709302 459186 709538
rect 459422 709302 459604 709538
rect 459004 709218 459604 709302
rect 459004 708982 459186 709218
rect 459422 708982 459604 709218
rect 455404 707658 456004 707680
rect 455404 707422 455586 707658
rect 455822 707422 456004 707658
rect 455404 707338 456004 707422
rect 455404 707102 455586 707338
rect 455822 707102 456004 707338
rect 444604 698018 444786 698254
rect 445022 698018 445204 698254
rect 444604 697934 445204 698018
rect 444604 697698 444786 697934
rect 445022 697698 445204 697934
rect 444604 662254 445204 697698
rect 444604 662018 444786 662254
rect 445022 662018 445204 662254
rect 444604 661934 445204 662018
rect 444604 661698 444786 661934
rect 445022 661698 445204 661934
rect 444604 626254 445204 661698
rect 444604 626018 444786 626254
rect 445022 626018 445204 626254
rect 444604 625934 445204 626018
rect 444604 625698 444786 625934
rect 445022 625698 445204 625934
rect 444604 590254 445204 625698
rect 444604 590018 444786 590254
rect 445022 590018 445204 590254
rect 444604 589934 445204 590018
rect 444604 589698 444786 589934
rect 445022 589698 445204 589934
rect 444604 554254 445204 589698
rect 444604 554018 444786 554254
rect 445022 554018 445204 554254
rect 444604 553934 445204 554018
rect 444604 553698 444786 553934
rect 445022 553698 445204 553934
rect 444604 518254 445204 553698
rect 444604 518018 444786 518254
rect 445022 518018 445204 518254
rect 444604 517934 445204 518018
rect 444604 517698 444786 517934
rect 445022 517698 445204 517934
rect 444604 482254 445204 517698
rect 444604 482018 444786 482254
rect 445022 482018 445204 482254
rect 444604 481934 445204 482018
rect 444604 481698 444786 481934
rect 445022 481698 445204 481934
rect 444604 446254 445204 481698
rect 444604 446018 444786 446254
rect 445022 446018 445204 446254
rect 444604 445934 445204 446018
rect 444604 445698 444786 445934
rect 445022 445698 445204 445934
rect 444604 410254 445204 445698
rect 444604 410018 444786 410254
rect 445022 410018 445204 410254
rect 444604 409934 445204 410018
rect 444604 409698 444786 409934
rect 445022 409698 445204 409934
rect 444604 374254 445204 409698
rect 444604 374018 444786 374254
rect 445022 374018 445204 374254
rect 444604 373934 445204 374018
rect 444604 373698 444786 373934
rect 445022 373698 445204 373934
rect 444604 338254 445204 373698
rect 444604 338018 444786 338254
rect 445022 338018 445204 338254
rect 444604 337934 445204 338018
rect 444604 337698 444786 337934
rect 445022 337698 445204 337934
rect 444604 302254 445204 337698
rect 444604 302018 444786 302254
rect 445022 302018 445204 302254
rect 444604 301934 445204 302018
rect 444604 301698 444786 301934
rect 445022 301698 445204 301934
rect 444604 266254 445204 301698
rect 444604 266018 444786 266254
rect 445022 266018 445204 266254
rect 444604 265934 445204 266018
rect 444604 265698 444786 265934
rect 445022 265698 445204 265934
rect 444604 230254 445204 265698
rect 444604 230018 444786 230254
rect 445022 230018 445204 230254
rect 444604 229934 445204 230018
rect 444604 229698 444786 229934
rect 445022 229698 445204 229934
rect 444604 194254 445204 229698
rect 444604 194018 444786 194254
rect 445022 194018 445204 194254
rect 444604 193934 445204 194018
rect 444604 193698 444786 193934
rect 445022 193698 445204 193934
rect 444604 158254 445204 193698
rect 444604 158018 444786 158254
rect 445022 158018 445204 158254
rect 444604 157934 445204 158018
rect 444604 157698 444786 157934
rect 445022 157698 445204 157934
rect 444604 122254 445204 157698
rect 444604 122018 444786 122254
rect 445022 122018 445204 122254
rect 444604 121934 445204 122018
rect 444604 121698 444786 121934
rect 445022 121698 445204 121934
rect 444604 86254 445204 121698
rect 444604 86018 444786 86254
rect 445022 86018 445204 86254
rect 444604 85934 445204 86018
rect 444604 85698 444786 85934
rect 445022 85698 445204 85934
rect 444604 50254 445204 85698
rect 444604 50018 444786 50254
rect 445022 50018 445204 50254
rect 444604 49934 445204 50018
rect 444604 49698 444786 49934
rect 445022 49698 445204 49934
rect 444604 14254 445204 49698
rect 444604 14018 444786 14254
rect 445022 14018 445204 14254
rect 444604 13934 445204 14018
rect 444604 13698 444786 13934
rect 445022 13698 445204 13934
rect 426604 -7162 426786 -6926
rect 427022 -7162 427204 -6926
rect 426604 -7246 427204 -7162
rect 426604 -7482 426786 -7246
rect 427022 -7482 427204 -7246
rect 426604 -7504 427204 -7482
rect 444604 -5986 445204 13698
rect 451804 705778 452404 705800
rect 451804 705542 451986 705778
rect 452222 705542 452404 705778
rect 451804 705458 452404 705542
rect 451804 705222 451986 705458
rect 452222 705222 452404 705458
rect 451804 669454 452404 705222
rect 451804 669218 451986 669454
rect 452222 669218 452404 669454
rect 451804 669134 452404 669218
rect 451804 668898 451986 669134
rect 452222 668898 452404 669134
rect 451804 633454 452404 668898
rect 451804 633218 451986 633454
rect 452222 633218 452404 633454
rect 451804 633134 452404 633218
rect 451804 632898 451986 633134
rect 452222 632898 452404 633134
rect 451804 597454 452404 632898
rect 451804 597218 451986 597454
rect 452222 597218 452404 597454
rect 451804 597134 452404 597218
rect 451804 596898 451986 597134
rect 452222 596898 452404 597134
rect 451804 561454 452404 596898
rect 451804 561218 451986 561454
rect 452222 561218 452404 561454
rect 451804 561134 452404 561218
rect 451804 560898 451986 561134
rect 452222 560898 452404 561134
rect 451804 525454 452404 560898
rect 451804 525218 451986 525454
rect 452222 525218 452404 525454
rect 451804 525134 452404 525218
rect 451804 524898 451986 525134
rect 452222 524898 452404 525134
rect 451804 489454 452404 524898
rect 451804 489218 451986 489454
rect 452222 489218 452404 489454
rect 451804 489134 452404 489218
rect 451804 488898 451986 489134
rect 452222 488898 452404 489134
rect 451804 453454 452404 488898
rect 451804 453218 451986 453454
rect 452222 453218 452404 453454
rect 451804 453134 452404 453218
rect 451804 452898 451986 453134
rect 452222 452898 452404 453134
rect 451804 417454 452404 452898
rect 451804 417218 451986 417454
rect 452222 417218 452404 417454
rect 451804 417134 452404 417218
rect 451804 416898 451986 417134
rect 452222 416898 452404 417134
rect 451804 381454 452404 416898
rect 451804 381218 451986 381454
rect 452222 381218 452404 381454
rect 451804 381134 452404 381218
rect 451804 380898 451986 381134
rect 452222 380898 452404 381134
rect 451804 345454 452404 380898
rect 451804 345218 451986 345454
rect 452222 345218 452404 345454
rect 451804 345134 452404 345218
rect 451804 344898 451986 345134
rect 452222 344898 452404 345134
rect 451804 309454 452404 344898
rect 451804 309218 451986 309454
rect 452222 309218 452404 309454
rect 451804 309134 452404 309218
rect 451804 308898 451986 309134
rect 452222 308898 452404 309134
rect 451804 273454 452404 308898
rect 451804 273218 451986 273454
rect 452222 273218 452404 273454
rect 451804 273134 452404 273218
rect 451804 272898 451986 273134
rect 452222 272898 452404 273134
rect 451804 237454 452404 272898
rect 451804 237218 451986 237454
rect 452222 237218 452404 237454
rect 451804 237134 452404 237218
rect 451804 236898 451986 237134
rect 452222 236898 452404 237134
rect 451804 201454 452404 236898
rect 451804 201218 451986 201454
rect 452222 201218 452404 201454
rect 451804 201134 452404 201218
rect 451804 200898 451986 201134
rect 452222 200898 452404 201134
rect 451804 165454 452404 200898
rect 451804 165218 451986 165454
rect 452222 165218 452404 165454
rect 451804 165134 452404 165218
rect 451804 164898 451986 165134
rect 452222 164898 452404 165134
rect 451804 129454 452404 164898
rect 451804 129218 451986 129454
rect 452222 129218 452404 129454
rect 451804 129134 452404 129218
rect 451804 128898 451986 129134
rect 452222 128898 452404 129134
rect 451804 93454 452404 128898
rect 451804 93218 451986 93454
rect 452222 93218 452404 93454
rect 451804 93134 452404 93218
rect 451804 92898 451986 93134
rect 452222 92898 452404 93134
rect 451804 57454 452404 92898
rect 451804 57218 451986 57454
rect 452222 57218 452404 57454
rect 451804 57134 452404 57218
rect 451804 56898 451986 57134
rect 452222 56898 452404 57134
rect 451804 21454 452404 56898
rect 451804 21218 451986 21454
rect 452222 21218 452404 21454
rect 451804 21134 452404 21218
rect 451804 20898 451986 21134
rect 452222 20898 452404 21134
rect 451804 -1286 452404 20898
rect 451804 -1522 451986 -1286
rect 452222 -1522 452404 -1286
rect 451804 -1606 452404 -1522
rect 451804 -1842 451986 -1606
rect 452222 -1842 452404 -1606
rect 451804 -1864 452404 -1842
rect 455404 673054 456004 707102
rect 455404 672818 455586 673054
rect 455822 672818 456004 673054
rect 455404 672734 456004 672818
rect 455404 672498 455586 672734
rect 455822 672498 456004 672734
rect 455404 637054 456004 672498
rect 455404 636818 455586 637054
rect 455822 636818 456004 637054
rect 455404 636734 456004 636818
rect 455404 636498 455586 636734
rect 455822 636498 456004 636734
rect 455404 601054 456004 636498
rect 455404 600818 455586 601054
rect 455822 600818 456004 601054
rect 455404 600734 456004 600818
rect 455404 600498 455586 600734
rect 455822 600498 456004 600734
rect 455404 565054 456004 600498
rect 455404 564818 455586 565054
rect 455822 564818 456004 565054
rect 455404 564734 456004 564818
rect 455404 564498 455586 564734
rect 455822 564498 456004 564734
rect 455404 529054 456004 564498
rect 455404 528818 455586 529054
rect 455822 528818 456004 529054
rect 455404 528734 456004 528818
rect 455404 528498 455586 528734
rect 455822 528498 456004 528734
rect 455404 493054 456004 528498
rect 455404 492818 455586 493054
rect 455822 492818 456004 493054
rect 455404 492734 456004 492818
rect 455404 492498 455586 492734
rect 455822 492498 456004 492734
rect 455404 457054 456004 492498
rect 455404 456818 455586 457054
rect 455822 456818 456004 457054
rect 455404 456734 456004 456818
rect 455404 456498 455586 456734
rect 455822 456498 456004 456734
rect 455404 421054 456004 456498
rect 455404 420818 455586 421054
rect 455822 420818 456004 421054
rect 455404 420734 456004 420818
rect 455404 420498 455586 420734
rect 455822 420498 456004 420734
rect 455404 385054 456004 420498
rect 455404 384818 455586 385054
rect 455822 384818 456004 385054
rect 455404 384734 456004 384818
rect 455404 384498 455586 384734
rect 455822 384498 456004 384734
rect 455404 349054 456004 384498
rect 455404 348818 455586 349054
rect 455822 348818 456004 349054
rect 455404 348734 456004 348818
rect 455404 348498 455586 348734
rect 455822 348498 456004 348734
rect 455404 313054 456004 348498
rect 455404 312818 455586 313054
rect 455822 312818 456004 313054
rect 455404 312734 456004 312818
rect 455404 312498 455586 312734
rect 455822 312498 456004 312734
rect 455404 277054 456004 312498
rect 455404 276818 455586 277054
rect 455822 276818 456004 277054
rect 455404 276734 456004 276818
rect 455404 276498 455586 276734
rect 455822 276498 456004 276734
rect 455404 241054 456004 276498
rect 455404 240818 455586 241054
rect 455822 240818 456004 241054
rect 455404 240734 456004 240818
rect 455404 240498 455586 240734
rect 455822 240498 456004 240734
rect 455404 205054 456004 240498
rect 455404 204818 455586 205054
rect 455822 204818 456004 205054
rect 455404 204734 456004 204818
rect 455404 204498 455586 204734
rect 455822 204498 456004 204734
rect 455404 169054 456004 204498
rect 455404 168818 455586 169054
rect 455822 168818 456004 169054
rect 455404 168734 456004 168818
rect 455404 168498 455586 168734
rect 455822 168498 456004 168734
rect 455404 133054 456004 168498
rect 455404 132818 455586 133054
rect 455822 132818 456004 133054
rect 455404 132734 456004 132818
rect 455404 132498 455586 132734
rect 455822 132498 456004 132734
rect 455404 97054 456004 132498
rect 455404 96818 455586 97054
rect 455822 96818 456004 97054
rect 455404 96734 456004 96818
rect 455404 96498 455586 96734
rect 455822 96498 456004 96734
rect 455404 61054 456004 96498
rect 455404 60818 455586 61054
rect 455822 60818 456004 61054
rect 455404 60734 456004 60818
rect 455404 60498 455586 60734
rect 455822 60498 456004 60734
rect 455404 25054 456004 60498
rect 455404 24818 455586 25054
rect 455822 24818 456004 25054
rect 455404 24734 456004 24818
rect 455404 24498 455586 24734
rect 455822 24498 456004 24734
rect 455404 -3166 456004 24498
rect 455404 -3402 455586 -3166
rect 455822 -3402 456004 -3166
rect 455404 -3486 456004 -3402
rect 455404 -3722 455586 -3486
rect 455822 -3722 456004 -3486
rect 455404 -3744 456004 -3722
rect 459004 676654 459604 708982
rect 459004 676418 459186 676654
rect 459422 676418 459604 676654
rect 459004 676334 459604 676418
rect 459004 676098 459186 676334
rect 459422 676098 459604 676334
rect 459004 640654 459604 676098
rect 459004 640418 459186 640654
rect 459422 640418 459604 640654
rect 459004 640334 459604 640418
rect 459004 640098 459186 640334
rect 459422 640098 459604 640334
rect 459004 604654 459604 640098
rect 459004 604418 459186 604654
rect 459422 604418 459604 604654
rect 459004 604334 459604 604418
rect 459004 604098 459186 604334
rect 459422 604098 459604 604334
rect 459004 568654 459604 604098
rect 459004 568418 459186 568654
rect 459422 568418 459604 568654
rect 459004 568334 459604 568418
rect 459004 568098 459186 568334
rect 459422 568098 459604 568334
rect 459004 532654 459604 568098
rect 459004 532418 459186 532654
rect 459422 532418 459604 532654
rect 459004 532334 459604 532418
rect 459004 532098 459186 532334
rect 459422 532098 459604 532334
rect 459004 496654 459604 532098
rect 459004 496418 459186 496654
rect 459422 496418 459604 496654
rect 459004 496334 459604 496418
rect 459004 496098 459186 496334
rect 459422 496098 459604 496334
rect 459004 460654 459604 496098
rect 459004 460418 459186 460654
rect 459422 460418 459604 460654
rect 459004 460334 459604 460418
rect 459004 460098 459186 460334
rect 459422 460098 459604 460334
rect 459004 424654 459604 460098
rect 459004 424418 459186 424654
rect 459422 424418 459604 424654
rect 459004 424334 459604 424418
rect 459004 424098 459186 424334
rect 459422 424098 459604 424334
rect 459004 388654 459604 424098
rect 459004 388418 459186 388654
rect 459422 388418 459604 388654
rect 459004 388334 459604 388418
rect 459004 388098 459186 388334
rect 459422 388098 459604 388334
rect 459004 352654 459604 388098
rect 459004 352418 459186 352654
rect 459422 352418 459604 352654
rect 459004 352334 459604 352418
rect 459004 352098 459186 352334
rect 459422 352098 459604 352334
rect 459004 316654 459604 352098
rect 459004 316418 459186 316654
rect 459422 316418 459604 316654
rect 459004 316334 459604 316418
rect 459004 316098 459186 316334
rect 459422 316098 459604 316334
rect 459004 280654 459604 316098
rect 459004 280418 459186 280654
rect 459422 280418 459604 280654
rect 459004 280334 459604 280418
rect 459004 280098 459186 280334
rect 459422 280098 459604 280334
rect 459004 244654 459604 280098
rect 459004 244418 459186 244654
rect 459422 244418 459604 244654
rect 459004 244334 459604 244418
rect 459004 244098 459186 244334
rect 459422 244098 459604 244334
rect 459004 208654 459604 244098
rect 459004 208418 459186 208654
rect 459422 208418 459604 208654
rect 459004 208334 459604 208418
rect 459004 208098 459186 208334
rect 459422 208098 459604 208334
rect 459004 172654 459604 208098
rect 459004 172418 459186 172654
rect 459422 172418 459604 172654
rect 459004 172334 459604 172418
rect 459004 172098 459186 172334
rect 459422 172098 459604 172334
rect 459004 136654 459604 172098
rect 459004 136418 459186 136654
rect 459422 136418 459604 136654
rect 459004 136334 459604 136418
rect 459004 136098 459186 136334
rect 459422 136098 459604 136334
rect 459004 100654 459604 136098
rect 459004 100418 459186 100654
rect 459422 100418 459604 100654
rect 459004 100334 459604 100418
rect 459004 100098 459186 100334
rect 459422 100098 459604 100334
rect 459004 64654 459604 100098
rect 459004 64418 459186 64654
rect 459422 64418 459604 64654
rect 459004 64334 459604 64418
rect 459004 64098 459186 64334
rect 459422 64098 459604 64334
rect 459004 28654 459604 64098
rect 459004 28418 459186 28654
rect 459422 28418 459604 28654
rect 459004 28334 459604 28418
rect 459004 28098 459186 28334
rect 459422 28098 459604 28334
rect 459004 -5046 459604 28098
rect 459004 -5282 459186 -5046
rect 459422 -5282 459604 -5046
rect 459004 -5366 459604 -5282
rect 459004 -5602 459186 -5366
rect 459422 -5602 459604 -5366
rect 459004 -5624 459604 -5602
rect 462604 680254 463204 710862
rect 480604 710478 481204 711440
rect 480604 710242 480786 710478
rect 481022 710242 481204 710478
rect 480604 710158 481204 710242
rect 480604 709922 480786 710158
rect 481022 709922 481204 710158
rect 477004 708598 477604 709560
rect 477004 708362 477186 708598
rect 477422 708362 477604 708598
rect 477004 708278 477604 708362
rect 477004 708042 477186 708278
rect 477422 708042 477604 708278
rect 473404 706718 474004 707680
rect 473404 706482 473586 706718
rect 473822 706482 474004 706718
rect 473404 706398 474004 706482
rect 473404 706162 473586 706398
rect 473822 706162 474004 706398
rect 462604 680018 462786 680254
rect 463022 680018 463204 680254
rect 462604 679934 463204 680018
rect 462604 679698 462786 679934
rect 463022 679698 463204 679934
rect 462604 644254 463204 679698
rect 462604 644018 462786 644254
rect 463022 644018 463204 644254
rect 462604 643934 463204 644018
rect 462604 643698 462786 643934
rect 463022 643698 463204 643934
rect 462604 608254 463204 643698
rect 462604 608018 462786 608254
rect 463022 608018 463204 608254
rect 462604 607934 463204 608018
rect 462604 607698 462786 607934
rect 463022 607698 463204 607934
rect 462604 572254 463204 607698
rect 462604 572018 462786 572254
rect 463022 572018 463204 572254
rect 462604 571934 463204 572018
rect 462604 571698 462786 571934
rect 463022 571698 463204 571934
rect 462604 536254 463204 571698
rect 462604 536018 462786 536254
rect 463022 536018 463204 536254
rect 462604 535934 463204 536018
rect 462604 535698 462786 535934
rect 463022 535698 463204 535934
rect 462604 500254 463204 535698
rect 462604 500018 462786 500254
rect 463022 500018 463204 500254
rect 462604 499934 463204 500018
rect 462604 499698 462786 499934
rect 463022 499698 463204 499934
rect 462604 464254 463204 499698
rect 462604 464018 462786 464254
rect 463022 464018 463204 464254
rect 462604 463934 463204 464018
rect 462604 463698 462786 463934
rect 463022 463698 463204 463934
rect 462604 428254 463204 463698
rect 462604 428018 462786 428254
rect 463022 428018 463204 428254
rect 462604 427934 463204 428018
rect 462604 427698 462786 427934
rect 463022 427698 463204 427934
rect 462604 392254 463204 427698
rect 462604 392018 462786 392254
rect 463022 392018 463204 392254
rect 462604 391934 463204 392018
rect 462604 391698 462786 391934
rect 463022 391698 463204 391934
rect 462604 356254 463204 391698
rect 462604 356018 462786 356254
rect 463022 356018 463204 356254
rect 462604 355934 463204 356018
rect 462604 355698 462786 355934
rect 463022 355698 463204 355934
rect 462604 320254 463204 355698
rect 462604 320018 462786 320254
rect 463022 320018 463204 320254
rect 462604 319934 463204 320018
rect 462604 319698 462786 319934
rect 463022 319698 463204 319934
rect 462604 284254 463204 319698
rect 462604 284018 462786 284254
rect 463022 284018 463204 284254
rect 462604 283934 463204 284018
rect 462604 283698 462786 283934
rect 463022 283698 463204 283934
rect 462604 248254 463204 283698
rect 462604 248018 462786 248254
rect 463022 248018 463204 248254
rect 462604 247934 463204 248018
rect 462604 247698 462786 247934
rect 463022 247698 463204 247934
rect 462604 212254 463204 247698
rect 462604 212018 462786 212254
rect 463022 212018 463204 212254
rect 462604 211934 463204 212018
rect 462604 211698 462786 211934
rect 463022 211698 463204 211934
rect 462604 176254 463204 211698
rect 462604 176018 462786 176254
rect 463022 176018 463204 176254
rect 462604 175934 463204 176018
rect 462604 175698 462786 175934
rect 463022 175698 463204 175934
rect 462604 140254 463204 175698
rect 462604 140018 462786 140254
rect 463022 140018 463204 140254
rect 462604 139934 463204 140018
rect 462604 139698 462786 139934
rect 463022 139698 463204 139934
rect 462604 104254 463204 139698
rect 462604 104018 462786 104254
rect 463022 104018 463204 104254
rect 462604 103934 463204 104018
rect 462604 103698 462786 103934
rect 463022 103698 463204 103934
rect 462604 68254 463204 103698
rect 462604 68018 462786 68254
rect 463022 68018 463204 68254
rect 462604 67934 463204 68018
rect 462604 67698 462786 67934
rect 463022 67698 463204 67934
rect 462604 32254 463204 67698
rect 462604 32018 462786 32254
rect 463022 32018 463204 32254
rect 462604 31934 463204 32018
rect 462604 31698 462786 31934
rect 463022 31698 463204 31934
rect 444604 -6222 444786 -5986
rect 445022 -6222 445204 -5986
rect 444604 -6306 445204 -6222
rect 444604 -6542 444786 -6306
rect 445022 -6542 445204 -6306
rect 444604 -7504 445204 -6542
rect 462604 -6926 463204 31698
rect 469804 704838 470404 705800
rect 469804 704602 469986 704838
rect 470222 704602 470404 704838
rect 469804 704518 470404 704602
rect 469804 704282 469986 704518
rect 470222 704282 470404 704518
rect 469804 687454 470404 704282
rect 469804 687218 469986 687454
rect 470222 687218 470404 687454
rect 469804 687134 470404 687218
rect 469804 686898 469986 687134
rect 470222 686898 470404 687134
rect 469804 651454 470404 686898
rect 469804 651218 469986 651454
rect 470222 651218 470404 651454
rect 469804 651134 470404 651218
rect 469804 650898 469986 651134
rect 470222 650898 470404 651134
rect 469804 615454 470404 650898
rect 469804 615218 469986 615454
rect 470222 615218 470404 615454
rect 469804 615134 470404 615218
rect 469804 614898 469986 615134
rect 470222 614898 470404 615134
rect 469804 579454 470404 614898
rect 469804 579218 469986 579454
rect 470222 579218 470404 579454
rect 469804 579134 470404 579218
rect 469804 578898 469986 579134
rect 470222 578898 470404 579134
rect 469804 543454 470404 578898
rect 469804 543218 469986 543454
rect 470222 543218 470404 543454
rect 469804 543134 470404 543218
rect 469804 542898 469986 543134
rect 470222 542898 470404 543134
rect 469804 507454 470404 542898
rect 469804 507218 469986 507454
rect 470222 507218 470404 507454
rect 469804 507134 470404 507218
rect 469804 506898 469986 507134
rect 470222 506898 470404 507134
rect 469804 471454 470404 506898
rect 469804 471218 469986 471454
rect 470222 471218 470404 471454
rect 469804 471134 470404 471218
rect 469804 470898 469986 471134
rect 470222 470898 470404 471134
rect 469804 435454 470404 470898
rect 469804 435218 469986 435454
rect 470222 435218 470404 435454
rect 469804 435134 470404 435218
rect 469804 434898 469986 435134
rect 470222 434898 470404 435134
rect 469804 399454 470404 434898
rect 469804 399218 469986 399454
rect 470222 399218 470404 399454
rect 469804 399134 470404 399218
rect 469804 398898 469986 399134
rect 470222 398898 470404 399134
rect 469804 363454 470404 398898
rect 469804 363218 469986 363454
rect 470222 363218 470404 363454
rect 469804 363134 470404 363218
rect 469804 362898 469986 363134
rect 470222 362898 470404 363134
rect 469804 327454 470404 362898
rect 469804 327218 469986 327454
rect 470222 327218 470404 327454
rect 469804 327134 470404 327218
rect 469804 326898 469986 327134
rect 470222 326898 470404 327134
rect 469804 291454 470404 326898
rect 469804 291218 469986 291454
rect 470222 291218 470404 291454
rect 469804 291134 470404 291218
rect 469804 290898 469986 291134
rect 470222 290898 470404 291134
rect 469804 255454 470404 290898
rect 469804 255218 469986 255454
rect 470222 255218 470404 255454
rect 469804 255134 470404 255218
rect 469804 254898 469986 255134
rect 470222 254898 470404 255134
rect 469804 219454 470404 254898
rect 469804 219218 469986 219454
rect 470222 219218 470404 219454
rect 469804 219134 470404 219218
rect 469804 218898 469986 219134
rect 470222 218898 470404 219134
rect 469804 183454 470404 218898
rect 469804 183218 469986 183454
rect 470222 183218 470404 183454
rect 469804 183134 470404 183218
rect 469804 182898 469986 183134
rect 470222 182898 470404 183134
rect 469804 147454 470404 182898
rect 469804 147218 469986 147454
rect 470222 147218 470404 147454
rect 469804 147134 470404 147218
rect 469804 146898 469986 147134
rect 470222 146898 470404 147134
rect 469804 111454 470404 146898
rect 469804 111218 469986 111454
rect 470222 111218 470404 111454
rect 469804 111134 470404 111218
rect 469804 110898 469986 111134
rect 470222 110898 470404 111134
rect 469804 75454 470404 110898
rect 469804 75218 469986 75454
rect 470222 75218 470404 75454
rect 469804 75134 470404 75218
rect 469804 74898 469986 75134
rect 470222 74898 470404 75134
rect 469804 39454 470404 74898
rect 469804 39218 469986 39454
rect 470222 39218 470404 39454
rect 469804 39134 470404 39218
rect 469804 38898 469986 39134
rect 470222 38898 470404 39134
rect 469804 3454 470404 38898
rect 469804 3218 469986 3454
rect 470222 3218 470404 3454
rect 469804 3134 470404 3218
rect 469804 2898 469986 3134
rect 470222 2898 470404 3134
rect 469804 -346 470404 2898
rect 469804 -582 469986 -346
rect 470222 -582 470404 -346
rect 469804 -666 470404 -582
rect 469804 -902 469986 -666
rect 470222 -902 470404 -666
rect 469804 -1864 470404 -902
rect 473404 691054 474004 706162
rect 473404 690818 473586 691054
rect 473822 690818 474004 691054
rect 473404 690734 474004 690818
rect 473404 690498 473586 690734
rect 473822 690498 474004 690734
rect 473404 655054 474004 690498
rect 473404 654818 473586 655054
rect 473822 654818 474004 655054
rect 473404 654734 474004 654818
rect 473404 654498 473586 654734
rect 473822 654498 474004 654734
rect 473404 619054 474004 654498
rect 473404 618818 473586 619054
rect 473822 618818 474004 619054
rect 473404 618734 474004 618818
rect 473404 618498 473586 618734
rect 473822 618498 474004 618734
rect 473404 583054 474004 618498
rect 473404 582818 473586 583054
rect 473822 582818 474004 583054
rect 473404 582734 474004 582818
rect 473404 582498 473586 582734
rect 473822 582498 474004 582734
rect 473404 547054 474004 582498
rect 473404 546818 473586 547054
rect 473822 546818 474004 547054
rect 473404 546734 474004 546818
rect 473404 546498 473586 546734
rect 473822 546498 474004 546734
rect 473404 511054 474004 546498
rect 473404 510818 473586 511054
rect 473822 510818 474004 511054
rect 473404 510734 474004 510818
rect 473404 510498 473586 510734
rect 473822 510498 474004 510734
rect 473404 475054 474004 510498
rect 473404 474818 473586 475054
rect 473822 474818 474004 475054
rect 473404 474734 474004 474818
rect 473404 474498 473586 474734
rect 473822 474498 474004 474734
rect 473404 439054 474004 474498
rect 473404 438818 473586 439054
rect 473822 438818 474004 439054
rect 473404 438734 474004 438818
rect 473404 438498 473586 438734
rect 473822 438498 474004 438734
rect 473404 403054 474004 438498
rect 473404 402818 473586 403054
rect 473822 402818 474004 403054
rect 473404 402734 474004 402818
rect 473404 402498 473586 402734
rect 473822 402498 474004 402734
rect 473404 367054 474004 402498
rect 473404 366818 473586 367054
rect 473822 366818 474004 367054
rect 473404 366734 474004 366818
rect 473404 366498 473586 366734
rect 473822 366498 474004 366734
rect 473404 331054 474004 366498
rect 473404 330818 473586 331054
rect 473822 330818 474004 331054
rect 473404 330734 474004 330818
rect 473404 330498 473586 330734
rect 473822 330498 474004 330734
rect 473404 295054 474004 330498
rect 473404 294818 473586 295054
rect 473822 294818 474004 295054
rect 473404 294734 474004 294818
rect 473404 294498 473586 294734
rect 473822 294498 474004 294734
rect 473404 259054 474004 294498
rect 473404 258818 473586 259054
rect 473822 258818 474004 259054
rect 473404 258734 474004 258818
rect 473404 258498 473586 258734
rect 473822 258498 474004 258734
rect 473404 223054 474004 258498
rect 473404 222818 473586 223054
rect 473822 222818 474004 223054
rect 473404 222734 474004 222818
rect 473404 222498 473586 222734
rect 473822 222498 474004 222734
rect 473404 187054 474004 222498
rect 473404 186818 473586 187054
rect 473822 186818 474004 187054
rect 473404 186734 474004 186818
rect 473404 186498 473586 186734
rect 473822 186498 474004 186734
rect 473404 151054 474004 186498
rect 473404 150818 473586 151054
rect 473822 150818 474004 151054
rect 473404 150734 474004 150818
rect 473404 150498 473586 150734
rect 473822 150498 474004 150734
rect 473404 115054 474004 150498
rect 473404 114818 473586 115054
rect 473822 114818 474004 115054
rect 473404 114734 474004 114818
rect 473404 114498 473586 114734
rect 473822 114498 474004 114734
rect 473404 79054 474004 114498
rect 473404 78818 473586 79054
rect 473822 78818 474004 79054
rect 473404 78734 474004 78818
rect 473404 78498 473586 78734
rect 473822 78498 474004 78734
rect 473404 43054 474004 78498
rect 473404 42818 473586 43054
rect 473822 42818 474004 43054
rect 473404 42734 474004 42818
rect 473404 42498 473586 42734
rect 473822 42498 474004 42734
rect 473404 7054 474004 42498
rect 473404 6818 473586 7054
rect 473822 6818 474004 7054
rect 473404 6734 474004 6818
rect 473404 6498 473586 6734
rect 473822 6498 474004 6734
rect 473404 -2226 474004 6498
rect 473404 -2462 473586 -2226
rect 473822 -2462 474004 -2226
rect 473404 -2546 474004 -2462
rect 473404 -2782 473586 -2546
rect 473822 -2782 474004 -2546
rect 473404 -3744 474004 -2782
rect 477004 694654 477604 708042
rect 477004 694418 477186 694654
rect 477422 694418 477604 694654
rect 477004 694334 477604 694418
rect 477004 694098 477186 694334
rect 477422 694098 477604 694334
rect 477004 658654 477604 694098
rect 477004 658418 477186 658654
rect 477422 658418 477604 658654
rect 477004 658334 477604 658418
rect 477004 658098 477186 658334
rect 477422 658098 477604 658334
rect 477004 622654 477604 658098
rect 477004 622418 477186 622654
rect 477422 622418 477604 622654
rect 477004 622334 477604 622418
rect 477004 622098 477186 622334
rect 477422 622098 477604 622334
rect 477004 586654 477604 622098
rect 477004 586418 477186 586654
rect 477422 586418 477604 586654
rect 477004 586334 477604 586418
rect 477004 586098 477186 586334
rect 477422 586098 477604 586334
rect 477004 550654 477604 586098
rect 477004 550418 477186 550654
rect 477422 550418 477604 550654
rect 477004 550334 477604 550418
rect 477004 550098 477186 550334
rect 477422 550098 477604 550334
rect 477004 514654 477604 550098
rect 477004 514418 477186 514654
rect 477422 514418 477604 514654
rect 477004 514334 477604 514418
rect 477004 514098 477186 514334
rect 477422 514098 477604 514334
rect 477004 478654 477604 514098
rect 477004 478418 477186 478654
rect 477422 478418 477604 478654
rect 477004 478334 477604 478418
rect 477004 478098 477186 478334
rect 477422 478098 477604 478334
rect 477004 442654 477604 478098
rect 477004 442418 477186 442654
rect 477422 442418 477604 442654
rect 477004 442334 477604 442418
rect 477004 442098 477186 442334
rect 477422 442098 477604 442334
rect 477004 406654 477604 442098
rect 477004 406418 477186 406654
rect 477422 406418 477604 406654
rect 477004 406334 477604 406418
rect 477004 406098 477186 406334
rect 477422 406098 477604 406334
rect 477004 370654 477604 406098
rect 477004 370418 477186 370654
rect 477422 370418 477604 370654
rect 477004 370334 477604 370418
rect 477004 370098 477186 370334
rect 477422 370098 477604 370334
rect 477004 334654 477604 370098
rect 477004 334418 477186 334654
rect 477422 334418 477604 334654
rect 477004 334334 477604 334418
rect 477004 334098 477186 334334
rect 477422 334098 477604 334334
rect 477004 298654 477604 334098
rect 477004 298418 477186 298654
rect 477422 298418 477604 298654
rect 477004 298334 477604 298418
rect 477004 298098 477186 298334
rect 477422 298098 477604 298334
rect 477004 262654 477604 298098
rect 477004 262418 477186 262654
rect 477422 262418 477604 262654
rect 477004 262334 477604 262418
rect 477004 262098 477186 262334
rect 477422 262098 477604 262334
rect 477004 226654 477604 262098
rect 477004 226418 477186 226654
rect 477422 226418 477604 226654
rect 477004 226334 477604 226418
rect 477004 226098 477186 226334
rect 477422 226098 477604 226334
rect 477004 190654 477604 226098
rect 477004 190418 477186 190654
rect 477422 190418 477604 190654
rect 477004 190334 477604 190418
rect 477004 190098 477186 190334
rect 477422 190098 477604 190334
rect 477004 154654 477604 190098
rect 477004 154418 477186 154654
rect 477422 154418 477604 154654
rect 477004 154334 477604 154418
rect 477004 154098 477186 154334
rect 477422 154098 477604 154334
rect 477004 118654 477604 154098
rect 477004 118418 477186 118654
rect 477422 118418 477604 118654
rect 477004 118334 477604 118418
rect 477004 118098 477186 118334
rect 477422 118098 477604 118334
rect 477004 82654 477604 118098
rect 477004 82418 477186 82654
rect 477422 82418 477604 82654
rect 477004 82334 477604 82418
rect 477004 82098 477186 82334
rect 477422 82098 477604 82334
rect 477004 46654 477604 82098
rect 477004 46418 477186 46654
rect 477422 46418 477604 46654
rect 477004 46334 477604 46418
rect 477004 46098 477186 46334
rect 477422 46098 477604 46334
rect 477004 10654 477604 46098
rect 477004 10418 477186 10654
rect 477422 10418 477604 10654
rect 477004 10334 477604 10418
rect 477004 10098 477186 10334
rect 477422 10098 477604 10334
rect 477004 -4106 477604 10098
rect 477004 -4342 477186 -4106
rect 477422 -4342 477604 -4106
rect 477004 -4426 477604 -4342
rect 477004 -4662 477186 -4426
rect 477422 -4662 477604 -4426
rect 477004 -5624 477604 -4662
rect 480604 698254 481204 709922
rect 498604 711418 499204 711440
rect 498604 711182 498786 711418
rect 499022 711182 499204 711418
rect 498604 711098 499204 711182
rect 498604 710862 498786 711098
rect 499022 710862 499204 711098
rect 495004 709538 495604 709560
rect 495004 709302 495186 709538
rect 495422 709302 495604 709538
rect 495004 709218 495604 709302
rect 495004 708982 495186 709218
rect 495422 708982 495604 709218
rect 491404 707658 492004 707680
rect 491404 707422 491586 707658
rect 491822 707422 492004 707658
rect 491404 707338 492004 707422
rect 491404 707102 491586 707338
rect 491822 707102 492004 707338
rect 480604 698018 480786 698254
rect 481022 698018 481204 698254
rect 480604 697934 481204 698018
rect 480604 697698 480786 697934
rect 481022 697698 481204 697934
rect 480604 662254 481204 697698
rect 480604 662018 480786 662254
rect 481022 662018 481204 662254
rect 480604 661934 481204 662018
rect 480604 661698 480786 661934
rect 481022 661698 481204 661934
rect 480604 626254 481204 661698
rect 480604 626018 480786 626254
rect 481022 626018 481204 626254
rect 480604 625934 481204 626018
rect 480604 625698 480786 625934
rect 481022 625698 481204 625934
rect 480604 590254 481204 625698
rect 480604 590018 480786 590254
rect 481022 590018 481204 590254
rect 480604 589934 481204 590018
rect 480604 589698 480786 589934
rect 481022 589698 481204 589934
rect 480604 554254 481204 589698
rect 480604 554018 480786 554254
rect 481022 554018 481204 554254
rect 480604 553934 481204 554018
rect 480604 553698 480786 553934
rect 481022 553698 481204 553934
rect 480604 518254 481204 553698
rect 480604 518018 480786 518254
rect 481022 518018 481204 518254
rect 480604 517934 481204 518018
rect 480604 517698 480786 517934
rect 481022 517698 481204 517934
rect 480604 482254 481204 517698
rect 480604 482018 480786 482254
rect 481022 482018 481204 482254
rect 480604 481934 481204 482018
rect 480604 481698 480786 481934
rect 481022 481698 481204 481934
rect 480604 446254 481204 481698
rect 480604 446018 480786 446254
rect 481022 446018 481204 446254
rect 480604 445934 481204 446018
rect 480604 445698 480786 445934
rect 481022 445698 481204 445934
rect 480604 410254 481204 445698
rect 480604 410018 480786 410254
rect 481022 410018 481204 410254
rect 480604 409934 481204 410018
rect 480604 409698 480786 409934
rect 481022 409698 481204 409934
rect 480604 374254 481204 409698
rect 480604 374018 480786 374254
rect 481022 374018 481204 374254
rect 480604 373934 481204 374018
rect 480604 373698 480786 373934
rect 481022 373698 481204 373934
rect 480604 338254 481204 373698
rect 480604 338018 480786 338254
rect 481022 338018 481204 338254
rect 480604 337934 481204 338018
rect 480604 337698 480786 337934
rect 481022 337698 481204 337934
rect 480604 302254 481204 337698
rect 480604 302018 480786 302254
rect 481022 302018 481204 302254
rect 480604 301934 481204 302018
rect 480604 301698 480786 301934
rect 481022 301698 481204 301934
rect 480604 266254 481204 301698
rect 480604 266018 480786 266254
rect 481022 266018 481204 266254
rect 480604 265934 481204 266018
rect 480604 265698 480786 265934
rect 481022 265698 481204 265934
rect 480604 230254 481204 265698
rect 480604 230018 480786 230254
rect 481022 230018 481204 230254
rect 480604 229934 481204 230018
rect 480604 229698 480786 229934
rect 481022 229698 481204 229934
rect 480604 194254 481204 229698
rect 480604 194018 480786 194254
rect 481022 194018 481204 194254
rect 480604 193934 481204 194018
rect 480604 193698 480786 193934
rect 481022 193698 481204 193934
rect 480604 158254 481204 193698
rect 480604 158018 480786 158254
rect 481022 158018 481204 158254
rect 480604 157934 481204 158018
rect 480604 157698 480786 157934
rect 481022 157698 481204 157934
rect 480604 122254 481204 157698
rect 480604 122018 480786 122254
rect 481022 122018 481204 122254
rect 480604 121934 481204 122018
rect 480604 121698 480786 121934
rect 481022 121698 481204 121934
rect 480604 86254 481204 121698
rect 480604 86018 480786 86254
rect 481022 86018 481204 86254
rect 480604 85934 481204 86018
rect 480604 85698 480786 85934
rect 481022 85698 481204 85934
rect 480604 50254 481204 85698
rect 480604 50018 480786 50254
rect 481022 50018 481204 50254
rect 480604 49934 481204 50018
rect 480604 49698 480786 49934
rect 481022 49698 481204 49934
rect 480604 14254 481204 49698
rect 480604 14018 480786 14254
rect 481022 14018 481204 14254
rect 480604 13934 481204 14018
rect 480604 13698 480786 13934
rect 481022 13698 481204 13934
rect 462604 -7162 462786 -6926
rect 463022 -7162 463204 -6926
rect 462604 -7246 463204 -7162
rect 462604 -7482 462786 -7246
rect 463022 -7482 463204 -7246
rect 462604 -7504 463204 -7482
rect 480604 -5986 481204 13698
rect 487804 705778 488404 705800
rect 487804 705542 487986 705778
rect 488222 705542 488404 705778
rect 487804 705458 488404 705542
rect 487804 705222 487986 705458
rect 488222 705222 488404 705458
rect 487804 669454 488404 705222
rect 487804 669218 487986 669454
rect 488222 669218 488404 669454
rect 487804 669134 488404 669218
rect 487804 668898 487986 669134
rect 488222 668898 488404 669134
rect 487804 633454 488404 668898
rect 487804 633218 487986 633454
rect 488222 633218 488404 633454
rect 487804 633134 488404 633218
rect 487804 632898 487986 633134
rect 488222 632898 488404 633134
rect 487804 597454 488404 632898
rect 487804 597218 487986 597454
rect 488222 597218 488404 597454
rect 487804 597134 488404 597218
rect 487804 596898 487986 597134
rect 488222 596898 488404 597134
rect 487804 561454 488404 596898
rect 487804 561218 487986 561454
rect 488222 561218 488404 561454
rect 487804 561134 488404 561218
rect 487804 560898 487986 561134
rect 488222 560898 488404 561134
rect 487804 525454 488404 560898
rect 487804 525218 487986 525454
rect 488222 525218 488404 525454
rect 487804 525134 488404 525218
rect 487804 524898 487986 525134
rect 488222 524898 488404 525134
rect 487804 489454 488404 524898
rect 487804 489218 487986 489454
rect 488222 489218 488404 489454
rect 487804 489134 488404 489218
rect 487804 488898 487986 489134
rect 488222 488898 488404 489134
rect 487804 453454 488404 488898
rect 487804 453218 487986 453454
rect 488222 453218 488404 453454
rect 487804 453134 488404 453218
rect 487804 452898 487986 453134
rect 488222 452898 488404 453134
rect 487804 417454 488404 452898
rect 487804 417218 487986 417454
rect 488222 417218 488404 417454
rect 487804 417134 488404 417218
rect 487804 416898 487986 417134
rect 488222 416898 488404 417134
rect 487804 381454 488404 416898
rect 487804 381218 487986 381454
rect 488222 381218 488404 381454
rect 487804 381134 488404 381218
rect 487804 380898 487986 381134
rect 488222 380898 488404 381134
rect 487804 345454 488404 380898
rect 487804 345218 487986 345454
rect 488222 345218 488404 345454
rect 487804 345134 488404 345218
rect 487804 344898 487986 345134
rect 488222 344898 488404 345134
rect 487804 309454 488404 344898
rect 487804 309218 487986 309454
rect 488222 309218 488404 309454
rect 487804 309134 488404 309218
rect 487804 308898 487986 309134
rect 488222 308898 488404 309134
rect 487804 273454 488404 308898
rect 487804 273218 487986 273454
rect 488222 273218 488404 273454
rect 487804 273134 488404 273218
rect 487804 272898 487986 273134
rect 488222 272898 488404 273134
rect 487804 237454 488404 272898
rect 487804 237218 487986 237454
rect 488222 237218 488404 237454
rect 487804 237134 488404 237218
rect 487804 236898 487986 237134
rect 488222 236898 488404 237134
rect 487804 201454 488404 236898
rect 487804 201218 487986 201454
rect 488222 201218 488404 201454
rect 487804 201134 488404 201218
rect 487804 200898 487986 201134
rect 488222 200898 488404 201134
rect 487804 165454 488404 200898
rect 487804 165218 487986 165454
rect 488222 165218 488404 165454
rect 487804 165134 488404 165218
rect 487804 164898 487986 165134
rect 488222 164898 488404 165134
rect 487804 129454 488404 164898
rect 487804 129218 487986 129454
rect 488222 129218 488404 129454
rect 487804 129134 488404 129218
rect 487804 128898 487986 129134
rect 488222 128898 488404 129134
rect 487804 93454 488404 128898
rect 487804 93218 487986 93454
rect 488222 93218 488404 93454
rect 487804 93134 488404 93218
rect 487804 92898 487986 93134
rect 488222 92898 488404 93134
rect 487804 57454 488404 92898
rect 487804 57218 487986 57454
rect 488222 57218 488404 57454
rect 487804 57134 488404 57218
rect 487804 56898 487986 57134
rect 488222 56898 488404 57134
rect 487804 21454 488404 56898
rect 487804 21218 487986 21454
rect 488222 21218 488404 21454
rect 487804 21134 488404 21218
rect 487804 20898 487986 21134
rect 488222 20898 488404 21134
rect 487804 -1286 488404 20898
rect 487804 -1522 487986 -1286
rect 488222 -1522 488404 -1286
rect 487804 -1606 488404 -1522
rect 487804 -1842 487986 -1606
rect 488222 -1842 488404 -1606
rect 487804 -1864 488404 -1842
rect 491404 673054 492004 707102
rect 491404 672818 491586 673054
rect 491822 672818 492004 673054
rect 491404 672734 492004 672818
rect 491404 672498 491586 672734
rect 491822 672498 492004 672734
rect 491404 637054 492004 672498
rect 491404 636818 491586 637054
rect 491822 636818 492004 637054
rect 491404 636734 492004 636818
rect 491404 636498 491586 636734
rect 491822 636498 492004 636734
rect 491404 601054 492004 636498
rect 491404 600818 491586 601054
rect 491822 600818 492004 601054
rect 491404 600734 492004 600818
rect 491404 600498 491586 600734
rect 491822 600498 492004 600734
rect 491404 565054 492004 600498
rect 491404 564818 491586 565054
rect 491822 564818 492004 565054
rect 491404 564734 492004 564818
rect 491404 564498 491586 564734
rect 491822 564498 492004 564734
rect 491404 529054 492004 564498
rect 491404 528818 491586 529054
rect 491822 528818 492004 529054
rect 491404 528734 492004 528818
rect 491404 528498 491586 528734
rect 491822 528498 492004 528734
rect 491404 493054 492004 528498
rect 491404 492818 491586 493054
rect 491822 492818 492004 493054
rect 491404 492734 492004 492818
rect 491404 492498 491586 492734
rect 491822 492498 492004 492734
rect 491404 457054 492004 492498
rect 491404 456818 491586 457054
rect 491822 456818 492004 457054
rect 491404 456734 492004 456818
rect 491404 456498 491586 456734
rect 491822 456498 492004 456734
rect 491404 421054 492004 456498
rect 491404 420818 491586 421054
rect 491822 420818 492004 421054
rect 491404 420734 492004 420818
rect 491404 420498 491586 420734
rect 491822 420498 492004 420734
rect 491404 385054 492004 420498
rect 491404 384818 491586 385054
rect 491822 384818 492004 385054
rect 491404 384734 492004 384818
rect 491404 384498 491586 384734
rect 491822 384498 492004 384734
rect 491404 349054 492004 384498
rect 491404 348818 491586 349054
rect 491822 348818 492004 349054
rect 491404 348734 492004 348818
rect 491404 348498 491586 348734
rect 491822 348498 492004 348734
rect 491404 313054 492004 348498
rect 491404 312818 491586 313054
rect 491822 312818 492004 313054
rect 491404 312734 492004 312818
rect 491404 312498 491586 312734
rect 491822 312498 492004 312734
rect 491404 277054 492004 312498
rect 491404 276818 491586 277054
rect 491822 276818 492004 277054
rect 491404 276734 492004 276818
rect 491404 276498 491586 276734
rect 491822 276498 492004 276734
rect 491404 241054 492004 276498
rect 491404 240818 491586 241054
rect 491822 240818 492004 241054
rect 491404 240734 492004 240818
rect 491404 240498 491586 240734
rect 491822 240498 492004 240734
rect 491404 205054 492004 240498
rect 491404 204818 491586 205054
rect 491822 204818 492004 205054
rect 491404 204734 492004 204818
rect 491404 204498 491586 204734
rect 491822 204498 492004 204734
rect 491404 169054 492004 204498
rect 491404 168818 491586 169054
rect 491822 168818 492004 169054
rect 491404 168734 492004 168818
rect 491404 168498 491586 168734
rect 491822 168498 492004 168734
rect 491404 133054 492004 168498
rect 491404 132818 491586 133054
rect 491822 132818 492004 133054
rect 491404 132734 492004 132818
rect 491404 132498 491586 132734
rect 491822 132498 492004 132734
rect 491404 97054 492004 132498
rect 491404 96818 491586 97054
rect 491822 96818 492004 97054
rect 491404 96734 492004 96818
rect 491404 96498 491586 96734
rect 491822 96498 492004 96734
rect 491404 61054 492004 96498
rect 491404 60818 491586 61054
rect 491822 60818 492004 61054
rect 491404 60734 492004 60818
rect 491404 60498 491586 60734
rect 491822 60498 492004 60734
rect 491404 25054 492004 60498
rect 491404 24818 491586 25054
rect 491822 24818 492004 25054
rect 491404 24734 492004 24818
rect 491404 24498 491586 24734
rect 491822 24498 492004 24734
rect 491404 -3166 492004 24498
rect 491404 -3402 491586 -3166
rect 491822 -3402 492004 -3166
rect 491404 -3486 492004 -3402
rect 491404 -3722 491586 -3486
rect 491822 -3722 492004 -3486
rect 491404 -3744 492004 -3722
rect 495004 676654 495604 708982
rect 495004 676418 495186 676654
rect 495422 676418 495604 676654
rect 495004 676334 495604 676418
rect 495004 676098 495186 676334
rect 495422 676098 495604 676334
rect 495004 640654 495604 676098
rect 495004 640418 495186 640654
rect 495422 640418 495604 640654
rect 495004 640334 495604 640418
rect 495004 640098 495186 640334
rect 495422 640098 495604 640334
rect 495004 604654 495604 640098
rect 495004 604418 495186 604654
rect 495422 604418 495604 604654
rect 495004 604334 495604 604418
rect 495004 604098 495186 604334
rect 495422 604098 495604 604334
rect 495004 568654 495604 604098
rect 495004 568418 495186 568654
rect 495422 568418 495604 568654
rect 495004 568334 495604 568418
rect 495004 568098 495186 568334
rect 495422 568098 495604 568334
rect 495004 532654 495604 568098
rect 495004 532418 495186 532654
rect 495422 532418 495604 532654
rect 495004 532334 495604 532418
rect 495004 532098 495186 532334
rect 495422 532098 495604 532334
rect 495004 496654 495604 532098
rect 495004 496418 495186 496654
rect 495422 496418 495604 496654
rect 495004 496334 495604 496418
rect 495004 496098 495186 496334
rect 495422 496098 495604 496334
rect 495004 460654 495604 496098
rect 495004 460418 495186 460654
rect 495422 460418 495604 460654
rect 495004 460334 495604 460418
rect 495004 460098 495186 460334
rect 495422 460098 495604 460334
rect 495004 424654 495604 460098
rect 495004 424418 495186 424654
rect 495422 424418 495604 424654
rect 495004 424334 495604 424418
rect 495004 424098 495186 424334
rect 495422 424098 495604 424334
rect 495004 388654 495604 424098
rect 495004 388418 495186 388654
rect 495422 388418 495604 388654
rect 495004 388334 495604 388418
rect 495004 388098 495186 388334
rect 495422 388098 495604 388334
rect 495004 352654 495604 388098
rect 495004 352418 495186 352654
rect 495422 352418 495604 352654
rect 495004 352334 495604 352418
rect 495004 352098 495186 352334
rect 495422 352098 495604 352334
rect 495004 316654 495604 352098
rect 495004 316418 495186 316654
rect 495422 316418 495604 316654
rect 495004 316334 495604 316418
rect 495004 316098 495186 316334
rect 495422 316098 495604 316334
rect 495004 280654 495604 316098
rect 495004 280418 495186 280654
rect 495422 280418 495604 280654
rect 495004 280334 495604 280418
rect 495004 280098 495186 280334
rect 495422 280098 495604 280334
rect 495004 244654 495604 280098
rect 495004 244418 495186 244654
rect 495422 244418 495604 244654
rect 495004 244334 495604 244418
rect 495004 244098 495186 244334
rect 495422 244098 495604 244334
rect 495004 208654 495604 244098
rect 495004 208418 495186 208654
rect 495422 208418 495604 208654
rect 495004 208334 495604 208418
rect 495004 208098 495186 208334
rect 495422 208098 495604 208334
rect 495004 172654 495604 208098
rect 495004 172418 495186 172654
rect 495422 172418 495604 172654
rect 495004 172334 495604 172418
rect 495004 172098 495186 172334
rect 495422 172098 495604 172334
rect 495004 136654 495604 172098
rect 495004 136418 495186 136654
rect 495422 136418 495604 136654
rect 495004 136334 495604 136418
rect 495004 136098 495186 136334
rect 495422 136098 495604 136334
rect 495004 100654 495604 136098
rect 495004 100418 495186 100654
rect 495422 100418 495604 100654
rect 495004 100334 495604 100418
rect 495004 100098 495186 100334
rect 495422 100098 495604 100334
rect 495004 64654 495604 100098
rect 495004 64418 495186 64654
rect 495422 64418 495604 64654
rect 495004 64334 495604 64418
rect 495004 64098 495186 64334
rect 495422 64098 495604 64334
rect 495004 28654 495604 64098
rect 495004 28418 495186 28654
rect 495422 28418 495604 28654
rect 495004 28334 495604 28418
rect 495004 28098 495186 28334
rect 495422 28098 495604 28334
rect 495004 -5046 495604 28098
rect 495004 -5282 495186 -5046
rect 495422 -5282 495604 -5046
rect 495004 -5366 495604 -5282
rect 495004 -5602 495186 -5366
rect 495422 -5602 495604 -5366
rect 495004 -5624 495604 -5602
rect 498604 680254 499204 710862
rect 516604 710478 517204 711440
rect 516604 710242 516786 710478
rect 517022 710242 517204 710478
rect 516604 710158 517204 710242
rect 516604 709922 516786 710158
rect 517022 709922 517204 710158
rect 513004 708598 513604 709560
rect 513004 708362 513186 708598
rect 513422 708362 513604 708598
rect 513004 708278 513604 708362
rect 513004 708042 513186 708278
rect 513422 708042 513604 708278
rect 509404 706718 510004 707680
rect 509404 706482 509586 706718
rect 509822 706482 510004 706718
rect 509404 706398 510004 706482
rect 509404 706162 509586 706398
rect 509822 706162 510004 706398
rect 498604 680018 498786 680254
rect 499022 680018 499204 680254
rect 498604 679934 499204 680018
rect 498604 679698 498786 679934
rect 499022 679698 499204 679934
rect 498604 644254 499204 679698
rect 498604 644018 498786 644254
rect 499022 644018 499204 644254
rect 498604 643934 499204 644018
rect 498604 643698 498786 643934
rect 499022 643698 499204 643934
rect 498604 608254 499204 643698
rect 498604 608018 498786 608254
rect 499022 608018 499204 608254
rect 498604 607934 499204 608018
rect 498604 607698 498786 607934
rect 499022 607698 499204 607934
rect 498604 572254 499204 607698
rect 498604 572018 498786 572254
rect 499022 572018 499204 572254
rect 498604 571934 499204 572018
rect 498604 571698 498786 571934
rect 499022 571698 499204 571934
rect 498604 536254 499204 571698
rect 498604 536018 498786 536254
rect 499022 536018 499204 536254
rect 498604 535934 499204 536018
rect 498604 535698 498786 535934
rect 499022 535698 499204 535934
rect 498604 500254 499204 535698
rect 498604 500018 498786 500254
rect 499022 500018 499204 500254
rect 498604 499934 499204 500018
rect 498604 499698 498786 499934
rect 499022 499698 499204 499934
rect 498604 464254 499204 499698
rect 498604 464018 498786 464254
rect 499022 464018 499204 464254
rect 498604 463934 499204 464018
rect 498604 463698 498786 463934
rect 499022 463698 499204 463934
rect 498604 428254 499204 463698
rect 498604 428018 498786 428254
rect 499022 428018 499204 428254
rect 498604 427934 499204 428018
rect 498604 427698 498786 427934
rect 499022 427698 499204 427934
rect 498604 392254 499204 427698
rect 498604 392018 498786 392254
rect 499022 392018 499204 392254
rect 498604 391934 499204 392018
rect 498604 391698 498786 391934
rect 499022 391698 499204 391934
rect 498604 356254 499204 391698
rect 498604 356018 498786 356254
rect 499022 356018 499204 356254
rect 498604 355934 499204 356018
rect 498604 355698 498786 355934
rect 499022 355698 499204 355934
rect 498604 320254 499204 355698
rect 498604 320018 498786 320254
rect 499022 320018 499204 320254
rect 498604 319934 499204 320018
rect 498604 319698 498786 319934
rect 499022 319698 499204 319934
rect 498604 284254 499204 319698
rect 498604 284018 498786 284254
rect 499022 284018 499204 284254
rect 498604 283934 499204 284018
rect 498604 283698 498786 283934
rect 499022 283698 499204 283934
rect 498604 248254 499204 283698
rect 498604 248018 498786 248254
rect 499022 248018 499204 248254
rect 498604 247934 499204 248018
rect 498604 247698 498786 247934
rect 499022 247698 499204 247934
rect 498604 212254 499204 247698
rect 498604 212018 498786 212254
rect 499022 212018 499204 212254
rect 498604 211934 499204 212018
rect 498604 211698 498786 211934
rect 499022 211698 499204 211934
rect 498604 176254 499204 211698
rect 498604 176018 498786 176254
rect 499022 176018 499204 176254
rect 498604 175934 499204 176018
rect 498604 175698 498786 175934
rect 499022 175698 499204 175934
rect 498604 140254 499204 175698
rect 498604 140018 498786 140254
rect 499022 140018 499204 140254
rect 498604 139934 499204 140018
rect 498604 139698 498786 139934
rect 499022 139698 499204 139934
rect 498604 104254 499204 139698
rect 498604 104018 498786 104254
rect 499022 104018 499204 104254
rect 498604 103934 499204 104018
rect 498604 103698 498786 103934
rect 499022 103698 499204 103934
rect 498604 68254 499204 103698
rect 498604 68018 498786 68254
rect 499022 68018 499204 68254
rect 498604 67934 499204 68018
rect 498604 67698 498786 67934
rect 499022 67698 499204 67934
rect 498604 32254 499204 67698
rect 498604 32018 498786 32254
rect 499022 32018 499204 32254
rect 498604 31934 499204 32018
rect 498604 31698 498786 31934
rect 499022 31698 499204 31934
rect 480604 -6222 480786 -5986
rect 481022 -6222 481204 -5986
rect 480604 -6306 481204 -6222
rect 480604 -6542 480786 -6306
rect 481022 -6542 481204 -6306
rect 480604 -7504 481204 -6542
rect 498604 -6926 499204 31698
rect 505804 704838 506404 705800
rect 505804 704602 505986 704838
rect 506222 704602 506404 704838
rect 505804 704518 506404 704602
rect 505804 704282 505986 704518
rect 506222 704282 506404 704518
rect 505804 687454 506404 704282
rect 505804 687218 505986 687454
rect 506222 687218 506404 687454
rect 505804 687134 506404 687218
rect 505804 686898 505986 687134
rect 506222 686898 506404 687134
rect 505804 651454 506404 686898
rect 505804 651218 505986 651454
rect 506222 651218 506404 651454
rect 505804 651134 506404 651218
rect 505804 650898 505986 651134
rect 506222 650898 506404 651134
rect 505804 615454 506404 650898
rect 505804 615218 505986 615454
rect 506222 615218 506404 615454
rect 505804 615134 506404 615218
rect 505804 614898 505986 615134
rect 506222 614898 506404 615134
rect 505804 579454 506404 614898
rect 505804 579218 505986 579454
rect 506222 579218 506404 579454
rect 505804 579134 506404 579218
rect 505804 578898 505986 579134
rect 506222 578898 506404 579134
rect 505804 543454 506404 578898
rect 505804 543218 505986 543454
rect 506222 543218 506404 543454
rect 505804 543134 506404 543218
rect 505804 542898 505986 543134
rect 506222 542898 506404 543134
rect 505804 507454 506404 542898
rect 505804 507218 505986 507454
rect 506222 507218 506404 507454
rect 505804 507134 506404 507218
rect 505804 506898 505986 507134
rect 506222 506898 506404 507134
rect 505804 471454 506404 506898
rect 505804 471218 505986 471454
rect 506222 471218 506404 471454
rect 505804 471134 506404 471218
rect 505804 470898 505986 471134
rect 506222 470898 506404 471134
rect 505804 435454 506404 470898
rect 505804 435218 505986 435454
rect 506222 435218 506404 435454
rect 505804 435134 506404 435218
rect 505804 434898 505986 435134
rect 506222 434898 506404 435134
rect 505804 399454 506404 434898
rect 505804 399218 505986 399454
rect 506222 399218 506404 399454
rect 505804 399134 506404 399218
rect 505804 398898 505986 399134
rect 506222 398898 506404 399134
rect 505804 363454 506404 398898
rect 505804 363218 505986 363454
rect 506222 363218 506404 363454
rect 505804 363134 506404 363218
rect 505804 362898 505986 363134
rect 506222 362898 506404 363134
rect 505804 327454 506404 362898
rect 505804 327218 505986 327454
rect 506222 327218 506404 327454
rect 505804 327134 506404 327218
rect 505804 326898 505986 327134
rect 506222 326898 506404 327134
rect 505804 291454 506404 326898
rect 505804 291218 505986 291454
rect 506222 291218 506404 291454
rect 505804 291134 506404 291218
rect 505804 290898 505986 291134
rect 506222 290898 506404 291134
rect 505804 255454 506404 290898
rect 505804 255218 505986 255454
rect 506222 255218 506404 255454
rect 505804 255134 506404 255218
rect 505804 254898 505986 255134
rect 506222 254898 506404 255134
rect 505804 219454 506404 254898
rect 505804 219218 505986 219454
rect 506222 219218 506404 219454
rect 505804 219134 506404 219218
rect 505804 218898 505986 219134
rect 506222 218898 506404 219134
rect 505804 183454 506404 218898
rect 505804 183218 505986 183454
rect 506222 183218 506404 183454
rect 505804 183134 506404 183218
rect 505804 182898 505986 183134
rect 506222 182898 506404 183134
rect 505804 147454 506404 182898
rect 505804 147218 505986 147454
rect 506222 147218 506404 147454
rect 505804 147134 506404 147218
rect 505804 146898 505986 147134
rect 506222 146898 506404 147134
rect 505804 111454 506404 146898
rect 505804 111218 505986 111454
rect 506222 111218 506404 111454
rect 505804 111134 506404 111218
rect 505804 110898 505986 111134
rect 506222 110898 506404 111134
rect 505804 75454 506404 110898
rect 505804 75218 505986 75454
rect 506222 75218 506404 75454
rect 505804 75134 506404 75218
rect 505804 74898 505986 75134
rect 506222 74898 506404 75134
rect 505804 39454 506404 74898
rect 505804 39218 505986 39454
rect 506222 39218 506404 39454
rect 505804 39134 506404 39218
rect 505804 38898 505986 39134
rect 506222 38898 506404 39134
rect 505804 3454 506404 38898
rect 505804 3218 505986 3454
rect 506222 3218 506404 3454
rect 505804 3134 506404 3218
rect 505804 2898 505986 3134
rect 506222 2898 506404 3134
rect 505804 -346 506404 2898
rect 505804 -582 505986 -346
rect 506222 -582 506404 -346
rect 505804 -666 506404 -582
rect 505804 -902 505986 -666
rect 506222 -902 506404 -666
rect 505804 -1864 506404 -902
rect 509404 691054 510004 706162
rect 509404 690818 509586 691054
rect 509822 690818 510004 691054
rect 509404 690734 510004 690818
rect 509404 690498 509586 690734
rect 509822 690498 510004 690734
rect 509404 655054 510004 690498
rect 509404 654818 509586 655054
rect 509822 654818 510004 655054
rect 509404 654734 510004 654818
rect 509404 654498 509586 654734
rect 509822 654498 510004 654734
rect 509404 619054 510004 654498
rect 509404 618818 509586 619054
rect 509822 618818 510004 619054
rect 509404 618734 510004 618818
rect 509404 618498 509586 618734
rect 509822 618498 510004 618734
rect 509404 583054 510004 618498
rect 509404 582818 509586 583054
rect 509822 582818 510004 583054
rect 509404 582734 510004 582818
rect 509404 582498 509586 582734
rect 509822 582498 510004 582734
rect 509404 547054 510004 582498
rect 509404 546818 509586 547054
rect 509822 546818 510004 547054
rect 509404 546734 510004 546818
rect 509404 546498 509586 546734
rect 509822 546498 510004 546734
rect 509404 511054 510004 546498
rect 509404 510818 509586 511054
rect 509822 510818 510004 511054
rect 509404 510734 510004 510818
rect 509404 510498 509586 510734
rect 509822 510498 510004 510734
rect 509404 475054 510004 510498
rect 509404 474818 509586 475054
rect 509822 474818 510004 475054
rect 509404 474734 510004 474818
rect 509404 474498 509586 474734
rect 509822 474498 510004 474734
rect 509404 439054 510004 474498
rect 509404 438818 509586 439054
rect 509822 438818 510004 439054
rect 509404 438734 510004 438818
rect 509404 438498 509586 438734
rect 509822 438498 510004 438734
rect 509404 403054 510004 438498
rect 509404 402818 509586 403054
rect 509822 402818 510004 403054
rect 509404 402734 510004 402818
rect 509404 402498 509586 402734
rect 509822 402498 510004 402734
rect 509404 367054 510004 402498
rect 509404 366818 509586 367054
rect 509822 366818 510004 367054
rect 509404 366734 510004 366818
rect 509404 366498 509586 366734
rect 509822 366498 510004 366734
rect 509404 331054 510004 366498
rect 509404 330818 509586 331054
rect 509822 330818 510004 331054
rect 509404 330734 510004 330818
rect 509404 330498 509586 330734
rect 509822 330498 510004 330734
rect 509404 295054 510004 330498
rect 509404 294818 509586 295054
rect 509822 294818 510004 295054
rect 509404 294734 510004 294818
rect 509404 294498 509586 294734
rect 509822 294498 510004 294734
rect 509404 259054 510004 294498
rect 509404 258818 509586 259054
rect 509822 258818 510004 259054
rect 509404 258734 510004 258818
rect 509404 258498 509586 258734
rect 509822 258498 510004 258734
rect 509404 223054 510004 258498
rect 509404 222818 509586 223054
rect 509822 222818 510004 223054
rect 509404 222734 510004 222818
rect 509404 222498 509586 222734
rect 509822 222498 510004 222734
rect 509404 187054 510004 222498
rect 509404 186818 509586 187054
rect 509822 186818 510004 187054
rect 509404 186734 510004 186818
rect 509404 186498 509586 186734
rect 509822 186498 510004 186734
rect 509404 151054 510004 186498
rect 509404 150818 509586 151054
rect 509822 150818 510004 151054
rect 509404 150734 510004 150818
rect 509404 150498 509586 150734
rect 509822 150498 510004 150734
rect 509404 115054 510004 150498
rect 509404 114818 509586 115054
rect 509822 114818 510004 115054
rect 509404 114734 510004 114818
rect 509404 114498 509586 114734
rect 509822 114498 510004 114734
rect 509404 79054 510004 114498
rect 509404 78818 509586 79054
rect 509822 78818 510004 79054
rect 509404 78734 510004 78818
rect 509404 78498 509586 78734
rect 509822 78498 510004 78734
rect 509404 43054 510004 78498
rect 509404 42818 509586 43054
rect 509822 42818 510004 43054
rect 509404 42734 510004 42818
rect 509404 42498 509586 42734
rect 509822 42498 510004 42734
rect 509404 7054 510004 42498
rect 509404 6818 509586 7054
rect 509822 6818 510004 7054
rect 509404 6734 510004 6818
rect 509404 6498 509586 6734
rect 509822 6498 510004 6734
rect 509404 -2226 510004 6498
rect 509404 -2462 509586 -2226
rect 509822 -2462 510004 -2226
rect 509404 -2546 510004 -2462
rect 509404 -2782 509586 -2546
rect 509822 -2782 510004 -2546
rect 509404 -3744 510004 -2782
rect 513004 694654 513604 708042
rect 513004 694418 513186 694654
rect 513422 694418 513604 694654
rect 513004 694334 513604 694418
rect 513004 694098 513186 694334
rect 513422 694098 513604 694334
rect 513004 658654 513604 694098
rect 513004 658418 513186 658654
rect 513422 658418 513604 658654
rect 513004 658334 513604 658418
rect 513004 658098 513186 658334
rect 513422 658098 513604 658334
rect 513004 622654 513604 658098
rect 513004 622418 513186 622654
rect 513422 622418 513604 622654
rect 513004 622334 513604 622418
rect 513004 622098 513186 622334
rect 513422 622098 513604 622334
rect 513004 586654 513604 622098
rect 513004 586418 513186 586654
rect 513422 586418 513604 586654
rect 513004 586334 513604 586418
rect 513004 586098 513186 586334
rect 513422 586098 513604 586334
rect 513004 550654 513604 586098
rect 513004 550418 513186 550654
rect 513422 550418 513604 550654
rect 513004 550334 513604 550418
rect 513004 550098 513186 550334
rect 513422 550098 513604 550334
rect 513004 514654 513604 550098
rect 513004 514418 513186 514654
rect 513422 514418 513604 514654
rect 513004 514334 513604 514418
rect 513004 514098 513186 514334
rect 513422 514098 513604 514334
rect 513004 478654 513604 514098
rect 513004 478418 513186 478654
rect 513422 478418 513604 478654
rect 513004 478334 513604 478418
rect 513004 478098 513186 478334
rect 513422 478098 513604 478334
rect 513004 442654 513604 478098
rect 513004 442418 513186 442654
rect 513422 442418 513604 442654
rect 513004 442334 513604 442418
rect 513004 442098 513186 442334
rect 513422 442098 513604 442334
rect 513004 406654 513604 442098
rect 513004 406418 513186 406654
rect 513422 406418 513604 406654
rect 513004 406334 513604 406418
rect 513004 406098 513186 406334
rect 513422 406098 513604 406334
rect 513004 370654 513604 406098
rect 513004 370418 513186 370654
rect 513422 370418 513604 370654
rect 513004 370334 513604 370418
rect 513004 370098 513186 370334
rect 513422 370098 513604 370334
rect 513004 334654 513604 370098
rect 513004 334418 513186 334654
rect 513422 334418 513604 334654
rect 513004 334334 513604 334418
rect 513004 334098 513186 334334
rect 513422 334098 513604 334334
rect 513004 298654 513604 334098
rect 513004 298418 513186 298654
rect 513422 298418 513604 298654
rect 513004 298334 513604 298418
rect 513004 298098 513186 298334
rect 513422 298098 513604 298334
rect 513004 262654 513604 298098
rect 513004 262418 513186 262654
rect 513422 262418 513604 262654
rect 513004 262334 513604 262418
rect 513004 262098 513186 262334
rect 513422 262098 513604 262334
rect 513004 226654 513604 262098
rect 513004 226418 513186 226654
rect 513422 226418 513604 226654
rect 513004 226334 513604 226418
rect 513004 226098 513186 226334
rect 513422 226098 513604 226334
rect 513004 190654 513604 226098
rect 513004 190418 513186 190654
rect 513422 190418 513604 190654
rect 513004 190334 513604 190418
rect 513004 190098 513186 190334
rect 513422 190098 513604 190334
rect 513004 154654 513604 190098
rect 513004 154418 513186 154654
rect 513422 154418 513604 154654
rect 513004 154334 513604 154418
rect 513004 154098 513186 154334
rect 513422 154098 513604 154334
rect 513004 118654 513604 154098
rect 513004 118418 513186 118654
rect 513422 118418 513604 118654
rect 513004 118334 513604 118418
rect 513004 118098 513186 118334
rect 513422 118098 513604 118334
rect 513004 82654 513604 118098
rect 513004 82418 513186 82654
rect 513422 82418 513604 82654
rect 513004 82334 513604 82418
rect 513004 82098 513186 82334
rect 513422 82098 513604 82334
rect 513004 46654 513604 82098
rect 513004 46418 513186 46654
rect 513422 46418 513604 46654
rect 513004 46334 513604 46418
rect 513004 46098 513186 46334
rect 513422 46098 513604 46334
rect 513004 10654 513604 46098
rect 513004 10418 513186 10654
rect 513422 10418 513604 10654
rect 513004 10334 513604 10418
rect 513004 10098 513186 10334
rect 513422 10098 513604 10334
rect 513004 -4106 513604 10098
rect 513004 -4342 513186 -4106
rect 513422 -4342 513604 -4106
rect 513004 -4426 513604 -4342
rect 513004 -4662 513186 -4426
rect 513422 -4662 513604 -4426
rect 513004 -5624 513604 -4662
rect 516604 698254 517204 709922
rect 534604 711418 535204 711440
rect 534604 711182 534786 711418
rect 535022 711182 535204 711418
rect 534604 711098 535204 711182
rect 534604 710862 534786 711098
rect 535022 710862 535204 711098
rect 531004 709538 531604 709560
rect 531004 709302 531186 709538
rect 531422 709302 531604 709538
rect 531004 709218 531604 709302
rect 531004 708982 531186 709218
rect 531422 708982 531604 709218
rect 527404 707658 528004 707680
rect 527404 707422 527586 707658
rect 527822 707422 528004 707658
rect 527404 707338 528004 707422
rect 527404 707102 527586 707338
rect 527822 707102 528004 707338
rect 516604 698018 516786 698254
rect 517022 698018 517204 698254
rect 516604 697934 517204 698018
rect 516604 697698 516786 697934
rect 517022 697698 517204 697934
rect 516604 662254 517204 697698
rect 516604 662018 516786 662254
rect 517022 662018 517204 662254
rect 516604 661934 517204 662018
rect 516604 661698 516786 661934
rect 517022 661698 517204 661934
rect 516604 626254 517204 661698
rect 516604 626018 516786 626254
rect 517022 626018 517204 626254
rect 516604 625934 517204 626018
rect 516604 625698 516786 625934
rect 517022 625698 517204 625934
rect 516604 590254 517204 625698
rect 516604 590018 516786 590254
rect 517022 590018 517204 590254
rect 516604 589934 517204 590018
rect 516604 589698 516786 589934
rect 517022 589698 517204 589934
rect 516604 554254 517204 589698
rect 516604 554018 516786 554254
rect 517022 554018 517204 554254
rect 516604 553934 517204 554018
rect 516604 553698 516786 553934
rect 517022 553698 517204 553934
rect 516604 518254 517204 553698
rect 516604 518018 516786 518254
rect 517022 518018 517204 518254
rect 516604 517934 517204 518018
rect 516604 517698 516786 517934
rect 517022 517698 517204 517934
rect 516604 482254 517204 517698
rect 516604 482018 516786 482254
rect 517022 482018 517204 482254
rect 516604 481934 517204 482018
rect 516604 481698 516786 481934
rect 517022 481698 517204 481934
rect 516604 446254 517204 481698
rect 516604 446018 516786 446254
rect 517022 446018 517204 446254
rect 516604 445934 517204 446018
rect 516604 445698 516786 445934
rect 517022 445698 517204 445934
rect 516604 410254 517204 445698
rect 516604 410018 516786 410254
rect 517022 410018 517204 410254
rect 516604 409934 517204 410018
rect 516604 409698 516786 409934
rect 517022 409698 517204 409934
rect 516604 374254 517204 409698
rect 516604 374018 516786 374254
rect 517022 374018 517204 374254
rect 516604 373934 517204 374018
rect 516604 373698 516786 373934
rect 517022 373698 517204 373934
rect 516604 338254 517204 373698
rect 516604 338018 516786 338254
rect 517022 338018 517204 338254
rect 516604 337934 517204 338018
rect 516604 337698 516786 337934
rect 517022 337698 517204 337934
rect 516604 302254 517204 337698
rect 516604 302018 516786 302254
rect 517022 302018 517204 302254
rect 516604 301934 517204 302018
rect 516604 301698 516786 301934
rect 517022 301698 517204 301934
rect 516604 266254 517204 301698
rect 516604 266018 516786 266254
rect 517022 266018 517204 266254
rect 516604 265934 517204 266018
rect 516604 265698 516786 265934
rect 517022 265698 517204 265934
rect 516604 230254 517204 265698
rect 516604 230018 516786 230254
rect 517022 230018 517204 230254
rect 516604 229934 517204 230018
rect 516604 229698 516786 229934
rect 517022 229698 517204 229934
rect 516604 194254 517204 229698
rect 516604 194018 516786 194254
rect 517022 194018 517204 194254
rect 516604 193934 517204 194018
rect 516604 193698 516786 193934
rect 517022 193698 517204 193934
rect 516604 158254 517204 193698
rect 516604 158018 516786 158254
rect 517022 158018 517204 158254
rect 516604 157934 517204 158018
rect 516604 157698 516786 157934
rect 517022 157698 517204 157934
rect 516604 122254 517204 157698
rect 516604 122018 516786 122254
rect 517022 122018 517204 122254
rect 516604 121934 517204 122018
rect 516604 121698 516786 121934
rect 517022 121698 517204 121934
rect 516604 86254 517204 121698
rect 516604 86018 516786 86254
rect 517022 86018 517204 86254
rect 516604 85934 517204 86018
rect 516604 85698 516786 85934
rect 517022 85698 517204 85934
rect 516604 50254 517204 85698
rect 516604 50018 516786 50254
rect 517022 50018 517204 50254
rect 516604 49934 517204 50018
rect 516604 49698 516786 49934
rect 517022 49698 517204 49934
rect 516604 14254 517204 49698
rect 516604 14018 516786 14254
rect 517022 14018 517204 14254
rect 516604 13934 517204 14018
rect 516604 13698 516786 13934
rect 517022 13698 517204 13934
rect 498604 -7162 498786 -6926
rect 499022 -7162 499204 -6926
rect 498604 -7246 499204 -7162
rect 498604 -7482 498786 -7246
rect 499022 -7482 499204 -7246
rect 498604 -7504 499204 -7482
rect 516604 -5986 517204 13698
rect 523804 705778 524404 705800
rect 523804 705542 523986 705778
rect 524222 705542 524404 705778
rect 523804 705458 524404 705542
rect 523804 705222 523986 705458
rect 524222 705222 524404 705458
rect 523804 669454 524404 705222
rect 523804 669218 523986 669454
rect 524222 669218 524404 669454
rect 523804 669134 524404 669218
rect 523804 668898 523986 669134
rect 524222 668898 524404 669134
rect 523804 633454 524404 668898
rect 523804 633218 523986 633454
rect 524222 633218 524404 633454
rect 523804 633134 524404 633218
rect 523804 632898 523986 633134
rect 524222 632898 524404 633134
rect 523804 597454 524404 632898
rect 523804 597218 523986 597454
rect 524222 597218 524404 597454
rect 523804 597134 524404 597218
rect 523804 596898 523986 597134
rect 524222 596898 524404 597134
rect 523804 561454 524404 596898
rect 523804 561218 523986 561454
rect 524222 561218 524404 561454
rect 523804 561134 524404 561218
rect 523804 560898 523986 561134
rect 524222 560898 524404 561134
rect 523804 525454 524404 560898
rect 523804 525218 523986 525454
rect 524222 525218 524404 525454
rect 523804 525134 524404 525218
rect 523804 524898 523986 525134
rect 524222 524898 524404 525134
rect 523804 489454 524404 524898
rect 523804 489218 523986 489454
rect 524222 489218 524404 489454
rect 523804 489134 524404 489218
rect 523804 488898 523986 489134
rect 524222 488898 524404 489134
rect 523804 453454 524404 488898
rect 523804 453218 523986 453454
rect 524222 453218 524404 453454
rect 523804 453134 524404 453218
rect 523804 452898 523986 453134
rect 524222 452898 524404 453134
rect 523804 417454 524404 452898
rect 523804 417218 523986 417454
rect 524222 417218 524404 417454
rect 523804 417134 524404 417218
rect 523804 416898 523986 417134
rect 524222 416898 524404 417134
rect 523804 381454 524404 416898
rect 523804 381218 523986 381454
rect 524222 381218 524404 381454
rect 523804 381134 524404 381218
rect 523804 380898 523986 381134
rect 524222 380898 524404 381134
rect 523804 345454 524404 380898
rect 523804 345218 523986 345454
rect 524222 345218 524404 345454
rect 523804 345134 524404 345218
rect 523804 344898 523986 345134
rect 524222 344898 524404 345134
rect 523804 309454 524404 344898
rect 523804 309218 523986 309454
rect 524222 309218 524404 309454
rect 523804 309134 524404 309218
rect 523804 308898 523986 309134
rect 524222 308898 524404 309134
rect 523804 273454 524404 308898
rect 523804 273218 523986 273454
rect 524222 273218 524404 273454
rect 523804 273134 524404 273218
rect 523804 272898 523986 273134
rect 524222 272898 524404 273134
rect 523804 237454 524404 272898
rect 523804 237218 523986 237454
rect 524222 237218 524404 237454
rect 523804 237134 524404 237218
rect 523804 236898 523986 237134
rect 524222 236898 524404 237134
rect 523804 201454 524404 236898
rect 523804 201218 523986 201454
rect 524222 201218 524404 201454
rect 523804 201134 524404 201218
rect 523804 200898 523986 201134
rect 524222 200898 524404 201134
rect 523804 165454 524404 200898
rect 523804 165218 523986 165454
rect 524222 165218 524404 165454
rect 523804 165134 524404 165218
rect 523804 164898 523986 165134
rect 524222 164898 524404 165134
rect 523804 129454 524404 164898
rect 523804 129218 523986 129454
rect 524222 129218 524404 129454
rect 523804 129134 524404 129218
rect 523804 128898 523986 129134
rect 524222 128898 524404 129134
rect 523804 93454 524404 128898
rect 523804 93218 523986 93454
rect 524222 93218 524404 93454
rect 523804 93134 524404 93218
rect 523804 92898 523986 93134
rect 524222 92898 524404 93134
rect 523804 57454 524404 92898
rect 523804 57218 523986 57454
rect 524222 57218 524404 57454
rect 523804 57134 524404 57218
rect 523804 56898 523986 57134
rect 524222 56898 524404 57134
rect 523804 21454 524404 56898
rect 523804 21218 523986 21454
rect 524222 21218 524404 21454
rect 523804 21134 524404 21218
rect 523804 20898 523986 21134
rect 524222 20898 524404 21134
rect 523804 -1286 524404 20898
rect 523804 -1522 523986 -1286
rect 524222 -1522 524404 -1286
rect 523804 -1606 524404 -1522
rect 523804 -1842 523986 -1606
rect 524222 -1842 524404 -1606
rect 523804 -1864 524404 -1842
rect 527404 673054 528004 707102
rect 527404 672818 527586 673054
rect 527822 672818 528004 673054
rect 527404 672734 528004 672818
rect 527404 672498 527586 672734
rect 527822 672498 528004 672734
rect 527404 637054 528004 672498
rect 527404 636818 527586 637054
rect 527822 636818 528004 637054
rect 527404 636734 528004 636818
rect 527404 636498 527586 636734
rect 527822 636498 528004 636734
rect 527404 601054 528004 636498
rect 527404 600818 527586 601054
rect 527822 600818 528004 601054
rect 527404 600734 528004 600818
rect 527404 600498 527586 600734
rect 527822 600498 528004 600734
rect 527404 565054 528004 600498
rect 527404 564818 527586 565054
rect 527822 564818 528004 565054
rect 527404 564734 528004 564818
rect 527404 564498 527586 564734
rect 527822 564498 528004 564734
rect 527404 529054 528004 564498
rect 527404 528818 527586 529054
rect 527822 528818 528004 529054
rect 527404 528734 528004 528818
rect 527404 528498 527586 528734
rect 527822 528498 528004 528734
rect 527404 493054 528004 528498
rect 527404 492818 527586 493054
rect 527822 492818 528004 493054
rect 527404 492734 528004 492818
rect 527404 492498 527586 492734
rect 527822 492498 528004 492734
rect 527404 457054 528004 492498
rect 527404 456818 527586 457054
rect 527822 456818 528004 457054
rect 527404 456734 528004 456818
rect 527404 456498 527586 456734
rect 527822 456498 528004 456734
rect 527404 421054 528004 456498
rect 527404 420818 527586 421054
rect 527822 420818 528004 421054
rect 527404 420734 528004 420818
rect 527404 420498 527586 420734
rect 527822 420498 528004 420734
rect 527404 385054 528004 420498
rect 527404 384818 527586 385054
rect 527822 384818 528004 385054
rect 527404 384734 528004 384818
rect 527404 384498 527586 384734
rect 527822 384498 528004 384734
rect 527404 349054 528004 384498
rect 527404 348818 527586 349054
rect 527822 348818 528004 349054
rect 527404 348734 528004 348818
rect 527404 348498 527586 348734
rect 527822 348498 528004 348734
rect 527404 313054 528004 348498
rect 527404 312818 527586 313054
rect 527822 312818 528004 313054
rect 527404 312734 528004 312818
rect 527404 312498 527586 312734
rect 527822 312498 528004 312734
rect 527404 277054 528004 312498
rect 527404 276818 527586 277054
rect 527822 276818 528004 277054
rect 527404 276734 528004 276818
rect 527404 276498 527586 276734
rect 527822 276498 528004 276734
rect 527404 241054 528004 276498
rect 527404 240818 527586 241054
rect 527822 240818 528004 241054
rect 527404 240734 528004 240818
rect 527404 240498 527586 240734
rect 527822 240498 528004 240734
rect 527404 205054 528004 240498
rect 527404 204818 527586 205054
rect 527822 204818 528004 205054
rect 527404 204734 528004 204818
rect 527404 204498 527586 204734
rect 527822 204498 528004 204734
rect 527404 169054 528004 204498
rect 527404 168818 527586 169054
rect 527822 168818 528004 169054
rect 527404 168734 528004 168818
rect 527404 168498 527586 168734
rect 527822 168498 528004 168734
rect 527404 133054 528004 168498
rect 527404 132818 527586 133054
rect 527822 132818 528004 133054
rect 527404 132734 528004 132818
rect 527404 132498 527586 132734
rect 527822 132498 528004 132734
rect 527404 97054 528004 132498
rect 527404 96818 527586 97054
rect 527822 96818 528004 97054
rect 527404 96734 528004 96818
rect 527404 96498 527586 96734
rect 527822 96498 528004 96734
rect 527404 61054 528004 96498
rect 527404 60818 527586 61054
rect 527822 60818 528004 61054
rect 527404 60734 528004 60818
rect 527404 60498 527586 60734
rect 527822 60498 528004 60734
rect 527404 25054 528004 60498
rect 527404 24818 527586 25054
rect 527822 24818 528004 25054
rect 527404 24734 528004 24818
rect 527404 24498 527586 24734
rect 527822 24498 528004 24734
rect 527404 -3166 528004 24498
rect 527404 -3402 527586 -3166
rect 527822 -3402 528004 -3166
rect 527404 -3486 528004 -3402
rect 527404 -3722 527586 -3486
rect 527822 -3722 528004 -3486
rect 527404 -3744 528004 -3722
rect 531004 676654 531604 708982
rect 531004 676418 531186 676654
rect 531422 676418 531604 676654
rect 531004 676334 531604 676418
rect 531004 676098 531186 676334
rect 531422 676098 531604 676334
rect 531004 640654 531604 676098
rect 531004 640418 531186 640654
rect 531422 640418 531604 640654
rect 531004 640334 531604 640418
rect 531004 640098 531186 640334
rect 531422 640098 531604 640334
rect 531004 604654 531604 640098
rect 531004 604418 531186 604654
rect 531422 604418 531604 604654
rect 531004 604334 531604 604418
rect 531004 604098 531186 604334
rect 531422 604098 531604 604334
rect 531004 568654 531604 604098
rect 531004 568418 531186 568654
rect 531422 568418 531604 568654
rect 531004 568334 531604 568418
rect 531004 568098 531186 568334
rect 531422 568098 531604 568334
rect 531004 532654 531604 568098
rect 531004 532418 531186 532654
rect 531422 532418 531604 532654
rect 531004 532334 531604 532418
rect 531004 532098 531186 532334
rect 531422 532098 531604 532334
rect 531004 496654 531604 532098
rect 531004 496418 531186 496654
rect 531422 496418 531604 496654
rect 531004 496334 531604 496418
rect 531004 496098 531186 496334
rect 531422 496098 531604 496334
rect 531004 460654 531604 496098
rect 531004 460418 531186 460654
rect 531422 460418 531604 460654
rect 531004 460334 531604 460418
rect 531004 460098 531186 460334
rect 531422 460098 531604 460334
rect 531004 424654 531604 460098
rect 531004 424418 531186 424654
rect 531422 424418 531604 424654
rect 531004 424334 531604 424418
rect 531004 424098 531186 424334
rect 531422 424098 531604 424334
rect 531004 388654 531604 424098
rect 531004 388418 531186 388654
rect 531422 388418 531604 388654
rect 531004 388334 531604 388418
rect 531004 388098 531186 388334
rect 531422 388098 531604 388334
rect 531004 352654 531604 388098
rect 531004 352418 531186 352654
rect 531422 352418 531604 352654
rect 531004 352334 531604 352418
rect 531004 352098 531186 352334
rect 531422 352098 531604 352334
rect 531004 316654 531604 352098
rect 531004 316418 531186 316654
rect 531422 316418 531604 316654
rect 531004 316334 531604 316418
rect 531004 316098 531186 316334
rect 531422 316098 531604 316334
rect 531004 280654 531604 316098
rect 531004 280418 531186 280654
rect 531422 280418 531604 280654
rect 531004 280334 531604 280418
rect 531004 280098 531186 280334
rect 531422 280098 531604 280334
rect 531004 244654 531604 280098
rect 531004 244418 531186 244654
rect 531422 244418 531604 244654
rect 531004 244334 531604 244418
rect 531004 244098 531186 244334
rect 531422 244098 531604 244334
rect 531004 208654 531604 244098
rect 531004 208418 531186 208654
rect 531422 208418 531604 208654
rect 531004 208334 531604 208418
rect 531004 208098 531186 208334
rect 531422 208098 531604 208334
rect 531004 172654 531604 208098
rect 531004 172418 531186 172654
rect 531422 172418 531604 172654
rect 531004 172334 531604 172418
rect 531004 172098 531186 172334
rect 531422 172098 531604 172334
rect 531004 136654 531604 172098
rect 531004 136418 531186 136654
rect 531422 136418 531604 136654
rect 531004 136334 531604 136418
rect 531004 136098 531186 136334
rect 531422 136098 531604 136334
rect 531004 100654 531604 136098
rect 531004 100418 531186 100654
rect 531422 100418 531604 100654
rect 531004 100334 531604 100418
rect 531004 100098 531186 100334
rect 531422 100098 531604 100334
rect 531004 64654 531604 100098
rect 531004 64418 531186 64654
rect 531422 64418 531604 64654
rect 531004 64334 531604 64418
rect 531004 64098 531186 64334
rect 531422 64098 531604 64334
rect 531004 28654 531604 64098
rect 531004 28418 531186 28654
rect 531422 28418 531604 28654
rect 531004 28334 531604 28418
rect 531004 28098 531186 28334
rect 531422 28098 531604 28334
rect 531004 -5046 531604 28098
rect 531004 -5282 531186 -5046
rect 531422 -5282 531604 -5046
rect 531004 -5366 531604 -5282
rect 531004 -5602 531186 -5366
rect 531422 -5602 531604 -5366
rect 531004 -5624 531604 -5602
rect 534604 680254 535204 710862
rect 552604 710478 553204 711440
rect 552604 710242 552786 710478
rect 553022 710242 553204 710478
rect 552604 710158 553204 710242
rect 552604 709922 552786 710158
rect 553022 709922 553204 710158
rect 549004 708598 549604 709560
rect 549004 708362 549186 708598
rect 549422 708362 549604 708598
rect 549004 708278 549604 708362
rect 549004 708042 549186 708278
rect 549422 708042 549604 708278
rect 545404 706718 546004 707680
rect 545404 706482 545586 706718
rect 545822 706482 546004 706718
rect 545404 706398 546004 706482
rect 545404 706162 545586 706398
rect 545822 706162 546004 706398
rect 534604 680018 534786 680254
rect 535022 680018 535204 680254
rect 534604 679934 535204 680018
rect 534604 679698 534786 679934
rect 535022 679698 535204 679934
rect 534604 644254 535204 679698
rect 534604 644018 534786 644254
rect 535022 644018 535204 644254
rect 534604 643934 535204 644018
rect 534604 643698 534786 643934
rect 535022 643698 535204 643934
rect 534604 608254 535204 643698
rect 534604 608018 534786 608254
rect 535022 608018 535204 608254
rect 534604 607934 535204 608018
rect 534604 607698 534786 607934
rect 535022 607698 535204 607934
rect 534604 572254 535204 607698
rect 534604 572018 534786 572254
rect 535022 572018 535204 572254
rect 534604 571934 535204 572018
rect 534604 571698 534786 571934
rect 535022 571698 535204 571934
rect 534604 536254 535204 571698
rect 534604 536018 534786 536254
rect 535022 536018 535204 536254
rect 534604 535934 535204 536018
rect 534604 535698 534786 535934
rect 535022 535698 535204 535934
rect 534604 500254 535204 535698
rect 534604 500018 534786 500254
rect 535022 500018 535204 500254
rect 534604 499934 535204 500018
rect 534604 499698 534786 499934
rect 535022 499698 535204 499934
rect 534604 464254 535204 499698
rect 534604 464018 534786 464254
rect 535022 464018 535204 464254
rect 534604 463934 535204 464018
rect 534604 463698 534786 463934
rect 535022 463698 535204 463934
rect 534604 428254 535204 463698
rect 534604 428018 534786 428254
rect 535022 428018 535204 428254
rect 534604 427934 535204 428018
rect 534604 427698 534786 427934
rect 535022 427698 535204 427934
rect 534604 392254 535204 427698
rect 534604 392018 534786 392254
rect 535022 392018 535204 392254
rect 534604 391934 535204 392018
rect 534604 391698 534786 391934
rect 535022 391698 535204 391934
rect 534604 356254 535204 391698
rect 534604 356018 534786 356254
rect 535022 356018 535204 356254
rect 534604 355934 535204 356018
rect 534604 355698 534786 355934
rect 535022 355698 535204 355934
rect 534604 320254 535204 355698
rect 534604 320018 534786 320254
rect 535022 320018 535204 320254
rect 534604 319934 535204 320018
rect 534604 319698 534786 319934
rect 535022 319698 535204 319934
rect 534604 284254 535204 319698
rect 534604 284018 534786 284254
rect 535022 284018 535204 284254
rect 534604 283934 535204 284018
rect 534604 283698 534786 283934
rect 535022 283698 535204 283934
rect 534604 248254 535204 283698
rect 534604 248018 534786 248254
rect 535022 248018 535204 248254
rect 534604 247934 535204 248018
rect 534604 247698 534786 247934
rect 535022 247698 535204 247934
rect 534604 212254 535204 247698
rect 534604 212018 534786 212254
rect 535022 212018 535204 212254
rect 534604 211934 535204 212018
rect 534604 211698 534786 211934
rect 535022 211698 535204 211934
rect 534604 176254 535204 211698
rect 534604 176018 534786 176254
rect 535022 176018 535204 176254
rect 534604 175934 535204 176018
rect 534604 175698 534786 175934
rect 535022 175698 535204 175934
rect 534604 140254 535204 175698
rect 534604 140018 534786 140254
rect 535022 140018 535204 140254
rect 534604 139934 535204 140018
rect 534604 139698 534786 139934
rect 535022 139698 535204 139934
rect 534604 104254 535204 139698
rect 534604 104018 534786 104254
rect 535022 104018 535204 104254
rect 534604 103934 535204 104018
rect 534604 103698 534786 103934
rect 535022 103698 535204 103934
rect 534604 68254 535204 103698
rect 534604 68018 534786 68254
rect 535022 68018 535204 68254
rect 534604 67934 535204 68018
rect 534604 67698 534786 67934
rect 535022 67698 535204 67934
rect 534604 32254 535204 67698
rect 534604 32018 534786 32254
rect 535022 32018 535204 32254
rect 534604 31934 535204 32018
rect 534604 31698 534786 31934
rect 535022 31698 535204 31934
rect 516604 -6222 516786 -5986
rect 517022 -6222 517204 -5986
rect 516604 -6306 517204 -6222
rect 516604 -6542 516786 -6306
rect 517022 -6542 517204 -6306
rect 516604 -7504 517204 -6542
rect 534604 -6926 535204 31698
rect 541804 704838 542404 705800
rect 541804 704602 541986 704838
rect 542222 704602 542404 704838
rect 541804 704518 542404 704602
rect 541804 704282 541986 704518
rect 542222 704282 542404 704518
rect 541804 687454 542404 704282
rect 541804 687218 541986 687454
rect 542222 687218 542404 687454
rect 541804 687134 542404 687218
rect 541804 686898 541986 687134
rect 542222 686898 542404 687134
rect 541804 651454 542404 686898
rect 541804 651218 541986 651454
rect 542222 651218 542404 651454
rect 541804 651134 542404 651218
rect 541804 650898 541986 651134
rect 542222 650898 542404 651134
rect 541804 615454 542404 650898
rect 541804 615218 541986 615454
rect 542222 615218 542404 615454
rect 541804 615134 542404 615218
rect 541804 614898 541986 615134
rect 542222 614898 542404 615134
rect 541804 579454 542404 614898
rect 541804 579218 541986 579454
rect 542222 579218 542404 579454
rect 541804 579134 542404 579218
rect 541804 578898 541986 579134
rect 542222 578898 542404 579134
rect 541804 543454 542404 578898
rect 541804 543218 541986 543454
rect 542222 543218 542404 543454
rect 541804 543134 542404 543218
rect 541804 542898 541986 543134
rect 542222 542898 542404 543134
rect 541804 507454 542404 542898
rect 541804 507218 541986 507454
rect 542222 507218 542404 507454
rect 541804 507134 542404 507218
rect 541804 506898 541986 507134
rect 542222 506898 542404 507134
rect 541804 471454 542404 506898
rect 541804 471218 541986 471454
rect 542222 471218 542404 471454
rect 541804 471134 542404 471218
rect 541804 470898 541986 471134
rect 542222 470898 542404 471134
rect 541804 435454 542404 470898
rect 541804 435218 541986 435454
rect 542222 435218 542404 435454
rect 541804 435134 542404 435218
rect 541804 434898 541986 435134
rect 542222 434898 542404 435134
rect 541804 399454 542404 434898
rect 541804 399218 541986 399454
rect 542222 399218 542404 399454
rect 541804 399134 542404 399218
rect 541804 398898 541986 399134
rect 542222 398898 542404 399134
rect 541804 363454 542404 398898
rect 541804 363218 541986 363454
rect 542222 363218 542404 363454
rect 541804 363134 542404 363218
rect 541804 362898 541986 363134
rect 542222 362898 542404 363134
rect 541804 327454 542404 362898
rect 541804 327218 541986 327454
rect 542222 327218 542404 327454
rect 541804 327134 542404 327218
rect 541804 326898 541986 327134
rect 542222 326898 542404 327134
rect 541804 291454 542404 326898
rect 541804 291218 541986 291454
rect 542222 291218 542404 291454
rect 541804 291134 542404 291218
rect 541804 290898 541986 291134
rect 542222 290898 542404 291134
rect 541804 255454 542404 290898
rect 541804 255218 541986 255454
rect 542222 255218 542404 255454
rect 541804 255134 542404 255218
rect 541804 254898 541986 255134
rect 542222 254898 542404 255134
rect 541804 219454 542404 254898
rect 541804 219218 541986 219454
rect 542222 219218 542404 219454
rect 541804 219134 542404 219218
rect 541804 218898 541986 219134
rect 542222 218898 542404 219134
rect 541804 183454 542404 218898
rect 541804 183218 541986 183454
rect 542222 183218 542404 183454
rect 541804 183134 542404 183218
rect 541804 182898 541986 183134
rect 542222 182898 542404 183134
rect 541804 147454 542404 182898
rect 541804 147218 541986 147454
rect 542222 147218 542404 147454
rect 541804 147134 542404 147218
rect 541804 146898 541986 147134
rect 542222 146898 542404 147134
rect 541804 111454 542404 146898
rect 541804 111218 541986 111454
rect 542222 111218 542404 111454
rect 541804 111134 542404 111218
rect 541804 110898 541986 111134
rect 542222 110898 542404 111134
rect 541804 75454 542404 110898
rect 541804 75218 541986 75454
rect 542222 75218 542404 75454
rect 541804 75134 542404 75218
rect 541804 74898 541986 75134
rect 542222 74898 542404 75134
rect 541804 39454 542404 74898
rect 541804 39218 541986 39454
rect 542222 39218 542404 39454
rect 541804 39134 542404 39218
rect 541804 38898 541986 39134
rect 542222 38898 542404 39134
rect 541804 3454 542404 38898
rect 541804 3218 541986 3454
rect 542222 3218 542404 3454
rect 541804 3134 542404 3218
rect 541804 2898 541986 3134
rect 542222 2898 542404 3134
rect 541804 -346 542404 2898
rect 541804 -582 541986 -346
rect 542222 -582 542404 -346
rect 541804 -666 542404 -582
rect 541804 -902 541986 -666
rect 542222 -902 542404 -666
rect 541804 -1864 542404 -902
rect 545404 691054 546004 706162
rect 545404 690818 545586 691054
rect 545822 690818 546004 691054
rect 545404 690734 546004 690818
rect 545404 690498 545586 690734
rect 545822 690498 546004 690734
rect 545404 655054 546004 690498
rect 545404 654818 545586 655054
rect 545822 654818 546004 655054
rect 545404 654734 546004 654818
rect 545404 654498 545586 654734
rect 545822 654498 546004 654734
rect 545404 619054 546004 654498
rect 545404 618818 545586 619054
rect 545822 618818 546004 619054
rect 545404 618734 546004 618818
rect 545404 618498 545586 618734
rect 545822 618498 546004 618734
rect 545404 583054 546004 618498
rect 545404 582818 545586 583054
rect 545822 582818 546004 583054
rect 545404 582734 546004 582818
rect 545404 582498 545586 582734
rect 545822 582498 546004 582734
rect 545404 547054 546004 582498
rect 545404 546818 545586 547054
rect 545822 546818 546004 547054
rect 545404 546734 546004 546818
rect 545404 546498 545586 546734
rect 545822 546498 546004 546734
rect 545404 511054 546004 546498
rect 545404 510818 545586 511054
rect 545822 510818 546004 511054
rect 545404 510734 546004 510818
rect 545404 510498 545586 510734
rect 545822 510498 546004 510734
rect 545404 475054 546004 510498
rect 545404 474818 545586 475054
rect 545822 474818 546004 475054
rect 545404 474734 546004 474818
rect 545404 474498 545586 474734
rect 545822 474498 546004 474734
rect 545404 439054 546004 474498
rect 545404 438818 545586 439054
rect 545822 438818 546004 439054
rect 545404 438734 546004 438818
rect 545404 438498 545586 438734
rect 545822 438498 546004 438734
rect 545404 403054 546004 438498
rect 545404 402818 545586 403054
rect 545822 402818 546004 403054
rect 545404 402734 546004 402818
rect 545404 402498 545586 402734
rect 545822 402498 546004 402734
rect 545404 367054 546004 402498
rect 545404 366818 545586 367054
rect 545822 366818 546004 367054
rect 545404 366734 546004 366818
rect 545404 366498 545586 366734
rect 545822 366498 546004 366734
rect 545404 331054 546004 366498
rect 545404 330818 545586 331054
rect 545822 330818 546004 331054
rect 545404 330734 546004 330818
rect 545404 330498 545586 330734
rect 545822 330498 546004 330734
rect 545404 295054 546004 330498
rect 545404 294818 545586 295054
rect 545822 294818 546004 295054
rect 545404 294734 546004 294818
rect 545404 294498 545586 294734
rect 545822 294498 546004 294734
rect 545404 259054 546004 294498
rect 545404 258818 545586 259054
rect 545822 258818 546004 259054
rect 545404 258734 546004 258818
rect 545404 258498 545586 258734
rect 545822 258498 546004 258734
rect 545404 223054 546004 258498
rect 545404 222818 545586 223054
rect 545822 222818 546004 223054
rect 545404 222734 546004 222818
rect 545404 222498 545586 222734
rect 545822 222498 546004 222734
rect 545404 187054 546004 222498
rect 545404 186818 545586 187054
rect 545822 186818 546004 187054
rect 545404 186734 546004 186818
rect 545404 186498 545586 186734
rect 545822 186498 546004 186734
rect 545404 151054 546004 186498
rect 545404 150818 545586 151054
rect 545822 150818 546004 151054
rect 545404 150734 546004 150818
rect 545404 150498 545586 150734
rect 545822 150498 546004 150734
rect 545404 115054 546004 150498
rect 545404 114818 545586 115054
rect 545822 114818 546004 115054
rect 545404 114734 546004 114818
rect 545404 114498 545586 114734
rect 545822 114498 546004 114734
rect 545404 79054 546004 114498
rect 545404 78818 545586 79054
rect 545822 78818 546004 79054
rect 545404 78734 546004 78818
rect 545404 78498 545586 78734
rect 545822 78498 546004 78734
rect 545404 43054 546004 78498
rect 545404 42818 545586 43054
rect 545822 42818 546004 43054
rect 545404 42734 546004 42818
rect 545404 42498 545586 42734
rect 545822 42498 546004 42734
rect 545404 7054 546004 42498
rect 545404 6818 545586 7054
rect 545822 6818 546004 7054
rect 545404 6734 546004 6818
rect 545404 6498 545586 6734
rect 545822 6498 546004 6734
rect 545404 -2226 546004 6498
rect 545404 -2462 545586 -2226
rect 545822 -2462 546004 -2226
rect 545404 -2546 546004 -2462
rect 545404 -2782 545586 -2546
rect 545822 -2782 546004 -2546
rect 545404 -3744 546004 -2782
rect 549004 694654 549604 708042
rect 549004 694418 549186 694654
rect 549422 694418 549604 694654
rect 549004 694334 549604 694418
rect 549004 694098 549186 694334
rect 549422 694098 549604 694334
rect 549004 658654 549604 694098
rect 549004 658418 549186 658654
rect 549422 658418 549604 658654
rect 549004 658334 549604 658418
rect 549004 658098 549186 658334
rect 549422 658098 549604 658334
rect 549004 622654 549604 658098
rect 549004 622418 549186 622654
rect 549422 622418 549604 622654
rect 549004 622334 549604 622418
rect 549004 622098 549186 622334
rect 549422 622098 549604 622334
rect 549004 586654 549604 622098
rect 549004 586418 549186 586654
rect 549422 586418 549604 586654
rect 549004 586334 549604 586418
rect 549004 586098 549186 586334
rect 549422 586098 549604 586334
rect 549004 550654 549604 586098
rect 549004 550418 549186 550654
rect 549422 550418 549604 550654
rect 549004 550334 549604 550418
rect 549004 550098 549186 550334
rect 549422 550098 549604 550334
rect 549004 514654 549604 550098
rect 549004 514418 549186 514654
rect 549422 514418 549604 514654
rect 549004 514334 549604 514418
rect 549004 514098 549186 514334
rect 549422 514098 549604 514334
rect 549004 478654 549604 514098
rect 549004 478418 549186 478654
rect 549422 478418 549604 478654
rect 549004 478334 549604 478418
rect 549004 478098 549186 478334
rect 549422 478098 549604 478334
rect 549004 442654 549604 478098
rect 549004 442418 549186 442654
rect 549422 442418 549604 442654
rect 549004 442334 549604 442418
rect 549004 442098 549186 442334
rect 549422 442098 549604 442334
rect 549004 406654 549604 442098
rect 549004 406418 549186 406654
rect 549422 406418 549604 406654
rect 549004 406334 549604 406418
rect 549004 406098 549186 406334
rect 549422 406098 549604 406334
rect 549004 370654 549604 406098
rect 549004 370418 549186 370654
rect 549422 370418 549604 370654
rect 549004 370334 549604 370418
rect 549004 370098 549186 370334
rect 549422 370098 549604 370334
rect 549004 334654 549604 370098
rect 549004 334418 549186 334654
rect 549422 334418 549604 334654
rect 549004 334334 549604 334418
rect 549004 334098 549186 334334
rect 549422 334098 549604 334334
rect 549004 298654 549604 334098
rect 549004 298418 549186 298654
rect 549422 298418 549604 298654
rect 549004 298334 549604 298418
rect 549004 298098 549186 298334
rect 549422 298098 549604 298334
rect 549004 262654 549604 298098
rect 549004 262418 549186 262654
rect 549422 262418 549604 262654
rect 549004 262334 549604 262418
rect 549004 262098 549186 262334
rect 549422 262098 549604 262334
rect 549004 226654 549604 262098
rect 549004 226418 549186 226654
rect 549422 226418 549604 226654
rect 549004 226334 549604 226418
rect 549004 226098 549186 226334
rect 549422 226098 549604 226334
rect 549004 190654 549604 226098
rect 549004 190418 549186 190654
rect 549422 190418 549604 190654
rect 549004 190334 549604 190418
rect 549004 190098 549186 190334
rect 549422 190098 549604 190334
rect 549004 154654 549604 190098
rect 549004 154418 549186 154654
rect 549422 154418 549604 154654
rect 549004 154334 549604 154418
rect 549004 154098 549186 154334
rect 549422 154098 549604 154334
rect 549004 118654 549604 154098
rect 549004 118418 549186 118654
rect 549422 118418 549604 118654
rect 549004 118334 549604 118418
rect 549004 118098 549186 118334
rect 549422 118098 549604 118334
rect 549004 82654 549604 118098
rect 549004 82418 549186 82654
rect 549422 82418 549604 82654
rect 549004 82334 549604 82418
rect 549004 82098 549186 82334
rect 549422 82098 549604 82334
rect 549004 46654 549604 82098
rect 549004 46418 549186 46654
rect 549422 46418 549604 46654
rect 549004 46334 549604 46418
rect 549004 46098 549186 46334
rect 549422 46098 549604 46334
rect 549004 10654 549604 46098
rect 549004 10418 549186 10654
rect 549422 10418 549604 10654
rect 549004 10334 549604 10418
rect 549004 10098 549186 10334
rect 549422 10098 549604 10334
rect 549004 -4106 549604 10098
rect 549004 -4342 549186 -4106
rect 549422 -4342 549604 -4106
rect 549004 -4426 549604 -4342
rect 549004 -4662 549186 -4426
rect 549422 -4662 549604 -4426
rect 549004 -5624 549604 -4662
rect 552604 698254 553204 709922
rect 570604 711418 571204 711440
rect 570604 711182 570786 711418
rect 571022 711182 571204 711418
rect 570604 711098 571204 711182
rect 570604 710862 570786 711098
rect 571022 710862 571204 711098
rect 567004 709538 567604 709560
rect 567004 709302 567186 709538
rect 567422 709302 567604 709538
rect 567004 709218 567604 709302
rect 567004 708982 567186 709218
rect 567422 708982 567604 709218
rect 563404 707658 564004 707680
rect 563404 707422 563586 707658
rect 563822 707422 564004 707658
rect 563404 707338 564004 707422
rect 563404 707102 563586 707338
rect 563822 707102 564004 707338
rect 552604 698018 552786 698254
rect 553022 698018 553204 698254
rect 552604 697934 553204 698018
rect 552604 697698 552786 697934
rect 553022 697698 553204 697934
rect 552604 662254 553204 697698
rect 552604 662018 552786 662254
rect 553022 662018 553204 662254
rect 552604 661934 553204 662018
rect 552604 661698 552786 661934
rect 553022 661698 553204 661934
rect 552604 626254 553204 661698
rect 552604 626018 552786 626254
rect 553022 626018 553204 626254
rect 552604 625934 553204 626018
rect 552604 625698 552786 625934
rect 553022 625698 553204 625934
rect 552604 590254 553204 625698
rect 552604 590018 552786 590254
rect 553022 590018 553204 590254
rect 552604 589934 553204 590018
rect 552604 589698 552786 589934
rect 553022 589698 553204 589934
rect 552604 554254 553204 589698
rect 552604 554018 552786 554254
rect 553022 554018 553204 554254
rect 552604 553934 553204 554018
rect 552604 553698 552786 553934
rect 553022 553698 553204 553934
rect 552604 518254 553204 553698
rect 552604 518018 552786 518254
rect 553022 518018 553204 518254
rect 552604 517934 553204 518018
rect 552604 517698 552786 517934
rect 553022 517698 553204 517934
rect 552604 482254 553204 517698
rect 552604 482018 552786 482254
rect 553022 482018 553204 482254
rect 552604 481934 553204 482018
rect 552604 481698 552786 481934
rect 553022 481698 553204 481934
rect 552604 446254 553204 481698
rect 552604 446018 552786 446254
rect 553022 446018 553204 446254
rect 552604 445934 553204 446018
rect 552604 445698 552786 445934
rect 553022 445698 553204 445934
rect 552604 410254 553204 445698
rect 552604 410018 552786 410254
rect 553022 410018 553204 410254
rect 552604 409934 553204 410018
rect 552604 409698 552786 409934
rect 553022 409698 553204 409934
rect 552604 374254 553204 409698
rect 552604 374018 552786 374254
rect 553022 374018 553204 374254
rect 552604 373934 553204 374018
rect 552604 373698 552786 373934
rect 553022 373698 553204 373934
rect 552604 338254 553204 373698
rect 552604 338018 552786 338254
rect 553022 338018 553204 338254
rect 552604 337934 553204 338018
rect 552604 337698 552786 337934
rect 553022 337698 553204 337934
rect 552604 302254 553204 337698
rect 552604 302018 552786 302254
rect 553022 302018 553204 302254
rect 552604 301934 553204 302018
rect 552604 301698 552786 301934
rect 553022 301698 553204 301934
rect 552604 266254 553204 301698
rect 552604 266018 552786 266254
rect 553022 266018 553204 266254
rect 552604 265934 553204 266018
rect 552604 265698 552786 265934
rect 553022 265698 553204 265934
rect 552604 230254 553204 265698
rect 552604 230018 552786 230254
rect 553022 230018 553204 230254
rect 552604 229934 553204 230018
rect 552604 229698 552786 229934
rect 553022 229698 553204 229934
rect 552604 194254 553204 229698
rect 552604 194018 552786 194254
rect 553022 194018 553204 194254
rect 552604 193934 553204 194018
rect 552604 193698 552786 193934
rect 553022 193698 553204 193934
rect 552604 158254 553204 193698
rect 552604 158018 552786 158254
rect 553022 158018 553204 158254
rect 552604 157934 553204 158018
rect 552604 157698 552786 157934
rect 553022 157698 553204 157934
rect 552604 122254 553204 157698
rect 552604 122018 552786 122254
rect 553022 122018 553204 122254
rect 552604 121934 553204 122018
rect 552604 121698 552786 121934
rect 553022 121698 553204 121934
rect 552604 86254 553204 121698
rect 552604 86018 552786 86254
rect 553022 86018 553204 86254
rect 552604 85934 553204 86018
rect 552604 85698 552786 85934
rect 553022 85698 553204 85934
rect 552604 50254 553204 85698
rect 552604 50018 552786 50254
rect 553022 50018 553204 50254
rect 552604 49934 553204 50018
rect 552604 49698 552786 49934
rect 553022 49698 553204 49934
rect 552604 14254 553204 49698
rect 552604 14018 552786 14254
rect 553022 14018 553204 14254
rect 552604 13934 553204 14018
rect 552604 13698 552786 13934
rect 553022 13698 553204 13934
rect 534604 -7162 534786 -6926
rect 535022 -7162 535204 -6926
rect 534604 -7246 535204 -7162
rect 534604 -7482 534786 -7246
rect 535022 -7482 535204 -7246
rect 534604 -7504 535204 -7482
rect 552604 -5986 553204 13698
rect 559804 705778 560404 705800
rect 559804 705542 559986 705778
rect 560222 705542 560404 705778
rect 559804 705458 560404 705542
rect 559804 705222 559986 705458
rect 560222 705222 560404 705458
rect 559804 669454 560404 705222
rect 559804 669218 559986 669454
rect 560222 669218 560404 669454
rect 559804 669134 560404 669218
rect 559804 668898 559986 669134
rect 560222 668898 560404 669134
rect 559804 633454 560404 668898
rect 559804 633218 559986 633454
rect 560222 633218 560404 633454
rect 559804 633134 560404 633218
rect 559804 632898 559986 633134
rect 560222 632898 560404 633134
rect 559804 597454 560404 632898
rect 559804 597218 559986 597454
rect 560222 597218 560404 597454
rect 559804 597134 560404 597218
rect 559804 596898 559986 597134
rect 560222 596898 560404 597134
rect 559804 561454 560404 596898
rect 559804 561218 559986 561454
rect 560222 561218 560404 561454
rect 559804 561134 560404 561218
rect 559804 560898 559986 561134
rect 560222 560898 560404 561134
rect 559804 525454 560404 560898
rect 559804 525218 559986 525454
rect 560222 525218 560404 525454
rect 559804 525134 560404 525218
rect 559804 524898 559986 525134
rect 560222 524898 560404 525134
rect 559804 489454 560404 524898
rect 559804 489218 559986 489454
rect 560222 489218 560404 489454
rect 559804 489134 560404 489218
rect 559804 488898 559986 489134
rect 560222 488898 560404 489134
rect 559804 453454 560404 488898
rect 559804 453218 559986 453454
rect 560222 453218 560404 453454
rect 559804 453134 560404 453218
rect 559804 452898 559986 453134
rect 560222 452898 560404 453134
rect 559804 417454 560404 452898
rect 559804 417218 559986 417454
rect 560222 417218 560404 417454
rect 559804 417134 560404 417218
rect 559804 416898 559986 417134
rect 560222 416898 560404 417134
rect 559804 381454 560404 416898
rect 559804 381218 559986 381454
rect 560222 381218 560404 381454
rect 559804 381134 560404 381218
rect 559804 380898 559986 381134
rect 560222 380898 560404 381134
rect 559804 345454 560404 380898
rect 559804 345218 559986 345454
rect 560222 345218 560404 345454
rect 559804 345134 560404 345218
rect 559804 344898 559986 345134
rect 560222 344898 560404 345134
rect 559804 309454 560404 344898
rect 559804 309218 559986 309454
rect 560222 309218 560404 309454
rect 559804 309134 560404 309218
rect 559804 308898 559986 309134
rect 560222 308898 560404 309134
rect 559804 273454 560404 308898
rect 559804 273218 559986 273454
rect 560222 273218 560404 273454
rect 559804 273134 560404 273218
rect 559804 272898 559986 273134
rect 560222 272898 560404 273134
rect 559804 237454 560404 272898
rect 559804 237218 559986 237454
rect 560222 237218 560404 237454
rect 559804 237134 560404 237218
rect 559804 236898 559986 237134
rect 560222 236898 560404 237134
rect 559804 201454 560404 236898
rect 559804 201218 559986 201454
rect 560222 201218 560404 201454
rect 559804 201134 560404 201218
rect 559804 200898 559986 201134
rect 560222 200898 560404 201134
rect 559804 165454 560404 200898
rect 559804 165218 559986 165454
rect 560222 165218 560404 165454
rect 559804 165134 560404 165218
rect 559804 164898 559986 165134
rect 560222 164898 560404 165134
rect 559804 129454 560404 164898
rect 559804 129218 559986 129454
rect 560222 129218 560404 129454
rect 559804 129134 560404 129218
rect 559804 128898 559986 129134
rect 560222 128898 560404 129134
rect 559804 93454 560404 128898
rect 559804 93218 559986 93454
rect 560222 93218 560404 93454
rect 559804 93134 560404 93218
rect 559804 92898 559986 93134
rect 560222 92898 560404 93134
rect 559804 57454 560404 92898
rect 559804 57218 559986 57454
rect 560222 57218 560404 57454
rect 559804 57134 560404 57218
rect 559804 56898 559986 57134
rect 560222 56898 560404 57134
rect 559804 21454 560404 56898
rect 559804 21218 559986 21454
rect 560222 21218 560404 21454
rect 559804 21134 560404 21218
rect 559804 20898 559986 21134
rect 560222 20898 560404 21134
rect 559804 -1286 560404 20898
rect 559804 -1522 559986 -1286
rect 560222 -1522 560404 -1286
rect 559804 -1606 560404 -1522
rect 559804 -1842 559986 -1606
rect 560222 -1842 560404 -1606
rect 559804 -1864 560404 -1842
rect 563404 673054 564004 707102
rect 563404 672818 563586 673054
rect 563822 672818 564004 673054
rect 563404 672734 564004 672818
rect 563404 672498 563586 672734
rect 563822 672498 564004 672734
rect 563404 637054 564004 672498
rect 563404 636818 563586 637054
rect 563822 636818 564004 637054
rect 563404 636734 564004 636818
rect 563404 636498 563586 636734
rect 563822 636498 564004 636734
rect 563404 601054 564004 636498
rect 563404 600818 563586 601054
rect 563822 600818 564004 601054
rect 563404 600734 564004 600818
rect 563404 600498 563586 600734
rect 563822 600498 564004 600734
rect 563404 565054 564004 600498
rect 563404 564818 563586 565054
rect 563822 564818 564004 565054
rect 563404 564734 564004 564818
rect 563404 564498 563586 564734
rect 563822 564498 564004 564734
rect 563404 529054 564004 564498
rect 563404 528818 563586 529054
rect 563822 528818 564004 529054
rect 563404 528734 564004 528818
rect 563404 528498 563586 528734
rect 563822 528498 564004 528734
rect 563404 493054 564004 528498
rect 563404 492818 563586 493054
rect 563822 492818 564004 493054
rect 563404 492734 564004 492818
rect 563404 492498 563586 492734
rect 563822 492498 564004 492734
rect 563404 457054 564004 492498
rect 563404 456818 563586 457054
rect 563822 456818 564004 457054
rect 563404 456734 564004 456818
rect 563404 456498 563586 456734
rect 563822 456498 564004 456734
rect 563404 421054 564004 456498
rect 563404 420818 563586 421054
rect 563822 420818 564004 421054
rect 563404 420734 564004 420818
rect 563404 420498 563586 420734
rect 563822 420498 564004 420734
rect 563404 385054 564004 420498
rect 563404 384818 563586 385054
rect 563822 384818 564004 385054
rect 563404 384734 564004 384818
rect 563404 384498 563586 384734
rect 563822 384498 564004 384734
rect 563404 349054 564004 384498
rect 563404 348818 563586 349054
rect 563822 348818 564004 349054
rect 563404 348734 564004 348818
rect 563404 348498 563586 348734
rect 563822 348498 564004 348734
rect 563404 313054 564004 348498
rect 563404 312818 563586 313054
rect 563822 312818 564004 313054
rect 563404 312734 564004 312818
rect 563404 312498 563586 312734
rect 563822 312498 564004 312734
rect 563404 277054 564004 312498
rect 563404 276818 563586 277054
rect 563822 276818 564004 277054
rect 563404 276734 564004 276818
rect 563404 276498 563586 276734
rect 563822 276498 564004 276734
rect 563404 241054 564004 276498
rect 563404 240818 563586 241054
rect 563822 240818 564004 241054
rect 563404 240734 564004 240818
rect 563404 240498 563586 240734
rect 563822 240498 564004 240734
rect 563404 205054 564004 240498
rect 563404 204818 563586 205054
rect 563822 204818 564004 205054
rect 563404 204734 564004 204818
rect 563404 204498 563586 204734
rect 563822 204498 564004 204734
rect 563404 169054 564004 204498
rect 563404 168818 563586 169054
rect 563822 168818 564004 169054
rect 563404 168734 564004 168818
rect 563404 168498 563586 168734
rect 563822 168498 564004 168734
rect 563404 133054 564004 168498
rect 563404 132818 563586 133054
rect 563822 132818 564004 133054
rect 563404 132734 564004 132818
rect 563404 132498 563586 132734
rect 563822 132498 564004 132734
rect 563404 97054 564004 132498
rect 563404 96818 563586 97054
rect 563822 96818 564004 97054
rect 563404 96734 564004 96818
rect 563404 96498 563586 96734
rect 563822 96498 564004 96734
rect 563404 61054 564004 96498
rect 563404 60818 563586 61054
rect 563822 60818 564004 61054
rect 563404 60734 564004 60818
rect 563404 60498 563586 60734
rect 563822 60498 564004 60734
rect 563404 25054 564004 60498
rect 563404 24818 563586 25054
rect 563822 24818 564004 25054
rect 563404 24734 564004 24818
rect 563404 24498 563586 24734
rect 563822 24498 564004 24734
rect 563404 -3166 564004 24498
rect 563404 -3402 563586 -3166
rect 563822 -3402 564004 -3166
rect 563404 -3486 564004 -3402
rect 563404 -3722 563586 -3486
rect 563822 -3722 564004 -3486
rect 563404 -3744 564004 -3722
rect 567004 676654 567604 708982
rect 567004 676418 567186 676654
rect 567422 676418 567604 676654
rect 567004 676334 567604 676418
rect 567004 676098 567186 676334
rect 567422 676098 567604 676334
rect 567004 640654 567604 676098
rect 567004 640418 567186 640654
rect 567422 640418 567604 640654
rect 567004 640334 567604 640418
rect 567004 640098 567186 640334
rect 567422 640098 567604 640334
rect 567004 604654 567604 640098
rect 567004 604418 567186 604654
rect 567422 604418 567604 604654
rect 567004 604334 567604 604418
rect 567004 604098 567186 604334
rect 567422 604098 567604 604334
rect 567004 568654 567604 604098
rect 567004 568418 567186 568654
rect 567422 568418 567604 568654
rect 567004 568334 567604 568418
rect 567004 568098 567186 568334
rect 567422 568098 567604 568334
rect 567004 532654 567604 568098
rect 567004 532418 567186 532654
rect 567422 532418 567604 532654
rect 567004 532334 567604 532418
rect 567004 532098 567186 532334
rect 567422 532098 567604 532334
rect 567004 496654 567604 532098
rect 567004 496418 567186 496654
rect 567422 496418 567604 496654
rect 567004 496334 567604 496418
rect 567004 496098 567186 496334
rect 567422 496098 567604 496334
rect 567004 460654 567604 496098
rect 567004 460418 567186 460654
rect 567422 460418 567604 460654
rect 567004 460334 567604 460418
rect 567004 460098 567186 460334
rect 567422 460098 567604 460334
rect 567004 424654 567604 460098
rect 567004 424418 567186 424654
rect 567422 424418 567604 424654
rect 567004 424334 567604 424418
rect 567004 424098 567186 424334
rect 567422 424098 567604 424334
rect 567004 388654 567604 424098
rect 567004 388418 567186 388654
rect 567422 388418 567604 388654
rect 567004 388334 567604 388418
rect 567004 388098 567186 388334
rect 567422 388098 567604 388334
rect 567004 352654 567604 388098
rect 567004 352418 567186 352654
rect 567422 352418 567604 352654
rect 567004 352334 567604 352418
rect 567004 352098 567186 352334
rect 567422 352098 567604 352334
rect 567004 316654 567604 352098
rect 567004 316418 567186 316654
rect 567422 316418 567604 316654
rect 567004 316334 567604 316418
rect 567004 316098 567186 316334
rect 567422 316098 567604 316334
rect 567004 280654 567604 316098
rect 567004 280418 567186 280654
rect 567422 280418 567604 280654
rect 567004 280334 567604 280418
rect 567004 280098 567186 280334
rect 567422 280098 567604 280334
rect 567004 244654 567604 280098
rect 567004 244418 567186 244654
rect 567422 244418 567604 244654
rect 567004 244334 567604 244418
rect 567004 244098 567186 244334
rect 567422 244098 567604 244334
rect 567004 208654 567604 244098
rect 567004 208418 567186 208654
rect 567422 208418 567604 208654
rect 567004 208334 567604 208418
rect 567004 208098 567186 208334
rect 567422 208098 567604 208334
rect 567004 172654 567604 208098
rect 567004 172418 567186 172654
rect 567422 172418 567604 172654
rect 567004 172334 567604 172418
rect 567004 172098 567186 172334
rect 567422 172098 567604 172334
rect 567004 136654 567604 172098
rect 567004 136418 567186 136654
rect 567422 136418 567604 136654
rect 567004 136334 567604 136418
rect 567004 136098 567186 136334
rect 567422 136098 567604 136334
rect 567004 100654 567604 136098
rect 567004 100418 567186 100654
rect 567422 100418 567604 100654
rect 567004 100334 567604 100418
rect 567004 100098 567186 100334
rect 567422 100098 567604 100334
rect 567004 64654 567604 100098
rect 567004 64418 567186 64654
rect 567422 64418 567604 64654
rect 567004 64334 567604 64418
rect 567004 64098 567186 64334
rect 567422 64098 567604 64334
rect 567004 28654 567604 64098
rect 567004 28418 567186 28654
rect 567422 28418 567604 28654
rect 567004 28334 567604 28418
rect 567004 28098 567186 28334
rect 567422 28098 567604 28334
rect 567004 -5046 567604 28098
rect 567004 -5282 567186 -5046
rect 567422 -5282 567604 -5046
rect 567004 -5366 567604 -5282
rect 567004 -5602 567186 -5366
rect 567422 -5602 567604 -5366
rect 567004 -5624 567604 -5602
rect 570604 680254 571204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 581404 706718 582004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 581404 706482 581586 706718
rect 581822 706482 582004 706718
rect 581404 706398 582004 706482
rect 581404 706162 581586 706398
rect 581822 706162 582004 706398
rect 570604 680018 570786 680254
rect 571022 680018 571204 680254
rect 570604 679934 571204 680018
rect 570604 679698 570786 679934
rect 571022 679698 571204 679934
rect 570604 644254 571204 679698
rect 570604 644018 570786 644254
rect 571022 644018 571204 644254
rect 570604 643934 571204 644018
rect 570604 643698 570786 643934
rect 571022 643698 571204 643934
rect 570604 608254 571204 643698
rect 570604 608018 570786 608254
rect 571022 608018 571204 608254
rect 570604 607934 571204 608018
rect 570604 607698 570786 607934
rect 571022 607698 571204 607934
rect 570604 572254 571204 607698
rect 570604 572018 570786 572254
rect 571022 572018 571204 572254
rect 570604 571934 571204 572018
rect 570604 571698 570786 571934
rect 571022 571698 571204 571934
rect 570604 536254 571204 571698
rect 570604 536018 570786 536254
rect 571022 536018 571204 536254
rect 570604 535934 571204 536018
rect 570604 535698 570786 535934
rect 571022 535698 571204 535934
rect 570604 500254 571204 535698
rect 570604 500018 570786 500254
rect 571022 500018 571204 500254
rect 570604 499934 571204 500018
rect 570604 499698 570786 499934
rect 571022 499698 571204 499934
rect 570604 464254 571204 499698
rect 570604 464018 570786 464254
rect 571022 464018 571204 464254
rect 570604 463934 571204 464018
rect 570604 463698 570786 463934
rect 571022 463698 571204 463934
rect 570604 428254 571204 463698
rect 570604 428018 570786 428254
rect 571022 428018 571204 428254
rect 570604 427934 571204 428018
rect 570604 427698 570786 427934
rect 571022 427698 571204 427934
rect 570604 392254 571204 427698
rect 570604 392018 570786 392254
rect 571022 392018 571204 392254
rect 570604 391934 571204 392018
rect 570604 391698 570786 391934
rect 571022 391698 571204 391934
rect 570604 356254 571204 391698
rect 570604 356018 570786 356254
rect 571022 356018 571204 356254
rect 570604 355934 571204 356018
rect 570604 355698 570786 355934
rect 571022 355698 571204 355934
rect 570604 320254 571204 355698
rect 570604 320018 570786 320254
rect 571022 320018 571204 320254
rect 570604 319934 571204 320018
rect 570604 319698 570786 319934
rect 571022 319698 571204 319934
rect 570604 284254 571204 319698
rect 570604 284018 570786 284254
rect 571022 284018 571204 284254
rect 570604 283934 571204 284018
rect 570604 283698 570786 283934
rect 571022 283698 571204 283934
rect 570604 248254 571204 283698
rect 570604 248018 570786 248254
rect 571022 248018 571204 248254
rect 570604 247934 571204 248018
rect 570604 247698 570786 247934
rect 571022 247698 571204 247934
rect 570604 212254 571204 247698
rect 570604 212018 570786 212254
rect 571022 212018 571204 212254
rect 570604 211934 571204 212018
rect 570604 211698 570786 211934
rect 571022 211698 571204 211934
rect 570604 176254 571204 211698
rect 570604 176018 570786 176254
rect 571022 176018 571204 176254
rect 570604 175934 571204 176018
rect 570604 175698 570786 175934
rect 571022 175698 571204 175934
rect 570604 140254 571204 175698
rect 570604 140018 570786 140254
rect 571022 140018 571204 140254
rect 570604 139934 571204 140018
rect 570604 139698 570786 139934
rect 571022 139698 571204 139934
rect 570604 104254 571204 139698
rect 570604 104018 570786 104254
rect 571022 104018 571204 104254
rect 570604 103934 571204 104018
rect 570604 103698 570786 103934
rect 571022 103698 571204 103934
rect 570604 68254 571204 103698
rect 570604 68018 570786 68254
rect 571022 68018 571204 68254
rect 570604 67934 571204 68018
rect 570604 67698 570786 67934
rect 571022 67698 571204 67934
rect 570604 32254 571204 67698
rect 570604 32018 570786 32254
rect 571022 32018 571204 32254
rect 570604 31934 571204 32018
rect 570604 31698 570786 31934
rect 571022 31698 571204 31934
rect 552604 -6222 552786 -5986
rect 553022 -6222 553204 -5986
rect 552604 -6306 553204 -6222
rect 552604 -6542 552786 -6306
rect 553022 -6542 553204 -6306
rect 552604 -7504 553204 -6542
rect 570604 -6926 571204 31698
rect 577804 704838 578404 705800
rect 577804 704602 577986 704838
rect 578222 704602 578404 704838
rect 577804 704518 578404 704602
rect 577804 704282 577986 704518
rect 578222 704282 578404 704518
rect 577804 687454 578404 704282
rect 577804 687218 577986 687454
rect 578222 687218 578404 687454
rect 577804 687134 578404 687218
rect 577804 686898 577986 687134
rect 578222 686898 578404 687134
rect 577804 651454 578404 686898
rect 577804 651218 577986 651454
rect 578222 651218 578404 651454
rect 577804 651134 578404 651218
rect 577804 650898 577986 651134
rect 578222 650898 578404 651134
rect 577804 615454 578404 650898
rect 577804 615218 577986 615454
rect 578222 615218 578404 615454
rect 577804 615134 578404 615218
rect 577804 614898 577986 615134
rect 578222 614898 578404 615134
rect 577804 579454 578404 614898
rect 577804 579218 577986 579454
rect 578222 579218 578404 579454
rect 577804 579134 578404 579218
rect 577804 578898 577986 579134
rect 578222 578898 578404 579134
rect 577804 543454 578404 578898
rect 577804 543218 577986 543454
rect 578222 543218 578404 543454
rect 577804 543134 578404 543218
rect 577804 542898 577986 543134
rect 578222 542898 578404 543134
rect 577804 507454 578404 542898
rect 577804 507218 577986 507454
rect 578222 507218 578404 507454
rect 577804 507134 578404 507218
rect 577804 506898 577986 507134
rect 578222 506898 578404 507134
rect 577804 471454 578404 506898
rect 577804 471218 577986 471454
rect 578222 471218 578404 471454
rect 577804 471134 578404 471218
rect 577804 470898 577986 471134
rect 578222 470898 578404 471134
rect 577804 435454 578404 470898
rect 577804 435218 577986 435454
rect 578222 435218 578404 435454
rect 577804 435134 578404 435218
rect 577804 434898 577986 435134
rect 578222 434898 578404 435134
rect 577804 399454 578404 434898
rect 577804 399218 577986 399454
rect 578222 399218 578404 399454
rect 577804 399134 578404 399218
rect 577804 398898 577986 399134
rect 578222 398898 578404 399134
rect 577804 363454 578404 398898
rect 577804 363218 577986 363454
rect 578222 363218 578404 363454
rect 577804 363134 578404 363218
rect 577804 362898 577986 363134
rect 578222 362898 578404 363134
rect 577804 327454 578404 362898
rect 577804 327218 577986 327454
rect 578222 327218 578404 327454
rect 577804 327134 578404 327218
rect 577804 326898 577986 327134
rect 578222 326898 578404 327134
rect 577804 291454 578404 326898
rect 577804 291218 577986 291454
rect 578222 291218 578404 291454
rect 577804 291134 578404 291218
rect 577804 290898 577986 291134
rect 578222 290898 578404 291134
rect 577804 255454 578404 290898
rect 577804 255218 577986 255454
rect 578222 255218 578404 255454
rect 577804 255134 578404 255218
rect 577804 254898 577986 255134
rect 578222 254898 578404 255134
rect 577804 219454 578404 254898
rect 577804 219218 577986 219454
rect 578222 219218 578404 219454
rect 577804 219134 578404 219218
rect 577804 218898 577986 219134
rect 578222 218898 578404 219134
rect 577804 183454 578404 218898
rect 577804 183218 577986 183454
rect 578222 183218 578404 183454
rect 577804 183134 578404 183218
rect 577804 182898 577986 183134
rect 578222 182898 578404 183134
rect 577804 147454 578404 182898
rect 577804 147218 577986 147454
rect 578222 147218 578404 147454
rect 577804 147134 578404 147218
rect 577804 146898 577986 147134
rect 578222 146898 578404 147134
rect 577804 111454 578404 146898
rect 577804 111218 577986 111454
rect 578222 111218 578404 111454
rect 577804 111134 578404 111218
rect 577804 110898 577986 111134
rect 578222 110898 578404 111134
rect 577804 75454 578404 110898
rect 577804 75218 577986 75454
rect 578222 75218 578404 75454
rect 577804 75134 578404 75218
rect 577804 74898 577986 75134
rect 578222 74898 578404 75134
rect 577804 39454 578404 74898
rect 577804 39218 577986 39454
rect 578222 39218 578404 39454
rect 577804 39134 578404 39218
rect 577804 38898 577986 39134
rect 578222 38898 578404 39134
rect 577804 3454 578404 38898
rect 577804 3218 577986 3454
rect 578222 3218 578404 3454
rect 577804 3134 578404 3218
rect 577804 2898 577986 3134
rect 578222 2898 578404 3134
rect 577804 -346 578404 2898
rect 577804 -582 577986 -346
rect 578222 -582 578404 -346
rect 577804 -666 578404 -582
rect 577804 -902 577986 -666
rect 578222 -902 578404 -666
rect 577804 -1864 578404 -902
rect 581404 691054 582004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 581404 690818 581586 691054
rect 581822 690818 582004 691054
rect 581404 690734 582004 690818
rect 581404 690498 581586 690734
rect 581822 690498 582004 690734
rect 581404 655054 582004 690498
rect 581404 654818 581586 655054
rect 581822 654818 582004 655054
rect 581404 654734 582004 654818
rect 581404 654498 581586 654734
rect 581822 654498 582004 654734
rect 581404 619054 582004 654498
rect 581404 618818 581586 619054
rect 581822 618818 582004 619054
rect 581404 618734 582004 618818
rect 581404 618498 581586 618734
rect 581822 618498 582004 618734
rect 581404 583054 582004 618498
rect 581404 582818 581586 583054
rect 581822 582818 582004 583054
rect 581404 582734 582004 582818
rect 581404 582498 581586 582734
rect 581822 582498 582004 582734
rect 581404 547054 582004 582498
rect 581404 546818 581586 547054
rect 581822 546818 582004 547054
rect 581404 546734 582004 546818
rect 581404 546498 581586 546734
rect 581822 546498 582004 546734
rect 581404 511054 582004 546498
rect 581404 510818 581586 511054
rect 581822 510818 582004 511054
rect 581404 510734 582004 510818
rect 581404 510498 581586 510734
rect 581822 510498 582004 510734
rect 581404 475054 582004 510498
rect 581404 474818 581586 475054
rect 581822 474818 582004 475054
rect 581404 474734 582004 474818
rect 581404 474498 581586 474734
rect 581822 474498 582004 474734
rect 581404 439054 582004 474498
rect 581404 438818 581586 439054
rect 581822 438818 582004 439054
rect 581404 438734 582004 438818
rect 581404 438498 581586 438734
rect 581822 438498 582004 438734
rect 581404 403054 582004 438498
rect 581404 402818 581586 403054
rect 581822 402818 582004 403054
rect 581404 402734 582004 402818
rect 581404 402498 581586 402734
rect 581822 402498 582004 402734
rect 581404 367054 582004 402498
rect 581404 366818 581586 367054
rect 581822 366818 582004 367054
rect 581404 366734 582004 366818
rect 581404 366498 581586 366734
rect 581822 366498 582004 366734
rect 581404 331054 582004 366498
rect 581404 330818 581586 331054
rect 581822 330818 582004 331054
rect 581404 330734 582004 330818
rect 581404 330498 581586 330734
rect 581822 330498 582004 330734
rect 581404 295054 582004 330498
rect 581404 294818 581586 295054
rect 581822 294818 582004 295054
rect 581404 294734 582004 294818
rect 581404 294498 581586 294734
rect 581822 294498 582004 294734
rect 581404 259054 582004 294498
rect 581404 258818 581586 259054
rect 581822 258818 582004 259054
rect 581404 258734 582004 258818
rect 581404 258498 581586 258734
rect 581822 258498 582004 258734
rect 581404 223054 582004 258498
rect 581404 222818 581586 223054
rect 581822 222818 582004 223054
rect 581404 222734 582004 222818
rect 581404 222498 581586 222734
rect 581822 222498 582004 222734
rect 581404 187054 582004 222498
rect 581404 186818 581586 187054
rect 581822 186818 582004 187054
rect 581404 186734 582004 186818
rect 581404 186498 581586 186734
rect 581822 186498 582004 186734
rect 581404 151054 582004 186498
rect 581404 150818 581586 151054
rect 581822 150818 582004 151054
rect 581404 150734 582004 150818
rect 581404 150498 581586 150734
rect 581822 150498 582004 150734
rect 581404 115054 582004 150498
rect 581404 114818 581586 115054
rect 581822 114818 582004 115054
rect 581404 114734 582004 114818
rect 581404 114498 581586 114734
rect 581822 114498 582004 114734
rect 581404 79054 582004 114498
rect 581404 78818 581586 79054
rect 581822 78818 582004 79054
rect 581404 78734 582004 78818
rect 581404 78498 581586 78734
rect 581822 78498 582004 78734
rect 581404 43054 582004 78498
rect 581404 42818 581586 43054
rect 581822 42818 582004 43054
rect 581404 42734 582004 42818
rect 581404 42498 581586 42734
rect 581822 42498 582004 42734
rect 581404 7054 582004 42498
rect 581404 6818 581586 7054
rect 581822 6818 582004 7054
rect 581404 6734 582004 6818
rect 581404 6498 581586 6734
rect 581822 6498 582004 6734
rect 581404 -2226 582004 6498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 687454 585920 704282
rect 585320 687218 585502 687454
rect 585738 687218 585920 687454
rect 585320 687134 585920 687218
rect 585320 686898 585502 687134
rect 585738 686898 585920 687134
rect 585320 651454 585920 686898
rect 585320 651218 585502 651454
rect 585738 651218 585920 651454
rect 585320 651134 585920 651218
rect 585320 650898 585502 651134
rect 585738 650898 585920 651134
rect 585320 615454 585920 650898
rect 585320 615218 585502 615454
rect 585738 615218 585920 615454
rect 585320 615134 585920 615218
rect 585320 614898 585502 615134
rect 585738 614898 585920 615134
rect 585320 579454 585920 614898
rect 585320 579218 585502 579454
rect 585738 579218 585920 579454
rect 585320 579134 585920 579218
rect 585320 578898 585502 579134
rect 585738 578898 585920 579134
rect 585320 543454 585920 578898
rect 585320 543218 585502 543454
rect 585738 543218 585920 543454
rect 585320 543134 585920 543218
rect 585320 542898 585502 543134
rect 585738 542898 585920 543134
rect 585320 507454 585920 542898
rect 585320 507218 585502 507454
rect 585738 507218 585920 507454
rect 585320 507134 585920 507218
rect 585320 506898 585502 507134
rect 585738 506898 585920 507134
rect 585320 471454 585920 506898
rect 585320 471218 585502 471454
rect 585738 471218 585920 471454
rect 585320 471134 585920 471218
rect 585320 470898 585502 471134
rect 585738 470898 585920 471134
rect 585320 435454 585920 470898
rect 585320 435218 585502 435454
rect 585738 435218 585920 435454
rect 585320 435134 585920 435218
rect 585320 434898 585502 435134
rect 585738 434898 585920 435134
rect 585320 399454 585920 434898
rect 585320 399218 585502 399454
rect 585738 399218 585920 399454
rect 585320 399134 585920 399218
rect 585320 398898 585502 399134
rect 585738 398898 585920 399134
rect 585320 363454 585920 398898
rect 585320 363218 585502 363454
rect 585738 363218 585920 363454
rect 585320 363134 585920 363218
rect 585320 362898 585502 363134
rect 585738 362898 585920 363134
rect 585320 327454 585920 362898
rect 585320 327218 585502 327454
rect 585738 327218 585920 327454
rect 585320 327134 585920 327218
rect 585320 326898 585502 327134
rect 585738 326898 585920 327134
rect 585320 291454 585920 326898
rect 585320 291218 585502 291454
rect 585738 291218 585920 291454
rect 585320 291134 585920 291218
rect 585320 290898 585502 291134
rect 585738 290898 585920 291134
rect 585320 255454 585920 290898
rect 585320 255218 585502 255454
rect 585738 255218 585920 255454
rect 585320 255134 585920 255218
rect 585320 254898 585502 255134
rect 585738 254898 585920 255134
rect 585320 219454 585920 254898
rect 585320 219218 585502 219454
rect 585738 219218 585920 219454
rect 585320 219134 585920 219218
rect 585320 218898 585502 219134
rect 585738 218898 585920 219134
rect 585320 183454 585920 218898
rect 585320 183218 585502 183454
rect 585738 183218 585920 183454
rect 585320 183134 585920 183218
rect 585320 182898 585502 183134
rect 585738 182898 585920 183134
rect 585320 147454 585920 182898
rect 585320 147218 585502 147454
rect 585738 147218 585920 147454
rect 585320 147134 585920 147218
rect 585320 146898 585502 147134
rect 585738 146898 585920 147134
rect 585320 111454 585920 146898
rect 585320 111218 585502 111454
rect 585738 111218 585920 111454
rect 585320 111134 585920 111218
rect 585320 110898 585502 111134
rect 585738 110898 585920 111134
rect 585320 75454 585920 110898
rect 585320 75218 585502 75454
rect 585738 75218 585920 75454
rect 585320 75134 585920 75218
rect 585320 74898 585502 75134
rect 585738 74898 585920 75134
rect 585320 39454 585920 74898
rect 585320 39218 585502 39454
rect 585738 39218 585920 39454
rect 585320 39134 585920 39218
rect 585320 38898 585502 39134
rect 585738 38898 585920 39134
rect 585320 3454 585920 38898
rect 585320 3218 585502 3454
rect 585738 3218 585920 3454
rect 585320 3134 585920 3218
rect 585320 2898 585502 3134
rect 585738 2898 585920 3134
rect 585320 -346 585920 2898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 669454 586860 705222
rect 586260 669218 586442 669454
rect 586678 669218 586860 669454
rect 586260 669134 586860 669218
rect 586260 668898 586442 669134
rect 586678 668898 586860 669134
rect 586260 633454 586860 668898
rect 586260 633218 586442 633454
rect 586678 633218 586860 633454
rect 586260 633134 586860 633218
rect 586260 632898 586442 633134
rect 586678 632898 586860 633134
rect 586260 597454 586860 632898
rect 586260 597218 586442 597454
rect 586678 597218 586860 597454
rect 586260 597134 586860 597218
rect 586260 596898 586442 597134
rect 586678 596898 586860 597134
rect 586260 561454 586860 596898
rect 586260 561218 586442 561454
rect 586678 561218 586860 561454
rect 586260 561134 586860 561218
rect 586260 560898 586442 561134
rect 586678 560898 586860 561134
rect 586260 525454 586860 560898
rect 586260 525218 586442 525454
rect 586678 525218 586860 525454
rect 586260 525134 586860 525218
rect 586260 524898 586442 525134
rect 586678 524898 586860 525134
rect 586260 489454 586860 524898
rect 586260 489218 586442 489454
rect 586678 489218 586860 489454
rect 586260 489134 586860 489218
rect 586260 488898 586442 489134
rect 586678 488898 586860 489134
rect 586260 453454 586860 488898
rect 586260 453218 586442 453454
rect 586678 453218 586860 453454
rect 586260 453134 586860 453218
rect 586260 452898 586442 453134
rect 586678 452898 586860 453134
rect 586260 417454 586860 452898
rect 586260 417218 586442 417454
rect 586678 417218 586860 417454
rect 586260 417134 586860 417218
rect 586260 416898 586442 417134
rect 586678 416898 586860 417134
rect 586260 381454 586860 416898
rect 586260 381218 586442 381454
rect 586678 381218 586860 381454
rect 586260 381134 586860 381218
rect 586260 380898 586442 381134
rect 586678 380898 586860 381134
rect 586260 345454 586860 380898
rect 586260 345218 586442 345454
rect 586678 345218 586860 345454
rect 586260 345134 586860 345218
rect 586260 344898 586442 345134
rect 586678 344898 586860 345134
rect 586260 309454 586860 344898
rect 586260 309218 586442 309454
rect 586678 309218 586860 309454
rect 586260 309134 586860 309218
rect 586260 308898 586442 309134
rect 586678 308898 586860 309134
rect 586260 273454 586860 308898
rect 586260 273218 586442 273454
rect 586678 273218 586860 273454
rect 586260 273134 586860 273218
rect 586260 272898 586442 273134
rect 586678 272898 586860 273134
rect 586260 237454 586860 272898
rect 586260 237218 586442 237454
rect 586678 237218 586860 237454
rect 586260 237134 586860 237218
rect 586260 236898 586442 237134
rect 586678 236898 586860 237134
rect 586260 201454 586860 236898
rect 586260 201218 586442 201454
rect 586678 201218 586860 201454
rect 586260 201134 586860 201218
rect 586260 200898 586442 201134
rect 586678 200898 586860 201134
rect 586260 165454 586860 200898
rect 586260 165218 586442 165454
rect 586678 165218 586860 165454
rect 586260 165134 586860 165218
rect 586260 164898 586442 165134
rect 586678 164898 586860 165134
rect 586260 129454 586860 164898
rect 586260 129218 586442 129454
rect 586678 129218 586860 129454
rect 586260 129134 586860 129218
rect 586260 128898 586442 129134
rect 586678 128898 586860 129134
rect 586260 93454 586860 128898
rect 586260 93218 586442 93454
rect 586678 93218 586860 93454
rect 586260 93134 586860 93218
rect 586260 92898 586442 93134
rect 586678 92898 586860 93134
rect 586260 57454 586860 92898
rect 586260 57218 586442 57454
rect 586678 57218 586860 57454
rect 586260 57134 586860 57218
rect 586260 56898 586442 57134
rect 586678 56898 586860 57134
rect 586260 21454 586860 56898
rect 586260 21218 586442 21454
rect 586678 21218 586860 21454
rect 586260 21134 586860 21218
rect 586260 20898 586442 21134
rect 586678 20898 586860 21134
rect 586260 -1286 586860 20898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 691054 587800 706162
rect 587200 690818 587382 691054
rect 587618 690818 587800 691054
rect 587200 690734 587800 690818
rect 587200 690498 587382 690734
rect 587618 690498 587800 690734
rect 587200 655054 587800 690498
rect 587200 654818 587382 655054
rect 587618 654818 587800 655054
rect 587200 654734 587800 654818
rect 587200 654498 587382 654734
rect 587618 654498 587800 654734
rect 587200 619054 587800 654498
rect 587200 618818 587382 619054
rect 587618 618818 587800 619054
rect 587200 618734 587800 618818
rect 587200 618498 587382 618734
rect 587618 618498 587800 618734
rect 587200 583054 587800 618498
rect 587200 582818 587382 583054
rect 587618 582818 587800 583054
rect 587200 582734 587800 582818
rect 587200 582498 587382 582734
rect 587618 582498 587800 582734
rect 587200 547054 587800 582498
rect 587200 546818 587382 547054
rect 587618 546818 587800 547054
rect 587200 546734 587800 546818
rect 587200 546498 587382 546734
rect 587618 546498 587800 546734
rect 587200 511054 587800 546498
rect 587200 510818 587382 511054
rect 587618 510818 587800 511054
rect 587200 510734 587800 510818
rect 587200 510498 587382 510734
rect 587618 510498 587800 510734
rect 587200 475054 587800 510498
rect 587200 474818 587382 475054
rect 587618 474818 587800 475054
rect 587200 474734 587800 474818
rect 587200 474498 587382 474734
rect 587618 474498 587800 474734
rect 587200 439054 587800 474498
rect 587200 438818 587382 439054
rect 587618 438818 587800 439054
rect 587200 438734 587800 438818
rect 587200 438498 587382 438734
rect 587618 438498 587800 438734
rect 587200 403054 587800 438498
rect 587200 402818 587382 403054
rect 587618 402818 587800 403054
rect 587200 402734 587800 402818
rect 587200 402498 587382 402734
rect 587618 402498 587800 402734
rect 587200 367054 587800 402498
rect 587200 366818 587382 367054
rect 587618 366818 587800 367054
rect 587200 366734 587800 366818
rect 587200 366498 587382 366734
rect 587618 366498 587800 366734
rect 587200 331054 587800 366498
rect 587200 330818 587382 331054
rect 587618 330818 587800 331054
rect 587200 330734 587800 330818
rect 587200 330498 587382 330734
rect 587618 330498 587800 330734
rect 587200 295054 587800 330498
rect 587200 294818 587382 295054
rect 587618 294818 587800 295054
rect 587200 294734 587800 294818
rect 587200 294498 587382 294734
rect 587618 294498 587800 294734
rect 587200 259054 587800 294498
rect 587200 258818 587382 259054
rect 587618 258818 587800 259054
rect 587200 258734 587800 258818
rect 587200 258498 587382 258734
rect 587618 258498 587800 258734
rect 587200 223054 587800 258498
rect 587200 222818 587382 223054
rect 587618 222818 587800 223054
rect 587200 222734 587800 222818
rect 587200 222498 587382 222734
rect 587618 222498 587800 222734
rect 587200 187054 587800 222498
rect 587200 186818 587382 187054
rect 587618 186818 587800 187054
rect 587200 186734 587800 186818
rect 587200 186498 587382 186734
rect 587618 186498 587800 186734
rect 587200 151054 587800 186498
rect 587200 150818 587382 151054
rect 587618 150818 587800 151054
rect 587200 150734 587800 150818
rect 587200 150498 587382 150734
rect 587618 150498 587800 150734
rect 587200 115054 587800 150498
rect 587200 114818 587382 115054
rect 587618 114818 587800 115054
rect 587200 114734 587800 114818
rect 587200 114498 587382 114734
rect 587618 114498 587800 114734
rect 587200 79054 587800 114498
rect 587200 78818 587382 79054
rect 587618 78818 587800 79054
rect 587200 78734 587800 78818
rect 587200 78498 587382 78734
rect 587618 78498 587800 78734
rect 587200 43054 587800 78498
rect 587200 42818 587382 43054
rect 587618 42818 587800 43054
rect 587200 42734 587800 42818
rect 587200 42498 587382 42734
rect 587618 42498 587800 42734
rect 587200 7054 587800 42498
rect 587200 6818 587382 7054
rect 587618 6818 587800 7054
rect 587200 6734 587800 6818
rect 587200 6498 587382 6734
rect 587618 6498 587800 6734
rect 581404 -2462 581586 -2226
rect 581822 -2462 582004 -2226
rect 581404 -2546 582004 -2462
rect 581404 -2782 581586 -2546
rect 581822 -2782 582004 -2546
rect 581404 -3744 582004 -2782
rect 587200 -2226 587800 6498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 673054 588740 707102
rect 588140 672818 588322 673054
rect 588558 672818 588740 673054
rect 588140 672734 588740 672818
rect 588140 672498 588322 672734
rect 588558 672498 588740 672734
rect 588140 637054 588740 672498
rect 588140 636818 588322 637054
rect 588558 636818 588740 637054
rect 588140 636734 588740 636818
rect 588140 636498 588322 636734
rect 588558 636498 588740 636734
rect 588140 601054 588740 636498
rect 588140 600818 588322 601054
rect 588558 600818 588740 601054
rect 588140 600734 588740 600818
rect 588140 600498 588322 600734
rect 588558 600498 588740 600734
rect 588140 565054 588740 600498
rect 588140 564818 588322 565054
rect 588558 564818 588740 565054
rect 588140 564734 588740 564818
rect 588140 564498 588322 564734
rect 588558 564498 588740 564734
rect 588140 529054 588740 564498
rect 588140 528818 588322 529054
rect 588558 528818 588740 529054
rect 588140 528734 588740 528818
rect 588140 528498 588322 528734
rect 588558 528498 588740 528734
rect 588140 493054 588740 528498
rect 588140 492818 588322 493054
rect 588558 492818 588740 493054
rect 588140 492734 588740 492818
rect 588140 492498 588322 492734
rect 588558 492498 588740 492734
rect 588140 457054 588740 492498
rect 588140 456818 588322 457054
rect 588558 456818 588740 457054
rect 588140 456734 588740 456818
rect 588140 456498 588322 456734
rect 588558 456498 588740 456734
rect 588140 421054 588740 456498
rect 588140 420818 588322 421054
rect 588558 420818 588740 421054
rect 588140 420734 588740 420818
rect 588140 420498 588322 420734
rect 588558 420498 588740 420734
rect 588140 385054 588740 420498
rect 588140 384818 588322 385054
rect 588558 384818 588740 385054
rect 588140 384734 588740 384818
rect 588140 384498 588322 384734
rect 588558 384498 588740 384734
rect 588140 349054 588740 384498
rect 588140 348818 588322 349054
rect 588558 348818 588740 349054
rect 588140 348734 588740 348818
rect 588140 348498 588322 348734
rect 588558 348498 588740 348734
rect 588140 313054 588740 348498
rect 588140 312818 588322 313054
rect 588558 312818 588740 313054
rect 588140 312734 588740 312818
rect 588140 312498 588322 312734
rect 588558 312498 588740 312734
rect 588140 277054 588740 312498
rect 588140 276818 588322 277054
rect 588558 276818 588740 277054
rect 588140 276734 588740 276818
rect 588140 276498 588322 276734
rect 588558 276498 588740 276734
rect 588140 241054 588740 276498
rect 588140 240818 588322 241054
rect 588558 240818 588740 241054
rect 588140 240734 588740 240818
rect 588140 240498 588322 240734
rect 588558 240498 588740 240734
rect 588140 205054 588740 240498
rect 588140 204818 588322 205054
rect 588558 204818 588740 205054
rect 588140 204734 588740 204818
rect 588140 204498 588322 204734
rect 588558 204498 588740 204734
rect 588140 169054 588740 204498
rect 588140 168818 588322 169054
rect 588558 168818 588740 169054
rect 588140 168734 588740 168818
rect 588140 168498 588322 168734
rect 588558 168498 588740 168734
rect 588140 133054 588740 168498
rect 588140 132818 588322 133054
rect 588558 132818 588740 133054
rect 588140 132734 588740 132818
rect 588140 132498 588322 132734
rect 588558 132498 588740 132734
rect 588140 97054 588740 132498
rect 588140 96818 588322 97054
rect 588558 96818 588740 97054
rect 588140 96734 588740 96818
rect 588140 96498 588322 96734
rect 588558 96498 588740 96734
rect 588140 61054 588740 96498
rect 588140 60818 588322 61054
rect 588558 60818 588740 61054
rect 588140 60734 588740 60818
rect 588140 60498 588322 60734
rect 588558 60498 588740 60734
rect 588140 25054 588740 60498
rect 588140 24818 588322 25054
rect 588558 24818 588740 25054
rect 588140 24734 588740 24818
rect 588140 24498 588322 24734
rect 588558 24498 588740 24734
rect 588140 -3166 588740 24498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 694654 589680 708042
rect 589080 694418 589262 694654
rect 589498 694418 589680 694654
rect 589080 694334 589680 694418
rect 589080 694098 589262 694334
rect 589498 694098 589680 694334
rect 589080 658654 589680 694098
rect 589080 658418 589262 658654
rect 589498 658418 589680 658654
rect 589080 658334 589680 658418
rect 589080 658098 589262 658334
rect 589498 658098 589680 658334
rect 589080 622654 589680 658098
rect 589080 622418 589262 622654
rect 589498 622418 589680 622654
rect 589080 622334 589680 622418
rect 589080 622098 589262 622334
rect 589498 622098 589680 622334
rect 589080 586654 589680 622098
rect 589080 586418 589262 586654
rect 589498 586418 589680 586654
rect 589080 586334 589680 586418
rect 589080 586098 589262 586334
rect 589498 586098 589680 586334
rect 589080 550654 589680 586098
rect 589080 550418 589262 550654
rect 589498 550418 589680 550654
rect 589080 550334 589680 550418
rect 589080 550098 589262 550334
rect 589498 550098 589680 550334
rect 589080 514654 589680 550098
rect 589080 514418 589262 514654
rect 589498 514418 589680 514654
rect 589080 514334 589680 514418
rect 589080 514098 589262 514334
rect 589498 514098 589680 514334
rect 589080 478654 589680 514098
rect 589080 478418 589262 478654
rect 589498 478418 589680 478654
rect 589080 478334 589680 478418
rect 589080 478098 589262 478334
rect 589498 478098 589680 478334
rect 589080 442654 589680 478098
rect 589080 442418 589262 442654
rect 589498 442418 589680 442654
rect 589080 442334 589680 442418
rect 589080 442098 589262 442334
rect 589498 442098 589680 442334
rect 589080 406654 589680 442098
rect 589080 406418 589262 406654
rect 589498 406418 589680 406654
rect 589080 406334 589680 406418
rect 589080 406098 589262 406334
rect 589498 406098 589680 406334
rect 589080 370654 589680 406098
rect 589080 370418 589262 370654
rect 589498 370418 589680 370654
rect 589080 370334 589680 370418
rect 589080 370098 589262 370334
rect 589498 370098 589680 370334
rect 589080 334654 589680 370098
rect 589080 334418 589262 334654
rect 589498 334418 589680 334654
rect 589080 334334 589680 334418
rect 589080 334098 589262 334334
rect 589498 334098 589680 334334
rect 589080 298654 589680 334098
rect 589080 298418 589262 298654
rect 589498 298418 589680 298654
rect 589080 298334 589680 298418
rect 589080 298098 589262 298334
rect 589498 298098 589680 298334
rect 589080 262654 589680 298098
rect 589080 262418 589262 262654
rect 589498 262418 589680 262654
rect 589080 262334 589680 262418
rect 589080 262098 589262 262334
rect 589498 262098 589680 262334
rect 589080 226654 589680 262098
rect 589080 226418 589262 226654
rect 589498 226418 589680 226654
rect 589080 226334 589680 226418
rect 589080 226098 589262 226334
rect 589498 226098 589680 226334
rect 589080 190654 589680 226098
rect 589080 190418 589262 190654
rect 589498 190418 589680 190654
rect 589080 190334 589680 190418
rect 589080 190098 589262 190334
rect 589498 190098 589680 190334
rect 589080 154654 589680 190098
rect 589080 154418 589262 154654
rect 589498 154418 589680 154654
rect 589080 154334 589680 154418
rect 589080 154098 589262 154334
rect 589498 154098 589680 154334
rect 589080 118654 589680 154098
rect 589080 118418 589262 118654
rect 589498 118418 589680 118654
rect 589080 118334 589680 118418
rect 589080 118098 589262 118334
rect 589498 118098 589680 118334
rect 589080 82654 589680 118098
rect 589080 82418 589262 82654
rect 589498 82418 589680 82654
rect 589080 82334 589680 82418
rect 589080 82098 589262 82334
rect 589498 82098 589680 82334
rect 589080 46654 589680 82098
rect 589080 46418 589262 46654
rect 589498 46418 589680 46654
rect 589080 46334 589680 46418
rect 589080 46098 589262 46334
rect 589498 46098 589680 46334
rect 589080 10654 589680 46098
rect 589080 10418 589262 10654
rect 589498 10418 589680 10654
rect 589080 10334 589680 10418
rect 589080 10098 589262 10334
rect 589498 10098 589680 10334
rect 589080 -4106 589680 10098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 676654 590620 708982
rect 590020 676418 590202 676654
rect 590438 676418 590620 676654
rect 590020 676334 590620 676418
rect 590020 676098 590202 676334
rect 590438 676098 590620 676334
rect 590020 640654 590620 676098
rect 590020 640418 590202 640654
rect 590438 640418 590620 640654
rect 590020 640334 590620 640418
rect 590020 640098 590202 640334
rect 590438 640098 590620 640334
rect 590020 604654 590620 640098
rect 590020 604418 590202 604654
rect 590438 604418 590620 604654
rect 590020 604334 590620 604418
rect 590020 604098 590202 604334
rect 590438 604098 590620 604334
rect 590020 568654 590620 604098
rect 590020 568418 590202 568654
rect 590438 568418 590620 568654
rect 590020 568334 590620 568418
rect 590020 568098 590202 568334
rect 590438 568098 590620 568334
rect 590020 532654 590620 568098
rect 590020 532418 590202 532654
rect 590438 532418 590620 532654
rect 590020 532334 590620 532418
rect 590020 532098 590202 532334
rect 590438 532098 590620 532334
rect 590020 496654 590620 532098
rect 590020 496418 590202 496654
rect 590438 496418 590620 496654
rect 590020 496334 590620 496418
rect 590020 496098 590202 496334
rect 590438 496098 590620 496334
rect 590020 460654 590620 496098
rect 590020 460418 590202 460654
rect 590438 460418 590620 460654
rect 590020 460334 590620 460418
rect 590020 460098 590202 460334
rect 590438 460098 590620 460334
rect 590020 424654 590620 460098
rect 590020 424418 590202 424654
rect 590438 424418 590620 424654
rect 590020 424334 590620 424418
rect 590020 424098 590202 424334
rect 590438 424098 590620 424334
rect 590020 388654 590620 424098
rect 590020 388418 590202 388654
rect 590438 388418 590620 388654
rect 590020 388334 590620 388418
rect 590020 388098 590202 388334
rect 590438 388098 590620 388334
rect 590020 352654 590620 388098
rect 590020 352418 590202 352654
rect 590438 352418 590620 352654
rect 590020 352334 590620 352418
rect 590020 352098 590202 352334
rect 590438 352098 590620 352334
rect 590020 316654 590620 352098
rect 590020 316418 590202 316654
rect 590438 316418 590620 316654
rect 590020 316334 590620 316418
rect 590020 316098 590202 316334
rect 590438 316098 590620 316334
rect 590020 280654 590620 316098
rect 590020 280418 590202 280654
rect 590438 280418 590620 280654
rect 590020 280334 590620 280418
rect 590020 280098 590202 280334
rect 590438 280098 590620 280334
rect 590020 244654 590620 280098
rect 590020 244418 590202 244654
rect 590438 244418 590620 244654
rect 590020 244334 590620 244418
rect 590020 244098 590202 244334
rect 590438 244098 590620 244334
rect 590020 208654 590620 244098
rect 590020 208418 590202 208654
rect 590438 208418 590620 208654
rect 590020 208334 590620 208418
rect 590020 208098 590202 208334
rect 590438 208098 590620 208334
rect 590020 172654 590620 208098
rect 590020 172418 590202 172654
rect 590438 172418 590620 172654
rect 590020 172334 590620 172418
rect 590020 172098 590202 172334
rect 590438 172098 590620 172334
rect 590020 136654 590620 172098
rect 590020 136418 590202 136654
rect 590438 136418 590620 136654
rect 590020 136334 590620 136418
rect 590020 136098 590202 136334
rect 590438 136098 590620 136334
rect 590020 100654 590620 136098
rect 590020 100418 590202 100654
rect 590438 100418 590620 100654
rect 590020 100334 590620 100418
rect 590020 100098 590202 100334
rect 590438 100098 590620 100334
rect 590020 64654 590620 100098
rect 590020 64418 590202 64654
rect 590438 64418 590620 64654
rect 590020 64334 590620 64418
rect 590020 64098 590202 64334
rect 590438 64098 590620 64334
rect 590020 28654 590620 64098
rect 590020 28418 590202 28654
rect 590438 28418 590620 28654
rect 590020 28334 590620 28418
rect 590020 28098 590202 28334
rect 590438 28098 590620 28334
rect 590020 -5046 590620 28098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 698254 591560 709922
rect 590960 698018 591142 698254
rect 591378 698018 591560 698254
rect 590960 697934 591560 698018
rect 590960 697698 591142 697934
rect 591378 697698 591560 697934
rect 590960 662254 591560 697698
rect 590960 662018 591142 662254
rect 591378 662018 591560 662254
rect 590960 661934 591560 662018
rect 590960 661698 591142 661934
rect 591378 661698 591560 661934
rect 590960 626254 591560 661698
rect 590960 626018 591142 626254
rect 591378 626018 591560 626254
rect 590960 625934 591560 626018
rect 590960 625698 591142 625934
rect 591378 625698 591560 625934
rect 590960 590254 591560 625698
rect 590960 590018 591142 590254
rect 591378 590018 591560 590254
rect 590960 589934 591560 590018
rect 590960 589698 591142 589934
rect 591378 589698 591560 589934
rect 590960 554254 591560 589698
rect 590960 554018 591142 554254
rect 591378 554018 591560 554254
rect 590960 553934 591560 554018
rect 590960 553698 591142 553934
rect 591378 553698 591560 553934
rect 590960 518254 591560 553698
rect 590960 518018 591142 518254
rect 591378 518018 591560 518254
rect 590960 517934 591560 518018
rect 590960 517698 591142 517934
rect 591378 517698 591560 517934
rect 590960 482254 591560 517698
rect 590960 482018 591142 482254
rect 591378 482018 591560 482254
rect 590960 481934 591560 482018
rect 590960 481698 591142 481934
rect 591378 481698 591560 481934
rect 590960 446254 591560 481698
rect 590960 446018 591142 446254
rect 591378 446018 591560 446254
rect 590960 445934 591560 446018
rect 590960 445698 591142 445934
rect 591378 445698 591560 445934
rect 590960 410254 591560 445698
rect 590960 410018 591142 410254
rect 591378 410018 591560 410254
rect 590960 409934 591560 410018
rect 590960 409698 591142 409934
rect 591378 409698 591560 409934
rect 590960 374254 591560 409698
rect 590960 374018 591142 374254
rect 591378 374018 591560 374254
rect 590960 373934 591560 374018
rect 590960 373698 591142 373934
rect 591378 373698 591560 373934
rect 590960 338254 591560 373698
rect 590960 338018 591142 338254
rect 591378 338018 591560 338254
rect 590960 337934 591560 338018
rect 590960 337698 591142 337934
rect 591378 337698 591560 337934
rect 590960 302254 591560 337698
rect 590960 302018 591142 302254
rect 591378 302018 591560 302254
rect 590960 301934 591560 302018
rect 590960 301698 591142 301934
rect 591378 301698 591560 301934
rect 590960 266254 591560 301698
rect 590960 266018 591142 266254
rect 591378 266018 591560 266254
rect 590960 265934 591560 266018
rect 590960 265698 591142 265934
rect 591378 265698 591560 265934
rect 590960 230254 591560 265698
rect 590960 230018 591142 230254
rect 591378 230018 591560 230254
rect 590960 229934 591560 230018
rect 590960 229698 591142 229934
rect 591378 229698 591560 229934
rect 590960 194254 591560 229698
rect 590960 194018 591142 194254
rect 591378 194018 591560 194254
rect 590960 193934 591560 194018
rect 590960 193698 591142 193934
rect 591378 193698 591560 193934
rect 590960 158254 591560 193698
rect 590960 158018 591142 158254
rect 591378 158018 591560 158254
rect 590960 157934 591560 158018
rect 590960 157698 591142 157934
rect 591378 157698 591560 157934
rect 590960 122254 591560 157698
rect 590960 122018 591142 122254
rect 591378 122018 591560 122254
rect 590960 121934 591560 122018
rect 590960 121698 591142 121934
rect 591378 121698 591560 121934
rect 590960 86254 591560 121698
rect 590960 86018 591142 86254
rect 591378 86018 591560 86254
rect 590960 85934 591560 86018
rect 590960 85698 591142 85934
rect 591378 85698 591560 85934
rect 590960 50254 591560 85698
rect 590960 50018 591142 50254
rect 591378 50018 591560 50254
rect 590960 49934 591560 50018
rect 590960 49698 591142 49934
rect 591378 49698 591560 49934
rect 590960 14254 591560 49698
rect 590960 14018 591142 14254
rect 591378 14018 591560 14254
rect 590960 13934 591560 14018
rect 590960 13698 591142 13934
rect 591378 13698 591560 13934
rect 590960 -5986 591560 13698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 680254 592500 710862
rect 591900 680018 592082 680254
rect 592318 680018 592500 680254
rect 591900 679934 592500 680018
rect 591900 679698 592082 679934
rect 592318 679698 592500 679934
rect 591900 644254 592500 679698
rect 591900 644018 592082 644254
rect 592318 644018 592500 644254
rect 591900 643934 592500 644018
rect 591900 643698 592082 643934
rect 592318 643698 592500 643934
rect 591900 608254 592500 643698
rect 591900 608018 592082 608254
rect 592318 608018 592500 608254
rect 591900 607934 592500 608018
rect 591900 607698 592082 607934
rect 592318 607698 592500 607934
rect 591900 572254 592500 607698
rect 591900 572018 592082 572254
rect 592318 572018 592500 572254
rect 591900 571934 592500 572018
rect 591900 571698 592082 571934
rect 592318 571698 592500 571934
rect 591900 536254 592500 571698
rect 591900 536018 592082 536254
rect 592318 536018 592500 536254
rect 591900 535934 592500 536018
rect 591900 535698 592082 535934
rect 592318 535698 592500 535934
rect 591900 500254 592500 535698
rect 591900 500018 592082 500254
rect 592318 500018 592500 500254
rect 591900 499934 592500 500018
rect 591900 499698 592082 499934
rect 592318 499698 592500 499934
rect 591900 464254 592500 499698
rect 591900 464018 592082 464254
rect 592318 464018 592500 464254
rect 591900 463934 592500 464018
rect 591900 463698 592082 463934
rect 592318 463698 592500 463934
rect 591900 428254 592500 463698
rect 591900 428018 592082 428254
rect 592318 428018 592500 428254
rect 591900 427934 592500 428018
rect 591900 427698 592082 427934
rect 592318 427698 592500 427934
rect 591900 392254 592500 427698
rect 591900 392018 592082 392254
rect 592318 392018 592500 392254
rect 591900 391934 592500 392018
rect 591900 391698 592082 391934
rect 592318 391698 592500 391934
rect 591900 356254 592500 391698
rect 591900 356018 592082 356254
rect 592318 356018 592500 356254
rect 591900 355934 592500 356018
rect 591900 355698 592082 355934
rect 592318 355698 592500 355934
rect 591900 320254 592500 355698
rect 591900 320018 592082 320254
rect 592318 320018 592500 320254
rect 591900 319934 592500 320018
rect 591900 319698 592082 319934
rect 592318 319698 592500 319934
rect 591900 284254 592500 319698
rect 591900 284018 592082 284254
rect 592318 284018 592500 284254
rect 591900 283934 592500 284018
rect 591900 283698 592082 283934
rect 592318 283698 592500 283934
rect 591900 248254 592500 283698
rect 591900 248018 592082 248254
rect 592318 248018 592500 248254
rect 591900 247934 592500 248018
rect 591900 247698 592082 247934
rect 592318 247698 592500 247934
rect 591900 212254 592500 247698
rect 591900 212018 592082 212254
rect 592318 212018 592500 212254
rect 591900 211934 592500 212018
rect 591900 211698 592082 211934
rect 592318 211698 592500 211934
rect 591900 176254 592500 211698
rect 591900 176018 592082 176254
rect 592318 176018 592500 176254
rect 591900 175934 592500 176018
rect 591900 175698 592082 175934
rect 592318 175698 592500 175934
rect 591900 140254 592500 175698
rect 591900 140018 592082 140254
rect 592318 140018 592500 140254
rect 591900 139934 592500 140018
rect 591900 139698 592082 139934
rect 592318 139698 592500 139934
rect 591900 104254 592500 139698
rect 591900 104018 592082 104254
rect 592318 104018 592500 104254
rect 591900 103934 592500 104018
rect 591900 103698 592082 103934
rect 592318 103698 592500 103934
rect 591900 68254 592500 103698
rect 591900 68018 592082 68254
rect 592318 68018 592500 68254
rect 591900 67934 592500 68018
rect 591900 67698 592082 67934
rect 592318 67698 592500 67934
rect 591900 32254 592500 67698
rect 591900 32018 592082 32254
rect 592318 32018 592500 32254
rect 591900 31934 592500 32018
rect 591900 31698 592082 31934
rect 592318 31698 592500 31934
rect 570604 -7162 570786 -6926
rect 571022 -7162 571204 -6926
rect 570604 -7246 571204 -7162
rect 570604 -7482 570786 -7246
rect 571022 -7482 571204 -7246
rect 570604 -7504 571204 -7482
rect 591900 -6926 592500 31698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 680018 -8158 680254
rect -8394 679698 -8158 679934
rect -8394 644018 -8158 644254
rect -8394 643698 -8158 643934
rect -8394 608018 -8158 608254
rect -8394 607698 -8158 607934
rect -8394 572018 -8158 572254
rect -8394 571698 -8158 571934
rect -8394 536018 -8158 536254
rect -8394 535698 -8158 535934
rect -8394 500018 -8158 500254
rect -8394 499698 -8158 499934
rect -8394 464018 -8158 464254
rect -8394 463698 -8158 463934
rect -8394 428018 -8158 428254
rect -8394 427698 -8158 427934
rect -8394 392018 -8158 392254
rect -8394 391698 -8158 391934
rect -8394 356018 -8158 356254
rect -8394 355698 -8158 355934
rect -8394 320018 -8158 320254
rect -8394 319698 -8158 319934
rect -8394 284018 -8158 284254
rect -8394 283698 -8158 283934
rect -8394 248018 -8158 248254
rect -8394 247698 -8158 247934
rect -8394 212018 -8158 212254
rect -8394 211698 -8158 211934
rect -8394 176018 -8158 176254
rect -8394 175698 -8158 175934
rect -8394 140018 -8158 140254
rect -8394 139698 -8158 139934
rect -8394 104018 -8158 104254
rect -8394 103698 -8158 103934
rect -8394 68018 -8158 68254
rect -8394 67698 -8158 67934
rect -8394 32018 -8158 32254
rect -8394 31698 -8158 31934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 12786 710242 13022 710478
rect 12786 709922 13022 710158
rect -7454 698018 -7218 698254
rect -7454 697698 -7218 697934
rect -7454 662018 -7218 662254
rect -7454 661698 -7218 661934
rect -7454 626018 -7218 626254
rect -7454 625698 -7218 625934
rect -7454 590018 -7218 590254
rect -7454 589698 -7218 589934
rect -7454 554018 -7218 554254
rect -7454 553698 -7218 553934
rect -7454 518018 -7218 518254
rect -7454 517698 -7218 517934
rect -7454 482018 -7218 482254
rect -7454 481698 -7218 481934
rect -7454 446018 -7218 446254
rect -7454 445698 -7218 445934
rect -7454 410018 -7218 410254
rect -7454 409698 -7218 409934
rect -7454 374018 -7218 374254
rect -7454 373698 -7218 373934
rect -7454 338018 -7218 338254
rect -7454 337698 -7218 337934
rect -7454 302018 -7218 302254
rect -7454 301698 -7218 301934
rect -7454 266018 -7218 266254
rect -7454 265698 -7218 265934
rect -7454 230018 -7218 230254
rect -7454 229698 -7218 229934
rect -7454 194018 -7218 194254
rect -7454 193698 -7218 193934
rect -7454 158018 -7218 158254
rect -7454 157698 -7218 157934
rect -7454 122018 -7218 122254
rect -7454 121698 -7218 121934
rect -7454 86018 -7218 86254
rect -7454 85698 -7218 85934
rect -7454 50018 -7218 50254
rect -7454 49698 -7218 49934
rect -7454 14018 -7218 14254
rect -7454 13698 -7218 13934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 676418 -6278 676654
rect -6514 676098 -6278 676334
rect -6514 640418 -6278 640654
rect -6514 640098 -6278 640334
rect -6514 604418 -6278 604654
rect -6514 604098 -6278 604334
rect -6514 568418 -6278 568654
rect -6514 568098 -6278 568334
rect -6514 532418 -6278 532654
rect -6514 532098 -6278 532334
rect -6514 496418 -6278 496654
rect -6514 496098 -6278 496334
rect -6514 460418 -6278 460654
rect -6514 460098 -6278 460334
rect -6514 424418 -6278 424654
rect -6514 424098 -6278 424334
rect -6514 388418 -6278 388654
rect -6514 388098 -6278 388334
rect -6514 352418 -6278 352654
rect -6514 352098 -6278 352334
rect -6514 316418 -6278 316654
rect -6514 316098 -6278 316334
rect -6514 280418 -6278 280654
rect -6514 280098 -6278 280334
rect -6514 244418 -6278 244654
rect -6514 244098 -6278 244334
rect -6514 208418 -6278 208654
rect -6514 208098 -6278 208334
rect -6514 172418 -6278 172654
rect -6514 172098 -6278 172334
rect -6514 136418 -6278 136654
rect -6514 136098 -6278 136334
rect -6514 100418 -6278 100654
rect -6514 100098 -6278 100334
rect -6514 64418 -6278 64654
rect -6514 64098 -6278 64334
rect -6514 28418 -6278 28654
rect -6514 28098 -6278 28334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 9186 708362 9422 708598
rect 9186 708042 9422 708278
rect -5574 694418 -5338 694654
rect -5574 694098 -5338 694334
rect -5574 658418 -5338 658654
rect -5574 658098 -5338 658334
rect -5574 622418 -5338 622654
rect -5574 622098 -5338 622334
rect -5574 586418 -5338 586654
rect -5574 586098 -5338 586334
rect -5574 550418 -5338 550654
rect -5574 550098 -5338 550334
rect -5574 514418 -5338 514654
rect -5574 514098 -5338 514334
rect -5574 478418 -5338 478654
rect -5574 478098 -5338 478334
rect -5574 442418 -5338 442654
rect -5574 442098 -5338 442334
rect -5574 406418 -5338 406654
rect -5574 406098 -5338 406334
rect -5574 370418 -5338 370654
rect -5574 370098 -5338 370334
rect -5574 334418 -5338 334654
rect -5574 334098 -5338 334334
rect -5574 298418 -5338 298654
rect -5574 298098 -5338 298334
rect -5574 262418 -5338 262654
rect -5574 262098 -5338 262334
rect -5574 226418 -5338 226654
rect -5574 226098 -5338 226334
rect -5574 190418 -5338 190654
rect -5574 190098 -5338 190334
rect -5574 154418 -5338 154654
rect -5574 154098 -5338 154334
rect -5574 118418 -5338 118654
rect -5574 118098 -5338 118334
rect -5574 82418 -5338 82654
rect -5574 82098 -5338 82334
rect -5574 46418 -5338 46654
rect -5574 46098 -5338 46334
rect -5574 10418 -5338 10654
rect -5574 10098 -5338 10334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 672818 -4398 673054
rect -4634 672498 -4398 672734
rect -4634 636818 -4398 637054
rect -4634 636498 -4398 636734
rect -4634 600818 -4398 601054
rect -4634 600498 -4398 600734
rect -4634 564818 -4398 565054
rect -4634 564498 -4398 564734
rect -4634 528818 -4398 529054
rect -4634 528498 -4398 528734
rect -4634 492818 -4398 493054
rect -4634 492498 -4398 492734
rect -4634 456818 -4398 457054
rect -4634 456498 -4398 456734
rect -4634 420818 -4398 421054
rect -4634 420498 -4398 420734
rect -4634 384818 -4398 385054
rect -4634 384498 -4398 384734
rect -4634 348818 -4398 349054
rect -4634 348498 -4398 348734
rect -4634 312818 -4398 313054
rect -4634 312498 -4398 312734
rect -4634 276818 -4398 277054
rect -4634 276498 -4398 276734
rect -4634 240818 -4398 241054
rect -4634 240498 -4398 240734
rect -4634 204818 -4398 205054
rect -4634 204498 -4398 204734
rect -4634 168818 -4398 169054
rect -4634 168498 -4398 168734
rect -4634 132818 -4398 133054
rect -4634 132498 -4398 132734
rect -4634 96818 -4398 97054
rect -4634 96498 -4398 96734
rect -4634 60818 -4398 61054
rect -4634 60498 -4398 60734
rect -4634 24818 -4398 25054
rect -4634 24498 -4398 24734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 5586 706482 5822 706718
rect 5586 706162 5822 706398
rect -3694 690818 -3458 691054
rect -3694 690498 -3458 690734
rect -3694 654818 -3458 655054
rect -3694 654498 -3458 654734
rect -3694 618818 -3458 619054
rect -3694 618498 -3458 618734
rect -3694 582818 -3458 583054
rect -3694 582498 -3458 582734
rect -3694 546818 -3458 547054
rect -3694 546498 -3458 546734
rect -3694 510818 -3458 511054
rect -3694 510498 -3458 510734
rect -3694 474818 -3458 475054
rect -3694 474498 -3458 474734
rect -3694 438818 -3458 439054
rect -3694 438498 -3458 438734
rect -3694 402818 -3458 403054
rect -3694 402498 -3458 402734
rect -3694 366818 -3458 367054
rect -3694 366498 -3458 366734
rect -3694 330818 -3458 331054
rect -3694 330498 -3458 330734
rect -3694 294818 -3458 295054
rect -3694 294498 -3458 294734
rect -3694 258818 -3458 259054
rect -3694 258498 -3458 258734
rect -3694 222818 -3458 223054
rect -3694 222498 -3458 222734
rect -3694 186818 -3458 187054
rect -3694 186498 -3458 186734
rect -3694 150818 -3458 151054
rect -3694 150498 -3458 150734
rect -3694 114818 -3458 115054
rect -3694 114498 -3458 114734
rect -3694 78818 -3458 79054
rect -3694 78498 -3458 78734
rect -3694 42818 -3458 43054
rect -3694 42498 -3458 42734
rect -3694 6818 -3458 7054
rect -3694 6498 -3458 6734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 669218 -2518 669454
rect -2754 668898 -2518 669134
rect -2754 633218 -2518 633454
rect -2754 632898 -2518 633134
rect -2754 597218 -2518 597454
rect -2754 596898 -2518 597134
rect -2754 561218 -2518 561454
rect -2754 560898 -2518 561134
rect -2754 525218 -2518 525454
rect -2754 524898 -2518 525134
rect -2754 489218 -2518 489454
rect -2754 488898 -2518 489134
rect -2754 453218 -2518 453454
rect -2754 452898 -2518 453134
rect -2754 417218 -2518 417454
rect -2754 416898 -2518 417134
rect -2754 381218 -2518 381454
rect -2754 380898 -2518 381134
rect -2754 345218 -2518 345454
rect -2754 344898 -2518 345134
rect -2754 309218 -2518 309454
rect -2754 308898 -2518 309134
rect -2754 273218 -2518 273454
rect -2754 272898 -2518 273134
rect -2754 237218 -2518 237454
rect -2754 236898 -2518 237134
rect -2754 201218 -2518 201454
rect -2754 200898 -2518 201134
rect -2754 165218 -2518 165454
rect -2754 164898 -2518 165134
rect -2754 129218 -2518 129454
rect -2754 128898 -2518 129134
rect -2754 93218 -2518 93454
rect -2754 92898 -2518 93134
rect -2754 57218 -2518 57454
rect -2754 56898 -2518 57134
rect -2754 21218 -2518 21454
rect -2754 20898 -2518 21134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 687218 -1578 687454
rect -1814 686898 -1578 687134
rect -1814 651218 -1578 651454
rect -1814 650898 -1578 651134
rect -1814 615218 -1578 615454
rect -1814 614898 -1578 615134
rect -1814 579218 -1578 579454
rect -1814 578898 -1578 579134
rect -1814 543218 -1578 543454
rect -1814 542898 -1578 543134
rect -1814 507218 -1578 507454
rect -1814 506898 -1578 507134
rect -1814 471218 -1578 471454
rect -1814 470898 -1578 471134
rect -1814 435218 -1578 435454
rect -1814 434898 -1578 435134
rect -1814 399218 -1578 399454
rect -1814 398898 -1578 399134
rect -1814 363218 -1578 363454
rect -1814 362898 -1578 363134
rect -1814 327218 -1578 327454
rect -1814 326898 -1578 327134
rect -1814 291218 -1578 291454
rect -1814 290898 -1578 291134
rect -1814 255218 -1578 255454
rect -1814 254898 -1578 255134
rect -1814 219218 -1578 219454
rect -1814 218898 -1578 219134
rect -1814 183218 -1578 183454
rect -1814 182898 -1578 183134
rect -1814 147218 -1578 147454
rect -1814 146898 -1578 147134
rect -1814 111218 -1578 111454
rect -1814 110898 -1578 111134
rect -1814 75218 -1578 75454
rect -1814 74898 -1578 75134
rect -1814 39218 -1578 39454
rect -1814 38898 -1578 39134
rect -1814 3218 -1578 3454
rect -1814 2898 -1578 3134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 1986 704602 2222 704838
rect 1986 704282 2222 704518
rect 1986 687218 2222 687454
rect 1986 686898 2222 687134
rect 5586 690818 5822 691054
rect 5586 690498 5822 690734
rect 1986 651218 2222 651454
rect 1986 650898 2222 651134
rect 1986 615218 2222 615454
rect 1986 614898 2222 615134
rect 1986 579218 2222 579454
rect 1986 578898 2222 579134
rect 1986 543218 2222 543454
rect 1986 542898 2222 543134
rect 1986 507218 2222 507454
rect 1986 506898 2222 507134
rect 1986 471218 2222 471454
rect 1986 470898 2222 471134
rect 1986 435218 2222 435454
rect 1986 434898 2222 435134
rect 5586 654818 5822 655054
rect 5586 654498 5822 654734
rect 5586 618818 5822 619054
rect 5586 618498 5822 618734
rect 5586 582818 5822 583054
rect 5586 582498 5822 582734
rect 5586 546818 5822 547054
rect 5586 546498 5822 546734
rect 5586 510818 5822 511054
rect 5586 510498 5822 510734
rect 5586 474818 5822 475054
rect 5586 474498 5822 474734
rect 5586 438818 5822 439054
rect 5586 438498 5822 438734
rect 1986 399218 2222 399454
rect 1986 398898 2222 399134
rect 1986 363218 2222 363454
rect 1986 362898 2222 363134
rect 1986 327218 2222 327454
rect 1986 326898 2222 327134
rect 1986 291218 2222 291454
rect 1986 290898 2222 291134
rect 1986 255218 2222 255454
rect 1986 254898 2222 255134
rect 1986 219218 2222 219454
rect 1986 218898 2222 219134
rect 1986 183218 2222 183454
rect 1986 182898 2222 183134
rect 1986 147218 2222 147454
rect 1986 146898 2222 147134
rect 1986 111218 2222 111454
rect 1986 110898 2222 111134
rect 1986 75218 2222 75454
rect 1986 74898 2222 75134
rect 1986 39218 2222 39454
rect 1986 38898 2222 39134
rect 1986 3218 2222 3454
rect 1986 2898 2222 3134
rect 1986 -582 2222 -346
rect 1986 -902 2222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 5586 402818 5822 403054
rect 5586 402498 5822 402734
rect 5586 366818 5822 367054
rect 5586 366498 5822 366734
rect 5586 330818 5822 331054
rect 5586 330498 5822 330734
rect 5586 294818 5822 295054
rect 5586 294498 5822 294734
rect 5586 258818 5822 259054
rect 5586 258498 5822 258734
rect 5586 222818 5822 223054
rect 5586 222498 5822 222734
rect 5586 186818 5822 187054
rect 5586 186498 5822 186734
rect 5586 150818 5822 151054
rect 5586 150498 5822 150734
rect 5586 114818 5822 115054
rect 5586 114498 5822 114734
rect 5586 78818 5822 79054
rect 5586 78498 5822 78734
rect 5586 42818 5822 43054
rect 5586 42498 5822 42734
rect 5586 6818 5822 7054
rect 5586 6498 5822 6734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 5586 -2462 5822 -2226
rect 5586 -2782 5822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 9186 694418 9422 694654
rect 9186 694098 9422 694334
rect 9186 658418 9422 658654
rect 9186 658098 9422 658334
rect 9186 622418 9422 622654
rect 9186 622098 9422 622334
rect 9186 586418 9422 586654
rect 9186 586098 9422 586334
rect 9186 550418 9422 550654
rect 9186 550098 9422 550334
rect 9186 514418 9422 514654
rect 9186 514098 9422 514334
rect 9186 478418 9422 478654
rect 9186 478098 9422 478334
rect 9186 442418 9422 442654
rect 9186 442098 9422 442334
rect 9186 406418 9422 406654
rect 9186 406098 9422 406334
rect 9186 370418 9422 370654
rect 9186 370098 9422 370334
rect 9186 334418 9422 334654
rect 9186 334098 9422 334334
rect 9186 298418 9422 298654
rect 9186 298098 9422 298334
rect 9186 262418 9422 262654
rect 9186 262098 9422 262334
rect 9186 226418 9422 226654
rect 9186 226098 9422 226334
rect 9186 190418 9422 190654
rect 9186 190098 9422 190334
rect 9186 154418 9422 154654
rect 9186 154098 9422 154334
rect 9186 118418 9422 118654
rect 9186 118098 9422 118334
rect 9186 82418 9422 82654
rect 9186 82098 9422 82334
rect 9186 46418 9422 46654
rect 9186 46098 9422 46334
rect 9186 10418 9422 10654
rect 9186 10098 9422 10334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 9186 -4342 9422 -4106
rect 9186 -4662 9422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 30786 711182 31022 711418
rect 30786 710862 31022 711098
rect 27186 709302 27422 709538
rect 27186 708982 27422 709218
rect 23586 707422 23822 707658
rect 23586 707102 23822 707338
rect 12786 698018 13022 698254
rect 12786 697698 13022 697934
rect 12786 662018 13022 662254
rect 12786 661698 13022 661934
rect 12786 626018 13022 626254
rect 12786 625698 13022 625934
rect 12786 590018 13022 590254
rect 12786 589698 13022 589934
rect 12786 554018 13022 554254
rect 12786 553698 13022 553934
rect 12786 518018 13022 518254
rect 12786 517698 13022 517934
rect 12786 482018 13022 482254
rect 12786 481698 13022 481934
rect 12786 446018 13022 446254
rect 12786 445698 13022 445934
rect 12786 410018 13022 410254
rect 12786 409698 13022 409934
rect 12786 374018 13022 374254
rect 12786 373698 13022 373934
rect 12786 338018 13022 338254
rect 12786 337698 13022 337934
rect 12786 302018 13022 302254
rect 12786 301698 13022 301934
rect 12786 266018 13022 266254
rect 12786 265698 13022 265934
rect 12786 230018 13022 230254
rect 12786 229698 13022 229934
rect 12786 194018 13022 194254
rect 12786 193698 13022 193934
rect 12786 158018 13022 158254
rect 12786 157698 13022 157934
rect 12786 122018 13022 122254
rect 12786 121698 13022 121934
rect 12786 86018 13022 86254
rect 12786 85698 13022 85934
rect 12786 50018 13022 50254
rect 12786 49698 13022 49934
rect 12786 14018 13022 14254
rect 12786 13698 13022 13934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 19986 705542 20222 705778
rect 19986 705222 20222 705458
rect 19986 669218 20222 669454
rect 19986 668898 20222 669134
rect 19986 633218 20222 633454
rect 19986 632898 20222 633134
rect 19986 597218 20222 597454
rect 19986 596898 20222 597134
rect 19986 561218 20222 561454
rect 19986 560898 20222 561134
rect 19986 525218 20222 525454
rect 19986 524898 20222 525134
rect 19986 489218 20222 489454
rect 19986 488898 20222 489134
rect 19986 453218 20222 453454
rect 19986 452898 20222 453134
rect 19986 417218 20222 417454
rect 19986 416898 20222 417134
rect 19986 381218 20222 381454
rect 19986 380898 20222 381134
rect 19986 345218 20222 345454
rect 19986 344898 20222 345134
rect 19986 309218 20222 309454
rect 19986 308898 20222 309134
rect 19986 273218 20222 273454
rect 19986 272898 20222 273134
rect 19986 237218 20222 237454
rect 19986 236898 20222 237134
rect 19986 201218 20222 201454
rect 19986 200898 20222 201134
rect 19986 165218 20222 165454
rect 19986 164898 20222 165134
rect 19986 129218 20222 129454
rect 19986 128898 20222 129134
rect 19986 93218 20222 93454
rect 19986 92898 20222 93134
rect 19986 57218 20222 57454
rect 19986 56898 20222 57134
rect 19986 21218 20222 21454
rect 19986 20898 20222 21134
rect 19986 -1522 20222 -1286
rect 19986 -1842 20222 -1606
rect 23586 672818 23822 673054
rect 23586 672498 23822 672734
rect 23586 636818 23822 637054
rect 23586 636498 23822 636734
rect 23586 600818 23822 601054
rect 23586 600498 23822 600734
rect 23586 564818 23822 565054
rect 23586 564498 23822 564734
rect 23586 528818 23822 529054
rect 23586 528498 23822 528734
rect 23586 492818 23822 493054
rect 23586 492498 23822 492734
rect 23586 456818 23822 457054
rect 23586 456498 23822 456734
rect 23586 420818 23822 421054
rect 23586 420498 23822 420734
rect 23586 384818 23822 385054
rect 23586 384498 23822 384734
rect 23586 348818 23822 349054
rect 23586 348498 23822 348734
rect 23586 312818 23822 313054
rect 23586 312498 23822 312734
rect 23586 276818 23822 277054
rect 23586 276498 23822 276734
rect 23586 240818 23822 241054
rect 23586 240498 23822 240734
rect 23586 204818 23822 205054
rect 23586 204498 23822 204734
rect 23586 168818 23822 169054
rect 23586 168498 23822 168734
rect 23586 132818 23822 133054
rect 23586 132498 23822 132734
rect 23586 96818 23822 97054
rect 23586 96498 23822 96734
rect 23586 60818 23822 61054
rect 23586 60498 23822 60734
rect 23586 24818 23822 25054
rect 23586 24498 23822 24734
rect 23586 -3402 23822 -3166
rect 23586 -3722 23822 -3486
rect 27186 676418 27422 676654
rect 27186 676098 27422 676334
rect 27186 640418 27422 640654
rect 27186 640098 27422 640334
rect 27186 604418 27422 604654
rect 27186 604098 27422 604334
rect 27186 568418 27422 568654
rect 27186 568098 27422 568334
rect 27186 532418 27422 532654
rect 27186 532098 27422 532334
rect 27186 496418 27422 496654
rect 27186 496098 27422 496334
rect 27186 460418 27422 460654
rect 27186 460098 27422 460334
rect 27186 424418 27422 424654
rect 27186 424098 27422 424334
rect 27186 388418 27422 388654
rect 27186 388098 27422 388334
rect 27186 352418 27422 352654
rect 27186 352098 27422 352334
rect 27186 316418 27422 316654
rect 27186 316098 27422 316334
rect 27186 280418 27422 280654
rect 27186 280098 27422 280334
rect 27186 244418 27422 244654
rect 27186 244098 27422 244334
rect 27186 208418 27422 208654
rect 27186 208098 27422 208334
rect 27186 172418 27422 172654
rect 27186 172098 27422 172334
rect 27186 136418 27422 136654
rect 27186 136098 27422 136334
rect 27186 100418 27422 100654
rect 27186 100098 27422 100334
rect 27186 64418 27422 64654
rect 27186 64098 27422 64334
rect 27186 28418 27422 28654
rect 27186 28098 27422 28334
rect 27186 -5282 27422 -5046
rect 27186 -5602 27422 -5366
rect 48786 710242 49022 710478
rect 48786 709922 49022 710158
rect 45186 708362 45422 708598
rect 45186 708042 45422 708278
rect 41586 706482 41822 706718
rect 41586 706162 41822 706398
rect 30786 680018 31022 680254
rect 30786 679698 31022 679934
rect 30786 644018 31022 644254
rect 30786 643698 31022 643934
rect 30786 608018 31022 608254
rect 30786 607698 31022 607934
rect 30786 572018 31022 572254
rect 30786 571698 31022 571934
rect 30786 536018 31022 536254
rect 30786 535698 31022 535934
rect 30786 500018 31022 500254
rect 30786 499698 31022 499934
rect 30786 464018 31022 464254
rect 30786 463698 31022 463934
rect 30786 428018 31022 428254
rect 30786 427698 31022 427934
rect 30786 392018 31022 392254
rect 30786 391698 31022 391934
rect 30786 356018 31022 356254
rect 30786 355698 31022 355934
rect 30786 320018 31022 320254
rect 30786 319698 31022 319934
rect 30786 284018 31022 284254
rect 30786 283698 31022 283934
rect 30786 248018 31022 248254
rect 30786 247698 31022 247934
rect 30786 212018 31022 212254
rect 30786 211698 31022 211934
rect 30786 176018 31022 176254
rect 30786 175698 31022 175934
rect 30786 140018 31022 140254
rect 30786 139698 31022 139934
rect 30786 104018 31022 104254
rect 30786 103698 31022 103934
rect 30786 68018 31022 68254
rect 30786 67698 31022 67934
rect 30786 32018 31022 32254
rect 30786 31698 31022 31934
rect 12786 -6222 13022 -5986
rect 12786 -6542 13022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 37986 704602 38222 704838
rect 37986 704282 38222 704518
rect 37986 687218 38222 687454
rect 37986 686898 38222 687134
rect 37986 651218 38222 651454
rect 37986 650898 38222 651134
rect 37986 615218 38222 615454
rect 37986 614898 38222 615134
rect 37986 579218 38222 579454
rect 37986 578898 38222 579134
rect 37986 543218 38222 543454
rect 37986 542898 38222 543134
rect 37986 507218 38222 507454
rect 37986 506898 38222 507134
rect 37986 471218 38222 471454
rect 37986 470898 38222 471134
rect 37986 435218 38222 435454
rect 37986 434898 38222 435134
rect 37986 399218 38222 399454
rect 37986 398898 38222 399134
rect 37986 363218 38222 363454
rect 37986 362898 38222 363134
rect 37986 327218 38222 327454
rect 37986 326898 38222 327134
rect 37986 291218 38222 291454
rect 37986 290898 38222 291134
rect 37986 255218 38222 255454
rect 37986 254898 38222 255134
rect 37986 219218 38222 219454
rect 37986 218898 38222 219134
rect 37986 183218 38222 183454
rect 37986 182898 38222 183134
rect 37986 147218 38222 147454
rect 37986 146898 38222 147134
rect 37986 111218 38222 111454
rect 37986 110898 38222 111134
rect 37986 75218 38222 75454
rect 37986 74898 38222 75134
rect 37986 39218 38222 39454
rect 37986 38898 38222 39134
rect 37986 3218 38222 3454
rect 37986 2898 38222 3134
rect 37986 -582 38222 -346
rect 37986 -902 38222 -666
rect 41586 690818 41822 691054
rect 41586 690498 41822 690734
rect 41586 654818 41822 655054
rect 41586 654498 41822 654734
rect 41586 618818 41822 619054
rect 41586 618498 41822 618734
rect 41586 582818 41822 583054
rect 41586 582498 41822 582734
rect 41586 546818 41822 547054
rect 41586 546498 41822 546734
rect 41586 510818 41822 511054
rect 41586 510498 41822 510734
rect 41586 474818 41822 475054
rect 41586 474498 41822 474734
rect 41586 438818 41822 439054
rect 41586 438498 41822 438734
rect 41586 402818 41822 403054
rect 41586 402498 41822 402734
rect 41586 366818 41822 367054
rect 41586 366498 41822 366734
rect 41586 330818 41822 331054
rect 41586 330498 41822 330734
rect 41586 294818 41822 295054
rect 41586 294498 41822 294734
rect 41586 258818 41822 259054
rect 41586 258498 41822 258734
rect 41586 222818 41822 223054
rect 41586 222498 41822 222734
rect 41586 186818 41822 187054
rect 41586 186498 41822 186734
rect 41586 150818 41822 151054
rect 41586 150498 41822 150734
rect 41586 114818 41822 115054
rect 41586 114498 41822 114734
rect 41586 78818 41822 79054
rect 41586 78498 41822 78734
rect 41586 42818 41822 43054
rect 41586 42498 41822 42734
rect 41586 6818 41822 7054
rect 41586 6498 41822 6734
rect 41586 -2462 41822 -2226
rect 41586 -2782 41822 -2546
rect 45186 694418 45422 694654
rect 45186 694098 45422 694334
rect 45186 658418 45422 658654
rect 45186 658098 45422 658334
rect 45186 622418 45422 622654
rect 45186 622098 45422 622334
rect 45186 586418 45422 586654
rect 45186 586098 45422 586334
rect 45186 550418 45422 550654
rect 45186 550098 45422 550334
rect 45186 514418 45422 514654
rect 45186 514098 45422 514334
rect 45186 478418 45422 478654
rect 45186 478098 45422 478334
rect 45186 442418 45422 442654
rect 45186 442098 45422 442334
rect 45186 406418 45422 406654
rect 45186 406098 45422 406334
rect 45186 370418 45422 370654
rect 45186 370098 45422 370334
rect 45186 334418 45422 334654
rect 45186 334098 45422 334334
rect 45186 298418 45422 298654
rect 45186 298098 45422 298334
rect 45186 262418 45422 262654
rect 45186 262098 45422 262334
rect 45186 226418 45422 226654
rect 45186 226098 45422 226334
rect 45186 190418 45422 190654
rect 45186 190098 45422 190334
rect 45186 154418 45422 154654
rect 45186 154098 45422 154334
rect 45186 118418 45422 118654
rect 45186 118098 45422 118334
rect 45186 82418 45422 82654
rect 45186 82098 45422 82334
rect 45186 46418 45422 46654
rect 45186 46098 45422 46334
rect 45186 10418 45422 10654
rect 45186 10098 45422 10334
rect 45186 -4342 45422 -4106
rect 45186 -4662 45422 -4426
rect 66786 711182 67022 711418
rect 66786 710862 67022 711098
rect 63186 709302 63422 709538
rect 63186 708982 63422 709218
rect 59586 707422 59822 707658
rect 59586 707102 59822 707338
rect 48786 698018 49022 698254
rect 48786 697698 49022 697934
rect 48786 662018 49022 662254
rect 48786 661698 49022 661934
rect 48786 626018 49022 626254
rect 48786 625698 49022 625934
rect 48786 590018 49022 590254
rect 48786 589698 49022 589934
rect 48786 554018 49022 554254
rect 48786 553698 49022 553934
rect 48786 518018 49022 518254
rect 48786 517698 49022 517934
rect 48786 482018 49022 482254
rect 48786 481698 49022 481934
rect 48786 446018 49022 446254
rect 48786 445698 49022 445934
rect 48786 410018 49022 410254
rect 48786 409698 49022 409934
rect 48786 374018 49022 374254
rect 48786 373698 49022 373934
rect 48786 338018 49022 338254
rect 48786 337698 49022 337934
rect 48786 302018 49022 302254
rect 48786 301698 49022 301934
rect 48786 266018 49022 266254
rect 48786 265698 49022 265934
rect 48786 230018 49022 230254
rect 48786 229698 49022 229934
rect 48786 194018 49022 194254
rect 48786 193698 49022 193934
rect 48786 158018 49022 158254
rect 48786 157698 49022 157934
rect 48786 122018 49022 122254
rect 48786 121698 49022 121934
rect 48786 86018 49022 86254
rect 48786 85698 49022 85934
rect 48786 50018 49022 50254
rect 48786 49698 49022 49934
rect 48786 14018 49022 14254
rect 48786 13698 49022 13934
rect 30786 -7162 31022 -6926
rect 30786 -7482 31022 -7246
rect 55986 705542 56222 705778
rect 55986 705222 56222 705458
rect 55986 669218 56222 669454
rect 55986 668898 56222 669134
rect 55986 633218 56222 633454
rect 55986 632898 56222 633134
rect 55986 597218 56222 597454
rect 55986 596898 56222 597134
rect 55986 561218 56222 561454
rect 55986 560898 56222 561134
rect 55986 525218 56222 525454
rect 55986 524898 56222 525134
rect 55986 489218 56222 489454
rect 55986 488898 56222 489134
rect 55986 453218 56222 453454
rect 55986 452898 56222 453134
rect 55986 417218 56222 417454
rect 55986 416898 56222 417134
rect 55986 381218 56222 381454
rect 55986 380898 56222 381134
rect 55986 345218 56222 345454
rect 55986 344898 56222 345134
rect 55986 309218 56222 309454
rect 55986 308898 56222 309134
rect 55986 273218 56222 273454
rect 55986 272898 56222 273134
rect 55986 237218 56222 237454
rect 55986 236898 56222 237134
rect 55986 201218 56222 201454
rect 55986 200898 56222 201134
rect 55986 165218 56222 165454
rect 55986 164898 56222 165134
rect 55986 129218 56222 129454
rect 55986 128898 56222 129134
rect 55986 93218 56222 93454
rect 55986 92898 56222 93134
rect 55986 57218 56222 57454
rect 55986 56898 56222 57134
rect 55986 21218 56222 21454
rect 55986 20898 56222 21134
rect 55986 -1522 56222 -1286
rect 55986 -1842 56222 -1606
rect 59586 672818 59822 673054
rect 59586 672498 59822 672734
rect 59586 636818 59822 637054
rect 59586 636498 59822 636734
rect 59586 600818 59822 601054
rect 59586 600498 59822 600734
rect 59586 564818 59822 565054
rect 59586 564498 59822 564734
rect 59586 528818 59822 529054
rect 59586 528498 59822 528734
rect 59586 492818 59822 493054
rect 59586 492498 59822 492734
rect 59586 456818 59822 457054
rect 59586 456498 59822 456734
rect 59586 420818 59822 421054
rect 59586 420498 59822 420734
rect 59586 384818 59822 385054
rect 59586 384498 59822 384734
rect 59586 348818 59822 349054
rect 59586 348498 59822 348734
rect 59586 312818 59822 313054
rect 59586 312498 59822 312734
rect 59586 276818 59822 277054
rect 59586 276498 59822 276734
rect 59586 240818 59822 241054
rect 59586 240498 59822 240734
rect 59586 204818 59822 205054
rect 59586 204498 59822 204734
rect 59586 168818 59822 169054
rect 59586 168498 59822 168734
rect 59586 132818 59822 133054
rect 59586 132498 59822 132734
rect 59586 96818 59822 97054
rect 59586 96498 59822 96734
rect 59586 60818 59822 61054
rect 59586 60498 59822 60734
rect 59586 24818 59822 25054
rect 59586 24498 59822 24734
rect 59586 -3402 59822 -3166
rect 59586 -3722 59822 -3486
rect 63186 676418 63422 676654
rect 63186 676098 63422 676334
rect 63186 640418 63422 640654
rect 63186 640098 63422 640334
rect 63186 604418 63422 604654
rect 63186 604098 63422 604334
rect 63186 568418 63422 568654
rect 63186 568098 63422 568334
rect 63186 532418 63422 532654
rect 63186 532098 63422 532334
rect 63186 496418 63422 496654
rect 63186 496098 63422 496334
rect 63186 460418 63422 460654
rect 63186 460098 63422 460334
rect 63186 424418 63422 424654
rect 63186 424098 63422 424334
rect 63186 388418 63422 388654
rect 63186 388098 63422 388334
rect 63186 352418 63422 352654
rect 63186 352098 63422 352334
rect 63186 316418 63422 316654
rect 63186 316098 63422 316334
rect 63186 280418 63422 280654
rect 63186 280098 63422 280334
rect 63186 244418 63422 244654
rect 63186 244098 63422 244334
rect 63186 208418 63422 208654
rect 63186 208098 63422 208334
rect 63186 172418 63422 172654
rect 63186 172098 63422 172334
rect 63186 136418 63422 136654
rect 63186 136098 63422 136334
rect 63186 100418 63422 100654
rect 63186 100098 63422 100334
rect 63186 64418 63422 64654
rect 63186 64098 63422 64334
rect 63186 28418 63422 28654
rect 63186 28098 63422 28334
rect 63186 -5282 63422 -5046
rect 63186 -5602 63422 -5366
rect 84786 710242 85022 710478
rect 84786 709922 85022 710158
rect 81186 708362 81422 708598
rect 81186 708042 81422 708278
rect 77586 706482 77822 706718
rect 77586 706162 77822 706398
rect 66786 680018 67022 680254
rect 66786 679698 67022 679934
rect 66786 644018 67022 644254
rect 66786 643698 67022 643934
rect 66786 608018 67022 608254
rect 66786 607698 67022 607934
rect 66786 572018 67022 572254
rect 66786 571698 67022 571934
rect 66786 536018 67022 536254
rect 66786 535698 67022 535934
rect 66786 500018 67022 500254
rect 66786 499698 67022 499934
rect 66786 464018 67022 464254
rect 66786 463698 67022 463934
rect 66786 428018 67022 428254
rect 66786 427698 67022 427934
rect 66786 392018 67022 392254
rect 66786 391698 67022 391934
rect 66786 356018 67022 356254
rect 66786 355698 67022 355934
rect 66786 320018 67022 320254
rect 66786 319698 67022 319934
rect 66786 284018 67022 284254
rect 66786 283698 67022 283934
rect 66786 248018 67022 248254
rect 66786 247698 67022 247934
rect 66786 212018 67022 212254
rect 66786 211698 67022 211934
rect 66786 176018 67022 176254
rect 66786 175698 67022 175934
rect 66786 140018 67022 140254
rect 66786 139698 67022 139934
rect 66786 104018 67022 104254
rect 66786 103698 67022 103934
rect 66786 68018 67022 68254
rect 66786 67698 67022 67934
rect 66786 32018 67022 32254
rect 66786 31698 67022 31934
rect 48786 -6222 49022 -5986
rect 48786 -6542 49022 -6306
rect 73986 704602 74222 704838
rect 73986 704282 74222 704518
rect 73986 687218 74222 687454
rect 73986 686898 74222 687134
rect 73986 651218 74222 651454
rect 73986 650898 74222 651134
rect 73986 615218 74222 615454
rect 73986 614898 74222 615134
rect 73986 579218 74222 579454
rect 73986 578898 74222 579134
rect 73986 543218 74222 543454
rect 73986 542898 74222 543134
rect 73986 507218 74222 507454
rect 73986 506898 74222 507134
rect 73986 471218 74222 471454
rect 73986 470898 74222 471134
rect 73986 435218 74222 435454
rect 73986 434898 74222 435134
rect 73986 399218 74222 399454
rect 73986 398898 74222 399134
rect 73986 363218 74222 363454
rect 73986 362898 74222 363134
rect 73986 327218 74222 327454
rect 73986 326898 74222 327134
rect 73986 291218 74222 291454
rect 73986 290898 74222 291134
rect 73986 255218 74222 255454
rect 73986 254898 74222 255134
rect 73986 219218 74222 219454
rect 73986 218898 74222 219134
rect 73986 183218 74222 183454
rect 73986 182898 74222 183134
rect 73986 147218 74222 147454
rect 73986 146898 74222 147134
rect 73986 111218 74222 111454
rect 73986 110898 74222 111134
rect 73986 75218 74222 75454
rect 73986 74898 74222 75134
rect 73986 39218 74222 39454
rect 73986 38898 74222 39134
rect 73986 3218 74222 3454
rect 73986 2898 74222 3134
rect 73986 -582 74222 -346
rect 73986 -902 74222 -666
rect 77586 690818 77822 691054
rect 77586 690498 77822 690734
rect 77586 654818 77822 655054
rect 77586 654498 77822 654734
rect 77586 618818 77822 619054
rect 77586 618498 77822 618734
rect 77586 582818 77822 583054
rect 77586 582498 77822 582734
rect 77586 546818 77822 547054
rect 77586 546498 77822 546734
rect 77586 510818 77822 511054
rect 77586 510498 77822 510734
rect 77586 474818 77822 475054
rect 77586 474498 77822 474734
rect 77586 438818 77822 439054
rect 77586 438498 77822 438734
rect 77586 402818 77822 403054
rect 77586 402498 77822 402734
rect 77586 366818 77822 367054
rect 77586 366498 77822 366734
rect 77586 330818 77822 331054
rect 77586 330498 77822 330734
rect 77586 294818 77822 295054
rect 77586 294498 77822 294734
rect 77586 258818 77822 259054
rect 77586 258498 77822 258734
rect 77586 222818 77822 223054
rect 77586 222498 77822 222734
rect 77586 186818 77822 187054
rect 77586 186498 77822 186734
rect 77586 150818 77822 151054
rect 77586 150498 77822 150734
rect 77586 114818 77822 115054
rect 77586 114498 77822 114734
rect 77586 78818 77822 79054
rect 77586 78498 77822 78734
rect 77586 42818 77822 43054
rect 77586 42498 77822 42734
rect 77586 6818 77822 7054
rect 77586 6498 77822 6734
rect 77586 -2462 77822 -2226
rect 77586 -2782 77822 -2546
rect 81186 694418 81422 694654
rect 81186 694098 81422 694334
rect 81186 658418 81422 658654
rect 81186 658098 81422 658334
rect 81186 622418 81422 622654
rect 81186 622098 81422 622334
rect 81186 586418 81422 586654
rect 81186 586098 81422 586334
rect 81186 550418 81422 550654
rect 81186 550098 81422 550334
rect 81186 514418 81422 514654
rect 81186 514098 81422 514334
rect 81186 478418 81422 478654
rect 81186 478098 81422 478334
rect 81186 442418 81422 442654
rect 81186 442098 81422 442334
rect 81186 406418 81422 406654
rect 81186 406098 81422 406334
rect 81186 370418 81422 370654
rect 81186 370098 81422 370334
rect 81186 334418 81422 334654
rect 81186 334098 81422 334334
rect 81186 298418 81422 298654
rect 81186 298098 81422 298334
rect 81186 262418 81422 262654
rect 81186 262098 81422 262334
rect 81186 226418 81422 226654
rect 81186 226098 81422 226334
rect 81186 190418 81422 190654
rect 81186 190098 81422 190334
rect 81186 154418 81422 154654
rect 81186 154098 81422 154334
rect 81186 118418 81422 118654
rect 81186 118098 81422 118334
rect 81186 82418 81422 82654
rect 81186 82098 81422 82334
rect 81186 46418 81422 46654
rect 81186 46098 81422 46334
rect 81186 10418 81422 10654
rect 81186 10098 81422 10334
rect 81186 -4342 81422 -4106
rect 81186 -4662 81422 -4426
rect 102786 711182 103022 711418
rect 102786 710862 103022 711098
rect 99186 709302 99422 709538
rect 99186 708982 99422 709218
rect 95586 707422 95822 707658
rect 95586 707102 95822 707338
rect 84786 698018 85022 698254
rect 84786 697698 85022 697934
rect 84786 662018 85022 662254
rect 84786 661698 85022 661934
rect 84786 626018 85022 626254
rect 84786 625698 85022 625934
rect 84786 590018 85022 590254
rect 84786 589698 85022 589934
rect 84786 554018 85022 554254
rect 84786 553698 85022 553934
rect 84786 518018 85022 518254
rect 84786 517698 85022 517934
rect 84786 482018 85022 482254
rect 84786 481698 85022 481934
rect 84786 446018 85022 446254
rect 84786 445698 85022 445934
rect 84786 410018 85022 410254
rect 84786 409698 85022 409934
rect 84786 374018 85022 374254
rect 84786 373698 85022 373934
rect 84786 338018 85022 338254
rect 84786 337698 85022 337934
rect 84786 302018 85022 302254
rect 84786 301698 85022 301934
rect 84786 266018 85022 266254
rect 84786 265698 85022 265934
rect 84786 230018 85022 230254
rect 84786 229698 85022 229934
rect 84786 194018 85022 194254
rect 84786 193698 85022 193934
rect 84786 158018 85022 158254
rect 84786 157698 85022 157934
rect 84786 122018 85022 122254
rect 84786 121698 85022 121934
rect 84786 86018 85022 86254
rect 84786 85698 85022 85934
rect 84786 50018 85022 50254
rect 84786 49698 85022 49934
rect 84786 14018 85022 14254
rect 84786 13698 85022 13934
rect 66786 -7162 67022 -6926
rect 66786 -7482 67022 -7246
rect 91986 705542 92222 705778
rect 91986 705222 92222 705458
rect 91986 669218 92222 669454
rect 91986 668898 92222 669134
rect 91986 633218 92222 633454
rect 91986 632898 92222 633134
rect 91986 597218 92222 597454
rect 91986 596898 92222 597134
rect 91986 561218 92222 561454
rect 91986 560898 92222 561134
rect 91986 525218 92222 525454
rect 91986 524898 92222 525134
rect 91986 489218 92222 489454
rect 91986 488898 92222 489134
rect 91986 453218 92222 453454
rect 91986 452898 92222 453134
rect 91986 417218 92222 417454
rect 91986 416898 92222 417134
rect 91986 381218 92222 381454
rect 91986 380898 92222 381134
rect 91986 345218 92222 345454
rect 91986 344898 92222 345134
rect 91986 309218 92222 309454
rect 91986 308898 92222 309134
rect 91986 273218 92222 273454
rect 91986 272898 92222 273134
rect 91986 237218 92222 237454
rect 91986 236898 92222 237134
rect 91986 201218 92222 201454
rect 91986 200898 92222 201134
rect 91986 165218 92222 165454
rect 91986 164898 92222 165134
rect 91986 129218 92222 129454
rect 91986 128898 92222 129134
rect 91986 93218 92222 93454
rect 91986 92898 92222 93134
rect 91986 57218 92222 57454
rect 91986 56898 92222 57134
rect 91986 21218 92222 21454
rect 91986 20898 92222 21134
rect 91986 -1522 92222 -1286
rect 91986 -1842 92222 -1606
rect 95586 672818 95822 673054
rect 95586 672498 95822 672734
rect 95586 636818 95822 637054
rect 95586 636498 95822 636734
rect 95586 600818 95822 601054
rect 95586 600498 95822 600734
rect 95586 564818 95822 565054
rect 95586 564498 95822 564734
rect 95586 528818 95822 529054
rect 95586 528498 95822 528734
rect 95586 492818 95822 493054
rect 95586 492498 95822 492734
rect 95586 456818 95822 457054
rect 95586 456498 95822 456734
rect 95586 420818 95822 421054
rect 95586 420498 95822 420734
rect 95586 384818 95822 385054
rect 95586 384498 95822 384734
rect 95586 348818 95822 349054
rect 95586 348498 95822 348734
rect 95586 312818 95822 313054
rect 95586 312498 95822 312734
rect 95586 276818 95822 277054
rect 95586 276498 95822 276734
rect 95586 240818 95822 241054
rect 95586 240498 95822 240734
rect 95586 204818 95822 205054
rect 95586 204498 95822 204734
rect 95586 168818 95822 169054
rect 95586 168498 95822 168734
rect 95586 132818 95822 133054
rect 95586 132498 95822 132734
rect 95586 96818 95822 97054
rect 95586 96498 95822 96734
rect 95586 60818 95822 61054
rect 95586 60498 95822 60734
rect 95586 24818 95822 25054
rect 95586 24498 95822 24734
rect 95586 -3402 95822 -3166
rect 95586 -3722 95822 -3486
rect 99186 676418 99422 676654
rect 99186 676098 99422 676334
rect 99186 640418 99422 640654
rect 99186 640098 99422 640334
rect 99186 604418 99422 604654
rect 99186 604098 99422 604334
rect 99186 568418 99422 568654
rect 99186 568098 99422 568334
rect 99186 532418 99422 532654
rect 99186 532098 99422 532334
rect 99186 496418 99422 496654
rect 99186 496098 99422 496334
rect 99186 460418 99422 460654
rect 99186 460098 99422 460334
rect 99186 424418 99422 424654
rect 99186 424098 99422 424334
rect 99186 388418 99422 388654
rect 99186 388098 99422 388334
rect 99186 352418 99422 352654
rect 99186 352098 99422 352334
rect 99186 316418 99422 316654
rect 99186 316098 99422 316334
rect 99186 280418 99422 280654
rect 99186 280098 99422 280334
rect 99186 244418 99422 244654
rect 99186 244098 99422 244334
rect 99186 208418 99422 208654
rect 99186 208098 99422 208334
rect 99186 172418 99422 172654
rect 99186 172098 99422 172334
rect 99186 136418 99422 136654
rect 99186 136098 99422 136334
rect 99186 100418 99422 100654
rect 99186 100098 99422 100334
rect 99186 64418 99422 64654
rect 99186 64098 99422 64334
rect 99186 28418 99422 28654
rect 99186 28098 99422 28334
rect 99186 -5282 99422 -5046
rect 99186 -5602 99422 -5366
rect 120786 710242 121022 710478
rect 120786 709922 121022 710158
rect 117186 708362 117422 708598
rect 117186 708042 117422 708278
rect 113586 706482 113822 706718
rect 113586 706162 113822 706398
rect 102786 680018 103022 680254
rect 102786 679698 103022 679934
rect 102786 644018 103022 644254
rect 102786 643698 103022 643934
rect 102786 608018 103022 608254
rect 102786 607698 103022 607934
rect 102786 572018 103022 572254
rect 102786 571698 103022 571934
rect 102786 536018 103022 536254
rect 102786 535698 103022 535934
rect 102786 500018 103022 500254
rect 102786 499698 103022 499934
rect 102786 464018 103022 464254
rect 102786 463698 103022 463934
rect 102786 428018 103022 428254
rect 102786 427698 103022 427934
rect 102786 392018 103022 392254
rect 102786 391698 103022 391934
rect 102786 356018 103022 356254
rect 102786 355698 103022 355934
rect 102786 320018 103022 320254
rect 102786 319698 103022 319934
rect 102786 284018 103022 284254
rect 102786 283698 103022 283934
rect 102786 248018 103022 248254
rect 102786 247698 103022 247934
rect 102786 212018 103022 212254
rect 102786 211698 103022 211934
rect 102786 176018 103022 176254
rect 102786 175698 103022 175934
rect 102786 140018 103022 140254
rect 102786 139698 103022 139934
rect 102786 104018 103022 104254
rect 102786 103698 103022 103934
rect 102786 68018 103022 68254
rect 102786 67698 103022 67934
rect 102786 32018 103022 32254
rect 102786 31698 103022 31934
rect 84786 -6222 85022 -5986
rect 84786 -6542 85022 -6306
rect 109986 704602 110222 704838
rect 109986 704282 110222 704518
rect 109986 687218 110222 687454
rect 109986 686898 110222 687134
rect 109986 651218 110222 651454
rect 109986 650898 110222 651134
rect 109986 615218 110222 615454
rect 109986 614898 110222 615134
rect 109986 579218 110222 579454
rect 109986 578898 110222 579134
rect 109986 543218 110222 543454
rect 109986 542898 110222 543134
rect 109986 507218 110222 507454
rect 109986 506898 110222 507134
rect 109986 471218 110222 471454
rect 109986 470898 110222 471134
rect 109986 435218 110222 435454
rect 109986 434898 110222 435134
rect 109986 399218 110222 399454
rect 109986 398898 110222 399134
rect 109986 363218 110222 363454
rect 109986 362898 110222 363134
rect 109986 327218 110222 327454
rect 109986 326898 110222 327134
rect 109986 291218 110222 291454
rect 109986 290898 110222 291134
rect 109986 255218 110222 255454
rect 109986 254898 110222 255134
rect 109986 219218 110222 219454
rect 109986 218898 110222 219134
rect 109986 183218 110222 183454
rect 109986 182898 110222 183134
rect 109986 147218 110222 147454
rect 109986 146898 110222 147134
rect 109986 111218 110222 111454
rect 109986 110898 110222 111134
rect 109986 75218 110222 75454
rect 109986 74898 110222 75134
rect 109986 39218 110222 39454
rect 109986 38898 110222 39134
rect 109986 3218 110222 3454
rect 109986 2898 110222 3134
rect 109986 -582 110222 -346
rect 109986 -902 110222 -666
rect 113586 690818 113822 691054
rect 113586 690498 113822 690734
rect 113586 654818 113822 655054
rect 113586 654498 113822 654734
rect 113586 618818 113822 619054
rect 113586 618498 113822 618734
rect 113586 582818 113822 583054
rect 113586 582498 113822 582734
rect 113586 546818 113822 547054
rect 113586 546498 113822 546734
rect 113586 510818 113822 511054
rect 113586 510498 113822 510734
rect 113586 474818 113822 475054
rect 113586 474498 113822 474734
rect 113586 438818 113822 439054
rect 113586 438498 113822 438734
rect 113586 402818 113822 403054
rect 113586 402498 113822 402734
rect 113586 366818 113822 367054
rect 113586 366498 113822 366734
rect 113586 330818 113822 331054
rect 113586 330498 113822 330734
rect 113586 294818 113822 295054
rect 113586 294498 113822 294734
rect 113586 258818 113822 259054
rect 113586 258498 113822 258734
rect 113586 222818 113822 223054
rect 113586 222498 113822 222734
rect 113586 186818 113822 187054
rect 113586 186498 113822 186734
rect 113586 150818 113822 151054
rect 113586 150498 113822 150734
rect 113586 114818 113822 115054
rect 113586 114498 113822 114734
rect 113586 78818 113822 79054
rect 113586 78498 113822 78734
rect 113586 42818 113822 43054
rect 113586 42498 113822 42734
rect 113586 6818 113822 7054
rect 113586 6498 113822 6734
rect 113586 -2462 113822 -2226
rect 113586 -2782 113822 -2546
rect 117186 694418 117422 694654
rect 117186 694098 117422 694334
rect 117186 658418 117422 658654
rect 117186 658098 117422 658334
rect 117186 622418 117422 622654
rect 117186 622098 117422 622334
rect 117186 586418 117422 586654
rect 117186 586098 117422 586334
rect 117186 550418 117422 550654
rect 117186 550098 117422 550334
rect 117186 514418 117422 514654
rect 117186 514098 117422 514334
rect 117186 478418 117422 478654
rect 117186 478098 117422 478334
rect 117186 442418 117422 442654
rect 117186 442098 117422 442334
rect 117186 406418 117422 406654
rect 117186 406098 117422 406334
rect 117186 370418 117422 370654
rect 117186 370098 117422 370334
rect 117186 334418 117422 334654
rect 117186 334098 117422 334334
rect 117186 298418 117422 298654
rect 117186 298098 117422 298334
rect 117186 262418 117422 262654
rect 117186 262098 117422 262334
rect 117186 226418 117422 226654
rect 117186 226098 117422 226334
rect 117186 190418 117422 190654
rect 117186 190098 117422 190334
rect 117186 154418 117422 154654
rect 117186 154098 117422 154334
rect 117186 118418 117422 118654
rect 117186 118098 117422 118334
rect 117186 82418 117422 82654
rect 117186 82098 117422 82334
rect 117186 46418 117422 46654
rect 117186 46098 117422 46334
rect 117186 10418 117422 10654
rect 117186 10098 117422 10334
rect 117186 -4342 117422 -4106
rect 117186 -4662 117422 -4426
rect 138786 711182 139022 711418
rect 138786 710862 139022 711098
rect 135186 709302 135422 709538
rect 135186 708982 135422 709218
rect 131586 707422 131822 707658
rect 131586 707102 131822 707338
rect 120786 698018 121022 698254
rect 120786 697698 121022 697934
rect 120786 662018 121022 662254
rect 120786 661698 121022 661934
rect 120786 626018 121022 626254
rect 120786 625698 121022 625934
rect 120786 590018 121022 590254
rect 120786 589698 121022 589934
rect 120786 554018 121022 554254
rect 120786 553698 121022 553934
rect 120786 518018 121022 518254
rect 120786 517698 121022 517934
rect 120786 482018 121022 482254
rect 120786 481698 121022 481934
rect 120786 446018 121022 446254
rect 120786 445698 121022 445934
rect 120786 410018 121022 410254
rect 120786 409698 121022 409934
rect 120786 374018 121022 374254
rect 120786 373698 121022 373934
rect 120786 338018 121022 338254
rect 120786 337698 121022 337934
rect 120786 302018 121022 302254
rect 120786 301698 121022 301934
rect 120786 266018 121022 266254
rect 120786 265698 121022 265934
rect 120786 230018 121022 230254
rect 120786 229698 121022 229934
rect 120786 194018 121022 194254
rect 120786 193698 121022 193934
rect 120786 158018 121022 158254
rect 120786 157698 121022 157934
rect 120786 122018 121022 122254
rect 120786 121698 121022 121934
rect 120786 86018 121022 86254
rect 120786 85698 121022 85934
rect 120786 50018 121022 50254
rect 120786 49698 121022 49934
rect 120786 14018 121022 14254
rect 120786 13698 121022 13934
rect 102786 -7162 103022 -6926
rect 102786 -7482 103022 -7246
rect 127986 705542 128222 705778
rect 127986 705222 128222 705458
rect 127986 669218 128222 669454
rect 127986 668898 128222 669134
rect 127986 633218 128222 633454
rect 127986 632898 128222 633134
rect 127986 597218 128222 597454
rect 127986 596898 128222 597134
rect 127986 561218 128222 561454
rect 127986 560898 128222 561134
rect 127986 525218 128222 525454
rect 127986 524898 128222 525134
rect 127986 489218 128222 489454
rect 127986 488898 128222 489134
rect 127986 453218 128222 453454
rect 127986 452898 128222 453134
rect 127986 417218 128222 417454
rect 127986 416898 128222 417134
rect 127986 381218 128222 381454
rect 127986 380898 128222 381134
rect 127986 345218 128222 345454
rect 127986 344898 128222 345134
rect 127986 309218 128222 309454
rect 127986 308898 128222 309134
rect 127986 273218 128222 273454
rect 127986 272898 128222 273134
rect 127986 237218 128222 237454
rect 127986 236898 128222 237134
rect 127986 201218 128222 201454
rect 127986 200898 128222 201134
rect 127986 165218 128222 165454
rect 127986 164898 128222 165134
rect 127986 129218 128222 129454
rect 127986 128898 128222 129134
rect 127986 93218 128222 93454
rect 127986 92898 128222 93134
rect 127986 57218 128222 57454
rect 127986 56898 128222 57134
rect 127986 21218 128222 21454
rect 127986 20898 128222 21134
rect 127986 -1522 128222 -1286
rect 127986 -1842 128222 -1606
rect 131586 672818 131822 673054
rect 131586 672498 131822 672734
rect 131586 636818 131822 637054
rect 131586 636498 131822 636734
rect 131586 600818 131822 601054
rect 131586 600498 131822 600734
rect 131586 564818 131822 565054
rect 131586 564498 131822 564734
rect 131586 528818 131822 529054
rect 131586 528498 131822 528734
rect 131586 492818 131822 493054
rect 131586 492498 131822 492734
rect 131586 456818 131822 457054
rect 131586 456498 131822 456734
rect 131586 420818 131822 421054
rect 131586 420498 131822 420734
rect 131586 384818 131822 385054
rect 131586 384498 131822 384734
rect 131586 348818 131822 349054
rect 131586 348498 131822 348734
rect 131586 312818 131822 313054
rect 131586 312498 131822 312734
rect 131586 276818 131822 277054
rect 131586 276498 131822 276734
rect 131586 240818 131822 241054
rect 131586 240498 131822 240734
rect 131586 204818 131822 205054
rect 131586 204498 131822 204734
rect 131586 168818 131822 169054
rect 131586 168498 131822 168734
rect 131586 132818 131822 133054
rect 131586 132498 131822 132734
rect 131586 96818 131822 97054
rect 131586 96498 131822 96734
rect 131586 60818 131822 61054
rect 131586 60498 131822 60734
rect 131586 24818 131822 25054
rect 131586 24498 131822 24734
rect 131586 -3402 131822 -3166
rect 131586 -3722 131822 -3486
rect 135186 676418 135422 676654
rect 135186 676098 135422 676334
rect 135186 640418 135422 640654
rect 135186 640098 135422 640334
rect 135186 604418 135422 604654
rect 135186 604098 135422 604334
rect 135186 568418 135422 568654
rect 135186 568098 135422 568334
rect 135186 532418 135422 532654
rect 135186 532098 135422 532334
rect 135186 496418 135422 496654
rect 135186 496098 135422 496334
rect 135186 460418 135422 460654
rect 135186 460098 135422 460334
rect 135186 424418 135422 424654
rect 135186 424098 135422 424334
rect 135186 388418 135422 388654
rect 135186 388098 135422 388334
rect 135186 352418 135422 352654
rect 135186 352098 135422 352334
rect 135186 316418 135422 316654
rect 135186 316098 135422 316334
rect 135186 280418 135422 280654
rect 135186 280098 135422 280334
rect 135186 244418 135422 244654
rect 135186 244098 135422 244334
rect 135186 208418 135422 208654
rect 135186 208098 135422 208334
rect 135186 172418 135422 172654
rect 135186 172098 135422 172334
rect 135186 136418 135422 136654
rect 135186 136098 135422 136334
rect 135186 100418 135422 100654
rect 135186 100098 135422 100334
rect 135186 64418 135422 64654
rect 135186 64098 135422 64334
rect 135186 28418 135422 28654
rect 135186 28098 135422 28334
rect 135186 -5282 135422 -5046
rect 135186 -5602 135422 -5366
rect 156786 710242 157022 710478
rect 156786 709922 157022 710158
rect 153186 708362 153422 708598
rect 153186 708042 153422 708278
rect 149586 706482 149822 706718
rect 149586 706162 149822 706398
rect 138786 680018 139022 680254
rect 138786 679698 139022 679934
rect 138786 644018 139022 644254
rect 138786 643698 139022 643934
rect 138786 608018 139022 608254
rect 138786 607698 139022 607934
rect 138786 572018 139022 572254
rect 138786 571698 139022 571934
rect 138786 536018 139022 536254
rect 138786 535698 139022 535934
rect 138786 500018 139022 500254
rect 138786 499698 139022 499934
rect 138786 464018 139022 464254
rect 138786 463698 139022 463934
rect 138786 428018 139022 428254
rect 138786 427698 139022 427934
rect 138786 392018 139022 392254
rect 138786 391698 139022 391934
rect 138786 356018 139022 356254
rect 138786 355698 139022 355934
rect 138786 320018 139022 320254
rect 138786 319698 139022 319934
rect 138786 284018 139022 284254
rect 138786 283698 139022 283934
rect 138786 248018 139022 248254
rect 138786 247698 139022 247934
rect 138786 212018 139022 212254
rect 138786 211698 139022 211934
rect 138786 176018 139022 176254
rect 138786 175698 139022 175934
rect 138786 140018 139022 140254
rect 138786 139698 139022 139934
rect 138786 104018 139022 104254
rect 138786 103698 139022 103934
rect 138786 68018 139022 68254
rect 138786 67698 139022 67934
rect 138786 32018 139022 32254
rect 138786 31698 139022 31934
rect 120786 -6222 121022 -5986
rect 120786 -6542 121022 -6306
rect 145986 704602 146222 704838
rect 145986 704282 146222 704518
rect 145986 687218 146222 687454
rect 145986 686898 146222 687134
rect 145986 651218 146222 651454
rect 145986 650898 146222 651134
rect 145986 615218 146222 615454
rect 145986 614898 146222 615134
rect 145986 579218 146222 579454
rect 145986 578898 146222 579134
rect 145986 543218 146222 543454
rect 145986 542898 146222 543134
rect 145986 507218 146222 507454
rect 145986 506898 146222 507134
rect 145986 471218 146222 471454
rect 145986 470898 146222 471134
rect 145986 435218 146222 435454
rect 145986 434898 146222 435134
rect 145986 399218 146222 399454
rect 145986 398898 146222 399134
rect 145986 363218 146222 363454
rect 145986 362898 146222 363134
rect 145986 327218 146222 327454
rect 145986 326898 146222 327134
rect 145986 291218 146222 291454
rect 145986 290898 146222 291134
rect 145986 255218 146222 255454
rect 145986 254898 146222 255134
rect 145986 219218 146222 219454
rect 145986 218898 146222 219134
rect 145986 183218 146222 183454
rect 145986 182898 146222 183134
rect 145986 147218 146222 147454
rect 145986 146898 146222 147134
rect 145986 111218 146222 111454
rect 145986 110898 146222 111134
rect 145986 75218 146222 75454
rect 145986 74898 146222 75134
rect 145986 39218 146222 39454
rect 145986 38898 146222 39134
rect 145986 3218 146222 3454
rect 145986 2898 146222 3134
rect 145986 -582 146222 -346
rect 145986 -902 146222 -666
rect 149586 690818 149822 691054
rect 149586 690498 149822 690734
rect 149586 654818 149822 655054
rect 149586 654498 149822 654734
rect 149586 618818 149822 619054
rect 149586 618498 149822 618734
rect 149586 582818 149822 583054
rect 149586 582498 149822 582734
rect 149586 546818 149822 547054
rect 149586 546498 149822 546734
rect 149586 510818 149822 511054
rect 149586 510498 149822 510734
rect 149586 474818 149822 475054
rect 149586 474498 149822 474734
rect 149586 438818 149822 439054
rect 149586 438498 149822 438734
rect 149586 402818 149822 403054
rect 149586 402498 149822 402734
rect 149586 366818 149822 367054
rect 149586 366498 149822 366734
rect 149586 330818 149822 331054
rect 149586 330498 149822 330734
rect 149586 294818 149822 295054
rect 149586 294498 149822 294734
rect 149586 258818 149822 259054
rect 149586 258498 149822 258734
rect 149586 222818 149822 223054
rect 149586 222498 149822 222734
rect 149586 186818 149822 187054
rect 149586 186498 149822 186734
rect 149586 150818 149822 151054
rect 149586 150498 149822 150734
rect 149586 114818 149822 115054
rect 149586 114498 149822 114734
rect 149586 78818 149822 79054
rect 149586 78498 149822 78734
rect 149586 42818 149822 43054
rect 149586 42498 149822 42734
rect 149586 6818 149822 7054
rect 149586 6498 149822 6734
rect 149586 -2462 149822 -2226
rect 149586 -2782 149822 -2546
rect 153186 694418 153422 694654
rect 153186 694098 153422 694334
rect 153186 658418 153422 658654
rect 153186 658098 153422 658334
rect 153186 622418 153422 622654
rect 153186 622098 153422 622334
rect 153186 586418 153422 586654
rect 153186 586098 153422 586334
rect 153186 550418 153422 550654
rect 153186 550098 153422 550334
rect 153186 514418 153422 514654
rect 153186 514098 153422 514334
rect 153186 478418 153422 478654
rect 153186 478098 153422 478334
rect 153186 442418 153422 442654
rect 153186 442098 153422 442334
rect 153186 406418 153422 406654
rect 153186 406098 153422 406334
rect 153186 370418 153422 370654
rect 153186 370098 153422 370334
rect 153186 334418 153422 334654
rect 153186 334098 153422 334334
rect 153186 298418 153422 298654
rect 153186 298098 153422 298334
rect 153186 262418 153422 262654
rect 153186 262098 153422 262334
rect 153186 226418 153422 226654
rect 153186 226098 153422 226334
rect 153186 190418 153422 190654
rect 153186 190098 153422 190334
rect 153186 154418 153422 154654
rect 153186 154098 153422 154334
rect 153186 118418 153422 118654
rect 153186 118098 153422 118334
rect 153186 82418 153422 82654
rect 153186 82098 153422 82334
rect 153186 46418 153422 46654
rect 153186 46098 153422 46334
rect 153186 10418 153422 10654
rect 153186 10098 153422 10334
rect 153186 -4342 153422 -4106
rect 153186 -4662 153422 -4426
rect 174786 711182 175022 711418
rect 174786 710862 175022 711098
rect 171186 709302 171422 709538
rect 171186 708982 171422 709218
rect 167586 707422 167822 707658
rect 167586 707102 167822 707338
rect 156786 698018 157022 698254
rect 156786 697698 157022 697934
rect 156786 662018 157022 662254
rect 156786 661698 157022 661934
rect 156786 626018 157022 626254
rect 156786 625698 157022 625934
rect 156786 590018 157022 590254
rect 156786 589698 157022 589934
rect 156786 554018 157022 554254
rect 156786 553698 157022 553934
rect 156786 518018 157022 518254
rect 156786 517698 157022 517934
rect 156786 482018 157022 482254
rect 156786 481698 157022 481934
rect 156786 446018 157022 446254
rect 156786 445698 157022 445934
rect 156786 410018 157022 410254
rect 156786 409698 157022 409934
rect 156786 374018 157022 374254
rect 156786 373698 157022 373934
rect 156786 338018 157022 338254
rect 156786 337698 157022 337934
rect 156786 302018 157022 302254
rect 156786 301698 157022 301934
rect 156786 266018 157022 266254
rect 156786 265698 157022 265934
rect 156786 230018 157022 230254
rect 156786 229698 157022 229934
rect 156786 194018 157022 194254
rect 156786 193698 157022 193934
rect 156786 158018 157022 158254
rect 156786 157698 157022 157934
rect 156786 122018 157022 122254
rect 156786 121698 157022 121934
rect 156786 86018 157022 86254
rect 156786 85698 157022 85934
rect 156786 50018 157022 50254
rect 156786 49698 157022 49934
rect 156786 14018 157022 14254
rect 156786 13698 157022 13934
rect 138786 -7162 139022 -6926
rect 138786 -7482 139022 -7246
rect 163986 705542 164222 705778
rect 163986 705222 164222 705458
rect 163986 669218 164222 669454
rect 163986 668898 164222 669134
rect 163986 633218 164222 633454
rect 163986 632898 164222 633134
rect 163986 597218 164222 597454
rect 163986 596898 164222 597134
rect 163986 561218 164222 561454
rect 163986 560898 164222 561134
rect 163986 525218 164222 525454
rect 163986 524898 164222 525134
rect 163986 489218 164222 489454
rect 163986 488898 164222 489134
rect 163986 453218 164222 453454
rect 163986 452898 164222 453134
rect 163986 417218 164222 417454
rect 163986 416898 164222 417134
rect 163986 381218 164222 381454
rect 163986 380898 164222 381134
rect 163986 345218 164222 345454
rect 163986 344898 164222 345134
rect 163986 309218 164222 309454
rect 163986 308898 164222 309134
rect 163986 273218 164222 273454
rect 163986 272898 164222 273134
rect 163986 237218 164222 237454
rect 163986 236898 164222 237134
rect 163986 201218 164222 201454
rect 163986 200898 164222 201134
rect 163986 165218 164222 165454
rect 163986 164898 164222 165134
rect 163986 129218 164222 129454
rect 163986 128898 164222 129134
rect 163986 93218 164222 93454
rect 163986 92898 164222 93134
rect 163986 57218 164222 57454
rect 163986 56898 164222 57134
rect 163986 21218 164222 21454
rect 163986 20898 164222 21134
rect 163986 -1522 164222 -1286
rect 163986 -1842 164222 -1606
rect 167586 672818 167822 673054
rect 167586 672498 167822 672734
rect 167586 636818 167822 637054
rect 167586 636498 167822 636734
rect 167586 600818 167822 601054
rect 167586 600498 167822 600734
rect 167586 564818 167822 565054
rect 167586 564498 167822 564734
rect 167586 528818 167822 529054
rect 167586 528498 167822 528734
rect 167586 492818 167822 493054
rect 167586 492498 167822 492734
rect 167586 456818 167822 457054
rect 167586 456498 167822 456734
rect 167586 420818 167822 421054
rect 167586 420498 167822 420734
rect 167586 384818 167822 385054
rect 167586 384498 167822 384734
rect 167586 348818 167822 349054
rect 167586 348498 167822 348734
rect 167586 312818 167822 313054
rect 167586 312498 167822 312734
rect 167586 276818 167822 277054
rect 167586 276498 167822 276734
rect 167586 240818 167822 241054
rect 167586 240498 167822 240734
rect 167586 204818 167822 205054
rect 167586 204498 167822 204734
rect 167586 168818 167822 169054
rect 167586 168498 167822 168734
rect 167586 132818 167822 133054
rect 167586 132498 167822 132734
rect 167586 96818 167822 97054
rect 167586 96498 167822 96734
rect 167586 60818 167822 61054
rect 167586 60498 167822 60734
rect 167586 24818 167822 25054
rect 167586 24498 167822 24734
rect 167586 -3402 167822 -3166
rect 167586 -3722 167822 -3486
rect 171186 676418 171422 676654
rect 171186 676098 171422 676334
rect 171186 640418 171422 640654
rect 171186 640098 171422 640334
rect 171186 604418 171422 604654
rect 171186 604098 171422 604334
rect 171186 568418 171422 568654
rect 171186 568098 171422 568334
rect 171186 532418 171422 532654
rect 171186 532098 171422 532334
rect 171186 496418 171422 496654
rect 171186 496098 171422 496334
rect 171186 460418 171422 460654
rect 171186 460098 171422 460334
rect 171186 424418 171422 424654
rect 171186 424098 171422 424334
rect 171186 388418 171422 388654
rect 171186 388098 171422 388334
rect 171186 352418 171422 352654
rect 171186 352098 171422 352334
rect 171186 316418 171422 316654
rect 171186 316098 171422 316334
rect 171186 280418 171422 280654
rect 171186 280098 171422 280334
rect 171186 244418 171422 244654
rect 171186 244098 171422 244334
rect 171186 208418 171422 208654
rect 171186 208098 171422 208334
rect 171186 172418 171422 172654
rect 171186 172098 171422 172334
rect 171186 136418 171422 136654
rect 171186 136098 171422 136334
rect 171186 100418 171422 100654
rect 171186 100098 171422 100334
rect 171186 64418 171422 64654
rect 171186 64098 171422 64334
rect 171186 28418 171422 28654
rect 171186 28098 171422 28334
rect 171186 -5282 171422 -5046
rect 171186 -5602 171422 -5366
rect 192786 710242 193022 710478
rect 192786 709922 193022 710158
rect 189186 708362 189422 708598
rect 189186 708042 189422 708278
rect 185586 706482 185822 706718
rect 185586 706162 185822 706398
rect 174786 680018 175022 680254
rect 174786 679698 175022 679934
rect 174786 644018 175022 644254
rect 174786 643698 175022 643934
rect 174786 608018 175022 608254
rect 174786 607698 175022 607934
rect 174786 572018 175022 572254
rect 174786 571698 175022 571934
rect 174786 536018 175022 536254
rect 174786 535698 175022 535934
rect 174786 500018 175022 500254
rect 174786 499698 175022 499934
rect 174786 464018 175022 464254
rect 174786 463698 175022 463934
rect 174786 428018 175022 428254
rect 174786 427698 175022 427934
rect 174786 392018 175022 392254
rect 174786 391698 175022 391934
rect 174786 356018 175022 356254
rect 174786 355698 175022 355934
rect 174786 320018 175022 320254
rect 174786 319698 175022 319934
rect 174786 284018 175022 284254
rect 174786 283698 175022 283934
rect 174786 248018 175022 248254
rect 174786 247698 175022 247934
rect 174786 212018 175022 212254
rect 174786 211698 175022 211934
rect 174786 176018 175022 176254
rect 174786 175698 175022 175934
rect 174786 140018 175022 140254
rect 174786 139698 175022 139934
rect 174786 104018 175022 104254
rect 174786 103698 175022 103934
rect 174786 68018 175022 68254
rect 174786 67698 175022 67934
rect 174786 32018 175022 32254
rect 174786 31698 175022 31934
rect 156786 -6222 157022 -5986
rect 156786 -6542 157022 -6306
rect 181986 704602 182222 704838
rect 181986 704282 182222 704518
rect 181986 687218 182222 687454
rect 181986 686898 182222 687134
rect 181986 651218 182222 651454
rect 181986 650898 182222 651134
rect 181986 615218 182222 615454
rect 181986 614898 182222 615134
rect 181986 579218 182222 579454
rect 181986 578898 182222 579134
rect 181986 543218 182222 543454
rect 181986 542898 182222 543134
rect 181986 507218 182222 507454
rect 181986 506898 182222 507134
rect 181986 471218 182222 471454
rect 181986 470898 182222 471134
rect 181986 435218 182222 435454
rect 181986 434898 182222 435134
rect 181986 399218 182222 399454
rect 181986 398898 182222 399134
rect 181986 363218 182222 363454
rect 181986 362898 182222 363134
rect 181986 327218 182222 327454
rect 181986 326898 182222 327134
rect 181986 291218 182222 291454
rect 181986 290898 182222 291134
rect 181986 255218 182222 255454
rect 181986 254898 182222 255134
rect 181986 219218 182222 219454
rect 181986 218898 182222 219134
rect 181986 183218 182222 183454
rect 181986 182898 182222 183134
rect 181986 147218 182222 147454
rect 181986 146898 182222 147134
rect 181986 111218 182222 111454
rect 181986 110898 182222 111134
rect 181986 75218 182222 75454
rect 181986 74898 182222 75134
rect 181986 39218 182222 39454
rect 181986 38898 182222 39134
rect 181986 3218 182222 3454
rect 181986 2898 182222 3134
rect 181986 -582 182222 -346
rect 181986 -902 182222 -666
rect 185586 690818 185822 691054
rect 185586 690498 185822 690734
rect 185586 654818 185822 655054
rect 185586 654498 185822 654734
rect 185586 618818 185822 619054
rect 185586 618498 185822 618734
rect 185586 582818 185822 583054
rect 185586 582498 185822 582734
rect 185586 546818 185822 547054
rect 185586 546498 185822 546734
rect 185586 510818 185822 511054
rect 185586 510498 185822 510734
rect 185586 474818 185822 475054
rect 185586 474498 185822 474734
rect 185586 438818 185822 439054
rect 185586 438498 185822 438734
rect 185586 402818 185822 403054
rect 185586 402498 185822 402734
rect 185586 366818 185822 367054
rect 185586 366498 185822 366734
rect 185586 330818 185822 331054
rect 185586 330498 185822 330734
rect 185586 294818 185822 295054
rect 185586 294498 185822 294734
rect 185586 258818 185822 259054
rect 185586 258498 185822 258734
rect 185586 222818 185822 223054
rect 185586 222498 185822 222734
rect 185586 186818 185822 187054
rect 185586 186498 185822 186734
rect 185586 150818 185822 151054
rect 185586 150498 185822 150734
rect 185586 114818 185822 115054
rect 185586 114498 185822 114734
rect 185586 78818 185822 79054
rect 185586 78498 185822 78734
rect 185586 42818 185822 43054
rect 185586 42498 185822 42734
rect 185586 6818 185822 7054
rect 185586 6498 185822 6734
rect 185586 -2462 185822 -2226
rect 185586 -2782 185822 -2546
rect 189186 694418 189422 694654
rect 189186 694098 189422 694334
rect 189186 658418 189422 658654
rect 189186 658098 189422 658334
rect 189186 622418 189422 622654
rect 189186 622098 189422 622334
rect 189186 586418 189422 586654
rect 189186 586098 189422 586334
rect 189186 550418 189422 550654
rect 189186 550098 189422 550334
rect 189186 514418 189422 514654
rect 189186 514098 189422 514334
rect 189186 478418 189422 478654
rect 189186 478098 189422 478334
rect 189186 442418 189422 442654
rect 189186 442098 189422 442334
rect 189186 406418 189422 406654
rect 189186 406098 189422 406334
rect 189186 370418 189422 370654
rect 189186 370098 189422 370334
rect 189186 334418 189422 334654
rect 189186 334098 189422 334334
rect 189186 298418 189422 298654
rect 189186 298098 189422 298334
rect 189186 262418 189422 262654
rect 189186 262098 189422 262334
rect 189186 226418 189422 226654
rect 189186 226098 189422 226334
rect 189186 190418 189422 190654
rect 189186 190098 189422 190334
rect 189186 154418 189422 154654
rect 189186 154098 189422 154334
rect 189186 118418 189422 118654
rect 189186 118098 189422 118334
rect 189186 82418 189422 82654
rect 189186 82098 189422 82334
rect 189186 46418 189422 46654
rect 189186 46098 189422 46334
rect 189186 10418 189422 10654
rect 189186 10098 189422 10334
rect 189186 -4342 189422 -4106
rect 189186 -4662 189422 -4426
rect 210786 711182 211022 711418
rect 210786 710862 211022 711098
rect 207186 709302 207422 709538
rect 207186 708982 207422 709218
rect 203586 707422 203822 707658
rect 203586 707102 203822 707338
rect 192786 698018 193022 698254
rect 192786 697698 193022 697934
rect 192786 662018 193022 662254
rect 192786 661698 193022 661934
rect 192786 626018 193022 626254
rect 192786 625698 193022 625934
rect 192786 590018 193022 590254
rect 192786 589698 193022 589934
rect 192786 554018 193022 554254
rect 192786 553698 193022 553934
rect 192786 518018 193022 518254
rect 192786 517698 193022 517934
rect 192786 482018 193022 482254
rect 192786 481698 193022 481934
rect 192786 446018 193022 446254
rect 192786 445698 193022 445934
rect 192786 410018 193022 410254
rect 192786 409698 193022 409934
rect 192786 374018 193022 374254
rect 192786 373698 193022 373934
rect 192786 338018 193022 338254
rect 192786 337698 193022 337934
rect 192786 302018 193022 302254
rect 192786 301698 193022 301934
rect 192786 266018 193022 266254
rect 192786 265698 193022 265934
rect 192786 230018 193022 230254
rect 192786 229698 193022 229934
rect 192786 194018 193022 194254
rect 192786 193698 193022 193934
rect 192786 158018 193022 158254
rect 192786 157698 193022 157934
rect 192786 122018 193022 122254
rect 192786 121698 193022 121934
rect 192786 86018 193022 86254
rect 192786 85698 193022 85934
rect 192786 50018 193022 50254
rect 192786 49698 193022 49934
rect 192786 14018 193022 14254
rect 192786 13698 193022 13934
rect 174786 -7162 175022 -6926
rect 174786 -7482 175022 -7246
rect 199986 705542 200222 705778
rect 199986 705222 200222 705458
rect 199986 669218 200222 669454
rect 199986 668898 200222 669134
rect 199986 633218 200222 633454
rect 199986 632898 200222 633134
rect 199986 597218 200222 597454
rect 199986 596898 200222 597134
rect 199986 561218 200222 561454
rect 199986 560898 200222 561134
rect 199986 525218 200222 525454
rect 199986 524898 200222 525134
rect 199986 489218 200222 489454
rect 199986 488898 200222 489134
rect 199986 453218 200222 453454
rect 199986 452898 200222 453134
rect 199986 417218 200222 417454
rect 199986 416898 200222 417134
rect 199986 381218 200222 381454
rect 199986 380898 200222 381134
rect 199986 345218 200222 345454
rect 199986 344898 200222 345134
rect 199986 309218 200222 309454
rect 199986 308898 200222 309134
rect 199986 273218 200222 273454
rect 199986 272898 200222 273134
rect 199986 237218 200222 237454
rect 199986 236898 200222 237134
rect 199986 201218 200222 201454
rect 199986 200898 200222 201134
rect 199986 165218 200222 165454
rect 199986 164898 200222 165134
rect 199986 129218 200222 129454
rect 199986 128898 200222 129134
rect 199986 93218 200222 93454
rect 199986 92898 200222 93134
rect 199986 57218 200222 57454
rect 199986 56898 200222 57134
rect 199986 21218 200222 21454
rect 199986 20898 200222 21134
rect 199986 -1522 200222 -1286
rect 199986 -1842 200222 -1606
rect 203586 672818 203822 673054
rect 203586 672498 203822 672734
rect 203586 636818 203822 637054
rect 203586 636498 203822 636734
rect 203586 600818 203822 601054
rect 203586 600498 203822 600734
rect 203586 564818 203822 565054
rect 203586 564498 203822 564734
rect 203586 528818 203822 529054
rect 203586 528498 203822 528734
rect 203586 492818 203822 493054
rect 203586 492498 203822 492734
rect 203586 456818 203822 457054
rect 203586 456498 203822 456734
rect 203586 420818 203822 421054
rect 203586 420498 203822 420734
rect 203586 384818 203822 385054
rect 203586 384498 203822 384734
rect 203586 348818 203822 349054
rect 203586 348498 203822 348734
rect 203586 312818 203822 313054
rect 203586 312498 203822 312734
rect 203586 276818 203822 277054
rect 203586 276498 203822 276734
rect 203586 240818 203822 241054
rect 203586 240498 203822 240734
rect 203586 204818 203822 205054
rect 203586 204498 203822 204734
rect 203586 168818 203822 169054
rect 203586 168498 203822 168734
rect 203586 132818 203822 133054
rect 203586 132498 203822 132734
rect 203586 96818 203822 97054
rect 203586 96498 203822 96734
rect 203586 60818 203822 61054
rect 203586 60498 203822 60734
rect 203586 24818 203822 25054
rect 203586 24498 203822 24734
rect 203586 -3402 203822 -3166
rect 203586 -3722 203822 -3486
rect 207186 676418 207422 676654
rect 207186 676098 207422 676334
rect 207186 640418 207422 640654
rect 207186 640098 207422 640334
rect 207186 604418 207422 604654
rect 207186 604098 207422 604334
rect 207186 568418 207422 568654
rect 207186 568098 207422 568334
rect 207186 532418 207422 532654
rect 207186 532098 207422 532334
rect 207186 496418 207422 496654
rect 207186 496098 207422 496334
rect 207186 460418 207422 460654
rect 207186 460098 207422 460334
rect 207186 424418 207422 424654
rect 207186 424098 207422 424334
rect 207186 388418 207422 388654
rect 207186 388098 207422 388334
rect 207186 352418 207422 352654
rect 207186 352098 207422 352334
rect 207186 316418 207422 316654
rect 207186 316098 207422 316334
rect 207186 280418 207422 280654
rect 207186 280098 207422 280334
rect 207186 244418 207422 244654
rect 207186 244098 207422 244334
rect 207186 208418 207422 208654
rect 207186 208098 207422 208334
rect 207186 172418 207422 172654
rect 207186 172098 207422 172334
rect 207186 136418 207422 136654
rect 207186 136098 207422 136334
rect 207186 100418 207422 100654
rect 207186 100098 207422 100334
rect 207186 64418 207422 64654
rect 207186 64098 207422 64334
rect 207186 28418 207422 28654
rect 207186 28098 207422 28334
rect 207186 -5282 207422 -5046
rect 207186 -5602 207422 -5366
rect 228786 710242 229022 710478
rect 228786 709922 229022 710158
rect 225186 708362 225422 708598
rect 225186 708042 225422 708278
rect 221586 706482 221822 706718
rect 221586 706162 221822 706398
rect 210786 680018 211022 680254
rect 210786 679698 211022 679934
rect 210786 644018 211022 644254
rect 210786 643698 211022 643934
rect 210786 608018 211022 608254
rect 210786 607698 211022 607934
rect 210786 572018 211022 572254
rect 210786 571698 211022 571934
rect 210786 536018 211022 536254
rect 210786 535698 211022 535934
rect 210786 500018 211022 500254
rect 210786 499698 211022 499934
rect 210786 464018 211022 464254
rect 210786 463698 211022 463934
rect 210786 428018 211022 428254
rect 210786 427698 211022 427934
rect 210786 392018 211022 392254
rect 210786 391698 211022 391934
rect 210786 356018 211022 356254
rect 210786 355698 211022 355934
rect 210786 320018 211022 320254
rect 210786 319698 211022 319934
rect 210786 284018 211022 284254
rect 210786 283698 211022 283934
rect 210786 248018 211022 248254
rect 210786 247698 211022 247934
rect 210786 212018 211022 212254
rect 210786 211698 211022 211934
rect 210786 176018 211022 176254
rect 210786 175698 211022 175934
rect 210786 140018 211022 140254
rect 210786 139698 211022 139934
rect 210786 104018 211022 104254
rect 210786 103698 211022 103934
rect 210786 68018 211022 68254
rect 210786 67698 211022 67934
rect 210786 32018 211022 32254
rect 210786 31698 211022 31934
rect 192786 -6222 193022 -5986
rect 192786 -6542 193022 -6306
rect 217986 704602 218222 704838
rect 217986 704282 218222 704518
rect 217986 687218 218222 687454
rect 217986 686898 218222 687134
rect 217986 651218 218222 651454
rect 217986 650898 218222 651134
rect 217986 615218 218222 615454
rect 217986 614898 218222 615134
rect 217986 579218 218222 579454
rect 217986 578898 218222 579134
rect 217986 543218 218222 543454
rect 217986 542898 218222 543134
rect 217986 507218 218222 507454
rect 217986 506898 218222 507134
rect 217986 471218 218222 471454
rect 217986 470898 218222 471134
rect 217986 435218 218222 435454
rect 217986 434898 218222 435134
rect 217986 399218 218222 399454
rect 217986 398898 218222 399134
rect 217986 363218 218222 363454
rect 217986 362898 218222 363134
rect 217986 327218 218222 327454
rect 217986 326898 218222 327134
rect 217986 291218 218222 291454
rect 217986 290898 218222 291134
rect 217986 255218 218222 255454
rect 217986 254898 218222 255134
rect 217986 219218 218222 219454
rect 217986 218898 218222 219134
rect 217986 183218 218222 183454
rect 217986 182898 218222 183134
rect 217986 147218 218222 147454
rect 217986 146898 218222 147134
rect 217986 111218 218222 111454
rect 217986 110898 218222 111134
rect 217986 75218 218222 75454
rect 217986 74898 218222 75134
rect 217986 39218 218222 39454
rect 217986 38898 218222 39134
rect 217986 3218 218222 3454
rect 217986 2898 218222 3134
rect 217986 -582 218222 -346
rect 217986 -902 218222 -666
rect 221586 690818 221822 691054
rect 221586 690498 221822 690734
rect 221586 654818 221822 655054
rect 221586 654498 221822 654734
rect 221586 618818 221822 619054
rect 221586 618498 221822 618734
rect 221586 582818 221822 583054
rect 221586 582498 221822 582734
rect 221586 546818 221822 547054
rect 221586 546498 221822 546734
rect 221586 510818 221822 511054
rect 221586 510498 221822 510734
rect 221586 474818 221822 475054
rect 221586 474498 221822 474734
rect 221586 438818 221822 439054
rect 221586 438498 221822 438734
rect 221586 402818 221822 403054
rect 221586 402498 221822 402734
rect 221586 366818 221822 367054
rect 221586 366498 221822 366734
rect 221586 330818 221822 331054
rect 221586 330498 221822 330734
rect 221586 294818 221822 295054
rect 221586 294498 221822 294734
rect 221586 258818 221822 259054
rect 221586 258498 221822 258734
rect 221586 222818 221822 223054
rect 221586 222498 221822 222734
rect 221586 186818 221822 187054
rect 221586 186498 221822 186734
rect 221586 150818 221822 151054
rect 221586 150498 221822 150734
rect 221586 114818 221822 115054
rect 221586 114498 221822 114734
rect 221586 78818 221822 79054
rect 221586 78498 221822 78734
rect 221586 42818 221822 43054
rect 221586 42498 221822 42734
rect 221586 6818 221822 7054
rect 221586 6498 221822 6734
rect 221586 -2462 221822 -2226
rect 221586 -2782 221822 -2546
rect 225186 694418 225422 694654
rect 225186 694098 225422 694334
rect 225186 658418 225422 658654
rect 225186 658098 225422 658334
rect 225186 622418 225422 622654
rect 225186 622098 225422 622334
rect 225186 586418 225422 586654
rect 225186 586098 225422 586334
rect 225186 550418 225422 550654
rect 225186 550098 225422 550334
rect 225186 514418 225422 514654
rect 225186 514098 225422 514334
rect 225186 478418 225422 478654
rect 225186 478098 225422 478334
rect 225186 442418 225422 442654
rect 225186 442098 225422 442334
rect 225186 406418 225422 406654
rect 225186 406098 225422 406334
rect 225186 370418 225422 370654
rect 225186 370098 225422 370334
rect 225186 334418 225422 334654
rect 225186 334098 225422 334334
rect 225186 298418 225422 298654
rect 225186 298098 225422 298334
rect 225186 262418 225422 262654
rect 225186 262098 225422 262334
rect 225186 226418 225422 226654
rect 225186 226098 225422 226334
rect 225186 190418 225422 190654
rect 225186 190098 225422 190334
rect 225186 154418 225422 154654
rect 225186 154098 225422 154334
rect 225186 118418 225422 118654
rect 225186 118098 225422 118334
rect 225186 82418 225422 82654
rect 225186 82098 225422 82334
rect 225186 46418 225422 46654
rect 225186 46098 225422 46334
rect 225186 10418 225422 10654
rect 225186 10098 225422 10334
rect 225186 -4342 225422 -4106
rect 225186 -4662 225422 -4426
rect 246786 711182 247022 711418
rect 246786 710862 247022 711098
rect 243186 709302 243422 709538
rect 243186 708982 243422 709218
rect 239586 707422 239822 707658
rect 239586 707102 239822 707338
rect 228786 698018 229022 698254
rect 228786 697698 229022 697934
rect 228786 662018 229022 662254
rect 228786 661698 229022 661934
rect 228786 626018 229022 626254
rect 228786 625698 229022 625934
rect 228786 590018 229022 590254
rect 228786 589698 229022 589934
rect 228786 554018 229022 554254
rect 228786 553698 229022 553934
rect 228786 518018 229022 518254
rect 228786 517698 229022 517934
rect 228786 482018 229022 482254
rect 228786 481698 229022 481934
rect 228786 446018 229022 446254
rect 228786 445698 229022 445934
rect 228786 410018 229022 410254
rect 235986 705542 236222 705778
rect 235986 705222 236222 705458
rect 235986 669218 236222 669454
rect 235986 668898 236222 669134
rect 235986 633218 236222 633454
rect 235986 632898 236222 633134
rect 235986 597218 236222 597454
rect 235986 596898 236222 597134
rect 235986 561218 236222 561454
rect 235986 560898 236222 561134
rect 235986 525218 236222 525454
rect 235986 524898 236222 525134
rect 235986 489218 236222 489454
rect 235986 488898 236222 489134
rect 235986 453218 236222 453454
rect 235986 452898 236222 453134
rect 235986 417218 236222 417454
rect 235986 416898 236222 417134
rect 239586 672818 239822 673054
rect 239586 672498 239822 672734
rect 239586 636818 239822 637054
rect 239586 636498 239822 636734
rect 239586 600818 239822 601054
rect 239586 600498 239822 600734
rect 239586 564818 239822 565054
rect 239586 564498 239822 564734
rect 239586 528818 239822 529054
rect 239586 528498 239822 528734
rect 239586 492818 239822 493054
rect 239586 492498 239822 492734
rect 239586 456818 239822 457054
rect 239586 456498 239822 456734
rect 239586 420818 239822 421054
rect 239586 420498 239822 420734
rect 243186 676418 243422 676654
rect 243186 676098 243422 676334
rect 243186 640418 243422 640654
rect 243186 640098 243422 640334
rect 243186 604418 243422 604654
rect 243186 604098 243422 604334
rect 243186 568418 243422 568654
rect 243186 568098 243422 568334
rect 243186 532418 243422 532654
rect 243186 532098 243422 532334
rect 243186 496418 243422 496654
rect 243186 496098 243422 496334
rect 243186 460418 243422 460654
rect 243186 460098 243422 460334
rect 243186 424418 243422 424654
rect 243186 424098 243422 424334
rect 264786 710242 265022 710478
rect 264786 709922 265022 710158
rect 261186 708362 261422 708598
rect 261186 708042 261422 708278
rect 257586 706482 257822 706718
rect 257586 706162 257822 706398
rect 246786 680018 247022 680254
rect 246786 679698 247022 679934
rect 246786 644018 247022 644254
rect 246786 643698 247022 643934
rect 246786 608018 247022 608254
rect 246786 607698 247022 607934
rect 246786 572018 247022 572254
rect 246786 571698 247022 571934
rect 246786 536018 247022 536254
rect 246786 535698 247022 535934
rect 246786 500018 247022 500254
rect 246786 499698 247022 499934
rect 246786 464018 247022 464254
rect 246786 463698 247022 463934
rect 246786 428018 247022 428254
rect 246786 427698 247022 427934
rect 253986 704602 254222 704838
rect 253986 704282 254222 704518
rect 253986 687218 254222 687454
rect 253986 686898 254222 687134
rect 253986 651218 254222 651454
rect 253986 650898 254222 651134
rect 253986 615218 254222 615454
rect 253986 614898 254222 615134
rect 253986 579218 254222 579454
rect 253986 578898 254222 579134
rect 253986 543218 254222 543454
rect 253986 542898 254222 543134
rect 253986 507218 254222 507454
rect 253986 506898 254222 507134
rect 253986 471218 254222 471454
rect 253986 470898 254222 471134
rect 253986 435218 254222 435454
rect 253986 434898 254222 435134
rect 257586 690818 257822 691054
rect 257586 690498 257822 690734
rect 257586 654818 257822 655054
rect 257586 654498 257822 654734
rect 257586 618818 257822 619054
rect 257586 618498 257822 618734
rect 257586 582818 257822 583054
rect 257586 582498 257822 582734
rect 257586 546818 257822 547054
rect 257586 546498 257822 546734
rect 257586 510818 257822 511054
rect 257586 510498 257822 510734
rect 257586 474818 257822 475054
rect 257586 474498 257822 474734
rect 257586 438818 257822 439054
rect 257586 438498 257822 438734
rect 261186 694418 261422 694654
rect 261186 694098 261422 694334
rect 261186 658418 261422 658654
rect 261186 658098 261422 658334
rect 261186 622418 261422 622654
rect 261186 622098 261422 622334
rect 261186 586418 261422 586654
rect 261186 586098 261422 586334
rect 261186 550418 261422 550654
rect 261186 550098 261422 550334
rect 261186 514418 261422 514654
rect 261186 514098 261422 514334
rect 261186 478418 261422 478654
rect 261186 478098 261422 478334
rect 261186 442418 261422 442654
rect 261186 442098 261422 442334
rect 282786 711182 283022 711418
rect 282786 710862 283022 711098
rect 279186 709302 279422 709538
rect 279186 708982 279422 709218
rect 275586 707422 275822 707658
rect 275586 707102 275822 707338
rect 264786 698018 265022 698254
rect 264786 697698 265022 697934
rect 264786 662018 265022 662254
rect 264786 661698 265022 661934
rect 264786 626018 265022 626254
rect 264786 625698 265022 625934
rect 264786 590018 265022 590254
rect 264786 589698 265022 589934
rect 264786 554018 265022 554254
rect 264786 553698 265022 553934
rect 264786 518018 265022 518254
rect 264786 517698 265022 517934
rect 264786 482018 265022 482254
rect 264786 481698 265022 481934
rect 264786 446018 265022 446254
rect 264786 445698 265022 445934
rect 271986 705542 272222 705778
rect 271986 705222 272222 705458
rect 271986 669218 272222 669454
rect 271986 668898 272222 669134
rect 271986 633218 272222 633454
rect 271986 632898 272222 633134
rect 271986 597218 272222 597454
rect 271986 596898 272222 597134
rect 271986 561218 272222 561454
rect 271986 560898 272222 561134
rect 271986 525218 272222 525454
rect 271986 524898 272222 525134
rect 271986 489218 272222 489454
rect 271986 488898 272222 489134
rect 271986 453218 272222 453454
rect 271986 452898 272222 453134
rect 271986 417218 272222 417454
rect 271986 416898 272222 417134
rect 275586 672818 275822 673054
rect 275586 672498 275822 672734
rect 275586 636818 275822 637054
rect 275586 636498 275822 636734
rect 275586 600818 275822 601054
rect 275586 600498 275822 600734
rect 275586 564818 275822 565054
rect 275586 564498 275822 564734
rect 275586 528818 275822 529054
rect 275586 528498 275822 528734
rect 275586 492818 275822 493054
rect 275586 492498 275822 492734
rect 275586 456818 275822 457054
rect 275586 456498 275822 456734
rect 275586 420818 275822 421054
rect 275586 420498 275822 420734
rect 279186 676418 279422 676654
rect 279186 676098 279422 676334
rect 279186 640418 279422 640654
rect 279186 640098 279422 640334
rect 279186 604418 279422 604654
rect 279186 604098 279422 604334
rect 279186 568418 279422 568654
rect 279186 568098 279422 568334
rect 279186 532418 279422 532654
rect 279186 532098 279422 532334
rect 279186 496418 279422 496654
rect 279186 496098 279422 496334
rect 279186 460418 279422 460654
rect 279186 460098 279422 460334
rect 279186 424418 279422 424654
rect 279186 424098 279422 424334
rect 300786 710242 301022 710478
rect 300786 709922 301022 710158
rect 297186 708362 297422 708598
rect 297186 708042 297422 708278
rect 293586 706482 293822 706718
rect 293586 706162 293822 706398
rect 282786 680018 283022 680254
rect 282786 679698 283022 679934
rect 282786 644018 283022 644254
rect 282786 643698 283022 643934
rect 282786 608018 283022 608254
rect 282786 607698 283022 607934
rect 282786 572018 283022 572254
rect 282786 571698 283022 571934
rect 282786 536018 283022 536254
rect 282786 535698 283022 535934
rect 282786 500018 283022 500254
rect 282786 499698 283022 499934
rect 282786 464018 283022 464254
rect 282786 463698 283022 463934
rect 282786 428018 283022 428254
rect 282786 427698 283022 427934
rect 289986 704602 290222 704838
rect 289986 704282 290222 704518
rect 289986 687218 290222 687454
rect 289986 686898 290222 687134
rect 289986 651218 290222 651454
rect 289986 650898 290222 651134
rect 289986 615218 290222 615454
rect 289986 614898 290222 615134
rect 289986 579218 290222 579454
rect 289986 578898 290222 579134
rect 289986 543218 290222 543454
rect 289986 542898 290222 543134
rect 289986 507218 290222 507454
rect 289986 506898 290222 507134
rect 289986 471218 290222 471454
rect 289986 470898 290222 471134
rect 289986 435218 290222 435454
rect 289986 434898 290222 435134
rect 293586 690818 293822 691054
rect 293586 690498 293822 690734
rect 293586 654818 293822 655054
rect 293586 654498 293822 654734
rect 293586 618818 293822 619054
rect 293586 618498 293822 618734
rect 293586 582818 293822 583054
rect 293586 582498 293822 582734
rect 293586 546818 293822 547054
rect 293586 546498 293822 546734
rect 293586 510818 293822 511054
rect 293586 510498 293822 510734
rect 293586 474818 293822 475054
rect 293586 474498 293822 474734
rect 293586 438818 293822 439054
rect 293586 438498 293822 438734
rect 297186 694418 297422 694654
rect 297186 694098 297422 694334
rect 297186 658418 297422 658654
rect 297186 658098 297422 658334
rect 297186 622418 297422 622654
rect 297186 622098 297422 622334
rect 297186 586418 297422 586654
rect 297186 586098 297422 586334
rect 297186 550418 297422 550654
rect 297186 550098 297422 550334
rect 297186 514418 297422 514654
rect 297186 514098 297422 514334
rect 297186 478418 297422 478654
rect 297186 478098 297422 478334
rect 297186 442418 297422 442654
rect 297186 442098 297422 442334
rect 318786 711182 319022 711418
rect 318786 710862 319022 711098
rect 315186 709302 315422 709538
rect 315186 708982 315422 709218
rect 311586 707422 311822 707658
rect 311586 707102 311822 707338
rect 300786 698018 301022 698254
rect 300786 697698 301022 697934
rect 300786 662018 301022 662254
rect 300786 661698 301022 661934
rect 300786 626018 301022 626254
rect 300786 625698 301022 625934
rect 300786 590018 301022 590254
rect 300786 589698 301022 589934
rect 300786 554018 301022 554254
rect 300786 553698 301022 553934
rect 300786 518018 301022 518254
rect 300786 517698 301022 517934
rect 300786 482018 301022 482254
rect 300786 481698 301022 481934
rect 300786 446018 301022 446254
rect 300786 445698 301022 445934
rect 307986 705542 308222 705778
rect 307986 705222 308222 705458
rect 307986 669218 308222 669454
rect 307986 668898 308222 669134
rect 307986 633218 308222 633454
rect 307986 632898 308222 633134
rect 307986 597218 308222 597454
rect 307986 596898 308222 597134
rect 307986 561218 308222 561454
rect 307986 560898 308222 561134
rect 307986 525218 308222 525454
rect 307986 524898 308222 525134
rect 307986 489218 308222 489454
rect 307986 488898 308222 489134
rect 307986 453218 308222 453454
rect 307986 452898 308222 453134
rect 307986 417218 308222 417454
rect 307986 416898 308222 417134
rect 228786 409698 229022 409934
rect 228786 374018 229022 374254
rect 228786 373698 229022 373934
rect 307986 381218 308222 381454
rect 307986 380898 308222 381134
rect 307986 345218 308222 345454
rect 307986 344898 308222 345134
rect 228786 338018 229022 338254
rect 228786 337698 229022 337934
rect 228786 302018 229022 302254
rect 228786 301698 229022 301934
rect 228786 266018 229022 266254
rect 228786 265698 229022 265934
rect 228786 230018 229022 230254
rect 228786 229698 229022 229934
rect 228786 194018 229022 194254
rect 228786 193698 229022 193934
rect 228786 158018 229022 158254
rect 228786 157698 229022 157934
rect 228786 122018 229022 122254
rect 228786 121698 229022 121934
rect 228786 86018 229022 86254
rect 228786 85698 229022 85934
rect 228786 50018 229022 50254
rect 228786 49698 229022 49934
rect 228786 14018 229022 14254
rect 228786 13698 229022 13934
rect 210786 -7162 211022 -6926
rect 210786 -7482 211022 -7246
rect 235986 309218 236222 309454
rect 235986 308898 236222 309134
rect 235986 273218 236222 273454
rect 235986 272898 236222 273134
rect 235986 237218 236222 237454
rect 235986 236898 236222 237134
rect 235986 201218 236222 201454
rect 235986 200898 236222 201134
rect 235986 165218 236222 165454
rect 235986 164898 236222 165134
rect 235986 129218 236222 129454
rect 235986 128898 236222 129134
rect 235986 93218 236222 93454
rect 235986 92898 236222 93134
rect 235986 57218 236222 57454
rect 235986 56898 236222 57134
rect 235986 21218 236222 21454
rect 235986 20898 236222 21134
rect 235986 -1522 236222 -1286
rect 235986 -1842 236222 -1606
rect 239586 312818 239822 313054
rect 239586 312498 239822 312734
rect 239586 276818 239822 277054
rect 239586 276498 239822 276734
rect 239586 240818 239822 241054
rect 239586 240498 239822 240734
rect 239586 204818 239822 205054
rect 239586 204498 239822 204734
rect 239586 168818 239822 169054
rect 239586 168498 239822 168734
rect 239586 132818 239822 133054
rect 239586 132498 239822 132734
rect 239586 96818 239822 97054
rect 239586 96498 239822 96734
rect 239586 60818 239822 61054
rect 239586 60498 239822 60734
rect 239586 24818 239822 25054
rect 239586 24498 239822 24734
rect 239586 -3402 239822 -3166
rect 239586 -3722 239822 -3486
rect 243186 316418 243422 316654
rect 243186 316098 243422 316334
rect 243186 280418 243422 280654
rect 243186 280098 243422 280334
rect 243186 244418 243422 244654
rect 243186 244098 243422 244334
rect 243186 208418 243422 208654
rect 243186 208098 243422 208334
rect 243186 172418 243422 172654
rect 243186 172098 243422 172334
rect 243186 136418 243422 136654
rect 243186 136098 243422 136334
rect 243186 100418 243422 100654
rect 243186 100098 243422 100334
rect 243186 64418 243422 64654
rect 243186 64098 243422 64334
rect 243186 28418 243422 28654
rect 243186 28098 243422 28334
rect 243186 -5282 243422 -5046
rect 243186 -5602 243422 -5366
rect 246786 320018 247022 320254
rect 246786 319698 247022 319934
rect 246786 284018 247022 284254
rect 246786 283698 247022 283934
rect 246786 248018 247022 248254
rect 246786 247698 247022 247934
rect 246786 212018 247022 212254
rect 246786 211698 247022 211934
rect 246786 176018 247022 176254
rect 246786 175698 247022 175934
rect 246786 140018 247022 140254
rect 246786 139698 247022 139934
rect 246786 104018 247022 104254
rect 246786 103698 247022 103934
rect 246786 68018 247022 68254
rect 246786 67698 247022 67934
rect 246786 32018 247022 32254
rect 246786 31698 247022 31934
rect 228786 -6222 229022 -5986
rect 228786 -6542 229022 -6306
rect 253986 327218 254222 327454
rect 253986 326898 254222 327134
rect 253986 291218 254222 291454
rect 253986 290898 254222 291134
rect 253986 255218 254222 255454
rect 253986 254898 254222 255134
rect 253986 219218 254222 219454
rect 253986 218898 254222 219134
rect 253986 183218 254222 183454
rect 253986 182898 254222 183134
rect 253986 147218 254222 147454
rect 253986 146898 254222 147134
rect 253986 111218 254222 111454
rect 253986 110898 254222 111134
rect 253986 75218 254222 75454
rect 253986 74898 254222 75134
rect 253986 39218 254222 39454
rect 253986 38898 254222 39134
rect 253986 3218 254222 3454
rect 253986 2898 254222 3134
rect 253986 -582 254222 -346
rect 253986 -902 254222 -666
rect 257586 330818 257822 331054
rect 257586 330498 257822 330734
rect 257586 294818 257822 295054
rect 257586 294498 257822 294734
rect 257586 258818 257822 259054
rect 257586 258498 257822 258734
rect 257586 222818 257822 223054
rect 257586 222498 257822 222734
rect 257586 186818 257822 187054
rect 257586 186498 257822 186734
rect 257586 150818 257822 151054
rect 257586 150498 257822 150734
rect 257586 114818 257822 115054
rect 257586 114498 257822 114734
rect 257586 78818 257822 79054
rect 257586 78498 257822 78734
rect 257586 42818 257822 43054
rect 257586 42498 257822 42734
rect 257586 6818 257822 7054
rect 257586 6498 257822 6734
rect 257586 -2462 257822 -2226
rect 257586 -2782 257822 -2546
rect 261186 334418 261422 334654
rect 261186 334098 261422 334334
rect 261186 298418 261422 298654
rect 261186 298098 261422 298334
rect 261186 262418 261422 262654
rect 261186 262098 261422 262334
rect 261186 226418 261422 226654
rect 261186 226098 261422 226334
rect 261186 190418 261422 190654
rect 261186 190098 261422 190334
rect 261186 154418 261422 154654
rect 261186 154098 261422 154334
rect 261186 118418 261422 118654
rect 261186 118098 261422 118334
rect 261186 82418 261422 82654
rect 261186 82098 261422 82334
rect 261186 46418 261422 46654
rect 261186 46098 261422 46334
rect 261186 10418 261422 10654
rect 261186 10098 261422 10334
rect 261186 -4342 261422 -4106
rect 261186 -4662 261422 -4426
rect 264786 302018 265022 302254
rect 264786 301698 265022 301934
rect 264786 266018 265022 266254
rect 264786 265698 265022 265934
rect 264786 230018 265022 230254
rect 264786 229698 265022 229934
rect 264786 194018 265022 194254
rect 264786 193698 265022 193934
rect 264786 158018 265022 158254
rect 264786 157698 265022 157934
rect 264786 122018 265022 122254
rect 264786 121698 265022 121934
rect 264786 86018 265022 86254
rect 264786 85698 265022 85934
rect 264786 50018 265022 50254
rect 264786 49698 265022 49934
rect 264786 14018 265022 14254
rect 264786 13698 265022 13934
rect 246786 -7162 247022 -6926
rect 246786 -7482 247022 -7246
rect 271986 309218 272222 309454
rect 271986 308898 272222 309134
rect 271986 273218 272222 273454
rect 271986 272898 272222 273134
rect 271986 237218 272222 237454
rect 271986 236898 272222 237134
rect 271986 201218 272222 201454
rect 271986 200898 272222 201134
rect 271986 165218 272222 165454
rect 271986 164898 272222 165134
rect 271986 129218 272222 129454
rect 271986 128898 272222 129134
rect 271986 93218 272222 93454
rect 271986 92898 272222 93134
rect 271986 57218 272222 57454
rect 271986 56898 272222 57134
rect 271986 21218 272222 21454
rect 271986 20898 272222 21134
rect 271986 -1522 272222 -1286
rect 271986 -1842 272222 -1606
rect 275586 312818 275822 313054
rect 275586 312498 275822 312734
rect 275586 276818 275822 277054
rect 275586 276498 275822 276734
rect 275586 240818 275822 241054
rect 275586 240498 275822 240734
rect 275586 204818 275822 205054
rect 275586 204498 275822 204734
rect 275586 168818 275822 169054
rect 275586 168498 275822 168734
rect 275586 132818 275822 133054
rect 275586 132498 275822 132734
rect 275586 96818 275822 97054
rect 275586 96498 275822 96734
rect 275586 60818 275822 61054
rect 275586 60498 275822 60734
rect 275586 24818 275822 25054
rect 275586 24498 275822 24734
rect 275586 -3402 275822 -3166
rect 275586 -3722 275822 -3486
rect 279186 316418 279422 316654
rect 279186 316098 279422 316334
rect 279186 280418 279422 280654
rect 279186 280098 279422 280334
rect 279186 244418 279422 244654
rect 279186 244098 279422 244334
rect 279186 208418 279422 208654
rect 279186 208098 279422 208334
rect 279186 172418 279422 172654
rect 279186 172098 279422 172334
rect 279186 136418 279422 136654
rect 279186 136098 279422 136334
rect 279186 100418 279422 100654
rect 279186 100098 279422 100334
rect 279186 64418 279422 64654
rect 279186 64098 279422 64334
rect 279186 28418 279422 28654
rect 279186 28098 279422 28334
rect 279186 -5282 279422 -5046
rect 279186 -5602 279422 -5366
rect 282786 320018 283022 320254
rect 282786 319698 283022 319934
rect 282786 284018 283022 284254
rect 282786 283698 283022 283934
rect 282786 248018 283022 248254
rect 282786 247698 283022 247934
rect 282786 212018 283022 212254
rect 282786 211698 283022 211934
rect 282786 176018 283022 176254
rect 282786 175698 283022 175934
rect 282786 140018 283022 140254
rect 282786 139698 283022 139934
rect 282786 104018 283022 104254
rect 282786 103698 283022 103934
rect 282786 68018 283022 68254
rect 282786 67698 283022 67934
rect 282786 32018 283022 32254
rect 282786 31698 283022 31934
rect 264786 -6222 265022 -5986
rect 264786 -6542 265022 -6306
rect 289986 327218 290222 327454
rect 289986 326898 290222 327134
rect 289986 291218 290222 291454
rect 289986 290898 290222 291134
rect 289986 255218 290222 255454
rect 289986 254898 290222 255134
rect 289986 219218 290222 219454
rect 289986 218898 290222 219134
rect 289986 183218 290222 183454
rect 289986 182898 290222 183134
rect 289986 147218 290222 147454
rect 289986 146898 290222 147134
rect 289986 111218 290222 111454
rect 289986 110898 290222 111134
rect 289986 75218 290222 75454
rect 289986 74898 290222 75134
rect 289986 39218 290222 39454
rect 289986 38898 290222 39134
rect 289986 3218 290222 3454
rect 289986 2898 290222 3134
rect 289986 -582 290222 -346
rect 289986 -902 290222 -666
rect 293586 330818 293822 331054
rect 293586 330498 293822 330734
rect 293586 294818 293822 295054
rect 293586 294498 293822 294734
rect 293586 258818 293822 259054
rect 293586 258498 293822 258734
rect 293586 222818 293822 223054
rect 293586 222498 293822 222734
rect 293586 186818 293822 187054
rect 293586 186498 293822 186734
rect 293586 150818 293822 151054
rect 293586 150498 293822 150734
rect 293586 114818 293822 115054
rect 293586 114498 293822 114734
rect 293586 78818 293822 79054
rect 293586 78498 293822 78734
rect 293586 42818 293822 43054
rect 293586 42498 293822 42734
rect 293586 6818 293822 7054
rect 293586 6498 293822 6734
rect 293586 -2462 293822 -2226
rect 293586 -2782 293822 -2546
rect 297186 334418 297422 334654
rect 297186 334098 297422 334334
rect 297186 298418 297422 298654
rect 297186 298098 297422 298334
rect 297186 262418 297422 262654
rect 297186 262098 297422 262334
rect 297186 226418 297422 226654
rect 297186 226098 297422 226334
rect 297186 190418 297422 190654
rect 297186 190098 297422 190334
rect 297186 154418 297422 154654
rect 297186 154098 297422 154334
rect 297186 118418 297422 118654
rect 297186 118098 297422 118334
rect 297186 82418 297422 82654
rect 297186 82098 297422 82334
rect 297186 46418 297422 46654
rect 297186 46098 297422 46334
rect 297186 10418 297422 10654
rect 297186 10098 297422 10334
rect 297186 -4342 297422 -4106
rect 297186 -4662 297422 -4426
rect 300786 302018 301022 302254
rect 300786 301698 301022 301934
rect 300786 266018 301022 266254
rect 300786 265698 301022 265934
rect 300786 230018 301022 230254
rect 300786 229698 301022 229934
rect 300786 194018 301022 194254
rect 300786 193698 301022 193934
rect 300786 158018 301022 158254
rect 300786 157698 301022 157934
rect 300786 122018 301022 122254
rect 300786 121698 301022 121934
rect 300786 86018 301022 86254
rect 300786 85698 301022 85934
rect 300786 50018 301022 50254
rect 300786 49698 301022 49934
rect 307986 309218 308222 309454
rect 307986 308898 308222 309134
rect 307986 273218 308222 273454
rect 307986 272898 308222 273134
rect 307986 237218 308222 237454
rect 307986 236898 308222 237134
rect 307986 201218 308222 201454
rect 307986 200898 308222 201134
rect 307986 165218 308222 165454
rect 307986 164898 308222 165134
rect 307986 129218 308222 129454
rect 307986 128898 308222 129134
rect 307986 93218 308222 93454
rect 307986 92898 308222 93134
rect 307986 57218 308222 57454
rect 307986 56898 308222 57134
rect 300786 14018 301022 14254
rect 300786 13698 301022 13934
rect 282786 -7162 283022 -6926
rect 282786 -7482 283022 -7246
rect 307986 21218 308222 21454
rect 307986 20898 308222 21134
rect 307986 -1522 308222 -1286
rect 307986 -1842 308222 -1606
rect 311586 672818 311822 673054
rect 311586 672498 311822 672734
rect 311586 636818 311822 637054
rect 311586 636498 311822 636734
rect 311586 600818 311822 601054
rect 311586 600498 311822 600734
rect 311586 564818 311822 565054
rect 311586 564498 311822 564734
rect 311586 528818 311822 529054
rect 311586 528498 311822 528734
rect 311586 492818 311822 493054
rect 311586 492498 311822 492734
rect 311586 456818 311822 457054
rect 311586 456498 311822 456734
rect 311586 420818 311822 421054
rect 311586 420498 311822 420734
rect 311586 384818 311822 385054
rect 311586 384498 311822 384734
rect 311586 348818 311822 349054
rect 311586 348498 311822 348734
rect 311586 312818 311822 313054
rect 311586 312498 311822 312734
rect 311586 276818 311822 277054
rect 311586 276498 311822 276734
rect 311586 240818 311822 241054
rect 311586 240498 311822 240734
rect 311586 204818 311822 205054
rect 311586 204498 311822 204734
rect 311586 168818 311822 169054
rect 311586 168498 311822 168734
rect 311586 132818 311822 133054
rect 311586 132498 311822 132734
rect 311586 96818 311822 97054
rect 311586 96498 311822 96734
rect 311586 60818 311822 61054
rect 311586 60498 311822 60734
rect 311586 24818 311822 25054
rect 311586 24498 311822 24734
rect 311586 -3402 311822 -3166
rect 311586 -3722 311822 -3486
rect 315186 676418 315422 676654
rect 315186 676098 315422 676334
rect 315186 640418 315422 640654
rect 315186 640098 315422 640334
rect 315186 604418 315422 604654
rect 315186 604098 315422 604334
rect 315186 568418 315422 568654
rect 315186 568098 315422 568334
rect 315186 532418 315422 532654
rect 315186 532098 315422 532334
rect 315186 496418 315422 496654
rect 315186 496098 315422 496334
rect 315186 460418 315422 460654
rect 315186 460098 315422 460334
rect 315186 424418 315422 424654
rect 315186 424098 315422 424334
rect 315186 388418 315422 388654
rect 315186 388098 315422 388334
rect 315186 352418 315422 352654
rect 315186 352098 315422 352334
rect 315186 316418 315422 316654
rect 315186 316098 315422 316334
rect 315186 280418 315422 280654
rect 315186 280098 315422 280334
rect 315186 244418 315422 244654
rect 315186 244098 315422 244334
rect 315186 208418 315422 208654
rect 315186 208098 315422 208334
rect 315186 172418 315422 172654
rect 315186 172098 315422 172334
rect 315186 136418 315422 136654
rect 315186 136098 315422 136334
rect 315186 100418 315422 100654
rect 315186 100098 315422 100334
rect 315186 64418 315422 64654
rect 315186 64098 315422 64334
rect 315186 28418 315422 28654
rect 315186 28098 315422 28334
rect 315186 -5282 315422 -5046
rect 315186 -5602 315422 -5366
rect 336786 710242 337022 710478
rect 336786 709922 337022 710158
rect 333186 708362 333422 708598
rect 333186 708042 333422 708278
rect 329586 706482 329822 706718
rect 329586 706162 329822 706398
rect 318786 680018 319022 680254
rect 318786 679698 319022 679934
rect 318786 644018 319022 644254
rect 318786 643698 319022 643934
rect 318786 608018 319022 608254
rect 318786 607698 319022 607934
rect 318786 572018 319022 572254
rect 318786 571698 319022 571934
rect 318786 536018 319022 536254
rect 318786 535698 319022 535934
rect 318786 500018 319022 500254
rect 318786 499698 319022 499934
rect 318786 464018 319022 464254
rect 318786 463698 319022 463934
rect 318786 428018 319022 428254
rect 318786 427698 319022 427934
rect 318786 392018 319022 392254
rect 318786 391698 319022 391934
rect 318786 356018 319022 356254
rect 318786 355698 319022 355934
rect 318786 320018 319022 320254
rect 318786 319698 319022 319934
rect 318786 284018 319022 284254
rect 318786 283698 319022 283934
rect 318786 248018 319022 248254
rect 318786 247698 319022 247934
rect 318786 212018 319022 212254
rect 318786 211698 319022 211934
rect 318786 176018 319022 176254
rect 318786 175698 319022 175934
rect 318786 140018 319022 140254
rect 318786 139698 319022 139934
rect 318786 104018 319022 104254
rect 318786 103698 319022 103934
rect 318786 68018 319022 68254
rect 318786 67698 319022 67934
rect 318786 32018 319022 32254
rect 318786 31698 319022 31934
rect 300786 -6222 301022 -5986
rect 300786 -6542 301022 -6306
rect 325986 704602 326222 704838
rect 325986 704282 326222 704518
rect 325986 687218 326222 687454
rect 325986 686898 326222 687134
rect 325986 651218 326222 651454
rect 325986 650898 326222 651134
rect 325986 615218 326222 615454
rect 325986 614898 326222 615134
rect 325986 579218 326222 579454
rect 325986 578898 326222 579134
rect 325986 543218 326222 543454
rect 325986 542898 326222 543134
rect 325986 507218 326222 507454
rect 325986 506898 326222 507134
rect 325986 471218 326222 471454
rect 325986 470898 326222 471134
rect 325986 435218 326222 435454
rect 325986 434898 326222 435134
rect 325986 399218 326222 399454
rect 325986 398898 326222 399134
rect 325986 363218 326222 363454
rect 325986 362898 326222 363134
rect 325986 327218 326222 327454
rect 325986 326898 326222 327134
rect 325986 291218 326222 291454
rect 325986 290898 326222 291134
rect 325986 255218 326222 255454
rect 325986 254898 326222 255134
rect 325986 219218 326222 219454
rect 325986 218898 326222 219134
rect 325986 183218 326222 183454
rect 325986 182898 326222 183134
rect 325986 147218 326222 147454
rect 325986 146898 326222 147134
rect 325986 111218 326222 111454
rect 325986 110898 326222 111134
rect 325986 75218 326222 75454
rect 325986 74898 326222 75134
rect 325986 39218 326222 39454
rect 325986 38898 326222 39134
rect 325986 3218 326222 3454
rect 325986 2898 326222 3134
rect 325986 -582 326222 -346
rect 325986 -902 326222 -666
rect 329586 690818 329822 691054
rect 329586 690498 329822 690734
rect 329586 654818 329822 655054
rect 329586 654498 329822 654734
rect 329586 618818 329822 619054
rect 329586 618498 329822 618734
rect 329586 582818 329822 583054
rect 329586 582498 329822 582734
rect 329586 546818 329822 547054
rect 329586 546498 329822 546734
rect 329586 510818 329822 511054
rect 329586 510498 329822 510734
rect 329586 474818 329822 475054
rect 329586 474498 329822 474734
rect 329586 438818 329822 439054
rect 329586 438498 329822 438734
rect 329586 402818 329822 403054
rect 329586 402498 329822 402734
rect 329586 366818 329822 367054
rect 329586 366498 329822 366734
rect 329586 330818 329822 331054
rect 329586 330498 329822 330734
rect 329586 294818 329822 295054
rect 329586 294498 329822 294734
rect 329586 258818 329822 259054
rect 329586 258498 329822 258734
rect 329586 222818 329822 223054
rect 329586 222498 329822 222734
rect 329586 186818 329822 187054
rect 329586 186498 329822 186734
rect 329586 150818 329822 151054
rect 329586 150498 329822 150734
rect 329586 114818 329822 115054
rect 329586 114498 329822 114734
rect 329586 78818 329822 79054
rect 329586 78498 329822 78734
rect 329586 42818 329822 43054
rect 329586 42498 329822 42734
rect 329586 6818 329822 7054
rect 329586 6498 329822 6734
rect 329586 -2462 329822 -2226
rect 329586 -2782 329822 -2546
rect 333186 694418 333422 694654
rect 333186 694098 333422 694334
rect 333186 658418 333422 658654
rect 333186 658098 333422 658334
rect 333186 622418 333422 622654
rect 333186 622098 333422 622334
rect 333186 586418 333422 586654
rect 333186 586098 333422 586334
rect 333186 550418 333422 550654
rect 333186 550098 333422 550334
rect 333186 514418 333422 514654
rect 333186 514098 333422 514334
rect 333186 478418 333422 478654
rect 333186 478098 333422 478334
rect 333186 442418 333422 442654
rect 333186 442098 333422 442334
rect 333186 406418 333422 406654
rect 333186 406098 333422 406334
rect 333186 370418 333422 370654
rect 333186 370098 333422 370334
rect 333186 334418 333422 334654
rect 333186 334098 333422 334334
rect 333186 298418 333422 298654
rect 333186 298098 333422 298334
rect 333186 262418 333422 262654
rect 333186 262098 333422 262334
rect 333186 226418 333422 226654
rect 333186 226098 333422 226334
rect 333186 190418 333422 190654
rect 333186 190098 333422 190334
rect 333186 154418 333422 154654
rect 333186 154098 333422 154334
rect 333186 118418 333422 118654
rect 333186 118098 333422 118334
rect 333186 82418 333422 82654
rect 333186 82098 333422 82334
rect 333186 46418 333422 46654
rect 333186 46098 333422 46334
rect 333186 10418 333422 10654
rect 333186 10098 333422 10334
rect 333186 -4342 333422 -4106
rect 333186 -4662 333422 -4426
rect 354786 711182 355022 711418
rect 354786 710862 355022 711098
rect 351186 709302 351422 709538
rect 351186 708982 351422 709218
rect 347586 707422 347822 707658
rect 347586 707102 347822 707338
rect 336786 698018 337022 698254
rect 336786 697698 337022 697934
rect 336786 662018 337022 662254
rect 336786 661698 337022 661934
rect 336786 626018 337022 626254
rect 336786 625698 337022 625934
rect 336786 590018 337022 590254
rect 336786 589698 337022 589934
rect 336786 554018 337022 554254
rect 336786 553698 337022 553934
rect 336786 518018 337022 518254
rect 336786 517698 337022 517934
rect 336786 482018 337022 482254
rect 336786 481698 337022 481934
rect 336786 446018 337022 446254
rect 336786 445698 337022 445934
rect 336786 410018 337022 410254
rect 336786 409698 337022 409934
rect 336786 374018 337022 374254
rect 336786 373698 337022 373934
rect 336786 338018 337022 338254
rect 336786 337698 337022 337934
rect 336786 302018 337022 302254
rect 336786 301698 337022 301934
rect 336786 266018 337022 266254
rect 336786 265698 337022 265934
rect 336786 230018 337022 230254
rect 336786 229698 337022 229934
rect 336786 194018 337022 194254
rect 336786 193698 337022 193934
rect 336786 158018 337022 158254
rect 336786 157698 337022 157934
rect 336786 122018 337022 122254
rect 336786 121698 337022 121934
rect 336786 86018 337022 86254
rect 336786 85698 337022 85934
rect 336786 50018 337022 50254
rect 336786 49698 337022 49934
rect 336786 14018 337022 14254
rect 336786 13698 337022 13934
rect 318786 -7162 319022 -6926
rect 318786 -7482 319022 -7246
rect 343986 705542 344222 705778
rect 343986 705222 344222 705458
rect 343986 669218 344222 669454
rect 343986 668898 344222 669134
rect 343986 633218 344222 633454
rect 343986 632898 344222 633134
rect 343986 597218 344222 597454
rect 343986 596898 344222 597134
rect 343986 561218 344222 561454
rect 343986 560898 344222 561134
rect 343986 525218 344222 525454
rect 343986 524898 344222 525134
rect 343986 489218 344222 489454
rect 343986 488898 344222 489134
rect 343986 453218 344222 453454
rect 343986 452898 344222 453134
rect 343986 417218 344222 417454
rect 343986 416898 344222 417134
rect 343986 381218 344222 381454
rect 343986 380898 344222 381134
rect 343986 345218 344222 345454
rect 343986 344898 344222 345134
rect 343986 309218 344222 309454
rect 343986 308898 344222 309134
rect 343986 273218 344222 273454
rect 343986 272898 344222 273134
rect 343986 237218 344222 237454
rect 343986 236898 344222 237134
rect 343986 201218 344222 201454
rect 343986 200898 344222 201134
rect 343986 165218 344222 165454
rect 343986 164898 344222 165134
rect 343986 129218 344222 129454
rect 343986 128898 344222 129134
rect 343986 93218 344222 93454
rect 343986 92898 344222 93134
rect 343986 57218 344222 57454
rect 343986 56898 344222 57134
rect 343986 21218 344222 21454
rect 343986 20898 344222 21134
rect 343986 -1522 344222 -1286
rect 343986 -1842 344222 -1606
rect 347586 672818 347822 673054
rect 347586 672498 347822 672734
rect 347586 636818 347822 637054
rect 347586 636498 347822 636734
rect 347586 600818 347822 601054
rect 347586 600498 347822 600734
rect 347586 564818 347822 565054
rect 347586 564498 347822 564734
rect 347586 528818 347822 529054
rect 347586 528498 347822 528734
rect 347586 492818 347822 493054
rect 347586 492498 347822 492734
rect 347586 456818 347822 457054
rect 347586 456498 347822 456734
rect 347586 420818 347822 421054
rect 347586 420498 347822 420734
rect 347586 384818 347822 385054
rect 347586 384498 347822 384734
rect 347586 348818 347822 349054
rect 347586 348498 347822 348734
rect 347586 312818 347822 313054
rect 347586 312498 347822 312734
rect 347586 276818 347822 277054
rect 347586 276498 347822 276734
rect 347586 240818 347822 241054
rect 347586 240498 347822 240734
rect 347586 204818 347822 205054
rect 347586 204498 347822 204734
rect 347586 168818 347822 169054
rect 347586 168498 347822 168734
rect 347586 132818 347822 133054
rect 347586 132498 347822 132734
rect 347586 96818 347822 97054
rect 347586 96498 347822 96734
rect 347586 60818 347822 61054
rect 347586 60498 347822 60734
rect 347586 24818 347822 25054
rect 347586 24498 347822 24734
rect 347586 -3402 347822 -3166
rect 347586 -3722 347822 -3486
rect 351186 676418 351422 676654
rect 351186 676098 351422 676334
rect 351186 640418 351422 640654
rect 351186 640098 351422 640334
rect 351186 604418 351422 604654
rect 351186 604098 351422 604334
rect 351186 568418 351422 568654
rect 351186 568098 351422 568334
rect 351186 532418 351422 532654
rect 351186 532098 351422 532334
rect 351186 496418 351422 496654
rect 351186 496098 351422 496334
rect 351186 460418 351422 460654
rect 351186 460098 351422 460334
rect 351186 424418 351422 424654
rect 351186 424098 351422 424334
rect 351186 388418 351422 388654
rect 351186 388098 351422 388334
rect 351186 352418 351422 352654
rect 351186 352098 351422 352334
rect 351186 316418 351422 316654
rect 351186 316098 351422 316334
rect 351186 280418 351422 280654
rect 351186 280098 351422 280334
rect 351186 244418 351422 244654
rect 351186 244098 351422 244334
rect 351186 208418 351422 208654
rect 351186 208098 351422 208334
rect 351186 172418 351422 172654
rect 351186 172098 351422 172334
rect 351186 136418 351422 136654
rect 351186 136098 351422 136334
rect 351186 100418 351422 100654
rect 351186 100098 351422 100334
rect 351186 64418 351422 64654
rect 351186 64098 351422 64334
rect 351186 28418 351422 28654
rect 351186 28098 351422 28334
rect 351186 -5282 351422 -5046
rect 351186 -5602 351422 -5366
rect 372786 710242 373022 710478
rect 372786 709922 373022 710158
rect 369186 708362 369422 708598
rect 369186 708042 369422 708278
rect 365586 706482 365822 706718
rect 365586 706162 365822 706398
rect 354786 680018 355022 680254
rect 354786 679698 355022 679934
rect 354786 644018 355022 644254
rect 354786 643698 355022 643934
rect 354786 608018 355022 608254
rect 354786 607698 355022 607934
rect 354786 572018 355022 572254
rect 354786 571698 355022 571934
rect 354786 536018 355022 536254
rect 354786 535698 355022 535934
rect 354786 500018 355022 500254
rect 354786 499698 355022 499934
rect 354786 464018 355022 464254
rect 354786 463698 355022 463934
rect 354786 428018 355022 428254
rect 354786 427698 355022 427934
rect 354786 392018 355022 392254
rect 354786 391698 355022 391934
rect 354786 356018 355022 356254
rect 354786 355698 355022 355934
rect 354786 320018 355022 320254
rect 354786 319698 355022 319934
rect 354786 284018 355022 284254
rect 354786 283698 355022 283934
rect 354786 248018 355022 248254
rect 354786 247698 355022 247934
rect 354786 212018 355022 212254
rect 354786 211698 355022 211934
rect 354786 176018 355022 176254
rect 354786 175698 355022 175934
rect 354786 140018 355022 140254
rect 354786 139698 355022 139934
rect 354786 104018 355022 104254
rect 354786 103698 355022 103934
rect 354786 68018 355022 68254
rect 354786 67698 355022 67934
rect 354786 32018 355022 32254
rect 354786 31698 355022 31934
rect 336786 -6222 337022 -5986
rect 336786 -6542 337022 -6306
rect 361986 704602 362222 704838
rect 361986 704282 362222 704518
rect 361986 687218 362222 687454
rect 361986 686898 362222 687134
rect 361986 651218 362222 651454
rect 361986 650898 362222 651134
rect 361986 615218 362222 615454
rect 361986 614898 362222 615134
rect 361986 579218 362222 579454
rect 361986 578898 362222 579134
rect 361986 543218 362222 543454
rect 361986 542898 362222 543134
rect 361986 507218 362222 507454
rect 361986 506898 362222 507134
rect 361986 471218 362222 471454
rect 361986 470898 362222 471134
rect 361986 435218 362222 435454
rect 361986 434898 362222 435134
rect 361986 399218 362222 399454
rect 361986 398898 362222 399134
rect 361986 363218 362222 363454
rect 361986 362898 362222 363134
rect 361986 327218 362222 327454
rect 361986 326898 362222 327134
rect 361986 291218 362222 291454
rect 361986 290898 362222 291134
rect 361986 255218 362222 255454
rect 361986 254898 362222 255134
rect 361986 219218 362222 219454
rect 361986 218898 362222 219134
rect 361986 183218 362222 183454
rect 361986 182898 362222 183134
rect 361986 147218 362222 147454
rect 361986 146898 362222 147134
rect 361986 111218 362222 111454
rect 361986 110898 362222 111134
rect 361986 75218 362222 75454
rect 361986 74898 362222 75134
rect 361986 39218 362222 39454
rect 361986 38898 362222 39134
rect 361986 3218 362222 3454
rect 361986 2898 362222 3134
rect 361986 -582 362222 -346
rect 361986 -902 362222 -666
rect 365586 690818 365822 691054
rect 365586 690498 365822 690734
rect 365586 654818 365822 655054
rect 365586 654498 365822 654734
rect 365586 618818 365822 619054
rect 365586 618498 365822 618734
rect 365586 582818 365822 583054
rect 365586 582498 365822 582734
rect 365586 546818 365822 547054
rect 365586 546498 365822 546734
rect 365586 510818 365822 511054
rect 365586 510498 365822 510734
rect 365586 474818 365822 475054
rect 365586 474498 365822 474734
rect 365586 438818 365822 439054
rect 365586 438498 365822 438734
rect 365586 402818 365822 403054
rect 365586 402498 365822 402734
rect 365586 366818 365822 367054
rect 365586 366498 365822 366734
rect 365586 330818 365822 331054
rect 365586 330498 365822 330734
rect 365586 294818 365822 295054
rect 365586 294498 365822 294734
rect 365586 258818 365822 259054
rect 365586 258498 365822 258734
rect 365586 222818 365822 223054
rect 365586 222498 365822 222734
rect 365586 186818 365822 187054
rect 365586 186498 365822 186734
rect 365586 150818 365822 151054
rect 365586 150498 365822 150734
rect 365586 114818 365822 115054
rect 365586 114498 365822 114734
rect 365586 78818 365822 79054
rect 365586 78498 365822 78734
rect 365586 42818 365822 43054
rect 365586 42498 365822 42734
rect 365586 6818 365822 7054
rect 365586 6498 365822 6734
rect 365586 -2462 365822 -2226
rect 365586 -2782 365822 -2546
rect 369186 694418 369422 694654
rect 369186 694098 369422 694334
rect 369186 658418 369422 658654
rect 369186 658098 369422 658334
rect 369186 622418 369422 622654
rect 369186 622098 369422 622334
rect 369186 586418 369422 586654
rect 369186 586098 369422 586334
rect 369186 550418 369422 550654
rect 369186 550098 369422 550334
rect 369186 514418 369422 514654
rect 369186 514098 369422 514334
rect 369186 478418 369422 478654
rect 369186 478098 369422 478334
rect 369186 442418 369422 442654
rect 369186 442098 369422 442334
rect 369186 406418 369422 406654
rect 369186 406098 369422 406334
rect 369186 370418 369422 370654
rect 369186 370098 369422 370334
rect 369186 334418 369422 334654
rect 369186 334098 369422 334334
rect 369186 298418 369422 298654
rect 369186 298098 369422 298334
rect 369186 262418 369422 262654
rect 369186 262098 369422 262334
rect 369186 226418 369422 226654
rect 369186 226098 369422 226334
rect 369186 190418 369422 190654
rect 369186 190098 369422 190334
rect 369186 154418 369422 154654
rect 369186 154098 369422 154334
rect 369186 118418 369422 118654
rect 369186 118098 369422 118334
rect 369186 82418 369422 82654
rect 369186 82098 369422 82334
rect 369186 46418 369422 46654
rect 369186 46098 369422 46334
rect 369186 10418 369422 10654
rect 369186 10098 369422 10334
rect 369186 -4342 369422 -4106
rect 369186 -4662 369422 -4426
rect 390786 711182 391022 711418
rect 390786 710862 391022 711098
rect 387186 709302 387422 709538
rect 387186 708982 387422 709218
rect 383586 707422 383822 707658
rect 383586 707102 383822 707338
rect 372786 698018 373022 698254
rect 372786 697698 373022 697934
rect 372786 662018 373022 662254
rect 372786 661698 373022 661934
rect 372786 626018 373022 626254
rect 372786 625698 373022 625934
rect 372786 590018 373022 590254
rect 372786 589698 373022 589934
rect 372786 554018 373022 554254
rect 372786 553698 373022 553934
rect 372786 518018 373022 518254
rect 372786 517698 373022 517934
rect 372786 482018 373022 482254
rect 372786 481698 373022 481934
rect 372786 446018 373022 446254
rect 372786 445698 373022 445934
rect 372786 410018 373022 410254
rect 372786 409698 373022 409934
rect 372786 374018 373022 374254
rect 372786 373698 373022 373934
rect 372786 338018 373022 338254
rect 372786 337698 373022 337934
rect 372786 302018 373022 302254
rect 372786 301698 373022 301934
rect 372786 266018 373022 266254
rect 372786 265698 373022 265934
rect 372786 230018 373022 230254
rect 372786 229698 373022 229934
rect 372786 194018 373022 194254
rect 372786 193698 373022 193934
rect 372786 158018 373022 158254
rect 372786 157698 373022 157934
rect 372786 122018 373022 122254
rect 372786 121698 373022 121934
rect 372786 86018 373022 86254
rect 372786 85698 373022 85934
rect 372786 50018 373022 50254
rect 372786 49698 373022 49934
rect 372786 14018 373022 14254
rect 372786 13698 373022 13934
rect 354786 -7162 355022 -6926
rect 354786 -7482 355022 -7246
rect 379986 705542 380222 705778
rect 379986 705222 380222 705458
rect 379986 669218 380222 669454
rect 379986 668898 380222 669134
rect 379986 633218 380222 633454
rect 379986 632898 380222 633134
rect 379986 597218 380222 597454
rect 379986 596898 380222 597134
rect 379986 561218 380222 561454
rect 379986 560898 380222 561134
rect 379986 525218 380222 525454
rect 379986 524898 380222 525134
rect 379986 489218 380222 489454
rect 379986 488898 380222 489134
rect 379986 453218 380222 453454
rect 379986 452898 380222 453134
rect 379986 417218 380222 417454
rect 379986 416898 380222 417134
rect 379986 381218 380222 381454
rect 379986 380898 380222 381134
rect 379986 345218 380222 345454
rect 379986 344898 380222 345134
rect 379986 309218 380222 309454
rect 379986 308898 380222 309134
rect 379986 273218 380222 273454
rect 379986 272898 380222 273134
rect 379986 237218 380222 237454
rect 379986 236898 380222 237134
rect 379986 201218 380222 201454
rect 379986 200898 380222 201134
rect 379986 165218 380222 165454
rect 379986 164898 380222 165134
rect 379986 129218 380222 129454
rect 379986 128898 380222 129134
rect 379986 93218 380222 93454
rect 379986 92898 380222 93134
rect 379986 57218 380222 57454
rect 379986 56898 380222 57134
rect 379986 21218 380222 21454
rect 379986 20898 380222 21134
rect 379986 -1522 380222 -1286
rect 379986 -1842 380222 -1606
rect 383586 672818 383822 673054
rect 383586 672498 383822 672734
rect 383586 636818 383822 637054
rect 383586 636498 383822 636734
rect 383586 600818 383822 601054
rect 383586 600498 383822 600734
rect 383586 564818 383822 565054
rect 383586 564498 383822 564734
rect 383586 528818 383822 529054
rect 383586 528498 383822 528734
rect 383586 492818 383822 493054
rect 383586 492498 383822 492734
rect 383586 456818 383822 457054
rect 383586 456498 383822 456734
rect 383586 420818 383822 421054
rect 383586 420498 383822 420734
rect 383586 384818 383822 385054
rect 383586 384498 383822 384734
rect 383586 348818 383822 349054
rect 383586 348498 383822 348734
rect 383586 312818 383822 313054
rect 383586 312498 383822 312734
rect 383586 276818 383822 277054
rect 383586 276498 383822 276734
rect 383586 240818 383822 241054
rect 383586 240498 383822 240734
rect 383586 204818 383822 205054
rect 383586 204498 383822 204734
rect 383586 168818 383822 169054
rect 383586 168498 383822 168734
rect 383586 132818 383822 133054
rect 383586 132498 383822 132734
rect 383586 96818 383822 97054
rect 383586 96498 383822 96734
rect 383586 60818 383822 61054
rect 383586 60498 383822 60734
rect 383586 24818 383822 25054
rect 383586 24498 383822 24734
rect 383586 -3402 383822 -3166
rect 383586 -3722 383822 -3486
rect 387186 676418 387422 676654
rect 387186 676098 387422 676334
rect 387186 640418 387422 640654
rect 387186 640098 387422 640334
rect 387186 604418 387422 604654
rect 387186 604098 387422 604334
rect 387186 568418 387422 568654
rect 387186 568098 387422 568334
rect 387186 532418 387422 532654
rect 387186 532098 387422 532334
rect 387186 496418 387422 496654
rect 387186 496098 387422 496334
rect 387186 460418 387422 460654
rect 387186 460098 387422 460334
rect 387186 424418 387422 424654
rect 387186 424098 387422 424334
rect 387186 388418 387422 388654
rect 387186 388098 387422 388334
rect 387186 352418 387422 352654
rect 387186 352098 387422 352334
rect 387186 316418 387422 316654
rect 387186 316098 387422 316334
rect 387186 280418 387422 280654
rect 387186 280098 387422 280334
rect 387186 244418 387422 244654
rect 387186 244098 387422 244334
rect 387186 208418 387422 208654
rect 387186 208098 387422 208334
rect 387186 172418 387422 172654
rect 387186 172098 387422 172334
rect 387186 136418 387422 136654
rect 387186 136098 387422 136334
rect 387186 100418 387422 100654
rect 387186 100098 387422 100334
rect 387186 64418 387422 64654
rect 387186 64098 387422 64334
rect 387186 28418 387422 28654
rect 387186 28098 387422 28334
rect 387186 -5282 387422 -5046
rect 387186 -5602 387422 -5366
rect 408786 710242 409022 710478
rect 408786 709922 409022 710158
rect 405186 708362 405422 708598
rect 405186 708042 405422 708278
rect 401586 706482 401822 706718
rect 401586 706162 401822 706398
rect 390786 680018 391022 680254
rect 390786 679698 391022 679934
rect 390786 644018 391022 644254
rect 390786 643698 391022 643934
rect 390786 608018 391022 608254
rect 390786 607698 391022 607934
rect 390786 572018 391022 572254
rect 390786 571698 391022 571934
rect 390786 536018 391022 536254
rect 390786 535698 391022 535934
rect 390786 500018 391022 500254
rect 390786 499698 391022 499934
rect 390786 464018 391022 464254
rect 390786 463698 391022 463934
rect 390786 428018 391022 428254
rect 390786 427698 391022 427934
rect 390786 392018 391022 392254
rect 390786 391698 391022 391934
rect 390786 356018 391022 356254
rect 390786 355698 391022 355934
rect 390786 320018 391022 320254
rect 390786 319698 391022 319934
rect 390786 284018 391022 284254
rect 390786 283698 391022 283934
rect 390786 248018 391022 248254
rect 390786 247698 391022 247934
rect 390786 212018 391022 212254
rect 390786 211698 391022 211934
rect 390786 176018 391022 176254
rect 390786 175698 391022 175934
rect 390786 140018 391022 140254
rect 390786 139698 391022 139934
rect 390786 104018 391022 104254
rect 390786 103698 391022 103934
rect 390786 68018 391022 68254
rect 390786 67698 391022 67934
rect 390786 32018 391022 32254
rect 390786 31698 391022 31934
rect 372786 -6222 373022 -5986
rect 372786 -6542 373022 -6306
rect 397986 704602 398222 704838
rect 397986 704282 398222 704518
rect 397986 687218 398222 687454
rect 397986 686898 398222 687134
rect 397986 651218 398222 651454
rect 397986 650898 398222 651134
rect 397986 615218 398222 615454
rect 397986 614898 398222 615134
rect 397986 579218 398222 579454
rect 397986 578898 398222 579134
rect 397986 543218 398222 543454
rect 397986 542898 398222 543134
rect 397986 507218 398222 507454
rect 397986 506898 398222 507134
rect 397986 471218 398222 471454
rect 397986 470898 398222 471134
rect 397986 435218 398222 435454
rect 397986 434898 398222 435134
rect 397986 399218 398222 399454
rect 397986 398898 398222 399134
rect 397986 363218 398222 363454
rect 397986 362898 398222 363134
rect 397986 327218 398222 327454
rect 397986 326898 398222 327134
rect 397986 291218 398222 291454
rect 397986 290898 398222 291134
rect 397986 255218 398222 255454
rect 397986 254898 398222 255134
rect 397986 219218 398222 219454
rect 397986 218898 398222 219134
rect 397986 183218 398222 183454
rect 397986 182898 398222 183134
rect 397986 147218 398222 147454
rect 397986 146898 398222 147134
rect 397986 111218 398222 111454
rect 397986 110898 398222 111134
rect 397986 75218 398222 75454
rect 397986 74898 398222 75134
rect 397986 39218 398222 39454
rect 397986 38898 398222 39134
rect 397986 3218 398222 3454
rect 397986 2898 398222 3134
rect 397986 -582 398222 -346
rect 397986 -902 398222 -666
rect 401586 690818 401822 691054
rect 401586 690498 401822 690734
rect 401586 654818 401822 655054
rect 401586 654498 401822 654734
rect 401586 618818 401822 619054
rect 401586 618498 401822 618734
rect 401586 582818 401822 583054
rect 401586 582498 401822 582734
rect 401586 546818 401822 547054
rect 401586 546498 401822 546734
rect 401586 510818 401822 511054
rect 401586 510498 401822 510734
rect 401586 474818 401822 475054
rect 401586 474498 401822 474734
rect 401586 438818 401822 439054
rect 401586 438498 401822 438734
rect 401586 402818 401822 403054
rect 401586 402498 401822 402734
rect 401586 366818 401822 367054
rect 401586 366498 401822 366734
rect 401586 330818 401822 331054
rect 401586 330498 401822 330734
rect 401586 294818 401822 295054
rect 401586 294498 401822 294734
rect 401586 258818 401822 259054
rect 401586 258498 401822 258734
rect 401586 222818 401822 223054
rect 401586 222498 401822 222734
rect 401586 186818 401822 187054
rect 401586 186498 401822 186734
rect 401586 150818 401822 151054
rect 401586 150498 401822 150734
rect 401586 114818 401822 115054
rect 401586 114498 401822 114734
rect 401586 78818 401822 79054
rect 401586 78498 401822 78734
rect 401586 42818 401822 43054
rect 401586 42498 401822 42734
rect 401586 6818 401822 7054
rect 401586 6498 401822 6734
rect 401586 -2462 401822 -2226
rect 401586 -2782 401822 -2546
rect 405186 694418 405422 694654
rect 405186 694098 405422 694334
rect 405186 658418 405422 658654
rect 405186 658098 405422 658334
rect 405186 622418 405422 622654
rect 405186 622098 405422 622334
rect 405186 586418 405422 586654
rect 405186 586098 405422 586334
rect 405186 550418 405422 550654
rect 405186 550098 405422 550334
rect 405186 514418 405422 514654
rect 405186 514098 405422 514334
rect 405186 478418 405422 478654
rect 405186 478098 405422 478334
rect 405186 442418 405422 442654
rect 405186 442098 405422 442334
rect 405186 406418 405422 406654
rect 405186 406098 405422 406334
rect 405186 370418 405422 370654
rect 405186 370098 405422 370334
rect 405186 334418 405422 334654
rect 405186 334098 405422 334334
rect 405186 298418 405422 298654
rect 405186 298098 405422 298334
rect 405186 262418 405422 262654
rect 405186 262098 405422 262334
rect 405186 226418 405422 226654
rect 405186 226098 405422 226334
rect 405186 190418 405422 190654
rect 405186 190098 405422 190334
rect 405186 154418 405422 154654
rect 405186 154098 405422 154334
rect 405186 118418 405422 118654
rect 405186 118098 405422 118334
rect 405186 82418 405422 82654
rect 405186 82098 405422 82334
rect 405186 46418 405422 46654
rect 405186 46098 405422 46334
rect 405186 10418 405422 10654
rect 405186 10098 405422 10334
rect 405186 -4342 405422 -4106
rect 405186 -4662 405422 -4426
rect 426786 711182 427022 711418
rect 426786 710862 427022 711098
rect 423186 709302 423422 709538
rect 423186 708982 423422 709218
rect 419586 707422 419822 707658
rect 419586 707102 419822 707338
rect 408786 698018 409022 698254
rect 408786 697698 409022 697934
rect 408786 662018 409022 662254
rect 408786 661698 409022 661934
rect 408786 626018 409022 626254
rect 408786 625698 409022 625934
rect 408786 590018 409022 590254
rect 408786 589698 409022 589934
rect 408786 554018 409022 554254
rect 408786 553698 409022 553934
rect 408786 518018 409022 518254
rect 408786 517698 409022 517934
rect 408786 482018 409022 482254
rect 408786 481698 409022 481934
rect 408786 446018 409022 446254
rect 408786 445698 409022 445934
rect 408786 410018 409022 410254
rect 408786 409698 409022 409934
rect 408786 374018 409022 374254
rect 408786 373698 409022 373934
rect 408786 338018 409022 338254
rect 408786 337698 409022 337934
rect 408786 302018 409022 302254
rect 408786 301698 409022 301934
rect 408786 266018 409022 266254
rect 408786 265698 409022 265934
rect 408786 230018 409022 230254
rect 408786 229698 409022 229934
rect 408786 194018 409022 194254
rect 408786 193698 409022 193934
rect 408786 158018 409022 158254
rect 408786 157698 409022 157934
rect 408786 122018 409022 122254
rect 408786 121698 409022 121934
rect 408786 86018 409022 86254
rect 408786 85698 409022 85934
rect 408786 50018 409022 50254
rect 408786 49698 409022 49934
rect 408786 14018 409022 14254
rect 408786 13698 409022 13934
rect 390786 -7162 391022 -6926
rect 390786 -7482 391022 -7246
rect 415986 705542 416222 705778
rect 415986 705222 416222 705458
rect 415986 669218 416222 669454
rect 415986 668898 416222 669134
rect 415986 633218 416222 633454
rect 415986 632898 416222 633134
rect 415986 597218 416222 597454
rect 415986 596898 416222 597134
rect 415986 561218 416222 561454
rect 415986 560898 416222 561134
rect 415986 525218 416222 525454
rect 415986 524898 416222 525134
rect 415986 489218 416222 489454
rect 415986 488898 416222 489134
rect 415986 453218 416222 453454
rect 415986 452898 416222 453134
rect 415986 417218 416222 417454
rect 415986 416898 416222 417134
rect 415986 381218 416222 381454
rect 415986 380898 416222 381134
rect 415986 345218 416222 345454
rect 415986 344898 416222 345134
rect 415986 309218 416222 309454
rect 415986 308898 416222 309134
rect 415986 273218 416222 273454
rect 415986 272898 416222 273134
rect 415986 237218 416222 237454
rect 415986 236898 416222 237134
rect 415986 201218 416222 201454
rect 415986 200898 416222 201134
rect 415986 165218 416222 165454
rect 415986 164898 416222 165134
rect 415986 129218 416222 129454
rect 415986 128898 416222 129134
rect 415986 93218 416222 93454
rect 415986 92898 416222 93134
rect 415986 57218 416222 57454
rect 415986 56898 416222 57134
rect 415986 21218 416222 21454
rect 415986 20898 416222 21134
rect 415986 -1522 416222 -1286
rect 415986 -1842 416222 -1606
rect 419586 672818 419822 673054
rect 419586 672498 419822 672734
rect 419586 636818 419822 637054
rect 419586 636498 419822 636734
rect 419586 600818 419822 601054
rect 419586 600498 419822 600734
rect 419586 564818 419822 565054
rect 419586 564498 419822 564734
rect 419586 528818 419822 529054
rect 419586 528498 419822 528734
rect 419586 492818 419822 493054
rect 419586 492498 419822 492734
rect 419586 456818 419822 457054
rect 419586 456498 419822 456734
rect 419586 420818 419822 421054
rect 419586 420498 419822 420734
rect 419586 384818 419822 385054
rect 419586 384498 419822 384734
rect 419586 348818 419822 349054
rect 419586 348498 419822 348734
rect 419586 312818 419822 313054
rect 419586 312498 419822 312734
rect 419586 276818 419822 277054
rect 419586 276498 419822 276734
rect 419586 240818 419822 241054
rect 419586 240498 419822 240734
rect 419586 204818 419822 205054
rect 419586 204498 419822 204734
rect 419586 168818 419822 169054
rect 419586 168498 419822 168734
rect 419586 132818 419822 133054
rect 419586 132498 419822 132734
rect 419586 96818 419822 97054
rect 419586 96498 419822 96734
rect 419586 60818 419822 61054
rect 419586 60498 419822 60734
rect 419586 24818 419822 25054
rect 419586 24498 419822 24734
rect 419586 -3402 419822 -3166
rect 419586 -3722 419822 -3486
rect 423186 676418 423422 676654
rect 423186 676098 423422 676334
rect 423186 640418 423422 640654
rect 423186 640098 423422 640334
rect 423186 604418 423422 604654
rect 423186 604098 423422 604334
rect 423186 568418 423422 568654
rect 423186 568098 423422 568334
rect 423186 532418 423422 532654
rect 423186 532098 423422 532334
rect 423186 496418 423422 496654
rect 423186 496098 423422 496334
rect 423186 460418 423422 460654
rect 423186 460098 423422 460334
rect 423186 424418 423422 424654
rect 423186 424098 423422 424334
rect 423186 388418 423422 388654
rect 423186 388098 423422 388334
rect 423186 352418 423422 352654
rect 423186 352098 423422 352334
rect 423186 316418 423422 316654
rect 423186 316098 423422 316334
rect 423186 280418 423422 280654
rect 423186 280098 423422 280334
rect 423186 244418 423422 244654
rect 423186 244098 423422 244334
rect 423186 208418 423422 208654
rect 423186 208098 423422 208334
rect 423186 172418 423422 172654
rect 423186 172098 423422 172334
rect 423186 136418 423422 136654
rect 423186 136098 423422 136334
rect 423186 100418 423422 100654
rect 423186 100098 423422 100334
rect 423186 64418 423422 64654
rect 423186 64098 423422 64334
rect 423186 28418 423422 28654
rect 423186 28098 423422 28334
rect 423186 -5282 423422 -5046
rect 423186 -5602 423422 -5366
rect 444786 710242 445022 710478
rect 444786 709922 445022 710158
rect 441186 708362 441422 708598
rect 441186 708042 441422 708278
rect 437586 706482 437822 706718
rect 437586 706162 437822 706398
rect 426786 680018 427022 680254
rect 426786 679698 427022 679934
rect 426786 644018 427022 644254
rect 426786 643698 427022 643934
rect 426786 608018 427022 608254
rect 426786 607698 427022 607934
rect 426786 572018 427022 572254
rect 426786 571698 427022 571934
rect 426786 536018 427022 536254
rect 426786 535698 427022 535934
rect 426786 500018 427022 500254
rect 426786 499698 427022 499934
rect 426786 464018 427022 464254
rect 426786 463698 427022 463934
rect 426786 428018 427022 428254
rect 426786 427698 427022 427934
rect 426786 392018 427022 392254
rect 426786 391698 427022 391934
rect 426786 356018 427022 356254
rect 426786 355698 427022 355934
rect 426786 320018 427022 320254
rect 426786 319698 427022 319934
rect 426786 284018 427022 284254
rect 426786 283698 427022 283934
rect 426786 248018 427022 248254
rect 426786 247698 427022 247934
rect 426786 212018 427022 212254
rect 426786 211698 427022 211934
rect 426786 176018 427022 176254
rect 426786 175698 427022 175934
rect 426786 140018 427022 140254
rect 426786 139698 427022 139934
rect 426786 104018 427022 104254
rect 426786 103698 427022 103934
rect 426786 68018 427022 68254
rect 426786 67698 427022 67934
rect 426786 32018 427022 32254
rect 426786 31698 427022 31934
rect 408786 -6222 409022 -5986
rect 408786 -6542 409022 -6306
rect 433986 704602 434222 704838
rect 433986 704282 434222 704518
rect 433986 687218 434222 687454
rect 433986 686898 434222 687134
rect 433986 651218 434222 651454
rect 433986 650898 434222 651134
rect 433986 615218 434222 615454
rect 433986 614898 434222 615134
rect 433986 579218 434222 579454
rect 433986 578898 434222 579134
rect 433986 543218 434222 543454
rect 433986 542898 434222 543134
rect 433986 507218 434222 507454
rect 433986 506898 434222 507134
rect 433986 471218 434222 471454
rect 433986 470898 434222 471134
rect 433986 435218 434222 435454
rect 433986 434898 434222 435134
rect 433986 399218 434222 399454
rect 433986 398898 434222 399134
rect 433986 363218 434222 363454
rect 433986 362898 434222 363134
rect 433986 327218 434222 327454
rect 433986 326898 434222 327134
rect 433986 291218 434222 291454
rect 433986 290898 434222 291134
rect 433986 255218 434222 255454
rect 433986 254898 434222 255134
rect 433986 219218 434222 219454
rect 433986 218898 434222 219134
rect 433986 183218 434222 183454
rect 433986 182898 434222 183134
rect 433986 147218 434222 147454
rect 433986 146898 434222 147134
rect 433986 111218 434222 111454
rect 433986 110898 434222 111134
rect 433986 75218 434222 75454
rect 433986 74898 434222 75134
rect 433986 39218 434222 39454
rect 433986 38898 434222 39134
rect 433986 3218 434222 3454
rect 433986 2898 434222 3134
rect 433986 -582 434222 -346
rect 433986 -902 434222 -666
rect 437586 690818 437822 691054
rect 437586 690498 437822 690734
rect 437586 654818 437822 655054
rect 437586 654498 437822 654734
rect 437586 618818 437822 619054
rect 437586 618498 437822 618734
rect 437586 582818 437822 583054
rect 437586 582498 437822 582734
rect 437586 546818 437822 547054
rect 437586 546498 437822 546734
rect 437586 510818 437822 511054
rect 437586 510498 437822 510734
rect 437586 474818 437822 475054
rect 437586 474498 437822 474734
rect 437586 438818 437822 439054
rect 437586 438498 437822 438734
rect 437586 402818 437822 403054
rect 437586 402498 437822 402734
rect 437586 366818 437822 367054
rect 437586 366498 437822 366734
rect 437586 330818 437822 331054
rect 437586 330498 437822 330734
rect 437586 294818 437822 295054
rect 437586 294498 437822 294734
rect 437586 258818 437822 259054
rect 437586 258498 437822 258734
rect 437586 222818 437822 223054
rect 437586 222498 437822 222734
rect 437586 186818 437822 187054
rect 437586 186498 437822 186734
rect 437586 150818 437822 151054
rect 437586 150498 437822 150734
rect 437586 114818 437822 115054
rect 437586 114498 437822 114734
rect 437586 78818 437822 79054
rect 437586 78498 437822 78734
rect 437586 42818 437822 43054
rect 437586 42498 437822 42734
rect 437586 6818 437822 7054
rect 437586 6498 437822 6734
rect 437586 -2462 437822 -2226
rect 437586 -2782 437822 -2546
rect 441186 694418 441422 694654
rect 441186 694098 441422 694334
rect 441186 658418 441422 658654
rect 441186 658098 441422 658334
rect 441186 622418 441422 622654
rect 441186 622098 441422 622334
rect 441186 586418 441422 586654
rect 441186 586098 441422 586334
rect 441186 550418 441422 550654
rect 441186 550098 441422 550334
rect 441186 514418 441422 514654
rect 441186 514098 441422 514334
rect 441186 478418 441422 478654
rect 441186 478098 441422 478334
rect 441186 442418 441422 442654
rect 441186 442098 441422 442334
rect 441186 406418 441422 406654
rect 441186 406098 441422 406334
rect 441186 370418 441422 370654
rect 441186 370098 441422 370334
rect 441186 334418 441422 334654
rect 441186 334098 441422 334334
rect 441186 298418 441422 298654
rect 441186 298098 441422 298334
rect 441186 262418 441422 262654
rect 441186 262098 441422 262334
rect 441186 226418 441422 226654
rect 441186 226098 441422 226334
rect 441186 190418 441422 190654
rect 441186 190098 441422 190334
rect 441186 154418 441422 154654
rect 441186 154098 441422 154334
rect 441186 118418 441422 118654
rect 441186 118098 441422 118334
rect 441186 82418 441422 82654
rect 441186 82098 441422 82334
rect 441186 46418 441422 46654
rect 441186 46098 441422 46334
rect 441186 10418 441422 10654
rect 441186 10098 441422 10334
rect 441186 -4342 441422 -4106
rect 441186 -4662 441422 -4426
rect 462786 711182 463022 711418
rect 462786 710862 463022 711098
rect 459186 709302 459422 709538
rect 459186 708982 459422 709218
rect 455586 707422 455822 707658
rect 455586 707102 455822 707338
rect 444786 698018 445022 698254
rect 444786 697698 445022 697934
rect 444786 662018 445022 662254
rect 444786 661698 445022 661934
rect 444786 626018 445022 626254
rect 444786 625698 445022 625934
rect 444786 590018 445022 590254
rect 444786 589698 445022 589934
rect 444786 554018 445022 554254
rect 444786 553698 445022 553934
rect 444786 518018 445022 518254
rect 444786 517698 445022 517934
rect 444786 482018 445022 482254
rect 444786 481698 445022 481934
rect 444786 446018 445022 446254
rect 444786 445698 445022 445934
rect 444786 410018 445022 410254
rect 444786 409698 445022 409934
rect 444786 374018 445022 374254
rect 444786 373698 445022 373934
rect 444786 338018 445022 338254
rect 444786 337698 445022 337934
rect 444786 302018 445022 302254
rect 444786 301698 445022 301934
rect 444786 266018 445022 266254
rect 444786 265698 445022 265934
rect 444786 230018 445022 230254
rect 444786 229698 445022 229934
rect 444786 194018 445022 194254
rect 444786 193698 445022 193934
rect 444786 158018 445022 158254
rect 444786 157698 445022 157934
rect 444786 122018 445022 122254
rect 444786 121698 445022 121934
rect 444786 86018 445022 86254
rect 444786 85698 445022 85934
rect 444786 50018 445022 50254
rect 444786 49698 445022 49934
rect 444786 14018 445022 14254
rect 444786 13698 445022 13934
rect 426786 -7162 427022 -6926
rect 426786 -7482 427022 -7246
rect 451986 705542 452222 705778
rect 451986 705222 452222 705458
rect 451986 669218 452222 669454
rect 451986 668898 452222 669134
rect 451986 633218 452222 633454
rect 451986 632898 452222 633134
rect 451986 597218 452222 597454
rect 451986 596898 452222 597134
rect 451986 561218 452222 561454
rect 451986 560898 452222 561134
rect 451986 525218 452222 525454
rect 451986 524898 452222 525134
rect 451986 489218 452222 489454
rect 451986 488898 452222 489134
rect 451986 453218 452222 453454
rect 451986 452898 452222 453134
rect 451986 417218 452222 417454
rect 451986 416898 452222 417134
rect 451986 381218 452222 381454
rect 451986 380898 452222 381134
rect 451986 345218 452222 345454
rect 451986 344898 452222 345134
rect 451986 309218 452222 309454
rect 451986 308898 452222 309134
rect 451986 273218 452222 273454
rect 451986 272898 452222 273134
rect 451986 237218 452222 237454
rect 451986 236898 452222 237134
rect 451986 201218 452222 201454
rect 451986 200898 452222 201134
rect 451986 165218 452222 165454
rect 451986 164898 452222 165134
rect 451986 129218 452222 129454
rect 451986 128898 452222 129134
rect 451986 93218 452222 93454
rect 451986 92898 452222 93134
rect 451986 57218 452222 57454
rect 451986 56898 452222 57134
rect 451986 21218 452222 21454
rect 451986 20898 452222 21134
rect 451986 -1522 452222 -1286
rect 451986 -1842 452222 -1606
rect 455586 672818 455822 673054
rect 455586 672498 455822 672734
rect 455586 636818 455822 637054
rect 455586 636498 455822 636734
rect 455586 600818 455822 601054
rect 455586 600498 455822 600734
rect 455586 564818 455822 565054
rect 455586 564498 455822 564734
rect 455586 528818 455822 529054
rect 455586 528498 455822 528734
rect 455586 492818 455822 493054
rect 455586 492498 455822 492734
rect 455586 456818 455822 457054
rect 455586 456498 455822 456734
rect 455586 420818 455822 421054
rect 455586 420498 455822 420734
rect 455586 384818 455822 385054
rect 455586 384498 455822 384734
rect 455586 348818 455822 349054
rect 455586 348498 455822 348734
rect 455586 312818 455822 313054
rect 455586 312498 455822 312734
rect 455586 276818 455822 277054
rect 455586 276498 455822 276734
rect 455586 240818 455822 241054
rect 455586 240498 455822 240734
rect 455586 204818 455822 205054
rect 455586 204498 455822 204734
rect 455586 168818 455822 169054
rect 455586 168498 455822 168734
rect 455586 132818 455822 133054
rect 455586 132498 455822 132734
rect 455586 96818 455822 97054
rect 455586 96498 455822 96734
rect 455586 60818 455822 61054
rect 455586 60498 455822 60734
rect 455586 24818 455822 25054
rect 455586 24498 455822 24734
rect 455586 -3402 455822 -3166
rect 455586 -3722 455822 -3486
rect 459186 676418 459422 676654
rect 459186 676098 459422 676334
rect 459186 640418 459422 640654
rect 459186 640098 459422 640334
rect 459186 604418 459422 604654
rect 459186 604098 459422 604334
rect 459186 568418 459422 568654
rect 459186 568098 459422 568334
rect 459186 532418 459422 532654
rect 459186 532098 459422 532334
rect 459186 496418 459422 496654
rect 459186 496098 459422 496334
rect 459186 460418 459422 460654
rect 459186 460098 459422 460334
rect 459186 424418 459422 424654
rect 459186 424098 459422 424334
rect 459186 388418 459422 388654
rect 459186 388098 459422 388334
rect 459186 352418 459422 352654
rect 459186 352098 459422 352334
rect 459186 316418 459422 316654
rect 459186 316098 459422 316334
rect 459186 280418 459422 280654
rect 459186 280098 459422 280334
rect 459186 244418 459422 244654
rect 459186 244098 459422 244334
rect 459186 208418 459422 208654
rect 459186 208098 459422 208334
rect 459186 172418 459422 172654
rect 459186 172098 459422 172334
rect 459186 136418 459422 136654
rect 459186 136098 459422 136334
rect 459186 100418 459422 100654
rect 459186 100098 459422 100334
rect 459186 64418 459422 64654
rect 459186 64098 459422 64334
rect 459186 28418 459422 28654
rect 459186 28098 459422 28334
rect 459186 -5282 459422 -5046
rect 459186 -5602 459422 -5366
rect 480786 710242 481022 710478
rect 480786 709922 481022 710158
rect 477186 708362 477422 708598
rect 477186 708042 477422 708278
rect 473586 706482 473822 706718
rect 473586 706162 473822 706398
rect 462786 680018 463022 680254
rect 462786 679698 463022 679934
rect 462786 644018 463022 644254
rect 462786 643698 463022 643934
rect 462786 608018 463022 608254
rect 462786 607698 463022 607934
rect 462786 572018 463022 572254
rect 462786 571698 463022 571934
rect 462786 536018 463022 536254
rect 462786 535698 463022 535934
rect 462786 500018 463022 500254
rect 462786 499698 463022 499934
rect 462786 464018 463022 464254
rect 462786 463698 463022 463934
rect 462786 428018 463022 428254
rect 462786 427698 463022 427934
rect 462786 392018 463022 392254
rect 462786 391698 463022 391934
rect 462786 356018 463022 356254
rect 462786 355698 463022 355934
rect 462786 320018 463022 320254
rect 462786 319698 463022 319934
rect 462786 284018 463022 284254
rect 462786 283698 463022 283934
rect 462786 248018 463022 248254
rect 462786 247698 463022 247934
rect 462786 212018 463022 212254
rect 462786 211698 463022 211934
rect 462786 176018 463022 176254
rect 462786 175698 463022 175934
rect 462786 140018 463022 140254
rect 462786 139698 463022 139934
rect 462786 104018 463022 104254
rect 462786 103698 463022 103934
rect 462786 68018 463022 68254
rect 462786 67698 463022 67934
rect 462786 32018 463022 32254
rect 462786 31698 463022 31934
rect 444786 -6222 445022 -5986
rect 444786 -6542 445022 -6306
rect 469986 704602 470222 704838
rect 469986 704282 470222 704518
rect 469986 687218 470222 687454
rect 469986 686898 470222 687134
rect 469986 651218 470222 651454
rect 469986 650898 470222 651134
rect 469986 615218 470222 615454
rect 469986 614898 470222 615134
rect 469986 579218 470222 579454
rect 469986 578898 470222 579134
rect 469986 543218 470222 543454
rect 469986 542898 470222 543134
rect 469986 507218 470222 507454
rect 469986 506898 470222 507134
rect 469986 471218 470222 471454
rect 469986 470898 470222 471134
rect 469986 435218 470222 435454
rect 469986 434898 470222 435134
rect 469986 399218 470222 399454
rect 469986 398898 470222 399134
rect 469986 363218 470222 363454
rect 469986 362898 470222 363134
rect 469986 327218 470222 327454
rect 469986 326898 470222 327134
rect 469986 291218 470222 291454
rect 469986 290898 470222 291134
rect 469986 255218 470222 255454
rect 469986 254898 470222 255134
rect 469986 219218 470222 219454
rect 469986 218898 470222 219134
rect 469986 183218 470222 183454
rect 469986 182898 470222 183134
rect 469986 147218 470222 147454
rect 469986 146898 470222 147134
rect 469986 111218 470222 111454
rect 469986 110898 470222 111134
rect 469986 75218 470222 75454
rect 469986 74898 470222 75134
rect 469986 39218 470222 39454
rect 469986 38898 470222 39134
rect 469986 3218 470222 3454
rect 469986 2898 470222 3134
rect 469986 -582 470222 -346
rect 469986 -902 470222 -666
rect 473586 690818 473822 691054
rect 473586 690498 473822 690734
rect 473586 654818 473822 655054
rect 473586 654498 473822 654734
rect 473586 618818 473822 619054
rect 473586 618498 473822 618734
rect 473586 582818 473822 583054
rect 473586 582498 473822 582734
rect 473586 546818 473822 547054
rect 473586 546498 473822 546734
rect 473586 510818 473822 511054
rect 473586 510498 473822 510734
rect 473586 474818 473822 475054
rect 473586 474498 473822 474734
rect 473586 438818 473822 439054
rect 473586 438498 473822 438734
rect 473586 402818 473822 403054
rect 473586 402498 473822 402734
rect 473586 366818 473822 367054
rect 473586 366498 473822 366734
rect 473586 330818 473822 331054
rect 473586 330498 473822 330734
rect 473586 294818 473822 295054
rect 473586 294498 473822 294734
rect 473586 258818 473822 259054
rect 473586 258498 473822 258734
rect 473586 222818 473822 223054
rect 473586 222498 473822 222734
rect 473586 186818 473822 187054
rect 473586 186498 473822 186734
rect 473586 150818 473822 151054
rect 473586 150498 473822 150734
rect 473586 114818 473822 115054
rect 473586 114498 473822 114734
rect 473586 78818 473822 79054
rect 473586 78498 473822 78734
rect 473586 42818 473822 43054
rect 473586 42498 473822 42734
rect 473586 6818 473822 7054
rect 473586 6498 473822 6734
rect 473586 -2462 473822 -2226
rect 473586 -2782 473822 -2546
rect 477186 694418 477422 694654
rect 477186 694098 477422 694334
rect 477186 658418 477422 658654
rect 477186 658098 477422 658334
rect 477186 622418 477422 622654
rect 477186 622098 477422 622334
rect 477186 586418 477422 586654
rect 477186 586098 477422 586334
rect 477186 550418 477422 550654
rect 477186 550098 477422 550334
rect 477186 514418 477422 514654
rect 477186 514098 477422 514334
rect 477186 478418 477422 478654
rect 477186 478098 477422 478334
rect 477186 442418 477422 442654
rect 477186 442098 477422 442334
rect 477186 406418 477422 406654
rect 477186 406098 477422 406334
rect 477186 370418 477422 370654
rect 477186 370098 477422 370334
rect 477186 334418 477422 334654
rect 477186 334098 477422 334334
rect 477186 298418 477422 298654
rect 477186 298098 477422 298334
rect 477186 262418 477422 262654
rect 477186 262098 477422 262334
rect 477186 226418 477422 226654
rect 477186 226098 477422 226334
rect 477186 190418 477422 190654
rect 477186 190098 477422 190334
rect 477186 154418 477422 154654
rect 477186 154098 477422 154334
rect 477186 118418 477422 118654
rect 477186 118098 477422 118334
rect 477186 82418 477422 82654
rect 477186 82098 477422 82334
rect 477186 46418 477422 46654
rect 477186 46098 477422 46334
rect 477186 10418 477422 10654
rect 477186 10098 477422 10334
rect 477186 -4342 477422 -4106
rect 477186 -4662 477422 -4426
rect 498786 711182 499022 711418
rect 498786 710862 499022 711098
rect 495186 709302 495422 709538
rect 495186 708982 495422 709218
rect 491586 707422 491822 707658
rect 491586 707102 491822 707338
rect 480786 698018 481022 698254
rect 480786 697698 481022 697934
rect 480786 662018 481022 662254
rect 480786 661698 481022 661934
rect 480786 626018 481022 626254
rect 480786 625698 481022 625934
rect 480786 590018 481022 590254
rect 480786 589698 481022 589934
rect 480786 554018 481022 554254
rect 480786 553698 481022 553934
rect 480786 518018 481022 518254
rect 480786 517698 481022 517934
rect 480786 482018 481022 482254
rect 480786 481698 481022 481934
rect 480786 446018 481022 446254
rect 480786 445698 481022 445934
rect 480786 410018 481022 410254
rect 480786 409698 481022 409934
rect 480786 374018 481022 374254
rect 480786 373698 481022 373934
rect 480786 338018 481022 338254
rect 480786 337698 481022 337934
rect 480786 302018 481022 302254
rect 480786 301698 481022 301934
rect 480786 266018 481022 266254
rect 480786 265698 481022 265934
rect 480786 230018 481022 230254
rect 480786 229698 481022 229934
rect 480786 194018 481022 194254
rect 480786 193698 481022 193934
rect 480786 158018 481022 158254
rect 480786 157698 481022 157934
rect 480786 122018 481022 122254
rect 480786 121698 481022 121934
rect 480786 86018 481022 86254
rect 480786 85698 481022 85934
rect 480786 50018 481022 50254
rect 480786 49698 481022 49934
rect 480786 14018 481022 14254
rect 480786 13698 481022 13934
rect 462786 -7162 463022 -6926
rect 462786 -7482 463022 -7246
rect 487986 705542 488222 705778
rect 487986 705222 488222 705458
rect 487986 669218 488222 669454
rect 487986 668898 488222 669134
rect 487986 633218 488222 633454
rect 487986 632898 488222 633134
rect 487986 597218 488222 597454
rect 487986 596898 488222 597134
rect 487986 561218 488222 561454
rect 487986 560898 488222 561134
rect 487986 525218 488222 525454
rect 487986 524898 488222 525134
rect 487986 489218 488222 489454
rect 487986 488898 488222 489134
rect 487986 453218 488222 453454
rect 487986 452898 488222 453134
rect 487986 417218 488222 417454
rect 487986 416898 488222 417134
rect 487986 381218 488222 381454
rect 487986 380898 488222 381134
rect 487986 345218 488222 345454
rect 487986 344898 488222 345134
rect 487986 309218 488222 309454
rect 487986 308898 488222 309134
rect 487986 273218 488222 273454
rect 487986 272898 488222 273134
rect 487986 237218 488222 237454
rect 487986 236898 488222 237134
rect 487986 201218 488222 201454
rect 487986 200898 488222 201134
rect 487986 165218 488222 165454
rect 487986 164898 488222 165134
rect 487986 129218 488222 129454
rect 487986 128898 488222 129134
rect 487986 93218 488222 93454
rect 487986 92898 488222 93134
rect 487986 57218 488222 57454
rect 487986 56898 488222 57134
rect 487986 21218 488222 21454
rect 487986 20898 488222 21134
rect 487986 -1522 488222 -1286
rect 487986 -1842 488222 -1606
rect 491586 672818 491822 673054
rect 491586 672498 491822 672734
rect 491586 636818 491822 637054
rect 491586 636498 491822 636734
rect 491586 600818 491822 601054
rect 491586 600498 491822 600734
rect 491586 564818 491822 565054
rect 491586 564498 491822 564734
rect 491586 528818 491822 529054
rect 491586 528498 491822 528734
rect 491586 492818 491822 493054
rect 491586 492498 491822 492734
rect 491586 456818 491822 457054
rect 491586 456498 491822 456734
rect 491586 420818 491822 421054
rect 491586 420498 491822 420734
rect 491586 384818 491822 385054
rect 491586 384498 491822 384734
rect 491586 348818 491822 349054
rect 491586 348498 491822 348734
rect 491586 312818 491822 313054
rect 491586 312498 491822 312734
rect 491586 276818 491822 277054
rect 491586 276498 491822 276734
rect 491586 240818 491822 241054
rect 491586 240498 491822 240734
rect 491586 204818 491822 205054
rect 491586 204498 491822 204734
rect 491586 168818 491822 169054
rect 491586 168498 491822 168734
rect 491586 132818 491822 133054
rect 491586 132498 491822 132734
rect 491586 96818 491822 97054
rect 491586 96498 491822 96734
rect 491586 60818 491822 61054
rect 491586 60498 491822 60734
rect 491586 24818 491822 25054
rect 491586 24498 491822 24734
rect 491586 -3402 491822 -3166
rect 491586 -3722 491822 -3486
rect 495186 676418 495422 676654
rect 495186 676098 495422 676334
rect 495186 640418 495422 640654
rect 495186 640098 495422 640334
rect 495186 604418 495422 604654
rect 495186 604098 495422 604334
rect 495186 568418 495422 568654
rect 495186 568098 495422 568334
rect 495186 532418 495422 532654
rect 495186 532098 495422 532334
rect 495186 496418 495422 496654
rect 495186 496098 495422 496334
rect 495186 460418 495422 460654
rect 495186 460098 495422 460334
rect 495186 424418 495422 424654
rect 495186 424098 495422 424334
rect 495186 388418 495422 388654
rect 495186 388098 495422 388334
rect 495186 352418 495422 352654
rect 495186 352098 495422 352334
rect 495186 316418 495422 316654
rect 495186 316098 495422 316334
rect 495186 280418 495422 280654
rect 495186 280098 495422 280334
rect 495186 244418 495422 244654
rect 495186 244098 495422 244334
rect 495186 208418 495422 208654
rect 495186 208098 495422 208334
rect 495186 172418 495422 172654
rect 495186 172098 495422 172334
rect 495186 136418 495422 136654
rect 495186 136098 495422 136334
rect 495186 100418 495422 100654
rect 495186 100098 495422 100334
rect 495186 64418 495422 64654
rect 495186 64098 495422 64334
rect 495186 28418 495422 28654
rect 495186 28098 495422 28334
rect 495186 -5282 495422 -5046
rect 495186 -5602 495422 -5366
rect 516786 710242 517022 710478
rect 516786 709922 517022 710158
rect 513186 708362 513422 708598
rect 513186 708042 513422 708278
rect 509586 706482 509822 706718
rect 509586 706162 509822 706398
rect 498786 680018 499022 680254
rect 498786 679698 499022 679934
rect 498786 644018 499022 644254
rect 498786 643698 499022 643934
rect 498786 608018 499022 608254
rect 498786 607698 499022 607934
rect 498786 572018 499022 572254
rect 498786 571698 499022 571934
rect 498786 536018 499022 536254
rect 498786 535698 499022 535934
rect 498786 500018 499022 500254
rect 498786 499698 499022 499934
rect 498786 464018 499022 464254
rect 498786 463698 499022 463934
rect 498786 428018 499022 428254
rect 498786 427698 499022 427934
rect 498786 392018 499022 392254
rect 498786 391698 499022 391934
rect 498786 356018 499022 356254
rect 498786 355698 499022 355934
rect 498786 320018 499022 320254
rect 498786 319698 499022 319934
rect 498786 284018 499022 284254
rect 498786 283698 499022 283934
rect 498786 248018 499022 248254
rect 498786 247698 499022 247934
rect 498786 212018 499022 212254
rect 498786 211698 499022 211934
rect 498786 176018 499022 176254
rect 498786 175698 499022 175934
rect 498786 140018 499022 140254
rect 498786 139698 499022 139934
rect 498786 104018 499022 104254
rect 498786 103698 499022 103934
rect 498786 68018 499022 68254
rect 498786 67698 499022 67934
rect 498786 32018 499022 32254
rect 498786 31698 499022 31934
rect 480786 -6222 481022 -5986
rect 480786 -6542 481022 -6306
rect 505986 704602 506222 704838
rect 505986 704282 506222 704518
rect 505986 687218 506222 687454
rect 505986 686898 506222 687134
rect 505986 651218 506222 651454
rect 505986 650898 506222 651134
rect 505986 615218 506222 615454
rect 505986 614898 506222 615134
rect 505986 579218 506222 579454
rect 505986 578898 506222 579134
rect 505986 543218 506222 543454
rect 505986 542898 506222 543134
rect 505986 507218 506222 507454
rect 505986 506898 506222 507134
rect 505986 471218 506222 471454
rect 505986 470898 506222 471134
rect 505986 435218 506222 435454
rect 505986 434898 506222 435134
rect 505986 399218 506222 399454
rect 505986 398898 506222 399134
rect 505986 363218 506222 363454
rect 505986 362898 506222 363134
rect 505986 327218 506222 327454
rect 505986 326898 506222 327134
rect 505986 291218 506222 291454
rect 505986 290898 506222 291134
rect 505986 255218 506222 255454
rect 505986 254898 506222 255134
rect 505986 219218 506222 219454
rect 505986 218898 506222 219134
rect 505986 183218 506222 183454
rect 505986 182898 506222 183134
rect 505986 147218 506222 147454
rect 505986 146898 506222 147134
rect 505986 111218 506222 111454
rect 505986 110898 506222 111134
rect 505986 75218 506222 75454
rect 505986 74898 506222 75134
rect 505986 39218 506222 39454
rect 505986 38898 506222 39134
rect 505986 3218 506222 3454
rect 505986 2898 506222 3134
rect 505986 -582 506222 -346
rect 505986 -902 506222 -666
rect 509586 690818 509822 691054
rect 509586 690498 509822 690734
rect 509586 654818 509822 655054
rect 509586 654498 509822 654734
rect 509586 618818 509822 619054
rect 509586 618498 509822 618734
rect 509586 582818 509822 583054
rect 509586 582498 509822 582734
rect 509586 546818 509822 547054
rect 509586 546498 509822 546734
rect 509586 510818 509822 511054
rect 509586 510498 509822 510734
rect 509586 474818 509822 475054
rect 509586 474498 509822 474734
rect 509586 438818 509822 439054
rect 509586 438498 509822 438734
rect 509586 402818 509822 403054
rect 509586 402498 509822 402734
rect 509586 366818 509822 367054
rect 509586 366498 509822 366734
rect 509586 330818 509822 331054
rect 509586 330498 509822 330734
rect 509586 294818 509822 295054
rect 509586 294498 509822 294734
rect 509586 258818 509822 259054
rect 509586 258498 509822 258734
rect 509586 222818 509822 223054
rect 509586 222498 509822 222734
rect 509586 186818 509822 187054
rect 509586 186498 509822 186734
rect 509586 150818 509822 151054
rect 509586 150498 509822 150734
rect 509586 114818 509822 115054
rect 509586 114498 509822 114734
rect 509586 78818 509822 79054
rect 509586 78498 509822 78734
rect 509586 42818 509822 43054
rect 509586 42498 509822 42734
rect 509586 6818 509822 7054
rect 509586 6498 509822 6734
rect 509586 -2462 509822 -2226
rect 509586 -2782 509822 -2546
rect 513186 694418 513422 694654
rect 513186 694098 513422 694334
rect 513186 658418 513422 658654
rect 513186 658098 513422 658334
rect 513186 622418 513422 622654
rect 513186 622098 513422 622334
rect 513186 586418 513422 586654
rect 513186 586098 513422 586334
rect 513186 550418 513422 550654
rect 513186 550098 513422 550334
rect 513186 514418 513422 514654
rect 513186 514098 513422 514334
rect 513186 478418 513422 478654
rect 513186 478098 513422 478334
rect 513186 442418 513422 442654
rect 513186 442098 513422 442334
rect 513186 406418 513422 406654
rect 513186 406098 513422 406334
rect 513186 370418 513422 370654
rect 513186 370098 513422 370334
rect 513186 334418 513422 334654
rect 513186 334098 513422 334334
rect 513186 298418 513422 298654
rect 513186 298098 513422 298334
rect 513186 262418 513422 262654
rect 513186 262098 513422 262334
rect 513186 226418 513422 226654
rect 513186 226098 513422 226334
rect 513186 190418 513422 190654
rect 513186 190098 513422 190334
rect 513186 154418 513422 154654
rect 513186 154098 513422 154334
rect 513186 118418 513422 118654
rect 513186 118098 513422 118334
rect 513186 82418 513422 82654
rect 513186 82098 513422 82334
rect 513186 46418 513422 46654
rect 513186 46098 513422 46334
rect 513186 10418 513422 10654
rect 513186 10098 513422 10334
rect 513186 -4342 513422 -4106
rect 513186 -4662 513422 -4426
rect 534786 711182 535022 711418
rect 534786 710862 535022 711098
rect 531186 709302 531422 709538
rect 531186 708982 531422 709218
rect 527586 707422 527822 707658
rect 527586 707102 527822 707338
rect 516786 698018 517022 698254
rect 516786 697698 517022 697934
rect 516786 662018 517022 662254
rect 516786 661698 517022 661934
rect 516786 626018 517022 626254
rect 516786 625698 517022 625934
rect 516786 590018 517022 590254
rect 516786 589698 517022 589934
rect 516786 554018 517022 554254
rect 516786 553698 517022 553934
rect 516786 518018 517022 518254
rect 516786 517698 517022 517934
rect 516786 482018 517022 482254
rect 516786 481698 517022 481934
rect 516786 446018 517022 446254
rect 516786 445698 517022 445934
rect 516786 410018 517022 410254
rect 516786 409698 517022 409934
rect 516786 374018 517022 374254
rect 516786 373698 517022 373934
rect 516786 338018 517022 338254
rect 516786 337698 517022 337934
rect 516786 302018 517022 302254
rect 516786 301698 517022 301934
rect 516786 266018 517022 266254
rect 516786 265698 517022 265934
rect 516786 230018 517022 230254
rect 516786 229698 517022 229934
rect 516786 194018 517022 194254
rect 516786 193698 517022 193934
rect 516786 158018 517022 158254
rect 516786 157698 517022 157934
rect 516786 122018 517022 122254
rect 516786 121698 517022 121934
rect 516786 86018 517022 86254
rect 516786 85698 517022 85934
rect 516786 50018 517022 50254
rect 516786 49698 517022 49934
rect 516786 14018 517022 14254
rect 516786 13698 517022 13934
rect 498786 -7162 499022 -6926
rect 498786 -7482 499022 -7246
rect 523986 705542 524222 705778
rect 523986 705222 524222 705458
rect 523986 669218 524222 669454
rect 523986 668898 524222 669134
rect 523986 633218 524222 633454
rect 523986 632898 524222 633134
rect 523986 597218 524222 597454
rect 523986 596898 524222 597134
rect 523986 561218 524222 561454
rect 523986 560898 524222 561134
rect 523986 525218 524222 525454
rect 523986 524898 524222 525134
rect 523986 489218 524222 489454
rect 523986 488898 524222 489134
rect 523986 453218 524222 453454
rect 523986 452898 524222 453134
rect 523986 417218 524222 417454
rect 523986 416898 524222 417134
rect 523986 381218 524222 381454
rect 523986 380898 524222 381134
rect 523986 345218 524222 345454
rect 523986 344898 524222 345134
rect 523986 309218 524222 309454
rect 523986 308898 524222 309134
rect 523986 273218 524222 273454
rect 523986 272898 524222 273134
rect 523986 237218 524222 237454
rect 523986 236898 524222 237134
rect 523986 201218 524222 201454
rect 523986 200898 524222 201134
rect 523986 165218 524222 165454
rect 523986 164898 524222 165134
rect 523986 129218 524222 129454
rect 523986 128898 524222 129134
rect 523986 93218 524222 93454
rect 523986 92898 524222 93134
rect 523986 57218 524222 57454
rect 523986 56898 524222 57134
rect 523986 21218 524222 21454
rect 523986 20898 524222 21134
rect 523986 -1522 524222 -1286
rect 523986 -1842 524222 -1606
rect 527586 672818 527822 673054
rect 527586 672498 527822 672734
rect 527586 636818 527822 637054
rect 527586 636498 527822 636734
rect 527586 600818 527822 601054
rect 527586 600498 527822 600734
rect 527586 564818 527822 565054
rect 527586 564498 527822 564734
rect 527586 528818 527822 529054
rect 527586 528498 527822 528734
rect 527586 492818 527822 493054
rect 527586 492498 527822 492734
rect 527586 456818 527822 457054
rect 527586 456498 527822 456734
rect 527586 420818 527822 421054
rect 527586 420498 527822 420734
rect 527586 384818 527822 385054
rect 527586 384498 527822 384734
rect 527586 348818 527822 349054
rect 527586 348498 527822 348734
rect 527586 312818 527822 313054
rect 527586 312498 527822 312734
rect 527586 276818 527822 277054
rect 527586 276498 527822 276734
rect 527586 240818 527822 241054
rect 527586 240498 527822 240734
rect 527586 204818 527822 205054
rect 527586 204498 527822 204734
rect 527586 168818 527822 169054
rect 527586 168498 527822 168734
rect 527586 132818 527822 133054
rect 527586 132498 527822 132734
rect 527586 96818 527822 97054
rect 527586 96498 527822 96734
rect 527586 60818 527822 61054
rect 527586 60498 527822 60734
rect 527586 24818 527822 25054
rect 527586 24498 527822 24734
rect 527586 -3402 527822 -3166
rect 527586 -3722 527822 -3486
rect 531186 676418 531422 676654
rect 531186 676098 531422 676334
rect 531186 640418 531422 640654
rect 531186 640098 531422 640334
rect 531186 604418 531422 604654
rect 531186 604098 531422 604334
rect 531186 568418 531422 568654
rect 531186 568098 531422 568334
rect 531186 532418 531422 532654
rect 531186 532098 531422 532334
rect 531186 496418 531422 496654
rect 531186 496098 531422 496334
rect 531186 460418 531422 460654
rect 531186 460098 531422 460334
rect 531186 424418 531422 424654
rect 531186 424098 531422 424334
rect 531186 388418 531422 388654
rect 531186 388098 531422 388334
rect 531186 352418 531422 352654
rect 531186 352098 531422 352334
rect 531186 316418 531422 316654
rect 531186 316098 531422 316334
rect 531186 280418 531422 280654
rect 531186 280098 531422 280334
rect 531186 244418 531422 244654
rect 531186 244098 531422 244334
rect 531186 208418 531422 208654
rect 531186 208098 531422 208334
rect 531186 172418 531422 172654
rect 531186 172098 531422 172334
rect 531186 136418 531422 136654
rect 531186 136098 531422 136334
rect 531186 100418 531422 100654
rect 531186 100098 531422 100334
rect 531186 64418 531422 64654
rect 531186 64098 531422 64334
rect 531186 28418 531422 28654
rect 531186 28098 531422 28334
rect 531186 -5282 531422 -5046
rect 531186 -5602 531422 -5366
rect 552786 710242 553022 710478
rect 552786 709922 553022 710158
rect 549186 708362 549422 708598
rect 549186 708042 549422 708278
rect 545586 706482 545822 706718
rect 545586 706162 545822 706398
rect 534786 680018 535022 680254
rect 534786 679698 535022 679934
rect 534786 644018 535022 644254
rect 534786 643698 535022 643934
rect 534786 608018 535022 608254
rect 534786 607698 535022 607934
rect 534786 572018 535022 572254
rect 534786 571698 535022 571934
rect 534786 536018 535022 536254
rect 534786 535698 535022 535934
rect 534786 500018 535022 500254
rect 534786 499698 535022 499934
rect 534786 464018 535022 464254
rect 534786 463698 535022 463934
rect 534786 428018 535022 428254
rect 534786 427698 535022 427934
rect 534786 392018 535022 392254
rect 534786 391698 535022 391934
rect 534786 356018 535022 356254
rect 534786 355698 535022 355934
rect 534786 320018 535022 320254
rect 534786 319698 535022 319934
rect 534786 284018 535022 284254
rect 534786 283698 535022 283934
rect 534786 248018 535022 248254
rect 534786 247698 535022 247934
rect 534786 212018 535022 212254
rect 534786 211698 535022 211934
rect 534786 176018 535022 176254
rect 534786 175698 535022 175934
rect 534786 140018 535022 140254
rect 534786 139698 535022 139934
rect 534786 104018 535022 104254
rect 534786 103698 535022 103934
rect 534786 68018 535022 68254
rect 534786 67698 535022 67934
rect 534786 32018 535022 32254
rect 534786 31698 535022 31934
rect 516786 -6222 517022 -5986
rect 516786 -6542 517022 -6306
rect 541986 704602 542222 704838
rect 541986 704282 542222 704518
rect 541986 687218 542222 687454
rect 541986 686898 542222 687134
rect 541986 651218 542222 651454
rect 541986 650898 542222 651134
rect 541986 615218 542222 615454
rect 541986 614898 542222 615134
rect 541986 579218 542222 579454
rect 541986 578898 542222 579134
rect 541986 543218 542222 543454
rect 541986 542898 542222 543134
rect 541986 507218 542222 507454
rect 541986 506898 542222 507134
rect 541986 471218 542222 471454
rect 541986 470898 542222 471134
rect 541986 435218 542222 435454
rect 541986 434898 542222 435134
rect 541986 399218 542222 399454
rect 541986 398898 542222 399134
rect 541986 363218 542222 363454
rect 541986 362898 542222 363134
rect 541986 327218 542222 327454
rect 541986 326898 542222 327134
rect 541986 291218 542222 291454
rect 541986 290898 542222 291134
rect 541986 255218 542222 255454
rect 541986 254898 542222 255134
rect 541986 219218 542222 219454
rect 541986 218898 542222 219134
rect 541986 183218 542222 183454
rect 541986 182898 542222 183134
rect 541986 147218 542222 147454
rect 541986 146898 542222 147134
rect 541986 111218 542222 111454
rect 541986 110898 542222 111134
rect 541986 75218 542222 75454
rect 541986 74898 542222 75134
rect 541986 39218 542222 39454
rect 541986 38898 542222 39134
rect 541986 3218 542222 3454
rect 541986 2898 542222 3134
rect 541986 -582 542222 -346
rect 541986 -902 542222 -666
rect 545586 690818 545822 691054
rect 545586 690498 545822 690734
rect 545586 654818 545822 655054
rect 545586 654498 545822 654734
rect 545586 618818 545822 619054
rect 545586 618498 545822 618734
rect 545586 582818 545822 583054
rect 545586 582498 545822 582734
rect 545586 546818 545822 547054
rect 545586 546498 545822 546734
rect 545586 510818 545822 511054
rect 545586 510498 545822 510734
rect 545586 474818 545822 475054
rect 545586 474498 545822 474734
rect 545586 438818 545822 439054
rect 545586 438498 545822 438734
rect 545586 402818 545822 403054
rect 545586 402498 545822 402734
rect 545586 366818 545822 367054
rect 545586 366498 545822 366734
rect 545586 330818 545822 331054
rect 545586 330498 545822 330734
rect 545586 294818 545822 295054
rect 545586 294498 545822 294734
rect 545586 258818 545822 259054
rect 545586 258498 545822 258734
rect 545586 222818 545822 223054
rect 545586 222498 545822 222734
rect 545586 186818 545822 187054
rect 545586 186498 545822 186734
rect 545586 150818 545822 151054
rect 545586 150498 545822 150734
rect 545586 114818 545822 115054
rect 545586 114498 545822 114734
rect 545586 78818 545822 79054
rect 545586 78498 545822 78734
rect 545586 42818 545822 43054
rect 545586 42498 545822 42734
rect 545586 6818 545822 7054
rect 545586 6498 545822 6734
rect 545586 -2462 545822 -2226
rect 545586 -2782 545822 -2546
rect 549186 694418 549422 694654
rect 549186 694098 549422 694334
rect 549186 658418 549422 658654
rect 549186 658098 549422 658334
rect 549186 622418 549422 622654
rect 549186 622098 549422 622334
rect 549186 586418 549422 586654
rect 549186 586098 549422 586334
rect 549186 550418 549422 550654
rect 549186 550098 549422 550334
rect 549186 514418 549422 514654
rect 549186 514098 549422 514334
rect 549186 478418 549422 478654
rect 549186 478098 549422 478334
rect 549186 442418 549422 442654
rect 549186 442098 549422 442334
rect 549186 406418 549422 406654
rect 549186 406098 549422 406334
rect 549186 370418 549422 370654
rect 549186 370098 549422 370334
rect 549186 334418 549422 334654
rect 549186 334098 549422 334334
rect 549186 298418 549422 298654
rect 549186 298098 549422 298334
rect 549186 262418 549422 262654
rect 549186 262098 549422 262334
rect 549186 226418 549422 226654
rect 549186 226098 549422 226334
rect 549186 190418 549422 190654
rect 549186 190098 549422 190334
rect 549186 154418 549422 154654
rect 549186 154098 549422 154334
rect 549186 118418 549422 118654
rect 549186 118098 549422 118334
rect 549186 82418 549422 82654
rect 549186 82098 549422 82334
rect 549186 46418 549422 46654
rect 549186 46098 549422 46334
rect 549186 10418 549422 10654
rect 549186 10098 549422 10334
rect 549186 -4342 549422 -4106
rect 549186 -4662 549422 -4426
rect 570786 711182 571022 711418
rect 570786 710862 571022 711098
rect 567186 709302 567422 709538
rect 567186 708982 567422 709218
rect 563586 707422 563822 707658
rect 563586 707102 563822 707338
rect 552786 698018 553022 698254
rect 552786 697698 553022 697934
rect 552786 662018 553022 662254
rect 552786 661698 553022 661934
rect 552786 626018 553022 626254
rect 552786 625698 553022 625934
rect 552786 590018 553022 590254
rect 552786 589698 553022 589934
rect 552786 554018 553022 554254
rect 552786 553698 553022 553934
rect 552786 518018 553022 518254
rect 552786 517698 553022 517934
rect 552786 482018 553022 482254
rect 552786 481698 553022 481934
rect 552786 446018 553022 446254
rect 552786 445698 553022 445934
rect 552786 410018 553022 410254
rect 552786 409698 553022 409934
rect 552786 374018 553022 374254
rect 552786 373698 553022 373934
rect 552786 338018 553022 338254
rect 552786 337698 553022 337934
rect 552786 302018 553022 302254
rect 552786 301698 553022 301934
rect 552786 266018 553022 266254
rect 552786 265698 553022 265934
rect 552786 230018 553022 230254
rect 552786 229698 553022 229934
rect 552786 194018 553022 194254
rect 552786 193698 553022 193934
rect 552786 158018 553022 158254
rect 552786 157698 553022 157934
rect 552786 122018 553022 122254
rect 552786 121698 553022 121934
rect 552786 86018 553022 86254
rect 552786 85698 553022 85934
rect 552786 50018 553022 50254
rect 552786 49698 553022 49934
rect 552786 14018 553022 14254
rect 552786 13698 553022 13934
rect 534786 -7162 535022 -6926
rect 534786 -7482 535022 -7246
rect 559986 705542 560222 705778
rect 559986 705222 560222 705458
rect 559986 669218 560222 669454
rect 559986 668898 560222 669134
rect 559986 633218 560222 633454
rect 559986 632898 560222 633134
rect 559986 597218 560222 597454
rect 559986 596898 560222 597134
rect 559986 561218 560222 561454
rect 559986 560898 560222 561134
rect 559986 525218 560222 525454
rect 559986 524898 560222 525134
rect 559986 489218 560222 489454
rect 559986 488898 560222 489134
rect 559986 453218 560222 453454
rect 559986 452898 560222 453134
rect 559986 417218 560222 417454
rect 559986 416898 560222 417134
rect 559986 381218 560222 381454
rect 559986 380898 560222 381134
rect 559986 345218 560222 345454
rect 559986 344898 560222 345134
rect 559986 309218 560222 309454
rect 559986 308898 560222 309134
rect 559986 273218 560222 273454
rect 559986 272898 560222 273134
rect 559986 237218 560222 237454
rect 559986 236898 560222 237134
rect 559986 201218 560222 201454
rect 559986 200898 560222 201134
rect 559986 165218 560222 165454
rect 559986 164898 560222 165134
rect 559986 129218 560222 129454
rect 559986 128898 560222 129134
rect 559986 93218 560222 93454
rect 559986 92898 560222 93134
rect 559986 57218 560222 57454
rect 559986 56898 560222 57134
rect 559986 21218 560222 21454
rect 559986 20898 560222 21134
rect 559986 -1522 560222 -1286
rect 559986 -1842 560222 -1606
rect 563586 672818 563822 673054
rect 563586 672498 563822 672734
rect 563586 636818 563822 637054
rect 563586 636498 563822 636734
rect 563586 600818 563822 601054
rect 563586 600498 563822 600734
rect 563586 564818 563822 565054
rect 563586 564498 563822 564734
rect 563586 528818 563822 529054
rect 563586 528498 563822 528734
rect 563586 492818 563822 493054
rect 563586 492498 563822 492734
rect 563586 456818 563822 457054
rect 563586 456498 563822 456734
rect 563586 420818 563822 421054
rect 563586 420498 563822 420734
rect 563586 384818 563822 385054
rect 563586 384498 563822 384734
rect 563586 348818 563822 349054
rect 563586 348498 563822 348734
rect 563586 312818 563822 313054
rect 563586 312498 563822 312734
rect 563586 276818 563822 277054
rect 563586 276498 563822 276734
rect 563586 240818 563822 241054
rect 563586 240498 563822 240734
rect 563586 204818 563822 205054
rect 563586 204498 563822 204734
rect 563586 168818 563822 169054
rect 563586 168498 563822 168734
rect 563586 132818 563822 133054
rect 563586 132498 563822 132734
rect 563586 96818 563822 97054
rect 563586 96498 563822 96734
rect 563586 60818 563822 61054
rect 563586 60498 563822 60734
rect 563586 24818 563822 25054
rect 563586 24498 563822 24734
rect 563586 -3402 563822 -3166
rect 563586 -3722 563822 -3486
rect 567186 676418 567422 676654
rect 567186 676098 567422 676334
rect 567186 640418 567422 640654
rect 567186 640098 567422 640334
rect 567186 604418 567422 604654
rect 567186 604098 567422 604334
rect 567186 568418 567422 568654
rect 567186 568098 567422 568334
rect 567186 532418 567422 532654
rect 567186 532098 567422 532334
rect 567186 496418 567422 496654
rect 567186 496098 567422 496334
rect 567186 460418 567422 460654
rect 567186 460098 567422 460334
rect 567186 424418 567422 424654
rect 567186 424098 567422 424334
rect 567186 388418 567422 388654
rect 567186 388098 567422 388334
rect 567186 352418 567422 352654
rect 567186 352098 567422 352334
rect 567186 316418 567422 316654
rect 567186 316098 567422 316334
rect 567186 280418 567422 280654
rect 567186 280098 567422 280334
rect 567186 244418 567422 244654
rect 567186 244098 567422 244334
rect 567186 208418 567422 208654
rect 567186 208098 567422 208334
rect 567186 172418 567422 172654
rect 567186 172098 567422 172334
rect 567186 136418 567422 136654
rect 567186 136098 567422 136334
rect 567186 100418 567422 100654
rect 567186 100098 567422 100334
rect 567186 64418 567422 64654
rect 567186 64098 567422 64334
rect 567186 28418 567422 28654
rect 567186 28098 567422 28334
rect 567186 -5282 567422 -5046
rect 567186 -5602 567422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 581586 706482 581822 706718
rect 581586 706162 581822 706398
rect 570786 680018 571022 680254
rect 570786 679698 571022 679934
rect 570786 644018 571022 644254
rect 570786 643698 571022 643934
rect 570786 608018 571022 608254
rect 570786 607698 571022 607934
rect 570786 572018 571022 572254
rect 570786 571698 571022 571934
rect 570786 536018 571022 536254
rect 570786 535698 571022 535934
rect 570786 500018 571022 500254
rect 570786 499698 571022 499934
rect 570786 464018 571022 464254
rect 570786 463698 571022 463934
rect 570786 428018 571022 428254
rect 570786 427698 571022 427934
rect 570786 392018 571022 392254
rect 570786 391698 571022 391934
rect 570786 356018 571022 356254
rect 570786 355698 571022 355934
rect 570786 320018 571022 320254
rect 570786 319698 571022 319934
rect 570786 284018 571022 284254
rect 570786 283698 571022 283934
rect 570786 248018 571022 248254
rect 570786 247698 571022 247934
rect 570786 212018 571022 212254
rect 570786 211698 571022 211934
rect 570786 176018 571022 176254
rect 570786 175698 571022 175934
rect 570786 140018 571022 140254
rect 570786 139698 571022 139934
rect 570786 104018 571022 104254
rect 570786 103698 571022 103934
rect 570786 68018 571022 68254
rect 570786 67698 571022 67934
rect 570786 32018 571022 32254
rect 570786 31698 571022 31934
rect 552786 -6222 553022 -5986
rect 552786 -6542 553022 -6306
rect 577986 704602 578222 704838
rect 577986 704282 578222 704518
rect 577986 687218 578222 687454
rect 577986 686898 578222 687134
rect 577986 651218 578222 651454
rect 577986 650898 578222 651134
rect 577986 615218 578222 615454
rect 577986 614898 578222 615134
rect 577986 579218 578222 579454
rect 577986 578898 578222 579134
rect 577986 543218 578222 543454
rect 577986 542898 578222 543134
rect 577986 507218 578222 507454
rect 577986 506898 578222 507134
rect 577986 471218 578222 471454
rect 577986 470898 578222 471134
rect 577986 435218 578222 435454
rect 577986 434898 578222 435134
rect 577986 399218 578222 399454
rect 577986 398898 578222 399134
rect 577986 363218 578222 363454
rect 577986 362898 578222 363134
rect 577986 327218 578222 327454
rect 577986 326898 578222 327134
rect 577986 291218 578222 291454
rect 577986 290898 578222 291134
rect 577986 255218 578222 255454
rect 577986 254898 578222 255134
rect 577986 219218 578222 219454
rect 577986 218898 578222 219134
rect 577986 183218 578222 183454
rect 577986 182898 578222 183134
rect 577986 147218 578222 147454
rect 577986 146898 578222 147134
rect 577986 111218 578222 111454
rect 577986 110898 578222 111134
rect 577986 75218 578222 75454
rect 577986 74898 578222 75134
rect 577986 39218 578222 39454
rect 577986 38898 578222 39134
rect 577986 3218 578222 3454
rect 577986 2898 578222 3134
rect 577986 -582 578222 -346
rect 577986 -902 578222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 581586 690818 581822 691054
rect 581586 690498 581822 690734
rect 581586 654818 581822 655054
rect 581586 654498 581822 654734
rect 581586 618818 581822 619054
rect 581586 618498 581822 618734
rect 581586 582818 581822 583054
rect 581586 582498 581822 582734
rect 581586 546818 581822 547054
rect 581586 546498 581822 546734
rect 581586 510818 581822 511054
rect 581586 510498 581822 510734
rect 581586 474818 581822 475054
rect 581586 474498 581822 474734
rect 581586 438818 581822 439054
rect 581586 438498 581822 438734
rect 581586 402818 581822 403054
rect 581586 402498 581822 402734
rect 581586 366818 581822 367054
rect 581586 366498 581822 366734
rect 581586 330818 581822 331054
rect 581586 330498 581822 330734
rect 581586 294818 581822 295054
rect 581586 294498 581822 294734
rect 581586 258818 581822 259054
rect 581586 258498 581822 258734
rect 581586 222818 581822 223054
rect 581586 222498 581822 222734
rect 581586 186818 581822 187054
rect 581586 186498 581822 186734
rect 581586 150818 581822 151054
rect 581586 150498 581822 150734
rect 581586 114818 581822 115054
rect 581586 114498 581822 114734
rect 581586 78818 581822 79054
rect 581586 78498 581822 78734
rect 581586 42818 581822 43054
rect 581586 42498 581822 42734
rect 581586 6818 581822 7054
rect 581586 6498 581822 6734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 687218 585738 687454
rect 585502 686898 585738 687134
rect 585502 651218 585738 651454
rect 585502 650898 585738 651134
rect 585502 615218 585738 615454
rect 585502 614898 585738 615134
rect 585502 579218 585738 579454
rect 585502 578898 585738 579134
rect 585502 543218 585738 543454
rect 585502 542898 585738 543134
rect 585502 507218 585738 507454
rect 585502 506898 585738 507134
rect 585502 471218 585738 471454
rect 585502 470898 585738 471134
rect 585502 435218 585738 435454
rect 585502 434898 585738 435134
rect 585502 399218 585738 399454
rect 585502 398898 585738 399134
rect 585502 363218 585738 363454
rect 585502 362898 585738 363134
rect 585502 327218 585738 327454
rect 585502 326898 585738 327134
rect 585502 291218 585738 291454
rect 585502 290898 585738 291134
rect 585502 255218 585738 255454
rect 585502 254898 585738 255134
rect 585502 219218 585738 219454
rect 585502 218898 585738 219134
rect 585502 183218 585738 183454
rect 585502 182898 585738 183134
rect 585502 147218 585738 147454
rect 585502 146898 585738 147134
rect 585502 111218 585738 111454
rect 585502 110898 585738 111134
rect 585502 75218 585738 75454
rect 585502 74898 585738 75134
rect 585502 39218 585738 39454
rect 585502 38898 585738 39134
rect 585502 3218 585738 3454
rect 585502 2898 585738 3134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 669218 586678 669454
rect 586442 668898 586678 669134
rect 586442 633218 586678 633454
rect 586442 632898 586678 633134
rect 586442 597218 586678 597454
rect 586442 596898 586678 597134
rect 586442 561218 586678 561454
rect 586442 560898 586678 561134
rect 586442 525218 586678 525454
rect 586442 524898 586678 525134
rect 586442 489218 586678 489454
rect 586442 488898 586678 489134
rect 586442 453218 586678 453454
rect 586442 452898 586678 453134
rect 586442 417218 586678 417454
rect 586442 416898 586678 417134
rect 586442 381218 586678 381454
rect 586442 380898 586678 381134
rect 586442 345218 586678 345454
rect 586442 344898 586678 345134
rect 586442 309218 586678 309454
rect 586442 308898 586678 309134
rect 586442 273218 586678 273454
rect 586442 272898 586678 273134
rect 586442 237218 586678 237454
rect 586442 236898 586678 237134
rect 586442 201218 586678 201454
rect 586442 200898 586678 201134
rect 586442 165218 586678 165454
rect 586442 164898 586678 165134
rect 586442 129218 586678 129454
rect 586442 128898 586678 129134
rect 586442 93218 586678 93454
rect 586442 92898 586678 93134
rect 586442 57218 586678 57454
rect 586442 56898 586678 57134
rect 586442 21218 586678 21454
rect 586442 20898 586678 21134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 690818 587618 691054
rect 587382 690498 587618 690734
rect 587382 654818 587618 655054
rect 587382 654498 587618 654734
rect 587382 618818 587618 619054
rect 587382 618498 587618 618734
rect 587382 582818 587618 583054
rect 587382 582498 587618 582734
rect 587382 546818 587618 547054
rect 587382 546498 587618 546734
rect 587382 510818 587618 511054
rect 587382 510498 587618 510734
rect 587382 474818 587618 475054
rect 587382 474498 587618 474734
rect 587382 438818 587618 439054
rect 587382 438498 587618 438734
rect 587382 402818 587618 403054
rect 587382 402498 587618 402734
rect 587382 366818 587618 367054
rect 587382 366498 587618 366734
rect 587382 330818 587618 331054
rect 587382 330498 587618 330734
rect 587382 294818 587618 295054
rect 587382 294498 587618 294734
rect 587382 258818 587618 259054
rect 587382 258498 587618 258734
rect 587382 222818 587618 223054
rect 587382 222498 587618 222734
rect 587382 186818 587618 187054
rect 587382 186498 587618 186734
rect 587382 150818 587618 151054
rect 587382 150498 587618 150734
rect 587382 114818 587618 115054
rect 587382 114498 587618 114734
rect 587382 78818 587618 79054
rect 587382 78498 587618 78734
rect 587382 42818 587618 43054
rect 587382 42498 587618 42734
rect 587382 6818 587618 7054
rect 587382 6498 587618 6734
rect 581586 -2462 581822 -2226
rect 581586 -2782 581822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 672818 588558 673054
rect 588322 672498 588558 672734
rect 588322 636818 588558 637054
rect 588322 636498 588558 636734
rect 588322 600818 588558 601054
rect 588322 600498 588558 600734
rect 588322 564818 588558 565054
rect 588322 564498 588558 564734
rect 588322 528818 588558 529054
rect 588322 528498 588558 528734
rect 588322 492818 588558 493054
rect 588322 492498 588558 492734
rect 588322 456818 588558 457054
rect 588322 456498 588558 456734
rect 588322 420818 588558 421054
rect 588322 420498 588558 420734
rect 588322 384818 588558 385054
rect 588322 384498 588558 384734
rect 588322 348818 588558 349054
rect 588322 348498 588558 348734
rect 588322 312818 588558 313054
rect 588322 312498 588558 312734
rect 588322 276818 588558 277054
rect 588322 276498 588558 276734
rect 588322 240818 588558 241054
rect 588322 240498 588558 240734
rect 588322 204818 588558 205054
rect 588322 204498 588558 204734
rect 588322 168818 588558 169054
rect 588322 168498 588558 168734
rect 588322 132818 588558 133054
rect 588322 132498 588558 132734
rect 588322 96818 588558 97054
rect 588322 96498 588558 96734
rect 588322 60818 588558 61054
rect 588322 60498 588558 60734
rect 588322 24818 588558 25054
rect 588322 24498 588558 24734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 694418 589498 694654
rect 589262 694098 589498 694334
rect 589262 658418 589498 658654
rect 589262 658098 589498 658334
rect 589262 622418 589498 622654
rect 589262 622098 589498 622334
rect 589262 586418 589498 586654
rect 589262 586098 589498 586334
rect 589262 550418 589498 550654
rect 589262 550098 589498 550334
rect 589262 514418 589498 514654
rect 589262 514098 589498 514334
rect 589262 478418 589498 478654
rect 589262 478098 589498 478334
rect 589262 442418 589498 442654
rect 589262 442098 589498 442334
rect 589262 406418 589498 406654
rect 589262 406098 589498 406334
rect 589262 370418 589498 370654
rect 589262 370098 589498 370334
rect 589262 334418 589498 334654
rect 589262 334098 589498 334334
rect 589262 298418 589498 298654
rect 589262 298098 589498 298334
rect 589262 262418 589498 262654
rect 589262 262098 589498 262334
rect 589262 226418 589498 226654
rect 589262 226098 589498 226334
rect 589262 190418 589498 190654
rect 589262 190098 589498 190334
rect 589262 154418 589498 154654
rect 589262 154098 589498 154334
rect 589262 118418 589498 118654
rect 589262 118098 589498 118334
rect 589262 82418 589498 82654
rect 589262 82098 589498 82334
rect 589262 46418 589498 46654
rect 589262 46098 589498 46334
rect 589262 10418 589498 10654
rect 589262 10098 589498 10334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 676418 590438 676654
rect 590202 676098 590438 676334
rect 590202 640418 590438 640654
rect 590202 640098 590438 640334
rect 590202 604418 590438 604654
rect 590202 604098 590438 604334
rect 590202 568418 590438 568654
rect 590202 568098 590438 568334
rect 590202 532418 590438 532654
rect 590202 532098 590438 532334
rect 590202 496418 590438 496654
rect 590202 496098 590438 496334
rect 590202 460418 590438 460654
rect 590202 460098 590438 460334
rect 590202 424418 590438 424654
rect 590202 424098 590438 424334
rect 590202 388418 590438 388654
rect 590202 388098 590438 388334
rect 590202 352418 590438 352654
rect 590202 352098 590438 352334
rect 590202 316418 590438 316654
rect 590202 316098 590438 316334
rect 590202 280418 590438 280654
rect 590202 280098 590438 280334
rect 590202 244418 590438 244654
rect 590202 244098 590438 244334
rect 590202 208418 590438 208654
rect 590202 208098 590438 208334
rect 590202 172418 590438 172654
rect 590202 172098 590438 172334
rect 590202 136418 590438 136654
rect 590202 136098 590438 136334
rect 590202 100418 590438 100654
rect 590202 100098 590438 100334
rect 590202 64418 590438 64654
rect 590202 64098 590438 64334
rect 590202 28418 590438 28654
rect 590202 28098 590438 28334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 698018 591378 698254
rect 591142 697698 591378 697934
rect 591142 662018 591378 662254
rect 591142 661698 591378 661934
rect 591142 626018 591378 626254
rect 591142 625698 591378 625934
rect 591142 590018 591378 590254
rect 591142 589698 591378 589934
rect 591142 554018 591378 554254
rect 591142 553698 591378 553934
rect 591142 518018 591378 518254
rect 591142 517698 591378 517934
rect 591142 482018 591378 482254
rect 591142 481698 591378 481934
rect 591142 446018 591378 446254
rect 591142 445698 591378 445934
rect 591142 410018 591378 410254
rect 591142 409698 591378 409934
rect 591142 374018 591378 374254
rect 591142 373698 591378 373934
rect 591142 338018 591378 338254
rect 591142 337698 591378 337934
rect 591142 302018 591378 302254
rect 591142 301698 591378 301934
rect 591142 266018 591378 266254
rect 591142 265698 591378 265934
rect 591142 230018 591378 230254
rect 591142 229698 591378 229934
rect 591142 194018 591378 194254
rect 591142 193698 591378 193934
rect 591142 158018 591378 158254
rect 591142 157698 591378 157934
rect 591142 122018 591378 122254
rect 591142 121698 591378 121934
rect 591142 86018 591378 86254
rect 591142 85698 591378 85934
rect 591142 50018 591378 50254
rect 591142 49698 591378 49934
rect 591142 14018 591378 14254
rect 591142 13698 591378 13934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 680018 592318 680254
rect 592082 679698 592318 679934
rect 592082 644018 592318 644254
rect 592082 643698 592318 643934
rect 592082 608018 592318 608254
rect 592082 607698 592318 607934
rect 592082 572018 592318 572254
rect 592082 571698 592318 571934
rect 592082 536018 592318 536254
rect 592082 535698 592318 535934
rect 592082 500018 592318 500254
rect 592082 499698 592318 499934
rect 592082 464018 592318 464254
rect 592082 463698 592318 463934
rect 592082 428018 592318 428254
rect 592082 427698 592318 427934
rect 592082 392018 592318 392254
rect 592082 391698 592318 391934
rect 592082 356018 592318 356254
rect 592082 355698 592318 355934
rect 592082 320018 592318 320254
rect 592082 319698 592318 319934
rect 592082 284018 592318 284254
rect 592082 283698 592318 283934
rect 592082 248018 592318 248254
rect 592082 247698 592318 247934
rect 592082 212018 592318 212254
rect 592082 211698 592318 211934
rect 592082 176018 592318 176254
rect 592082 175698 592318 175934
rect 592082 140018 592318 140254
rect 592082 139698 592318 139934
rect 592082 104018 592318 104254
rect 592082 103698 592318 103934
rect 592082 68018 592318 68254
rect 592082 67698 592318 67934
rect 592082 32018 592318 32254
rect 592082 31698 592318 31934
rect 570786 -7162 571022 -6926
rect 570786 -7482 571022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 30786 711418
rect 31022 711182 66786 711418
rect 67022 711182 102786 711418
rect 103022 711182 138786 711418
rect 139022 711182 174786 711418
rect 175022 711182 210786 711418
rect 211022 711182 246786 711418
rect 247022 711182 282786 711418
rect 283022 711182 318786 711418
rect 319022 711182 354786 711418
rect 355022 711182 390786 711418
rect 391022 711182 426786 711418
rect 427022 711182 462786 711418
rect 463022 711182 498786 711418
rect 499022 711182 534786 711418
rect 535022 711182 570786 711418
rect 571022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 30786 711098
rect 31022 710862 66786 711098
rect 67022 710862 102786 711098
rect 103022 710862 138786 711098
rect 139022 710862 174786 711098
rect 175022 710862 210786 711098
rect 211022 710862 246786 711098
rect 247022 710862 282786 711098
rect 283022 710862 318786 711098
rect 319022 710862 354786 711098
rect 355022 710862 390786 711098
rect 391022 710862 426786 711098
rect 427022 710862 462786 711098
rect 463022 710862 498786 711098
rect 499022 710862 534786 711098
rect 535022 710862 570786 711098
rect 571022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 12786 710478
rect 13022 710242 48786 710478
rect 49022 710242 84786 710478
rect 85022 710242 120786 710478
rect 121022 710242 156786 710478
rect 157022 710242 192786 710478
rect 193022 710242 228786 710478
rect 229022 710242 264786 710478
rect 265022 710242 300786 710478
rect 301022 710242 336786 710478
rect 337022 710242 372786 710478
rect 373022 710242 408786 710478
rect 409022 710242 444786 710478
rect 445022 710242 480786 710478
rect 481022 710242 516786 710478
rect 517022 710242 552786 710478
rect 553022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 12786 710158
rect 13022 709922 48786 710158
rect 49022 709922 84786 710158
rect 85022 709922 120786 710158
rect 121022 709922 156786 710158
rect 157022 709922 192786 710158
rect 193022 709922 228786 710158
rect 229022 709922 264786 710158
rect 265022 709922 300786 710158
rect 301022 709922 336786 710158
rect 337022 709922 372786 710158
rect 373022 709922 408786 710158
rect 409022 709922 444786 710158
rect 445022 709922 480786 710158
rect 481022 709922 516786 710158
rect 517022 709922 552786 710158
rect 553022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 27186 709538
rect 27422 709302 63186 709538
rect 63422 709302 99186 709538
rect 99422 709302 135186 709538
rect 135422 709302 171186 709538
rect 171422 709302 207186 709538
rect 207422 709302 243186 709538
rect 243422 709302 279186 709538
rect 279422 709302 315186 709538
rect 315422 709302 351186 709538
rect 351422 709302 387186 709538
rect 387422 709302 423186 709538
rect 423422 709302 459186 709538
rect 459422 709302 495186 709538
rect 495422 709302 531186 709538
rect 531422 709302 567186 709538
rect 567422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 27186 709218
rect 27422 708982 63186 709218
rect 63422 708982 99186 709218
rect 99422 708982 135186 709218
rect 135422 708982 171186 709218
rect 171422 708982 207186 709218
rect 207422 708982 243186 709218
rect 243422 708982 279186 709218
rect 279422 708982 315186 709218
rect 315422 708982 351186 709218
rect 351422 708982 387186 709218
rect 387422 708982 423186 709218
rect 423422 708982 459186 709218
rect 459422 708982 495186 709218
rect 495422 708982 531186 709218
rect 531422 708982 567186 709218
rect 567422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 9186 708598
rect 9422 708362 45186 708598
rect 45422 708362 81186 708598
rect 81422 708362 117186 708598
rect 117422 708362 153186 708598
rect 153422 708362 189186 708598
rect 189422 708362 225186 708598
rect 225422 708362 261186 708598
rect 261422 708362 297186 708598
rect 297422 708362 333186 708598
rect 333422 708362 369186 708598
rect 369422 708362 405186 708598
rect 405422 708362 441186 708598
rect 441422 708362 477186 708598
rect 477422 708362 513186 708598
rect 513422 708362 549186 708598
rect 549422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 9186 708278
rect 9422 708042 45186 708278
rect 45422 708042 81186 708278
rect 81422 708042 117186 708278
rect 117422 708042 153186 708278
rect 153422 708042 189186 708278
rect 189422 708042 225186 708278
rect 225422 708042 261186 708278
rect 261422 708042 297186 708278
rect 297422 708042 333186 708278
rect 333422 708042 369186 708278
rect 369422 708042 405186 708278
rect 405422 708042 441186 708278
rect 441422 708042 477186 708278
rect 477422 708042 513186 708278
rect 513422 708042 549186 708278
rect 549422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 23586 707658
rect 23822 707422 59586 707658
rect 59822 707422 95586 707658
rect 95822 707422 131586 707658
rect 131822 707422 167586 707658
rect 167822 707422 203586 707658
rect 203822 707422 239586 707658
rect 239822 707422 275586 707658
rect 275822 707422 311586 707658
rect 311822 707422 347586 707658
rect 347822 707422 383586 707658
rect 383822 707422 419586 707658
rect 419822 707422 455586 707658
rect 455822 707422 491586 707658
rect 491822 707422 527586 707658
rect 527822 707422 563586 707658
rect 563822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 23586 707338
rect 23822 707102 59586 707338
rect 59822 707102 95586 707338
rect 95822 707102 131586 707338
rect 131822 707102 167586 707338
rect 167822 707102 203586 707338
rect 203822 707102 239586 707338
rect 239822 707102 275586 707338
rect 275822 707102 311586 707338
rect 311822 707102 347586 707338
rect 347822 707102 383586 707338
rect 383822 707102 419586 707338
rect 419822 707102 455586 707338
rect 455822 707102 491586 707338
rect 491822 707102 527586 707338
rect 527822 707102 563586 707338
rect 563822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 5586 706718
rect 5822 706482 41586 706718
rect 41822 706482 77586 706718
rect 77822 706482 113586 706718
rect 113822 706482 149586 706718
rect 149822 706482 185586 706718
rect 185822 706482 221586 706718
rect 221822 706482 257586 706718
rect 257822 706482 293586 706718
rect 293822 706482 329586 706718
rect 329822 706482 365586 706718
rect 365822 706482 401586 706718
rect 401822 706482 437586 706718
rect 437822 706482 473586 706718
rect 473822 706482 509586 706718
rect 509822 706482 545586 706718
rect 545822 706482 581586 706718
rect 581822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 5586 706398
rect 5822 706162 41586 706398
rect 41822 706162 77586 706398
rect 77822 706162 113586 706398
rect 113822 706162 149586 706398
rect 149822 706162 185586 706398
rect 185822 706162 221586 706398
rect 221822 706162 257586 706398
rect 257822 706162 293586 706398
rect 293822 706162 329586 706398
rect 329822 706162 365586 706398
rect 365822 706162 401586 706398
rect 401822 706162 437586 706398
rect 437822 706162 473586 706398
rect 473822 706162 509586 706398
rect 509822 706162 545586 706398
rect 545822 706162 581586 706398
rect 581822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 19986 705778
rect 20222 705542 55986 705778
rect 56222 705542 91986 705778
rect 92222 705542 127986 705778
rect 128222 705542 163986 705778
rect 164222 705542 199986 705778
rect 200222 705542 235986 705778
rect 236222 705542 271986 705778
rect 272222 705542 307986 705778
rect 308222 705542 343986 705778
rect 344222 705542 379986 705778
rect 380222 705542 415986 705778
rect 416222 705542 451986 705778
rect 452222 705542 487986 705778
rect 488222 705542 523986 705778
rect 524222 705542 559986 705778
rect 560222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 19986 705458
rect 20222 705222 55986 705458
rect 56222 705222 91986 705458
rect 92222 705222 127986 705458
rect 128222 705222 163986 705458
rect 164222 705222 199986 705458
rect 200222 705222 235986 705458
rect 236222 705222 271986 705458
rect 272222 705222 307986 705458
rect 308222 705222 343986 705458
rect 344222 705222 379986 705458
rect 380222 705222 415986 705458
rect 416222 705222 451986 705458
rect 452222 705222 487986 705458
rect 488222 705222 523986 705458
rect 524222 705222 559986 705458
rect 560222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 1986 704838
rect 2222 704602 37986 704838
rect 38222 704602 73986 704838
rect 74222 704602 109986 704838
rect 110222 704602 145986 704838
rect 146222 704602 181986 704838
rect 182222 704602 217986 704838
rect 218222 704602 253986 704838
rect 254222 704602 289986 704838
rect 290222 704602 325986 704838
rect 326222 704602 361986 704838
rect 362222 704602 397986 704838
rect 398222 704602 433986 704838
rect 434222 704602 469986 704838
rect 470222 704602 505986 704838
rect 506222 704602 541986 704838
rect 542222 704602 577986 704838
rect 578222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 1986 704518
rect 2222 704282 37986 704518
rect 38222 704282 73986 704518
rect 74222 704282 109986 704518
rect 110222 704282 145986 704518
rect 146222 704282 181986 704518
rect 182222 704282 217986 704518
rect 218222 704282 253986 704518
rect 254222 704282 289986 704518
rect 290222 704282 325986 704518
rect 326222 704282 361986 704518
rect 362222 704282 397986 704518
rect 398222 704282 433986 704518
rect 434222 704282 469986 704518
rect 470222 704282 505986 704518
rect 506222 704282 541986 704518
rect 542222 704282 577986 704518
rect 578222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect -7636 698276 -7036 698278
rect 12604 698276 13204 698278
rect 48604 698276 49204 698278
rect 84604 698276 85204 698278
rect 120604 698276 121204 698278
rect 156604 698276 157204 698278
rect 192604 698276 193204 698278
rect 228604 698276 229204 698278
rect 264604 698276 265204 698278
rect 300604 698276 301204 698278
rect 336604 698276 337204 698278
rect 372604 698276 373204 698278
rect 408604 698276 409204 698278
rect 444604 698276 445204 698278
rect 480604 698276 481204 698278
rect 516604 698276 517204 698278
rect 552604 698276 553204 698278
rect 590960 698276 591560 698278
rect -8576 698254 592500 698276
rect -8576 698018 -7454 698254
rect -7218 698018 12786 698254
rect 13022 698018 48786 698254
rect 49022 698018 84786 698254
rect 85022 698018 120786 698254
rect 121022 698018 156786 698254
rect 157022 698018 192786 698254
rect 193022 698018 228786 698254
rect 229022 698018 264786 698254
rect 265022 698018 300786 698254
rect 301022 698018 336786 698254
rect 337022 698018 372786 698254
rect 373022 698018 408786 698254
rect 409022 698018 444786 698254
rect 445022 698018 480786 698254
rect 481022 698018 516786 698254
rect 517022 698018 552786 698254
rect 553022 698018 591142 698254
rect 591378 698018 592500 698254
rect -8576 697934 592500 698018
rect -8576 697698 -7454 697934
rect -7218 697698 12786 697934
rect 13022 697698 48786 697934
rect 49022 697698 84786 697934
rect 85022 697698 120786 697934
rect 121022 697698 156786 697934
rect 157022 697698 192786 697934
rect 193022 697698 228786 697934
rect 229022 697698 264786 697934
rect 265022 697698 300786 697934
rect 301022 697698 336786 697934
rect 337022 697698 372786 697934
rect 373022 697698 408786 697934
rect 409022 697698 444786 697934
rect 445022 697698 480786 697934
rect 481022 697698 516786 697934
rect 517022 697698 552786 697934
rect 553022 697698 591142 697934
rect 591378 697698 592500 697934
rect -8576 697676 592500 697698
rect -7636 697674 -7036 697676
rect 12604 697674 13204 697676
rect 48604 697674 49204 697676
rect 84604 697674 85204 697676
rect 120604 697674 121204 697676
rect 156604 697674 157204 697676
rect 192604 697674 193204 697676
rect 228604 697674 229204 697676
rect 264604 697674 265204 697676
rect 300604 697674 301204 697676
rect 336604 697674 337204 697676
rect 372604 697674 373204 697676
rect 408604 697674 409204 697676
rect 444604 697674 445204 697676
rect 480604 697674 481204 697676
rect 516604 697674 517204 697676
rect 552604 697674 553204 697676
rect 590960 697674 591560 697676
rect -5756 694676 -5156 694678
rect 9004 694676 9604 694678
rect 45004 694676 45604 694678
rect 81004 694676 81604 694678
rect 117004 694676 117604 694678
rect 153004 694676 153604 694678
rect 189004 694676 189604 694678
rect 225004 694676 225604 694678
rect 261004 694676 261604 694678
rect 297004 694676 297604 694678
rect 333004 694676 333604 694678
rect 369004 694676 369604 694678
rect 405004 694676 405604 694678
rect 441004 694676 441604 694678
rect 477004 694676 477604 694678
rect 513004 694676 513604 694678
rect 549004 694676 549604 694678
rect 589080 694676 589680 694678
rect -6696 694654 590620 694676
rect -6696 694418 -5574 694654
rect -5338 694418 9186 694654
rect 9422 694418 45186 694654
rect 45422 694418 81186 694654
rect 81422 694418 117186 694654
rect 117422 694418 153186 694654
rect 153422 694418 189186 694654
rect 189422 694418 225186 694654
rect 225422 694418 261186 694654
rect 261422 694418 297186 694654
rect 297422 694418 333186 694654
rect 333422 694418 369186 694654
rect 369422 694418 405186 694654
rect 405422 694418 441186 694654
rect 441422 694418 477186 694654
rect 477422 694418 513186 694654
rect 513422 694418 549186 694654
rect 549422 694418 589262 694654
rect 589498 694418 590620 694654
rect -6696 694334 590620 694418
rect -6696 694098 -5574 694334
rect -5338 694098 9186 694334
rect 9422 694098 45186 694334
rect 45422 694098 81186 694334
rect 81422 694098 117186 694334
rect 117422 694098 153186 694334
rect 153422 694098 189186 694334
rect 189422 694098 225186 694334
rect 225422 694098 261186 694334
rect 261422 694098 297186 694334
rect 297422 694098 333186 694334
rect 333422 694098 369186 694334
rect 369422 694098 405186 694334
rect 405422 694098 441186 694334
rect 441422 694098 477186 694334
rect 477422 694098 513186 694334
rect 513422 694098 549186 694334
rect 549422 694098 589262 694334
rect 589498 694098 590620 694334
rect -6696 694076 590620 694098
rect -5756 694074 -5156 694076
rect 9004 694074 9604 694076
rect 45004 694074 45604 694076
rect 81004 694074 81604 694076
rect 117004 694074 117604 694076
rect 153004 694074 153604 694076
rect 189004 694074 189604 694076
rect 225004 694074 225604 694076
rect 261004 694074 261604 694076
rect 297004 694074 297604 694076
rect 333004 694074 333604 694076
rect 369004 694074 369604 694076
rect 405004 694074 405604 694076
rect 441004 694074 441604 694076
rect 477004 694074 477604 694076
rect 513004 694074 513604 694076
rect 549004 694074 549604 694076
rect 589080 694074 589680 694076
rect -3876 691076 -3276 691078
rect 5404 691076 6004 691078
rect 41404 691076 42004 691078
rect 77404 691076 78004 691078
rect 113404 691076 114004 691078
rect 149404 691076 150004 691078
rect 185404 691076 186004 691078
rect 221404 691076 222004 691078
rect 257404 691076 258004 691078
rect 293404 691076 294004 691078
rect 329404 691076 330004 691078
rect 365404 691076 366004 691078
rect 401404 691076 402004 691078
rect 437404 691076 438004 691078
rect 473404 691076 474004 691078
rect 509404 691076 510004 691078
rect 545404 691076 546004 691078
rect 581404 691076 582004 691078
rect 587200 691076 587800 691078
rect -4816 691054 588740 691076
rect -4816 690818 -3694 691054
rect -3458 690818 5586 691054
rect 5822 690818 41586 691054
rect 41822 690818 77586 691054
rect 77822 690818 113586 691054
rect 113822 690818 149586 691054
rect 149822 690818 185586 691054
rect 185822 690818 221586 691054
rect 221822 690818 257586 691054
rect 257822 690818 293586 691054
rect 293822 690818 329586 691054
rect 329822 690818 365586 691054
rect 365822 690818 401586 691054
rect 401822 690818 437586 691054
rect 437822 690818 473586 691054
rect 473822 690818 509586 691054
rect 509822 690818 545586 691054
rect 545822 690818 581586 691054
rect 581822 690818 587382 691054
rect 587618 690818 588740 691054
rect -4816 690734 588740 690818
rect -4816 690498 -3694 690734
rect -3458 690498 5586 690734
rect 5822 690498 41586 690734
rect 41822 690498 77586 690734
rect 77822 690498 113586 690734
rect 113822 690498 149586 690734
rect 149822 690498 185586 690734
rect 185822 690498 221586 690734
rect 221822 690498 257586 690734
rect 257822 690498 293586 690734
rect 293822 690498 329586 690734
rect 329822 690498 365586 690734
rect 365822 690498 401586 690734
rect 401822 690498 437586 690734
rect 437822 690498 473586 690734
rect 473822 690498 509586 690734
rect 509822 690498 545586 690734
rect 545822 690498 581586 690734
rect 581822 690498 587382 690734
rect 587618 690498 588740 690734
rect -4816 690476 588740 690498
rect -3876 690474 -3276 690476
rect 5404 690474 6004 690476
rect 41404 690474 42004 690476
rect 77404 690474 78004 690476
rect 113404 690474 114004 690476
rect 149404 690474 150004 690476
rect 185404 690474 186004 690476
rect 221404 690474 222004 690476
rect 257404 690474 258004 690476
rect 293404 690474 294004 690476
rect 329404 690474 330004 690476
rect 365404 690474 366004 690476
rect 401404 690474 402004 690476
rect 437404 690474 438004 690476
rect 473404 690474 474004 690476
rect 509404 690474 510004 690476
rect 545404 690474 546004 690476
rect 581404 690474 582004 690476
rect 587200 690474 587800 690476
rect -1996 687476 -1396 687478
rect 1804 687476 2404 687478
rect 37804 687476 38404 687478
rect 73804 687476 74404 687478
rect 109804 687476 110404 687478
rect 145804 687476 146404 687478
rect 181804 687476 182404 687478
rect 217804 687476 218404 687478
rect 253804 687476 254404 687478
rect 289804 687476 290404 687478
rect 325804 687476 326404 687478
rect 361804 687476 362404 687478
rect 397804 687476 398404 687478
rect 433804 687476 434404 687478
rect 469804 687476 470404 687478
rect 505804 687476 506404 687478
rect 541804 687476 542404 687478
rect 577804 687476 578404 687478
rect 585320 687476 585920 687478
rect -2936 687454 586860 687476
rect -2936 687218 -1814 687454
rect -1578 687218 1986 687454
rect 2222 687218 37986 687454
rect 38222 687218 73986 687454
rect 74222 687218 109986 687454
rect 110222 687218 145986 687454
rect 146222 687218 181986 687454
rect 182222 687218 217986 687454
rect 218222 687218 253986 687454
rect 254222 687218 289986 687454
rect 290222 687218 325986 687454
rect 326222 687218 361986 687454
rect 362222 687218 397986 687454
rect 398222 687218 433986 687454
rect 434222 687218 469986 687454
rect 470222 687218 505986 687454
rect 506222 687218 541986 687454
rect 542222 687218 577986 687454
rect 578222 687218 585502 687454
rect 585738 687218 586860 687454
rect -2936 687134 586860 687218
rect -2936 686898 -1814 687134
rect -1578 686898 1986 687134
rect 2222 686898 37986 687134
rect 38222 686898 73986 687134
rect 74222 686898 109986 687134
rect 110222 686898 145986 687134
rect 146222 686898 181986 687134
rect 182222 686898 217986 687134
rect 218222 686898 253986 687134
rect 254222 686898 289986 687134
rect 290222 686898 325986 687134
rect 326222 686898 361986 687134
rect 362222 686898 397986 687134
rect 398222 686898 433986 687134
rect 434222 686898 469986 687134
rect 470222 686898 505986 687134
rect 506222 686898 541986 687134
rect 542222 686898 577986 687134
rect 578222 686898 585502 687134
rect 585738 686898 586860 687134
rect -2936 686876 586860 686898
rect -1996 686874 -1396 686876
rect 1804 686874 2404 686876
rect 37804 686874 38404 686876
rect 73804 686874 74404 686876
rect 109804 686874 110404 686876
rect 145804 686874 146404 686876
rect 181804 686874 182404 686876
rect 217804 686874 218404 686876
rect 253804 686874 254404 686876
rect 289804 686874 290404 686876
rect 325804 686874 326404 686876
rect 361804 686874 362404 686876
rect 397804 686874 398404 686876
rect 433804 686874 434404 686876
rect 469804 686874 470404 686876
rect 505804 686874 506404 686876
rect 541804 686874 542404 686876
rect 577804 686874 578404 686876
rect 585320 686874 585920 686876
rect -8576 680276 -7976 680278
rect 30604 680276 31204 680278
rect 66604 680276 67204 680278
rect 102604 680276 103204 680278
rect 138604 680276 139204 680278
rect 174604 680276 175204 680278
rect 210604 680276 211204 680278
rect 246604 680276 247204 680278
rect 282604 680276 283204 680278
rect 318604 680276 319204 680278
rect 354604 680276 355204 680278
rect 390604 680276 391204 680278
rect 426604 680276 427204 680278
rect 462604 680276 463204 680278
rect 498604 680276 499204 680278
rect 534604 680276 535204 680278
rect 570604 680276 571204 680278
rect 591900 680276 592500 680278
rect -8576 680254 592500 680276
rect -8576 680018 -8394 680254
rect -8158 680018 30786 680254
rect 31022 680018 66786 680254
rect 67022 680018 102786 680254
rect 103022 680018 138786 680254
rect 139022 680018 174786 680254
rect 175022 680018 210786 680254
rect 211022 680018 246786 680254
rect 247022 680018 282786 680254
rect 283022 680018 318786 680254
rect 319022 680018 354786 680254
rect 355022 680018 390786 680254
rect 391022 680018 426786 680254
rect 427022 680018 462786 680254
rect 463022 680018 498786 680254
rect 499022 680018 534786 680254
rect 535022 680018 570786 680254
rect 571022 680018 592082 680254
rect 592318 680018 592500 680254
rect -8576 679934 592500 680018
rect -8576 679698 -8394 679934
rect -8158 679698 30786 679934
rect 31022 679698 66786 679934
rect 67022 679698 102786 679934
rect 103022 679698 138786 679934
rect 139022 679698 174786 679934
rect 175022 679698 210786 679934
rect 211022 679698 246786 679934
rect 247022 679698 282786 679934
rect 283022 679698 318786 679934
rect 319022 679698 354786 679934
rect 355022 679698 390786 679934
rect 391022 679698 426786 679934
rect 427022 679698 462786 679934
rect 463022 679698 498786 679934
rect 499022 679698 534786 679934
rect 535022 679698 570786 679934
rect 571022 679698 592082 679934
rect 592318 679698 592500 679934
rect -8576 679676 592500 679698
rect -8576 679674 -7976 679676
rect 30604 679674 31204 679676
rect 66604 679674 67204 679676
rect 102604 679674 103204 679676
rect 138604 679674 139204 679676
rect 174604 679674 175204 679676
rect 210604 679674 211204 679676
rect 246604 679674 247204 679676
rect 282604 679674 283204 679676
rect 318604 679674 319204 679676
rect 354604 679674 355204 679676
rect 390604 679674 391204 679676
rect 426604 679674 427204 679676
rect 462604 679674 463204 679676
rect 498604 679674 499204 679676
rect 534604 679674 535204 679676
rect 570604 679674 571204 679676
rect 591900 679674 592500 679676
rect -6696 676676 -6096 676678
rect 27004 676676 27604 676678
rect 63004 676676 63604 676678
rect 99004 676676 99604 676678
rect 135004 676676 135604 676678
rect 171004 676676 171604 676678
rect 207004 676676 207604 676678
rect 243004 676676 243604 676678
rect 279004 676676 279604 676678
rect 315004 676676 315604 676678
rect 351004 676676 351604 676678
rect 387004 676676 387604 676678
rect 423004 676676 423604 676678
rect 459004 676676 459604 676678
rect 495004 676676 495604 676678
rect 531004 676676 531604 676678
rect 567004 676676 567604 676678
rect 590020 676676 590620 676678
rect -6696 676654 590620 676676
rect -6696 676418 -6514 676654
rect -6278 676418 27186 676654
rect 27422 676418 63186 676654
rect 63422 676418 99186 676654
rect 99422 676418 135186 676654
rect 135422 676418 171186 676654
rect 171422 676418 207186 676654
rect 207422 676418 243186 676654
rect 243422 676418 279186 676654
rect 279422 676418 315186 676654
rect 315422 676418 351186 676654
rect 351422 676418 387186 676654
rect 387422 676418 423186 676654
rect 423422 676418 459186 676654
rect 459422 676418 495186 676654
rect 495422 676418 531186 676654
rect 531422 676418 567186 676654
rect 567422 676418 590202 676654
rect 590438 676418 590620 676654
rect -6696 676334 590620 676418
rect -6696 676098 -6514 676334
rect -6278 676098 27186 676334
rect 27422 676098 63186 676334
rect 63422 676098 99186 676334
rect 99422 676098 135186 676334
rect 135422 676098 171186 676334
rect 171422 676098 207186 676334
rect 207422 676098 243186 676334
rect 243422 676098 279186 676334
rect 279422 676098 315186 676334
rect 315422 676098 351186 676334
rect 351422 676098 387186 676334
rect 387422 676098 423186 676334
rect 423422 676098 459186 676334
rect 459422 676098 495186 676334
rect 495422 676098 531186 676334
rect 531422 676098 567186 676334
rect 567422 676098 590202 676334
rect 590438 676098 590620 676334
rect -6696 676076 590620 676098
rect -6696 676074 -6096 676076
rect 27004 676074 27604 676076
rect 63004 676074 63604 676076
rect 99004 676074 99604 676076
rect 135004 676074 135604 676076
rect 171004 676074 171604 676076
rect 207004 676074 207604 676076
rect 243004 676074 243604 676076
rect 279004 676074 279604 676076
rect 315004 676074 315604 676076
rect 351004 676074 351604 676076
rect 387004 676074 387604 676076
rect 423004 676074 423604 676076
rect 459004 676074 459604 676076
rect 495004 676074 495604 676076
rect 531004 676074 531604 676076
rect 567004 676074 567604 676076
rect 590020 676074 590620 676076
rect -4816 673076 -4216 673078
rect 23404 673076 24004 673078
rect 59404 673076 60004 673078
rect 95404 673076 96004 673078
rect 131404 673076 132004 673078
rect 167404 673076 168004 673078
rect 203404 673076 204004 673078
rect 239404 673076 240004 673078
rect 275404 673076 276004 673078
rect 311404 673076 312004 673078
rect 347404 673076 348004 673078
rect 383404 673076 384004 673078
rect 419404 673076 420004 673078
rect 455404 673076 456004 673078
rect 491404 673076 492004 673078
rect 527404 673076 528004 673078
rect 563404 673076 564004 673078
rect 588140 673076 588740 673078
rect -4816 673054 588740 673076
rect -4816 672818 -4634 673054
rect -4398 672818 23586 673054
rect 23822 672818 59586 673054
rect 59822 672818 95586 673054
rect 95822 672818 131586 673054
rect 131822 672818 167586 673054
rect 167822 672818 203586 673054
rect 203822 672818 239586 673054
rect 239822 672818 275586 673054
rect 275822 672818 311586 673054
rect 311822 672818 347586 673054
rect 347822 672818 383586 673054
rect 383822 672818 419586 673054
rect 419822 672818 455586 673054
rect 455822 672818 491586 673054
rect 491822 672818 527586 673054
rect 527822 672818 563586 673054
rect 563822 672818 588322 673054
rect 588558 672818 588740 673054
rect -4816 672734 588740 672818
rect -4816 672498 -4634 672734
rect -4398 672498 23586 672734
rect 23822 672498 59586 672734
rect 59822 672498 95586 672734
rect 95822 672498 131586 672734
rect 131822 672498 167586 672734
rect 167822 672498 203586 672734
rect 203822 672498 239586 672734
rect 239822 672498 275586 672734
rect 275822 672498 311586 672734
rect 311822 672498 347586 672734
rect 347822 672498 383586 672734
rect 383822 672498 419586 672734
rect 419822 672498 455586 672734
rect 455822 672498 491586 672734
rect 491822 672498 527586 672734
rect 527822 672498 563586 672734
rect 563822 672498 588322 672734
rect 588558 672498 588740 672734
rect -4816 672476 588740 672498
rect -4816 672474 -4216 672476
rect 23404 672474 24004 672476
rect 59404 672474 60004 672476
rect 95404 672474 96004 672476
rect 131404 672474 132004 672476
rect 167404 672474 168004 672476
rect 203404 672474 204004 672476
rect 239404 672474 240004 672476
rect 275404 672474 276004 672476
rect 311404 672474 312004 672476
rect 347404 672474 348004 672476
rect 383404 672474 384004 672476
rect 419404 672474 420004 672476
rect 455404 672474 456004 672476
rect 491404 672474 492004 672476
rect 527404 672474 528004 672476
rect 563404 672474 564004 672476
rect 588140 672474 588740 672476
rect -2936 669476 -2336 669478
rect 19804 669476 20404 669478
rect 55804 669476 56404 669478
rect 91804 669476 92404 669478
rect 127804 669476 128404 669478
rect 163804 669476 164404 669478
rect 199804 669476 200404 669478
rect 235804 669476 236404 669478
rect 271804 669476 272404 669478
rect 307804 669476 308404 669478
rect 343804 669476 344404 669478
rect 379804 669476 380404 669478
rect 415804 669476 416404 669478
rect 451804 669476 452404 669478
rect 487804 669476 488404 669478
rect 523804 669476 524404 669478
rect 559804 669476 560404 669478
rect 586260 669476 586860 669478
rect -2936 669454 586860 669476
rect -2936 669218 -2754 669454
rect -2518 669218 19986 669454
rect 20222 669218 55986 669454
rect 56222 669218 91986 669454
rect 92222 669218 127986 669454
rect 128222 669218 163986 669454
rect 164222 669218 199986 669454
rect 200222 669218 235986 669454
rect 236222 669218 271986 669454
rect 272222 669218 307986 669454
rect 308222 669218 343986 669454
rect 344222 669218 379986 669454
rect 380222 669218 415986 669454
rect 416222 669218 451986 669454
rect 452222 669218 487986 669454
rect 488222 669218 523986 669454
rect 524222 669218 559986 669454
rect 560222 669218 586442 669454
rect 586678 669218 586860 669454
rect -2936 669134 586860 669218
rect -2936 668898 -2754 669134
rect -2518 668898 19986 669134
rect 20222 668898 55986 669134
rect 56222 668898 91986 669134
rect 92222 668898 127986 669134
rect 128222 668898 163986 669134
rect 164222 668898 199986 669134
rect 200222 668898 235986 669134
rect 236222 668898 271986 669134
rect 272222 668898 307986 669134
rect 308222 668898 343986 669134
rect 344222 668898 379986 669134
rect 380222 668898 415986 669134
rect 416222 668898 451986 669134
rect 452222 668898 487986 669134
rect 488222 668898 523986 669134
rect 524222 668898 559986 669134
rect 560222 668898 586442 669134
rect 586678 668898 586860 669134
rect -2936 668876 586860 668898
rect -2936 668874 -2336 668876
rect 19804 668874 20404 668876
rect 55804 668874 56404 668876
rect 91804 668874 92404 668876
rect 127804 668874 128404 668876
rect 163804 668874 164404 668876
rect 199804 668874 200404 668876
rect 235804 668874 236404 668876
rect 271804 668874 272404 668876
rect 307804 668874 308404 668876
rect 343804 668874 344404 668876
rect 379804 668874 380404 668876
rect 415804 668874 416404 668876
rect 451804 668874 452404 668876
rect 487804 668874 488404 668876
rect 523804 668874 524404 668876
rect 559804 668874 560404 668876
rect 586260 668874 586860 668876
rect -7636 662276 -7036 662278
rect 12604 662276 13204 662278
rect 48604 662276 49204 662278
rect 84604 662276 85204 662278
rect 120604 662276 121204 662278
rect 156604 662276 157204 662278
rect 192604 662276 193204 662278
rect 228604 662276 229204 662278
rect 264604 662276 265204 662278
rect 300604 662276 301204 662278
rect 336604 662276 337204 662278
rect 372604 662276 373204 662278
rect 408604 662276 409204 662278
rect 444604 662276 445204 662278
rect 480604 662276 481204 662278
rect 516604 662276 517204 662278
rect 552604 662276 553204 662278
rect 590960 662276 591560 662278
rect -8576 662254 592500 662276
rect -8576 662018 -7454 662254
rect -7218 662018 12786 662254
rect 13022 662018 48786 662254
rect 49022 662018 84786 662254
rect 85022 662018 120786 662254
rect 121022 662018 156786 662254
rect 157022 662018 192786 662254
rect 193022 662018 228786 662254
rect 229022 662018 264786 662254
rect 265022 662018 300786 662254
rect 301022 662018 336786 662254
rect 337022 662018 372786 662254
rect 373022 662018 408786 662254
rect 409022 662018 444786 662254
rect 445022 662018 480786 662254
rect 481022 662018 516786 662254
rect 517022 662018 552786 662254
rect 553022 662018 591142 662254
rect 591378 662018 592500 662254
rect -8576 661934 592500 662018
rect -8576 661698 -7454 661934
rect -7218 661698 12786 661934
rect 13022 661698 48786 661934
rect 49022 661698 84786 661934
rect 85022 661698 120786 661934
rect 121022 661698 156786 661934
rect 157022 661698 192786 661934
rect 193022 661698 228786 661934
rect 229022 661698 264786 661934
rect 265022 661698 300786 661934
rect 301022 661698 336786 661934
rect 337022 661698 372786 661934
rect 373022 661698 408786 661934
rect 409022 661698 444786 661934
rect 445022 661698 480786 661934
rect 481022 661698 516786 661934
rect 517022 661698 552786 661934
rect 553022 661698 591142 661934
rect 591378 661698 592500 661934
rect -8576 661676 592500 661698
rect -7636 661674 -7036 661676
rect 12604 661674 13204 661676
rect 48604 661674 49204 661676
rect 84604 661674 85204 661676
rect 120604 661674 121204 661676
rect 156604 661674 157204 661676
rect 192604 661674 193204 661676
rect 228604 661674 229204 661676
rect 264604 661674 265204 661676
rect 300604 661674 301204 661676
rect 336604 661674 337204 661676
rect 372604 661674 373204 661676
rect 408604 661674 409204 661676
rect 444604 661674 445204 661676
rect 480604 661674 481204 661676
rect 516604 661674 517204 661676
rect 552604 661674 553204 661676
rect 590960 661674 591560 661676
rect -5756 658676 -5156 658678
rect 9004 658676 9604 658678
rect 45004 658676 45604 658678
rect 81004 658676 81604 658678
rect 117004 658676 117604 658678
rect 153004 658676 153604 658678
rect 189004 658676 189604 658678
rect 225004 658676 225604 658678
rect 261004 658676 261604 658678
rect 297004 658676 297604 658678
rect 333004 658676 333604 658678
rect 369004 658676 369604 658678
rect 405004 658676 405604 658678
rect 441004 658676 441604 658678
rect 477004 658676 477604 658678
rect 513004 658676 513604 658678
rect 549004 658676 549604 658678
rect 589080 658676 589680 658678
rect -6696 658654 590620 658676
rect -6696 658418 -5574 658654
rect -5338 658418 9186 658654
rect 9422 658418 45186 658654
rect 45422 658418 81186 658654
rect 81422 658418 117186 658654
rect 117422 658418 153186 658654
rect 153422 658418 189186 658654
rect 189422 658418 225186 658654
rect 225422 658418 261186 658654
rect 261422 658418 297186 658654
rect 297422 658418 333186 658654
rect 333422 658418 369186 658654
rect 369422 658418 405186 658654
rect 405422 658418 441186 658654
rect 441422 658418 477186 658654
rect 477422 658418 513186 658654
rect 513422 658418 549186 658654
rect 549422 658418 589262 658654
rect 589498 658418 590620 658654
rect -6696 658334 590620 658418
rect -6696 658098 -5574 658334
rect -5338 658098 9186 658334
rect 9422 658098 45186 658334
rect 45422 658098 81186 658334
rect 81422 658098 117186 658334
rect 117422 658098 153186 658334
rect 153422 658098 189186 658334
rect 189422 658098 225186 658334
rect 225422 658098 261186 658334
rect 261422 658098 297186 658334
rect 297422 658098 333186 658334
rect 333422 658098 369186 658334
rect 369422 658098 405186 658334
rect 405422 658098 441186 658334
rect 441422 658098 477186 658334
rect 477422 658098 513186 658334
rect 513422 658098 549186 658334
rect 549422 658098 589262 658334
rect 589498 658098 590620 658334
rect -6696 658076 590620 658098
rect -5756 658074 -5156 658076
rect 9004 658074 9604 658076
rect 45004 658074 45604 658076
rect 81004 658074 81604 658076
rect 117004 658074 117604 658076
rect 153004 658074 153604 658076
rect 189004 658074 189604 658076
rect 225004 658074 225604 658076
rect 261004 658074 261604 658076
rect 297004 658074 297604 658076
rect 333004 658074 333604 658076
rect 369004 658074 369604 658076
rect 405004 658074 405604 658076
rect 441004 658074 441604 658076
rect 477004 658074 477604 658076
rect 513004 658074 513604 658076
rect 549004 658074 549604 658076
rect 589080 658074 589680 658076
rect -3876 655076 -3276 655078
rect 5404 655076 6004 655078
rect 41404 655076 42004 655078
rect 77404 655076 78004 655078
rect 113404 655076 114004 655078
rect 149404 655076 150004 655078
rect 185404 655076 186004 655078
rect 221404 655076 222004 655078
rect 257404 655076 258004 655078
rect 293404 655076 294004 655078
rect 329404 655076 330004 655078
rect 365404 655076 366004 655078
rect 401404 655076 402004 655078
rect 437404 655076 438004 655078
rect 473404 655076 474004 655078
rect 509404 655076 510004 655078
rect 545404 655076 546004 655078
rect 581404 655076 582004 655078
rect 587200 655076 587800 655078
rect -4816 655054 588740 655076
rect -4816 654818 -3694 655054
rect -3458 654818 5586 655054
rect 5822 654818 41586 655054
rect 41822 654818 77586 655054
rect 77822 654818 113586 655054
rect 113822 654818 149586 655054
rect 149822 654818 185586 655054
rect 185822 654818 221586 655054
rect 221822 654818 257586 655054
rect 257822 654818 293586 655054
rect 293822 654818 329586 655054
rect 329822 654818 365586 655054
rect 365822 654818 401586 655054
rect 401822 654818 437586 655054
rect 437822 654818 473586 655054
rect 473822 654818 509586 655054
rect 509822 654818 545586 655054
rect 545822 654818 581586 655054
rect 581822 654818 587382 655054
rect 587618 654818 588740 655054
rect -4816 654734 588740 654818
rect -4816 654498 -3694 654734
rect -3458 654498 5586 654734
rect 5822 654498 41586 654734
rect 41822 654498 77586 654734
rect 77822 654498 113586 654734
rect 113822 654498 149586 654734
rect 149822 654498 185586 654734
rect 185822 654498 221586 654734
rect 221822 654498 257586 654734
rect 257822 654498 293586 654734
rect 293822 654498 329586 654734
rect 329822 654498 365586 654734
rect 365822 654498 401586 654734
rect 401822 654498 437586 654734
rect 437822 654498 473586 654734
rect 473822 654498 509586 654734
rect 509822 654498 545586 654734
rect 545822 654498 581586 654734
rect 581822 654498 587382 654734
rect 587618 654498 588740 654734
rect -4816 654476 588740 654498
rect -3876 654474 -3276 654476
rect 5404 654474 6004 654476
rect 41404 654474 42004 654476
rect 77404 654474 78004 654476
rect 113404 654474 114004 654476
rect 149404 654474 150004 654476
rect 185404 654474 186004 654476
rect 221404 654474 222004 654476
rect 257404 654474 258004 654476
rect 293404 654474 294004 654476
rect 329404 654474 330004 654476
rect 365404 654474 366004 654476
rect 401404 654474 402004 654476
rect 437404 654474 438004 654476
rect 473404 654474 474004 654476
rect 509404 654474 510004 654476
rect 545404 654474 546004 654476
rect 581404 654474 582004 654476
rect 587200 654474 587800 654476
rect -1996 651476 -1396 651478
rect 1804 651476 2404 651478
rect 37804 651476 38404 651478
rect 73804 651476 74404 651478
rect 109804 651476 110404 651478
rect 145804 651476 146404 651478
rect 181804 651476 182404 651478
rect 217804 651476 218404 651478
rect 253804 651476 254404 651478
rect 289804 651476 290404 651478
rect 325804 651476 326404 651478
rect 361804 651476 362404 651478
rect 397804 651476 398404 651478
rect 433804 651476 434404 651478
rect 469804 651476 470404 651478
rect 505804 651476 506404 651478
rect 541804 651476 542404 651478
rect 577804 651476 578404 651478
rect 585320 651476 585920 651478
rect -2936 651454 586860 651476
rect -2936 651218 -1814 651454
rect -1578 651218 1986 651454
rect 2222 651218 37986 651454
rect 38222 651218 73986 651454
rect 74222 651218 109986 651454
rect 110222 651218 145986 651454
rect 146222 651218 181986 651454
rect 182222 651218 217986 651454
rect 218222 651218 253986 651454
rect 254222 651218 289986 651454
rect 290222 651218 325986 651454
rect 326222 651218 361986 651454
rect 362222 651218 397986 651454
rect 398222 651218 433986 651454
rect 434222 651218 469986 651454
rect 470222 651218 505986 651454
rect 506222 651218 541986 651454
rect 542222 651218 577986 651454
rect 578222 651218 585502 651454
rect 585738 651218 586860 651454
rect -2936 651134 586860 651218
rect -2936 650898 -1814 651134
rect -1578 650898 1986 651134
rect 2222 650898 37986 651134
rect 38222 650898 73986 651134
rect 74222 650898 109986 651134
rect 110222 650898 145986 651134
rect 146222 650898 181986 651134
rect 182222 650898 217986 651134
rect 218222 650898 253986 651134
rect 254222 650898 289986 651134
rect 290222 650898 325986 651134
rect 326222 650898 361986 651134
rect 362222 650898 397986 651134
rect 398222 650898 433986 651134
rect 434222 650898 469986 651134
rect 470222 650898 505986 651134
rect 506222 650898 541986 651134
rect 542222 650898 577986 651134
rect 578222 650898 585502 651134
rect 585738 650898 586860 651134
rect -2936 650876 586860 650898
rect -1996 650874 -1396 650876
rect 1804 650874 2404 650876
rect 37804 650874 38404 650876
rect 73804 650874 74404 650876
rect 109804 650874 110404 650876
rect 145804 650874 146404 650876
rect 181804 650874 182404 650876
rect 217804 650874 218404 650876
rect 253804 650874 254404 650876
rect 289804 650874 290404 650876
rect 325804 650874 326404 650876
rect 361804 650874 362404 650876
rect 397804 650874 398404 650876
rect 433804 650874 434404 650876
rect 469804 650874 470404 650876
rect 505804 650874 506404 650876
rect 541804 650874 542404 650876
rect 577804 650874 578404 650876
rect 585320 650874 585920 650876
rect -8576 644276 -7976 644278
rect 30604 644276 31204 644278
rect 66604 644276 67204 644278
rect 102604 644276 103204 644278
rect 138604 644276 139204 644278
rect 174604 644276 175204 644278
rect 210604 644276 211204 644278
rect 246604 644276 247204 644278
rect 282604 644276 283204 644278
rect 318604 644276 319204 644278
rect 354604 644276 355204 644278
rect 390604 644276 391204 644278
rect 426604 644276 427204 644278
rect 462604 644276 463204 644278
rect 498604 644276 499204 644278
rect 534604 644276 535204 644278
rect 570604 644276 571204 644278
rect 591900 644276 592500 644278
rect -8576 644254 592500 644276
rect -8576 644018 -8394 644254
rect -8158 644018 30786 644254
rect 31022 644018 66786 644254
rect 67022 644018 102786 644254
rect 103022 644018 138786 644254
rect 139022 644018 174786 644254
rect 175022 644018 210786 644254
rect 211022 644018 246786 644254
rect 247022 644018 282786 644254
rect 283022 644018 318786 644254
rect 319022 644018 354786 644254
rect 355022 644018 390786 644254
rect 391022 644018 426786 644254
rect 427022 644018 462786 644254
rect 463022 644018 498786 644254
rect 499022 644018 534786 644254
rect 535022 644018 570786 644254
rect 571022 644018 592082 644254
rect 592318 644018 592500 644254
rect -8576 643934 592500 644018
rect -8576 643698 -8394 643934
rect -8158 643698 30786 643934
rect 31022 643698 66786 643934
rect 67022 643698 102786 643934
rect 103022 643698 138786 643934
rect 139022 643698 174786 643934
rect 175022 643698 210786 643934
rect 211022 643698 246786 643934
rect 247022 643698 282786 643934
rect 283022 643698 318786 643934
rect 319022 643698 354786 643934
rect 355022 643698 390786 643934
rect 391022 643698 426786 643934
rect 427022 643698 462786 643934
rect 463022 643698 498786 643934
rect 499022 643698 534786 643934
rect 535022 643698 570786 643934
rect 571022 643698 592082 643934
rect 592318 643698 592500 643934
rect -8576 643676 592500 643698
rect -8576 643674 -7976 643676
rect 30604 643674 31204 643676
rect 66604 643674 67204 643676
rect 102604 643674 103204 643676
rect 138604 643674 139204 643676
rect 174604 643674 175204 643676
rect 210604 643674 211204 643676
rect 246604 643674 247204 643676
rect 282604 643674 283204 643676
rect 318604 643674 319204 643676
rect 354604 643674 355204 643676
rect 390604 643674 391204 643676
rect 426604 643674 427204 643676
rect 462604 643674 463204 643676
rect 498604 643674 499204 643676
rect 534604 643674 535204 643676
rect 570604 643674 571204 643676
rect 591900 643674 592500 643676
rect -6696 640676 -6096 640678
rect 27004 640676 27604 640678
rect 63004 640676 63604 640678
rect 99004 640676 99604 640678
rect 135004 640676 135604 640678
rect 171004 640676 171604 640678
rect 207004 640676 207604 640678
rect 243004 640676 243604 640678
rect 279004 640676 279604 640678
rect 315004 640676 315604 640678
rect 351004 640676 351604 640678
rect 387004 640676 387604 640678
rect 423004 640676 423604 640678
rect 459004 640676 459604 640678
rect 495004 640676 495604 640678
rect 531004 640676 531604 640678
rect 567004 640676 567604 640678
rect 590020 640676 590620 640678
rect -6696 640654 590620 640676
rect -6696 640418 -6514 640654
rect -6278 640418 27186 640654
rect 27422 640418 63186 640654
rect 63422 640418 99186 640654
rect 99422 640418 135186 640654
rect 135422 640418 171186 640654
rect 171422 640418 207186 640654
rect 207422 640418 243186 640654
rect 243422 640418 279186 640654
rect 279422 640418 315186 640654
rect 315422 640418 351186 640654
rect 351422 640418 387186 640654
rect 387422 640418 423186 640654
rect 423422 640418 459186 640654
rect 459422 640418 495186 640654
rect 495422 640418 531186 640654
rect 531422 640418 567186 640654
rect 567422 640418 590202 640654
rect 590438 640418 590620 640654
rect -6696 640334 590620 640418
rect -6696 640098 -6514 640334
rect -6278 640098 27186 640334
rect 27422 640098 63186 640334
rect 63422 640098 99186 640334
rect 99422 640098 135186 640334
rect 135422 640098 171186 640334
rect 171422 640098 207186 640334
rect 207422 640098 243186 640334
rect 243422 640098 279186 640334
rect 279422 640098 315186 640334
rect 315422 640098 351186 640334
rect 351422 640098 387186 640334
rect 387422 640098 423186 640334
rect 423422 640098 459186 640334
rect 459422 640098 495186 640334
rect 495422 640098 531186 640334
rect 531422 640098 567186 640334
rect 567422 640098 590202 640334
rect 590438 640098 590620 640334
rect -6696 640076 590620 640098
rect -6696 640074 -6096 640076
rect 27004 640074 27604 640076
rect 63004 640074 63604 640076
rect 99004 640074 99604 640076
rect 135004 640074 135604 640076
rect 171004 640074 171604 640076
rect 207004 640074 207604 640076
rect 243004 640074 243604 640076
rect 279004 640074 279604 640076
rect 315004 640074 315604 640076
rect 351004 640074 351604 640076
rect 387004 640074 387604 640076
rect 423004 640074 423604 640076
rect 459004 640074 459604 640076
rect 495004 640074 495604 640076
rect 531004 640074 531604 640076
rect 567004 640074 567604 640076
rect 590020 640074 590620 640076
rect -4816 637076 -4216 637078
rect 23404 637076 24004 637078
rect 59404 637076 60004 637078
rect 95404 637076 96004 637078
rect 131404 637076 132004 637078
rect 167404 637076 168004 637078
rect 203404 637076 204004 637078
rect 239404 637076 240004 637078
rect 275404 637076 276004 637078
rect 311404 637076 312004 637078
rect 347404 637076 348004 637078
rect 383404 637076 384004 637078
rect 419404 637076 420004 637078
rect 455404 637076 456004 637078
rect 491404 637076 492004 637078
rect 527404 637076 528004 637078
rect 563404 637076 564004 637078
rect 588140 637076 588740 637078
rect -4816 637054 588740 637076
rect -4816 636818 -4634 637054
rect -4398 636818 23586 637054
rect 23822 636818 59586 637054
rect 59822 636818 95586 637054
rect 95822 636818 131586 637054
rect 131822 636818 167586 637054
rect 167822 636818 203586 637054
rect 203822 636818 239586 637054
rect 239822 636818 275586 637054
rect 275822 636818 311586 637054
rect 311822 636818 347586 637054
rect 347822 636818 383586 637054
rect 383822 636818 419586 637054
rect 419822 636818 455586 637054
rect 455822 636818 491586 637054
rect 491822 636818 527586 637054
rect 527822 636818 563586 637054
rect 563822 636818 588322 637054
rect 588558 636818 588740 637054
rect -4816 636734 588740 636818
rect -4816 636498 -4634 636734
rect -4398 636498 23586 636734
rect 23822 636498 59586 636734
rect 59822 636498 95586 636734
rect 95822 636498 131586 636734
rect 131822 636498 167586 636734
rect 167822 636498 203586 636734
rect 203822 636498 239586 636734
rect 239822 636498 275586 636734
rect 275822 636498 311586 636734
rect 311822 636498 347586 636734
rect 347822 636498 383586 636734
rect 383822 636498 419586 636734
rect 419822 636498 455586 636734
rect 455822 636498 491586 636734
rect 491822 636498 527586 636734
rect 527822 636498 563586 636734
rect 563822 636498 588322 636734
rect 588558 636498 588740 636734
rect -4816 636476 588740 636498
rect -4816 636474 -4216 636476
rect 23404 636474 24004 636476
rect 59404 636474 60004 636476
rect 95404 636474 96004 636476
rect 131404 636474 132004 636476
rect 167404 636474 168004 636476
rect 203404 636474 204004 636476
rect 239404 636474 240004 636476
rect 275404 636474 276004 636476
rect 311404 636474 312004 636476
rect 347404 636474 348004 636476
rect 383404 636474 384004 636476
rect 419404 636474 420004 636476
rect 455404 636474 456004 636476
rect 491404 636474 492004 636476
rect 527404 636474 528004 636476
rect 563404 636474 564004 636476
rect 588140 636474 588740 636476
rect -2936 633476 -2336 633478
rect 19804 633476 20404 633478
rect 55804 633476 56404 633478
rect 91804 633476 92404 633478
rect 127804 633476 128404 633478
rect 163804 633476 164404 633478
rect 199804 633476 200404 633478
rect 235804 633476 236404 633478
rect 271804 633476 272404 633478
rect 307804 633476 308404 633478
rect 343804 633476 344404 633478
rect 379804 633476 380404 633478
rect 415804 633476 416404 633478
rect 451804 633476 452404 633478
rect 487804 633476 488404 633478
rect 523804 633476 524404 633478
rect 559804 633476 560404 633478
rect 586260 633476 586860 633478
rect -2936 633454 586860 633476
rect -2936 633218 -2754 633454
rect -2518 633218 19986 633454
rect 20222 633218 55986 633454
rect 56222 633218 91986 633454
rect 92222 633218 127986 633454
rect 128222 633218 163986 633454
rect 164222 633218 199986 633454
rect 200222 633218 235986 633454
rect 236222 633218 271986 633454
rect 272222 633218 307986 633454
rect 308222 633218 343986 633454
rect 344222 633218 379986 633454
rect 380222 633218 415986 633454
rect 416222 633218 451986 633454
rect 452222 633218 487986 633454
rect 488222 633218 523986 633454
rect 524222 633218 559986 633454
rect 560222 633218 586442 633454
rect 586678 633218 586860 633454
rect -2936 633134 586860 633218
rect -2936 632898 -2754 633134
rect -2518 632898 19986 633134
rect 20222 632898 55986 633134
rect 56222 632898 91986 633134
rect 92222 632898 127986 633134
rect 128222 632898 163986 633134
rect 164222 632898 199986 633134
rect 200222 632898 235986 633134
rect 236222 632898 271986 633134
rect 272222 632898 307986 633134
rect 308222 632898 343986 633134
rect 344222 632898 379986 633134
rect 380222 632898 415986 633134
rect 416222 632898 451986 633134
rect 452222 632898 487986 633134
rect 488222 632898 523986 633134
rect 524222 632898 559986 633134
rect 560222 632898 586442 633134
rect 586678 632898 586860 633134
rect -2936 632876 586860 632898
rect -2936 632874 -2336 632876
rect 19804 632874 20404 632876
rect 55804 632874 56404 632876
rect 91804 632874 92404 632876
rect 127804 632874 128404 632876
rect 163804 632874 164404 632876
rect 199804 632874 200404 632876
rect 235804 632874 236404 632876
rect 271804 632874 272404 632876
rect 307804 632874 308404 632876
rect 343804 632874 344404 632876
rect 379804 632874 380404 632876
rect 415804 632874 416404 632876
rect 451804 632874 452404 632876
rect 487804 632874 488404 632876
rect 523804 632874 524404 632876
rect 559804 632874 560404 632876
rect 586260 632874 586860 632876
rect -7636 626276 -7036 626278
rect 12604 626276 13204 626278
rect 48604 626276 49204 626278
rect 84604 626276 85204 626278
rect 120604 626276 121204 626278
rect 156604 626276 157204 626278
rect 192604 626276 193204 626278
rect 228604 626276 229204 626278
rect 264604 626276 265204 626278
rect 300604 626276 301204 626278
rect 336604 626276 337204 626278
rect 372604 626276 373204 626278
rect 408604 626276 409204 626278
rect 444604 626276 445204 626278
rect 480604 626276 481204 626278
rect 516604 626276 517204 626278
rect 552604 626276 553204 626278
rect 590960 626276 591560 626278
rect -8576 626254 592500 626276
rect -8576 626018 -7454 626254
rect -7218 626018 12786 626254
rect 13022 626018 48786 626254
rect 49022 626018 84786 626254
rect 85022 626018 120786 626254
rect 121022 626018 156786 626254
rect 157022 626018 192786 626254
rect 193022 626018 228786 626254
rect 229022 626018 264786 626254
rect 265022 626018 300786 626254
rect 301022 626018 336786 626254
rect 337022 626018 372786 626254
rect 373022 626018 408786 626254
rect 409022 626018 444786 626254
rect 445022 626018 480786 626254
rect 481022 626018 516786 626254
rect 517022 626018 552786 626254
rect 553022 626018 591142 626254
rect 591378 626018 592500 626254
rect -8576 625934 592500 626018
rect -8576 625698 -7454 625934
rect -7218 625698 12786 625934
rect 13022 625698 48786 625934
rect 49022 625698 84786 625934
rect 85022 625698 120786 625934
rect 121022 625698 156786 625934
rect 157022 625698 192786 625934
rect 193022 625698 228786 625934
rect 229022 625698 264786 625934
rect 265022 625698 300786 625934
rect 301022 625698 336786 625934
rect 337022 625698 372786 625934
rect 373022 625698 408786 625934
rect 409022 625698 444786 625934
rect 445022 625698 480786 625934
rect 481022 625698 516786 625934
rect 517022 625698 552786 625934
rect 553022 625698 591142 625934
rect 591378 625698 592500 625934
rect -8576 625676 592500 625698
rect -7636 625674 -7036 625676
rect 12604 625674 13204 625676
rect 48604 625674 49204 625676
rect 84604 625674 85204 625676
rect 120604 625674 121204 625676
rect 156604 625674 157204 625676
rect 192604 625674 193204 625676
rect 228604 625674 229204 625676
rect 264604 625674 265204 625676
rect 300604 625674 301204 625676
rect 336604 625674 337204 625676
rect 372604 625674 373204 625676
rect 408604 625674 409204 625676
rect 444604 625674 445204 625676
rect 480604 625674 481204 625676
rect 516604 625674 517204 625676
rect 552604 625674 553204 625676
rect 590960 625674 591560 625676
rect -5756 622676 -5156 622678
rect 9004 622676 9604 622678
rect 45004 622676 45604 622678
rect 81004 622676 81604 622678
rect 117004 622676 117604 622678
rect 153004 622676 153604 622678
rect 189004 622676 189604 622678
rect 225004 622676 225604 622678
rect 261004 622676 261604 622678
rect 297004 622676 297604 622678
rect 333004 622676 333604 622678
rect 369004 622676 369604 622678
rect 405004 622676 405604 622678
rect 441004 622676 441604 622678
rect 477004 622676 477604 622678
rect 513004 622676 513604 622678
rect 549004 622676 549604 622678
rect 589080 622676 589680 622678
rect -6696 622654 590620 622676
rect -6696 622418 -5574 622654
rect -5338 622418 9186 622654
rect 9422 622418 45186 622654
rect 45422 622418 81186 622654
rect 81422 622418 117186 622654
rect 117422 622418 153186 622654
rect 153422 622418 189186 622654
rect 189422 622418 225186 622654
rect 225422 622418 261186 622654
rect 261422 622418 297186 622654
rect 297422 622418 333186 622654
rect 333422 622418 369186 622654
rect 369422 622418 405186 622654
rect 405422 622418 441186 622654
rect 441422 622418 477186 622654
rect 477422 622418 513186 622654
rect 513422 622418 549186 622654
rect 549422 622418 589262 622654
rect 589498 622418 590620 622654
rect -6696 622334 590620 622418
rect -6696 622098 -5574 622334
rect -5338 622098 9186 622334
rect 9422 622098 45186 622334
rect 45422 622098 81186 622334
rect 81422 622098 117186 622334
rect 117422 622098 153186 622334
rect 153422 622098 189186 622334
rect 189422 622098 225186 622334
rect 225422 622098 261186 622334
rect 261422 622098 297186 622334
rect 297422 622098 333186 622334
rect 333422 622098 369186 622334
rect 369422 622098 405186 622334
rect 405422 622098 441186 622334
rect 441422 622098 477186 622334
rect 477422 622098 513186 622334
rect 513422 622098 549186 622334
rect 549422 622098 589262 622334
rect 589498 622098 590620 622334
rect -6696 622076 590620 622098
rect -5756 622074 -5156 622076
rect 9004 622074 9604 622076
rect 45004 622074 45604 622076
rect 81004 622074 81604 622076
rect 117004 622074 117604 622076
rect 153004 622074 153604 622076
rect 189004 622074 189604 622076
rect 225004 622074 225604 622076
rect 261004 622074 261604 622076
rect 297004 622074 297604 622076
rect 333004 622074 333604 622076
rect 369004 622074 369604 622076
rect 405004 622074 405604 622076
rect 441004 622074 441604 622076
rect 477004 622074 477604 622076
rect 513004 622074 513604 622076
rect 549004 622074 549604 622076
rect 589080 622074 589680 622076
rect -3876 619076 -3276 619078
rect 5404 619076 6004 619078
rect 41404 619076 42004 619078
rect 77404 619076 78004 619078
rect 113404 619076 114004 619078
rect 149404 619076 150004 619078
rect 185404 619076 186004 619078
rect 221404 619076 222004 619078
rect 257404 619076 258004 619078
rect 293404 619076 294004 619078
rect 329404 619076 330004 619078
rect 365404 619076 366004 619078
rect 401404 619076 402004 619078
rect 437404 619076 438004 619078
rect 473404 619076 474004 619078
rect 509404 619076 510004 619078
rect 545404 619076 546004 619078
rect 581404 619076 582004 619078
rect 587200 619076 587800 619078
rect -4816 619054 588740 619076
rect -4816 618818 -3694 619054
rect -3458 618818 5586 619054
rect 5822 618818 41586 619054
rect 41822 618818 77586 619054
rect 77822 618818 113586 619054
rect 113822 618818 149586 619054
rect 149822 618818 185586 619054
rect 185822 618818 221586 619054
rect 221822 618818 257586 619054
rect 257822 618818 293586 619054
rect 293822 618818 329586 619054
rect 329822 618818 365586 619054
rect 365822 618818 401586 619054
rect 401822 618818 437586 619054
rect 437822 618818 473586 619054
rect 473822 618818 509586 619054
rect 509822 618818 545586 619054
rect 545822 618818 581586 619054
rect 581822 618818 587382 619054
rect 587618 618818 588740 619054
rect -4816 618734 588740 618818
rect -4816 618498 -3694 618734
rect -3458 618498 5586 618734
rect 5822 618498 41586 618734
rect 41822 618498 77586 618734
rect 77822 618498 113586 618734
rect 113822 618498 149586 618734
rect 149822 618498 185586 618734
rect 185822 618498 221586 618734
rect 221822 618498 257586 618734
rect 257822 618498 293586 618734
rect 293822 618498 329586 618734
rect 329822 618498 365586 618734
rect 365822 618498 401586 618734
rect 401822 618498 437586 618734
rect 437822 618498 473586 618734
rect 473822 618498 509586 618734
rect 509822 618498 545586 618734
rect 545822 618498 581586 618734
rect 581822 618498 587382 618734
rect 587618 618498 588740 618734
rect -4816 618476 588740 618498
rect -3876 618474 -3276 618476
rect 5404 618474 6004 618476
rect 41404 618474 42004 618476
rect 77404 618474 78004 618476
rect 113404 618474 114004 618476
rect 149404 618474 150004 618476
rect 185404 618474 186004 618476
rect 221404 618474 222004 618476
rect 257404 618474 258004 618476
rect 293404 618474 294004 618476
rect 329404 618474 330004 618476
rect 365404 618474 366004 618476
rect 401404 618474 402004 618476
rect 437404 618474 438004 618476
rect 473404 618474 474004 618476
rect 509404 618474 510004 618476
rect 545404 618474 546004 618476
rect 581404 618474 582004 618476
rect 587200 618474 587800 618476
rect -1996 615476 -1396 615478
rect 1804 615476 2404 615478
rect 37804 615476 38404 615478
rect 73804 615476 74404 615478
rect 109804 615476 110404 615478
rect 145804 615476 146404 615478
rect 181804 615476 182404 615478
rect 217804 615476 218404 615478
rect 253804 615476 254404 615478
rect 289804 615476 290404 615478
rect 325804 615476 326404 615478
rect 361804 615476 362404 615478
rect 397804 615476 398404 615478
rect 433804 615476 434404 615478
rect 469804 615476 470404 615478
rect 505804 615476 506404 615478
rect 541804 615476 542404 615478
rect 577804 615476 578404 615478
rect 585320 615476 585920 615478
rect -2936 615454 586860 615476
rect -2936 615218 -1814 615454
rect -1578 615218 1986 615454
rect 2222 615218 37986 615454
rect 38222 615218 73986 615454
rect 74222 615218 109986 615454
rect 110222 615218 145986 615454
rect 146222 615218 181986 615454
rect 182222 615218 217986 615454
rect 218222 615218 253986 615454
rect 254222 615218 289986 615454
rect 290222 615218 325986 615454
rect 326222 615218 361986 615454
rect 362222 615218 397986 615454
rect 398222 615218 433986 615454
rect 434222 615218 469986 615454
rect 470222 615218 505986 615454
rect 506222 615218 541986 615454
rect 542222 615218 577986 615454
rect 578222 615218 585502 615454
rect 585738 615218 586860 615454
rect -2936 615134 586860 615218
rect -2936 614898 -1814 615134
rect -1578 614898 1986 615134
rect 2222 614898 37986 615134
rect 38222 614898 73986 615134
rect 74222 614898 109986 615134
rect 110222 614898 145986 615134
rect 146222 614898 181986 615134
rect 182222 614898 217986 615134
rect 218222 614898 253986 615134
rect 254222 614898 289986 615134
rect 290222 614898 325986 615134
rect 326222 614898 361986 615134
rect 362222 614898 397986 615134
rect 398222 614898 433986 615134
rect 434222 614898 469986 615134
rect 470222 614898 505986 615134
rect 506222 614898 541986 615134
rect 542222 614898 577986 615134
rect 578222 614898 585502 615134
rect 585738 614898 586860 615134
rect -2936 614876 586860 614898
rect -1996 614874 -1396 614876
rect 1804 614874 2404 614876
rect 37804 614874 38404 614876
rect 73804 614874 74404 614876
rect 109804 614874 110404 614876
rect 145804 614874 146404 614876
rect 181804 614874 182404 614876
rect 217804 614874 218404 614876
rect 253804 614874 254404 614876
rect 289804 614874 290404 614876
rect 325804 614874 326404 614876
rect 361804 614874 362404 614876
rect 397804 614874 398404 614876
rect 433804 614874 434404 614876
rect 469804 614874 470404 614876
rect 505804 614874 506404 614876
rect 541804 614874 542404 614876
rect 577804 614874 578404 614876
rect 585320 614874 585920 614876
rect -8576 608276 -7976 608278
rect 30604 608276 31204 608278
rect 66604 608276 67204 608278
rect 102604 608276 103204 608278
rect 138604 608276 139204 608278
rect 174604 608276 175204 608278
rect 210604 608276 211204 608278
rect 246604 608276 247204 608278
rect 282604 608276 283204 608278
rect 318604 608276 319204 608278
rect 354604 608276 355204 608278
rect 390604 608276 391204 608278
rect 426604 608276 427204 608278
rect 462604 608276 463204 608278
rect 498604 608276 499204 608278
rect 534604 608276 535204 608278
rect 570604 608276 571204 608278
rect 591900 608276 592500 608278
rect -8576 608254 592500 608276
rect -8576 608018 -8394 608254
rect -8158 608018 30786 608254
rect 31022 608018 66786 608254
rect 67022 608018 102786 608254
rect 103022 608018 138786 608254
rect 139022 608018 174786 608254
rect 175022 608018 210786 608254
rect 211022 608018 246786 608254
rect 247022 608018 282786 608254
rect 283022 608018 318786 608254
rect 319022 608018 354786 608254
rect 355022 608018 390786 608254
rect 391022 608018 426786 608254
rect 427022 608018 462786 608254
rect 463022 608018 498786 608254
rect 499022 608018 534786 608254
rect 535022 608018 570786 608254
rect 571022 608018 592082 608254
rect 592318 608018 592500 608254
rect -8576 607934 592500 608018
rect -8576 607698 -8394 607934
rect -8158 607698 30786 607934
rect 31022 607698 66786 607934
rect 67022 607698 102786 607934
rect 103022 607698 138786 607934
rect 139022 607698 174786 607934
rect 175022 607698 210786 607934
rect 211022 607698 246786 607934
rect 247022 607698 282786 607934
rect 283022 607698 318786 607934
rect 319022 607698 354786 607934
rect 355022 607698 390786 607934
rect 391022 607698 426786 607934
rect 427022 607698 462786 607934
rect 463022 607698 498786 607934
rect 499022 607698 534786 607934
rect 535022 607698 570786 607934
rect 571022 607698 592082 607934
rect 592318 607698 592500 607934
rect -8576 607676 592500 607698
rect -8576 607674 -7976 607676
rect 30604 607674 31204 607676
rect 66604 607674 67204 607676
rect 102604 607674 103204 607676
rect 138604 607674 139204 607676
rect 174604 607674 175204 607676
rect 210604 607674 211204 607676
rect 246604 607674 247204 607676
rect 282604 607674 283204 607676
rect 318604 607674 319204 607676
rect 354604 607674 355204 607676
rect 390604 607674 391204 607676
rect 426604 607674 427204 607676
rect 462604 607674 463204 607676
rect 498604 607674 499204 607676
rect 534604 607674 535204 607676
rect 570604 607674 571204 607676
rect 591900 607674 592500 607676
rect -6696 604676 -6096 604678
rect 27004 604676 27604 604678
rect 63004 604676 63604 604678
rect 99004 604676 99604 604678
rect 135004 604676 135604 604678
rect 171004 604676 171604 604678
rect 207004 604676 207604 604678
rect 243004 604676 243604 604678
rect 279004 604676 279604 604678
rect 315004 604676 315604 604678
rect 351004 604676 351604 604678
rect 387004 604676 387604 604678
rect 423004 604676 423604 604678
rect 459004 604676 459604 604678
rect 495004 604676 495604 604678
rect 531004 604676 531604 604678
rect 567004 604676 567604 604678
rect 590020 604676 590620 604678
rect -6696 604654 590620 604676
rect -6696 604418 -6514 604654
rect -6278 604418 27186 604654
rect 27422 604418 63186 604654
rect 63422 604418 99186 604654
rect 99422 604418 135186 604654
rect 135422 604418 171186 604654
rect 171422 604418 207186 604654
rect 207422 604418 243186 604654
rect 243422 604418 279186 604654
rect 279422 604418 315186 604654
rect 315422 604418 351186 604654
rect 351422 604418 387186 604654
rect 387422 604418 423186 604654
rect 423422 604418 459186 604654
rect 459422 604418 495186 604654
rect 495422 604418 531186 604654
rect 531422 604418 567186 604654
rect 567422 604418 590202 604654
rect 590438 604418 590620 604654
rect -6696 604334 590620 604418
rect -6696 604098 -6514 604334
rect -6278 604098 27186 604334
rect 27422 604098 63186 604334
rect 63422 604098 99186 604334
rect 99422 604098 135186 604334
rect 135422 604098 171186 604334
rect 171422 604098 207186 604334
rect 207422 604098 243186 604334
rect 243422 604098 279186 604334
rect 279422 604098 315186 604334
rect 315422 604098 351186 604334
rect 351422 604098 387186 604334
rect 387422 604098 423186 604334
rect 423422 604098 459186 604334
rect 459422 604098 495186 604334
rect 495422 604098 531186 604334
rect 531422 604098 567186 604334
rect 567422 604098 590202 604334
rect 590438 604098 590620 604334
rect -6696 604076 590620 604098
rect -6696 604074 -6096 604076
rect 27004 604074 27604 604076
rect 63004 604074 63604 604076
rect 99004 604074 99604 604076
rect 135004 604074 135604 604076
rect 171004 604074 171604 604076
rect 207004 604074 207604 604076
rect 243004 604074 243604 604076
rect 279004 604074 279604 604076
rect 315004 604074 315604 604076
rect 351004 604074 351604 604076
rect 387004 604074 387604 604076
rect 423004 604074 423604 604076
rect 459004 604074 459604 604076
rect 495004 604074 495604 604076
rect 531004 604074 531604 604076
rect 567004 604074 567604 604076
rect 590020 604074 590620 604076
rect -4816 601076 -4216 601078
rect 23404 601076 24004 601078
rect 59404 601076 60004 601078
rect 95404 601076 96004 601078
rect 131404 601076 132004 601078
rect 167404 601076 168004 601078
rect 203404 601076 204004 601078
rect 239404 601076 240004 601078
rect 275404 601076 276004 601078
rect 311404 601076 312004 601078
rect 347404 601076 348004 601078
rect 383404 601076 384004 601078
rect 419404 601076 420004 601078
rect 455404 601076 456004 601078
rect 491404 601076 492004 601078
rect 527404 601076 528004 601078
rect 563404 601076 564004 601078
rect 588140 601076 588740 601078
rect -4816 601054 588740 601076
rect -4816 600818 -4634 601054
rect -4398 600818 23586 601054
rect 23822 600818 59586 601054
rect 59822 600818 95586 601054
rect 95822 600818 131586 601054
rect 131822 600818 167586 601054
rect 167822 600818 203586 601054
rect 203822 600818 239586 601054
rect 239822 600818 275586 601054
rect 275822 600818 311586 601054
rect 311822 600818 347586 601054
rect 347822 600818 383586 601054
rect 383822 600818 419586 601054
rect 419822 600818 455586 601054
rect 455822 600818 491586 601054
rect 491822 600818 527586 601054
rect 527822 600818 563586 601054
rect 563822 600818 588322 601054
rect 588558 600818 588740 601054
rect -4816 600734 588740 600818
rect -4816 600498 -4634 600734
rect -4398 600498 23586 600734
rect 23822 600498 59586 600734
rect 59822 600498 95586 600734
rect 95822 600498 131586 600734
rect 131822 600498 167586 600734
rect 167822 600498 203586 600734
rect 203822 600498 239586 600734
rect 239822 600498 275586 600734
rect 275822 600498 311586 600734
rect 311822 600498 347586 600734
rect 347822 600498 383586 600734
rect 383822 600498 419586 600734
rect 419822 600498 455586 600734
rect 455822 600498 491586 600734
rect 491822 600498 527586 600734
rect 527822 600498 563586 600734
rect 563822 600498 588322 600734
rect 588558 600498 588740 600734
rect -4816 600476 588740 600498
rect -4816 600474 -4216 600476
rect 23404 600474 24004 600476
rect 59404 600474 60004 600476
rect 95404 600474 96004 600476
rect 131404 600474 132004 600476
rect 167404 600474 168004 600476
rect 203404 600474 204004 600476
rect 239404 600474 240004 600476
rect 275404 600474 276004 600476
rect 311404 600474 312004 600476
rect 347404 600474 348004 600476
rect 383404 600474 384004 600476
rect 419404 600474 420004 600476
rect 455404 600474 456004 600476
rect 491404 600474 492004 600476
rect 527404 600474 528004 600476
rect 563404 600474 564004 600476
rect 588140 600474 588740 600476
rect -2936 597476 -2336 597478
rect 19804 597476 20404 597478
rect 55804 597476 56404 597478
rect 91804 597476 92404 597478
rect 127804 597476 128404 597478
rect 163804 597476 164404 597478
rect 199804 597476 200404 597478
rect 235804 597476 236404 597478
rect 271804 597476 272404 597478
rect 307804 597476 308404 597478
rect 343804 597476 344404 597478
rect 379804 597476 380404 597478
rect 415804 597476 416404 597478
rect 451804 597476 452404 597478
rect 487804 597476 488404 597478
rect 523804 597476 524404 597478
rect 559804 597476 560404 597478
rect 586260 597476 586860 597478
rect -2936 597454 586860 597476
rect -2936 597218 -2754 597454
rect -2518 597218 19986 597454
rect 20222 597218 55986 597454
rect 56222 597218 91986 597454
rect 92222 597218 127986 597454
rect 128222 597218 163986 597454
rect 164222 597218 199986 597454
rect 200222 597218 235986 597454
rect 236222 597218 271986 597454
rect 272222 597218 307986 597454
rect 308222 597218 343986 597454
rect 344222 597218 379986 597454
rect 380222 597218 415986 597454
rect 416222 597218 451986 597454
rect 452222 597218 487986 597454
rect 488222 597218 523986 597454
rect 524222 597218 559986 597454
rect 560222 597218 586442 597454
rect 586678 597218 586860 597454
rect -2936 597134 586860 597218
rect -2936 596898 -2754 597134
rect -2518 596898 19986 597134
rect 20222 596898 55986 597134
rect 56222 596898 91986 597134
rect 92222 596898 127986 597134
rect 128222 596898 163986 597134
rect 164222 596898 199986 597134
rect 200222 596898 235986 597134
rect 236222 596898 271986 597134
rect 272222 596898 307986 597134
rect 308222 596898 343986 597134
rect 344222 596898 379986 597134
rect 380222 596898 415986 597134
rect 416222 596898 451986 597134
rect 452222 596898 487986 597134
rect 488222 596898 523986 597134
rect 524222 596898 559986 597134
rect 560222 596898 586442 597134
rect 586678 596898 586860 597134
rect -2936 596876 586860 596898
rect -2936 596874 -2336 596876
rect 19804 596874 20404 596876
rect 55804 596874 56404 596876
rect 91804 596874 92404 596876
rect 127804 596874 128404 596876
rect 163804 596874 164404 596876
rect 199804 596874 200404 596876
rect 235804 596874 236404 596876
rect 271804 596874 272404 596876
rect 307804 596874 308404 596876
rect 343804 596874 344404 596876
rect 379804 596874 380404 596876
rect 415804 596874 416404 596876
rect 451804 596874 452404 596876
rect 487804 596874 488404 596876
rect 523804 596874 524404 596876
rect 559804 596874 560404 596876
rect 586260 596874 586860 596876
rect -7636 590276 -7036 590278
rect 12604 590276 13204 590278
rect 48604 590276 49204 590278
rect 84604 590276 85204 590278
rect 120604 590276 121204 590278
rect 156604 590276 157204 590278
rect 192604 590276 193204 590278
rect 228604 590276 229204 590278
rect 264604 590276 265204 590278
rect 300604 590276 301204 590278
rect 336604 590276 337204 590278
rect 372604 590276 373204 590278
rect 408604 590276 409204 590278
rect 444604 590276 445204 590278
rect 480604 590276 481204 590278
rect 516604 590276 517204 590278
rect 552604 590276 553204 590278
rect 590960 590276 591560 590278
rect -8576 590254 592500 590276
rect -8576 590018 -7454 590254
rect -7218 590018 12786 590254
rect 13022 590018 48786 590254
rect 49022 590018 84786 590254
rect 85022 590018 120786 590254
rect 121022 590018 156786 590254
rect 157022 590018 192786 590254
rect 193022 590018 228786 590254
rect 229022 590018 264786 590254
rect 265022 590018 300786 590254
rect 301022 590018 336786 590254
rect 337022 590018 372786 590254
rect 373022 590018 408786 590254
rect 409022 590018 444786 590254
rect 445022 590018 480786 590254
rect 481022 590018 516786 590254
rect 517022 590018 552786 590254
rect 553022 590018 591142 590254
rect 591378 590018 592500 590254
rect -8576 589934 592500 590018
rect -8576 589698 -7454 589934
rect -7218 589698 12786 589934
rect 13022 589698 48786 589934
rect 49022 589698 84786 589934
rect 85022 589698 120786 589934
rect 121022 589698 156786 589934
rect 157022 589698 192786 589934
rect 193022 589698 228786 589934
rect 229022 589698 264786 589934
rect 265022 589698 300786 589934
rect 301022 589698 336786 589934
rect 337022 589698 372786 589934
rect 373022 589698 408786 589934
rect 409022 589698 444786 589934
rect 445022 589698 480786 589934
rect 481022 589698 516786 589934
rect 517022 589698 552786 589934
rect 553022 589698 591142 589934
rect 591378 589698 592500 589934
rect -8576 589676 592500 589698
rect -7636 589674 -7036 589676
rect 12604 589674 13204 589676
rect 48604 589674 49204 589676
rect 84604 589674 85204 589676
rect 120604 589674 121204 589676
rect 156604 589674 157204 589676
rect 192604 589674 193204 589676
rect 228604 589674 229204 589676
rect 264604 589674 265204 589676
rect 300604 589674 301204 589676
rect 336604 589674 337204 589676
rect 372604 589674 373204 589676
rect 408604 589674 409204 589676
rect 444604 589674 445204 589676
rect 480604 589674 481204 589676
rect 516604 589674 517204 589676
rect 552604 589674 553204 589676
rect 590960 589674 591560 589676
rect -5756 586676 -5156 586678
rect 9004 586676 9604 586678
rect 45004 586676 45604 586678
rect 81004 586676 81604 586678
rect 117004 586676 117604 586678
rect 153004 586676 153604 586678
rect 189004 586676 189604 586678
rect 225004 586676 225604 586678
rect 261004 586676 261604 586678
rect 297004 586676 297604 586678
rect 333004 586676 333604 586678
rect 369004 586676 369604 586678
rect 405004 586676 405604 586678
rect 441004 586676 441604 586678
rect 477004 586676 477604 586678
rect 513004 586676 513604 586678
rect 549004 586676 549604 586678
rect 589080 586676 589680 586678
rect -6696 586654 590620 586676
rect -6696 586418 -5574 586654
rect -5338 586418 9186 586654
rect 9422 586418 45186 586654
rect 45422 586418 81186 586654
rect 81422 586418 117186 586654
rect 117422 586418 153186 586654
rect 153422 586418 189186 586654
rect 189422 586418 225186 586654
rect 225422 586418 261186 586654
rect 261422 586418 297186 586654
rect 297422 586418 333186 586654
rect 333422 586418 369186 586654
rect 369422 586418 405186 586654
rect 405422 586418 441186 586654
rect 441422 586418 477186 586654
rect 477422 586418 513186 586654
rect 513422 586418 549186 586654
rect 549422 586418 589262 586654
rect 589498 586418 590620 586654
rect -6696 586334 590620 586418
rect -6696 586098 -5574 586334
rect -5338 586098 9186 586334
rect 9422 586098 45186 586334
rect 45422 586098 81186 586334
rect 81422 586098 117186 586334
rect 117422 586098 153186 586334
rect 153422 586098 189186 586334
rect 189422 586098 225186 586334
rect 225422 586098 261186 586334
rect 261422 586098 297186 586334
rect 297422 586098 333186 586334
rect 333422 586098 369186 586334
rect 369422 586098 405186 586334
rect 405422 586098 441186 586334
rect 441422 586098 477186 586334
rect 477422 586098 513186 586334
rect 513422 586098 549186 586334
rect 549422 586098 589262 586334
rect 589498 586098 590620 586334
rect -6696 586076 590620 586098
rect -5756 586074 -5156 586076
rect 9004 586074 9604 586076
rect 45004 586074 45604 586076
rect 81004 586074 81604 586076
rect 117004 586074 117604 586076
rect 153004 586074 153604 586076
rect 189004 586074 189604 586076
rect 225004 586074 225604 586076
rect 261004 586074 261604 586076
rect 297004 586074 297604 586076
rect 333004 586074 333604 586076
rect 369004 586074 369604 586076
rect 405004 586074 405604 586076
rect 441004 586074 441604 586076
rect 477004 586074 477604 586076
rect 513004 586074 513604 586076
rect 549004 586074 549604 586076
rect 589080 586074 589680 586076
rect -3876 583076 -3276 583078
rect 5404 583076 6004 583078
rect 41404 583076 42004 583078
rect 77404 583076 78004 583078
rect 113404 583076 114004 583078
rect 149404 583076 150004 583078
rect 185404 583076 186004 583078
rect 221404 583076 222004 583078
rect 257404 583076 258004 583078
rect 293404 583076 294004 583078
rect 329404 583076 330004 583078
rect 365404 583076 366004 583078
rect 401404 583076 402004 583078
rect 437404 583076 438004 583078
rect 473404 583076 474004 583078
rect 509404 583076 510004 583078
rect 545404 583076 546004 583078
rect 581404 583076 582004 583078
rect 587200 583076 587800 583078
rect -4816 583054 588740 583076
rect -4816 582818 -3694 583054
rect -3458 582818 5586 583054
rect 5822 582818 41586 583054
rect 41822 582818 77586 583054
rect 77822 582818 113586 583054
rect 113822 582818 149586 583054
rect 149822 582818 185586 583054
rect 185822 582818 221586 583054
rect 221822 582818 257586 583054
rect 257822 582818 293586 583054
rect 293822 582818 329586 583054
rect 329822 582818 365586 583054
rect 365822 582818 401586 583054
rect 401822 582818 437586 583054
rect 437822 582818 473586 583054
rect 473822 582818 509586 583054
rect 509822 582818 545586 583054
rect 545822 582818 581586 583054
rect 581822 582818 587382 583054
rect 587618 582818 588740 583054
rect -4816 582734 588740 582818
rect -4816 582498 -3694 582734
rect -3458 582498 5586 582734
rect 5822 582498 41586 582734
rect 41822 582498 77586 582734
rect 77822 582498 113586 582734
rect 113822 582498 149586 582734
rect 149822 582498 185586 582734
rect 185822 582498 221586 582734
rect 221822 582498 257586 582734
rect 257822 582498 293586 582734
rect 293822 582498 329586 582734
rect 329822 582498 365586 582734
rect 365822 582498 401586 582734
rect 401822 582498 437586 582734
rect 437822 582498 473586 582734
rect 473822 582498 509586 582734
rect 509822 582498 545586 582734
rect 545822 582498 581586 582734
rect 581822 582498 587382 582734
rect 587618 582498 588740 582734
rect -4816 582476 588740 582498
rect -3876 582474 -3276 582476
rect 5404 582474 6004 582476
rect 41404 582474 42004 582476
rect 77404 582474 78004 582476
rect 113404 582474 114004 582476
rect 149404 582474 150004 582476
rect 185404 582474 186004 582476
rect 221404 582474 222004 582476
rect 257404 582474 258004 582476
rect 293404 582474 294004 582476
rect 329404 582474 330004 582476
rect 365404 582474 366004 582476
rect 401404 582474 402004 582476
rect 437404 582474 438004 582476
rect 473404 582474 474004 582476
rect 509404 582474 510004 582476
rect 545404 582474 546004 582476
rect 581404 582474 582004 582476
rect 587200 582474 587800 582476
rect -1996 579476 -1396 579478
rect 1804 579476 2404 579478
rect 37804 579476 38404 579478
rect 73804 579476 74404 579478
rect 109804 579476 110404 579478
rect 145804 579476 146404 579478
rect 181804 579476 182404 579478
rect 217804 579476 218404 579478
rect 253804 579476 254404 579478
rect 289804 579476 290404 579478
rect 325804 579476 326404 579478
rect 361804 579476 362404 579478
rect 397804 579476 398404 579478
rect 433804 579476 434404 579478
rect 469804 579476 470404 579478
rect 505804 579476 506404 579478
rect 541804 579476 542404 579478
rect 577804 579476 578404 579478
rect 585320 579476 585920 579478
rect -2936 579454 586860 579476
rect -2936 579218 -1814 579454
rect -1578 579218 1986 579454
rect 2222 579218 37986 579454
rect 38222 579218 73986 579454
rect 74222 579218 109986 579454
rect 110222 579218 145986 579454
rect 146222 579218 181986 579454
rect 182222 579218 217986 579454
rect 218222 579218 253986 579454
rect 254222 579218 289986 579454
rect 290222 579218 325986 579454
rect 326222 579218 361986 579454
rect 362222 579218 397986 579454
rect 398222 579218 433986 579454
rect 434222 579218 469986 579454
rect 470222 579218 505986 579454
rect 506222 579218 541986 579454
rect 542222 579218 577986 579454
rect 578222 579218 585502 579454
rect 585738 579218 586860 579454
rect -2936 579134 586860 579218
rect -2936 578898 -1814 579134
rect -1578 578898 1986 579134
rect 2222 578898 37986 579134
rect 38222 578898 73986 579134
rect 74222 578898 109986 579134
rect 110222 578898 145986 579134
rect 146222 578898 181986 579134
rect 182222 578898 217986 579134
rect 218222 578898 253986 579134
rect 254222 578898 289986 579134
rect 290222 578898 325986 579134
rect 326222 578898 361986 579134
rect 362222 578898 397986 579134
rect 398222 578898 433986 579134
rect 434222 578898 469986 579134
rect 470222 578898 505986 579134
rect 506222 578898 541986 579134
rect 542222 578898 577986 579134
rect 578222 578898 585502 579134
rect 585738 578898 586860 579134
rect -2936 578876 586860 578898
rect -1996 578874 -1396 578876
rect 1804 578874 2404 578876
rect 37804 578874 38404 578876
rect 73804 578874 74404 578876
rect 109804 578874 110404 578876
rect 145804 578874 146404 578876
rect 181804 578874 182404 578876
rect 217804 578874 218404 578876
rect 253804 578874 254404 578876
rect 289804 578874 290404 578876
rect 325804 578874 326404 578876
rect 361804 578874 362404 578876
rect 397804 578874 398404 578876
rect 433804 578874 434404 578876
rect 469804 578874 470404 578876
rect 505804 578874 506404 578876
rect 541804 578874 542404 578876
rect 577804 578874 578404 578876
rect 585320 578874 585920 578876
rect -8576 572276 -7976 572278
rect 30604 572276 31204 572278
rect 66604 572276 67204 572278
rect 102604 572276 103204 572278
rect 138604 572276 139204 572278
rect 174604 572276 175204 572278
rect 210604 572276 211204 572278
rect 246604 572276 247204 572278
rect 282604 572276 283204 572278
rect 318604 572276 319204 572278
rect 354604 572276 355204 572278
rect 390604 572276 391204 572278
rect 426604 572276 427204 572278
rect 462604 572276 463204 572278
rect 498604 572276 499204 572278
rect 534604 572276 535204 572278
rect 570604 572276 571204 572278
rect 591900 572276 592500 572278
rect -8576 572254 592500 572276
rect -8576 572018 -8394 572254
rect -8158 572018 30786 572254
rect 31022 572018 66786 572254
rect 67022 572018 102786 572254
rect 103022 572018 138786 572254
rect 139022 572018 174786 572254
rect 175022 572018 210786 572254
rect 211022 572018 246786 572254
rect 247022 572018 282786 572254
rect 283022 572018 318786 572254
rect 319022 572018 354786 572254
rect 355022 572018 390786 572254
rect 391022 572018 426786 572254
rect 427022 572018 462786 572254
rect 463022 572018 498786 572254
rect 499022 572018 534786 572254
rect 535022 572018 570786 572254
rect 571022 572018 592082 572254
rect 592318 572018 592500 572254
rect -8576 571934 592500 572018
rect -8576 571698 -8394 571934
rect -8158 571698 30786 571934
rect 31022 571698 66786 571934
rect 67022 571698 102786 571934
rect 103022 571698 138786 571934
rect 139022 571698 174786 571934
rect 175022 571698 210786 571934
rect 211022 571698 246786 571934
rect 247022 571698 282786 571934
rect 283022 571698 318786 571934
rect 319022 571698 354786 571934
rect 355022 571698 390786 571934
rect 391022 571698 426786 571934
rect 427022 571698 462786 571934
rect 463022 571698 498786 571934
rect 499022 571698 534786 571934
rect 535022 571698 570786 571934
rect 571022 571698 592082 571934
rect 592318 571698 592500 571934
rect -8576 571676 592500 571698
rect -8576 571674 -7976 571676
rect 30604 571674 31204 571676
rect 66604 571674 67204 571676
rect 102604 571674 103204 571676
rect 138604 571674 139204 571676
rect 174604 571674 175204 571676
rect 210604 571674 211204 571676
rect 246604 571674 247204 571676
rect 282604 571674 283204 571676
rect 318604 571674 319204 571676
rect 354604 571674 355204 571676
rect 390604 571674 391204 571676
rect 426604 571674 427204 571676
rect 462604 571674 463204 571676
rect 498604 571674 499204 571676
rect 534604 571674 535204 571676
rect 570604 571674 571204 571676
rect 591900 571674 592500 571676
rect -6696 568676 -6096 568678
rect 27004 568676 27604 568678
rect 63004 568676 63604 568678
rect 99004 568676 99604 568678
rect 135004 568676 135604 568678
rect 171004 568676 171604 568678
rect 207004 568676 207604 568678
rect 243004 568676 243604 568678
rect 279004 568676 279604 568678
rect 315004 568676 315604 568678
rect 351004 568676 351604 568678
rect 387004 568676 387604 568678
rect 423004 568676 423604 568678
rect 459004 568676 459604 568678
rect 495004 568676 495604 568678
rect 531004 568676 531604 568678
rect 567004 568676 567604 568678
rect 590020 568676 590620 568678
rect -6696 568654 590620 568676
rect -6696 568418 -6514 568654
rect -6278 568418 27186 568654
rect 27422 568418 63186 568654
rect 63422 568418 99186 568654
rect 99422 568418 135186 568654
rect 135422 568418 171186 568654
rect 171422 568418 207186 568654
rect 207422 568418 243186 568654
rect 243422 568418 279186 568654
rect 279422 568418 315186 568654
rect 315422 568418 351186 568654
rect 351422 568418 387186 568654
rect 387422 568418 423186 568654
rect 423422 568418 459186 568654
rect 459422 568418 495186 568654
rect 495422 568418 531186 568654
rect 531422 568418 567186 568654
rect 567422 568418 590202 568654
rect 590438 568418 590620 568654
rect -6696 568334 590620 568418
rect -6696 568098 -6514 568334
rect -6278 568098 27186 568334
rect 27422 568098 63186 568334
rect 63422 568098 99186 568334
rect 99422 568098 135186 568334
rect 135422 568098 171186 568334
rect 171422 568098 207186 568334
rect 207422 568098 243186 568334
rect 243422 568098 279186 568334
rect 279422 568098 315186 568334
rect 315422 568098 351186 568334
rect 351422 568098 387186 568334
rect 387422 568098 423186 568334
rect 423422 568098 459186 568334
rect 459422 568098 495186 568334
rect 495422 568098 531186 568334
rect 531422 568098 567186 568334
rect 567422 568098 590202 568334
rect 590438 568098 590620 568334
rect -6696 568076 590620 568098
rect -6696 568074 -6096 568076
rect 27004 568074 27604 568076
rect 63004 568074 63604 568076
rect 99004 568074 99604 568076
rect 135004 568074 135604 568076
rect 171004 568074 171604 568076
rect 207004 568074 207604 568076
rect 243004 568074 243604 568076
rect 279004 568074 279604 568076
rect 315004 568074 315604 568076
rect 351004 568074 351604 568076
rect 387004 568074 387604 568076
rect 423004 568074 423604 568076
rect 459004 568074 459604 568076
rect 495004 568074 495604 568076
rect 531004 568074 531604 568076
rect 567004 568074 567604 568076
rect 590020 568074 590620 568076
rect -4816 565076 -4216 565078
rect 23404 565076 24004 565078
rect 59404 565076 60004 565078
rect 95404 565076 96004 565078
rect 131404 565076 132004 565078
rect 167404 565076 168004 565078
rect 203404 565076 204004 565078
rect 239404 565076 240004 565078
rect 275404 565076 276004 565078
rect 311404 565076 312004 565078
rect 347404 565076 348004 565078
rect 383404 565076 384004 565078
rect 419404 565076 420004 565078
rect 455404 565076 456004 565078
rect 491404 565076 492004 565078
rect 527404 565076 528004 565078
rect 563404 565076 564004 565078
rect 588140 565076 588740 565078
rect -4816 565054 588740 565076
rect -4816 564818 -4634 565054
rect -4398 564818 23586 565054
rect 23822 564818 59586 565054
rect 59822 564818 95586 565054
rect 95822 564818 131586 565054
rect 131822 564818 167586 565054
rect 167822 564818 203586 565054
rect 203822 564818 239586 565054
rect 239822 564818 275586 565054
rect 275822 564818 311586 565054
rect 311822 564818 347586 565054
rect 347822 564818 383586 565054
rect 383822 564818 419586 565054
rect 419822 564818 455586 565054
rect 455822 564818 491586 565054
rect 491822 564818 527586 565054
rect 527822 564818 563586 565054
rect 563822 564818 588322 565054
rect 588558 564818 588740 565054
rect -4816 564734 588740 564818
rect -4816 564498 -4634 564734
rect -4398 564498 23586 564734
rect 23822 564498 59586 564734
rect 59822 564498 95586 564734
rect 95822 564498 131586 564734
rect 131822 564498 167586 564734
rect 167822 564498 203586 564734
rect 203822 564498 239586 564734
rect 239822 564498 275586 564734
rect 275822 564498 311586 564734
rect 311822 564498 347586 564734
rect 347822 564498 383586 564734
rect 383822 564498 419586 564734
rect 419822 564498 455586 564734
rect 455822 564498 491586 564734
rect 491822 564498 527586 564734
rect 527822 564498 563586 564734
rect 563822 564498 588322 564734
rect 588558 564498 588740 564734
rect -4816 564476 588740 564498
rect -4816 564474 -4216 564476
rect 23404 564474 24004 564476
rect 59404 564474 60004 564476
rect 95404 564474 96004 564476
rect 131404 564474 132004 564476
rect 167404 564474 168004 564476
rect 203404 564474 204004 564476
rect 239404 564474 240004 564476
rect 275404 564474 276004 564476
rect 311404 564474 312004 564476
rect 347404 564474 348004 564476
rect 383404 564474 384004 564476
rect 419404 564474 420004 564476
rect 455404 564474 456004 564476
rect 491404 564474 492004 564476
rect 527404 564474 528004 564476
rect 563404 564474 564004 564476
rect 588140 564474 588740 564476
rect -2936 561476 -2336 561478
rect 19804 561476 20404 561478
rect 55804 561476 56404 561478
rect 91804 561476 92404 561478
rect 127804 561476 128404 561478
rect 163804 561476 164404 561478
rect 199804 561476 200404 561478
rect 235804 561476 236404 561478
rect 271804 561476 272404 561478
rect 307804 561476 308404 561478
rect 343804 561476 344404 561478
rect 379804 561476 380404 561478
rect 415804 561476 416404 561478
rect 451804 561476 452404 561478
rect 487804 561476 488404 561478
rect 523804 561476 524404 561478
rect 559804 561476 560404 561478
rect 586260 561476 586860 561478
rect -2936 561454 586860 561476
rect -2936 561218 -2754 561454
rect -2518 561218 19986 561454
rect 20222 561218 55986 561454
rect 56222 561218 91986 561454
rect 92222 561218 127986 561454
rect 128222 561218 163986 561454
rect 164222 561218 199986 561454
rect 200222 561218 235986 561454
rect 236222 561218 271986 561454
rect 272222 561218 307986 561454
rect 308222 561218 343986 561454
rect 344222 561218 379986 561454
rect 380222 561218 415986 561454
rect 416222 561218 451986 561454
rect 452222 561218 487986 561454
rect 488222 561218 523986 561454
rect 524222 561218 559986 561454
rect 560222 561218 586442 561454
rect 586678 561218 586860 561454
rect -2936 561134 586860 561218
rect -2936 560898 -2754 561134
rect -2518 560898 19986 561134
rect 20222 560898 55986 561134
rect 56222 560898 91986 561134
rect 92222 560898 127986 561134
rect 128222 560898 163986 561134
rect 164222 560898 199986 561134
rect 200222 560898 235986 561134
rect 236222 560898 271986 561134
rect 272222 560898 307986 561134
rect 308222 560898 343986 561134
rect 344222 560898 379986 561134
rect 380222 560898 415986 561134
rect 416222 560898 451986 561134
rect 452222 560898 487986 561134
rect 488222 560898 523986 561134
rect 524222 560898 559986 561134
rect 560222 560898 586442 561134
rect 586678 560898 586860 561134
rect -2936 560876 586860 560898
rect -2936 560874 -2336 560876
rect 19804 560874 20404 560876
rect 55804 560874 56404 560876
rect 91804 560874 92404 560876
rect 127804 560874 128404 560876
rect 163804 560874 164404 560876
rect 199804 560874 200404 560876
rect 235804 560874 236404 560876
rect 271804 560874 272404 560876
rect 307804 560874 308404 560876
rect 343804 560874 344404 560876
rect 379804 560874 380404 560876
rect 415804 560874 416404 560876
rect 451804 560874 452404 560876
rect 487804 560874 488404 560876
rect 523804 560874 524404 560876
rect 559804 560874 560404 560876
rect 586260 560874 586860 560876
rect -7636 554276 -7036 554278
rect 12604 554276 13204 554278
rect 48604 554276 49204 554278
rect 84604 554276 85204 554278
rect 120604 554276 121204 554278
rect 156604 554276 157204 554278
rect 192604 554276 193204 554278
rect 228604 554276 229204 554278
rect 264604 554276 265204 554278
rect 300604 554276 301204 554278
rect 336604 554276 337204 554278
rect 372604 554276 373204 554278
rect 408604 554276 409204 554278
rect 444604 554276 445204 554278
rect 480604 554276 481204 554278
rect 516604 554276 517204 554278
rect 552604 554276 553204 554278
rect 590960 554276 591560 554278
rect -8576 554254 592500 554276
rect -8576 554018 -7454 554254
rect -7218 554018 12786 554254
rect 13022 554018 48786 554254
rect 49022 554018 84786 554254
rect 85022 554018 120786 554254
rect 121022 554018 156786 554254
rect 157022 554018 192786 554254
rect 193022 554018 228786 554254
rect 229022 554018 264786 554254
rect 265022 554018 300786 554254
rect 301022 554018 336786 554254
rect 337022 554018 372786 554254
rect 373022 554018 408786 554254
rect 409022 554018 444786 554254
rect 445022 554018 480786 554254
rect 481022 554018 516786 554254
rect 517022 554018 552786 554254
rect 553022 554018 591142 554254
rect 591378 554018 592500 554254
rect -8576 553934 592500 554018
rect -8576 553698 -7454 553934
rect -7218 553698 12786 553934
rect 13022 553698 48786 553934
rect 49022 553698 84786 553934
rect 85022 553698 120786 553934
rect 121022 553698 156786 553934
rect 157022 553698 192786 553934
rect 193022 553698 228786 553934
rect 229022 553698 264786 553934
rect 265022 553698 300786 553934
rect 301022 553698 336786 553934
rect 337022 553698 372786 553934
rect 373022 553698 408786 553934
rect 409022 553698 444786 553934
rect 445022 553698 480786 553934
rect 481022 553698 516786 553934
rect 517022 553698 552786 553934
rect 553022 553698 591142 553934
rect 591378 553698 592500 553934
rect -8576 553676 592500 553698
rect -7636 553674 -7036 553676
rect 12604 553674 13204 553676
rect 48604 553674 49204 553676
rect 84604 553674 85204 553676
rect 120604 553674 121204 553676
rect 156604 553674 157204 553676
rect 192604 553674 193204 553676
rect 228604 553674 229204 553676
rect 264604 553674 265204 553676
rect 300604 553674 301204 553676
rect 336604 553674 337204 553676
rect 372604 553674 373204 553676
rect 408604 553674 409204 553676
rect 444604 553674 445204 553676
rect 480604 553674 481204 553676
rect 516604 553674 517204 553676
rect 552604 553674 553204 553676
rect 590960 553674 591560 553676
rect -5756 550676 -5156 550678
rect 9004 550676 9604 550678
rect 45004 550676 45604 550678
rect 81004 550676 81604 550678
rect 117004 550676 117604 550678
rect 153004 550676 153604 550678
rect 189004 550676 189604 550678
rect 225004 550676 225604 550678
rect 261004 550676 261604 550678
rect 297004 550676 297604 550678
rect 333004 550676 333604 550678
rect 369004 550676 369604 550678
rect 405004 550676 405604 550678
rect 441004 550676 441604 550678
rect 477004 550676 477604 550678
rect 513004 550676 513604 550678
rect 549004 550676 549604 550678
rect 589080 550676 589680 550678
rect -6696 550654 590620 550676
rect -6696 550418 -5574 550654
rect -5338 550418 9186 550654
rect 9422 550418 45186 550654
rect 45422 550418 81186 550654
rect 81422 550418 117186 550654
rect 117422 550418 153186 550654
rect 153422 550418 189186 550654
rect 189422 550418 225186 550654
rect 225422 550418 261186 550654
rect 261422 550418 297186 550654
rect 297422 550418 333186 550654
rect 333422 550418 369186 550654
rect 369422 550418 405186 550654
rect 405422 550418 441186 550654
rect 441422 550418 477186 550654
rect 477422 550418 513186 550654
rect 513422 550418 549186 550654
rect 549422 550418 589262 550654
rect 589498 550418 590620 550654
rect -6696 550334 590620 550418
rect -6696 550098 -5574 550334
rect -5338 550098 9186 550334
rect 9422 550098 45186 550334
rect 45422 550098 81186 550334
rect 81422 550098 117186 550334
rect 117422 550098 153186 550334
rect 153422 550098 189186 550334
rect 189422 550098 225186 550334
rect 225422 550098 261186 550334
rect 261422 550098 297186 550334
rect 297422 550098 333186 550334
rect 333422 550098 369186 550334
rect 369422 550098 405186 550334
rect 405422 550098 441186 550334
rect 441422 550098 477186 550334
rect 477422 550098 513186 550334
rect 513422 550098 549186 550334
rect 549422 550098 589262 550334
rect 589498 550098 590620 550334
rect -6696 550076 590620 550098
rect -5756 550074 -5156 550076
rect 9004 550074 9604 550076
rect 45004 550074 45604 550076
rect 81004 550074 81604 550076
rect 117004 550074 117604 550076
rect 153004 550074 153604 550076
rect 189004 550074 189604 550076
rect 225004 550074 225604 550076
rect 261004 550074 261604 550076
rect 297004 550074 297604 550076
rect 333004 550074 333604 550076
rect 369004 550074 369604 550076
rect 405004 550074 405604 550076
rect 441004 550074 441604 550076
rect 477004 550074 477604 550076
rect 513004 550074 513604 550076
rect 549004 550074 549604 550076
rect 589080 550074 589680 550076
rect -3876 547076 -3276 547078
rect 5404 547076 6004 547078
rect 41404 547076 42004 547078
rect 77404 547076 78004 547078
rect 113404 547076 114004 547078
rect 149404 547076 150004 547078
rect 185404 547076 186004 547078
rect 221404 547076 222004 547078
rect 257404 547076 258004 547078
rect 293404 547076 294004 547078
rect 329404 547076 330004 547078
rect 365404 547076 366004 547078
rect 401404 547076 402004 547078
rect 437404 547076 438004 547078
rect 473404 547076 474004 547078
rect 509404 547076 510004 547078
rect 545404 547076 546004 547078
rect 581404 547076 582004 547078
rect 587200 547076 587800 547078
rect -4816 547054 588740 547076
rect -4816 546818 -3694 547054
rect -3458 546818 5586 547054
rect 5822 546818 41586 547054
rect 41822 546818 77586 547054
rect 77822 546818 113586 547054
rect 113822 546818 149586 547054
rect 149822 546818 185586 547054
rect 185822 546818 221586 547054
rect 221822 546818 257586 547054
rect 257822 546818 293586 547054
rect 293822 546818 329586 547054
rect 329822 546818 365586 547054
rect 365822 546818 401586 547054
rect 401822 546818 437586 547054
rect 437822 546818 473586 547054
rect 473822 546818 509586 547054
rect 509822 546818 545586 547054
rect 545822 546818 581586 547054
rect 581822 546818 587382 547054
rect 587618 546818 588740 547054
rect -4816 546734 588740 546818
rect -4816 546498 -3694 546734
rect -3458 546498 5586 546734
rect 5822 546498 41586 546734
rect 41822 546498 77586 546734
rect 77822 546498 113586 546734
rect 113822 546498 149586 546734
rect 149822 546498 185586 546734
rect 185822 546498 221586 546734
rect 221822 546498 257586 546734
rect 257822 546498 293586 546734
rect 293822 546498 329586 546734
rect 329822 546498 365586 546734
rect 365822 546498 401586 546734
rect 401822 546498 437586 546734
rect 437822 546498 473586 546734
rect 473822 546498 509586 546734
rect 509822 546498 545586 546734
rect 545822 546498 581586 546734
rect 581822 546498 587382 546734
rect 587618 546498 588740 546734
rect -4816 546476 588740 546498
rect -3876 546474 -3276 546476
rect 5404 546474 6004 546476
rect 41404 546474 42004 546476
rect 77404 546474 78004 546476
rect 113404 546474 114004 546476
rect 149404 546474 150004 546476
rect 185404 546474 186004 546476
rect 221404 546474 222004 546476
rect 257404 546474 258004 546476
rect 293404 546474 294004 546476
rect 329404 546474 330004 546476
rect 365404 546474 366004 546476
rect 401404 546474 402004 546476
rect 437404 546474 438004 546476
rect 473404 546474 474004 546476
rect 509404 546474 510004 546476
rect 545404 546474 546004 546476
rect 581404 546474 582004 546476
rect 587200 546474 587800 546476
rect -1996 543476 -1396 543478
rect 1804 543476 2404 543478
rect 37804 543476 38404 543478
rect 73804 543476 74404 543478
rect 109804 543476 110404 543478
rect 145804 543476 146404 543478
rect 181804 543476 182404 543478
rect 217804 543476 218404 543478
rect 253804 543476 254404 543478
rect 289804 543476 290404 543478
rect 325804 543476 326404 543478
rect 361804 543476 362404 543478
rect 397804 543476 398404 543478
rect 433804 543476 434404 543478
rect 469804 543476 470404 543478
rect 505804 543476 506404 543478
rect 541804 543476 542404 543478
rect 577804 543476 578404 543478
rect 585320 543476 585920 543478
rect -2936 543454 586860 543476
rect -2936 543218 -1814 543454
rect -1578 543218 1986 543454
rect 2222 543218 37986 543454
rect 38222 543218 73986 543454
rect 74222 543218 109986 543454
rect 110222 543218 145986 543454
rect 146222 543218 181986 543454
rect 182222 543218 217986 543454
rect 218222 543218 253986 543454
rect 254222 543218 289986 543454
rect 290222 543218 325986 543454
rect 326222 543218 361986 543454
rect 362222 543218 397986 543454
rect 398222 543218 433986 543454
rect 434222 543218 469986 543454
rect 470222 543218 505986 543454
rect 506222 543218 541986 543454
rect 542222 543218 577986 543454
rect 578222 543218 585502 543454
rect 585738 543218 586860 543454
rect -2936 543134 586860 543218
rect -2936 542898 -1814 543134
rect -1578 542898 1986 543134
rect 2222 542898 37986 543134
rect 38222 542898 73986 543134
rect 74222 542898 109986 543134
rect 110222 542898 145986 543134
rect 146222 542898 181986 543134
rect 182222 542898 217986 543134
rect 218222 542898 253986 543134
rect 254222 542898 289986 543134
rect 290222 542898 325986 543134
rect 326222 542898 361986 543134
rect 362222 542898 397986 543134
rect 398222 542898 433986 543134
rect 434222 542898 469986 543134
rect 470222 542898 505986 543134
rect 506222 542898 541986 543134
rect 542222 542898 577986 543134
rect 578222 542898 585502 543134
rect 585738 542898 586860 543134
rect -2936 542876 586860 542898
rect -1996 542874 -1396 542876
rect 1804 542874 2404 542876
rect 37804 542874 38404 542876
rect 73804 542874 74404 542876
rect 109804 542874 110404 542876
rect 145804 542874 146404 542876
rect 181804 542874 182404 542876
rect 217804 542874 218404 542876
rect 253804 542874 254404 542876
rect 289804 542874 290404 542876
rect 325804 542874 326404 542876
rect 361804 542874 362404 542876
rect 397804 542874 398404 542876
rect 433804 542874 434404 542876
rect 469804 542874 470404 542876
rect 505804 542874 506404 542876
rect 541804 542874 542404 542876
rect 577804 542874 578404 542876
rect 585320 542874 585920 542876
rect -8576 536276 -7976 536278
rect 30604 536276 31204 536278
rect 66604 536276 67204 536278
rect 102604 536276 103204 536278
rect 138604 536276 139204 536278
rect 174604 536276 175204 536278
rect 210604 536276 211204 536278
rect 246604 536276 247204 536278
rect 282604 536276 283204 536278
rect 318604 536276 319204 536278
rect 354604 536276 355204 536278
rect 390604 536276 391204 536278
rect 426604 536276 427204 536278
rect 462604 536276 463204 536278
rect 498604 536276 499204 536278
rect 534604 536276 535204 536278
rect 570604 536276 571204 536278
rect 591900 536276 592500 536278
rect -8576 536254 592500 536276
rect -8576 536018 -8394 536254
rect -8158 536018 30786 536254
rect 31022 536018 66786 536254
rect 67022 536018 102786 536254
rect 103022 536018 138786 536254
rect 139022 536018 174786 536254
rect 175022 536018 210786 536254
rect 211022 536018 246786 536254
rect 247022 536018 282786 536254
rect 283022 536018 318786 536254
rect 319022 536018 354786 536254
rect 355022 536018 390786 536254
rect 391022 536018 426786 536254
rect 427022 536018 462786 536254
rect 463022 536018 498786 536254
rect 499022 536018 534786 536254
rect 535022 536018 570786 536254
rect 571022 536018 592082 536254
rect 592318 536018 592500 536254
rect -8576 535934 592500 536018
rect -8576 535698 -8394 535934
rect -8158 535698 30786 535934
rect 31022 535698 66786 535934
rect 67022 535698 102786 535934
rect 103022 535698 138786 535934
rect 139022 535698 174786 535934
rect 175022 535698 210786 535934
rect 211022 535698 246786 535934
rect 247022 535698 282786 535934
rect 283022 535698 318786 535934
rect 319022 535698 354786 535934
rect 355022 535698 390786 535934
rect 391022 535698 426786 535934
rect 427022 535698 462786 535934
rect 463022 535698 498786 535934
rect 499022 535698 534786 535934
rect 535022 535698 570786 535934
rect 571022 535698 592082 535934
rect 592318 535698 592500 535934
rect -8576 535676 592500 535698
rect -8576 535674 -7976 535676
rect 30604 535674 31204 535676
rect 66604 535674 67204 535676
rect 102604 535674 103204 535676
rect 138604 535674 139204 535676
rect 174604 535674 175204 535676
rect 210604 535674 211204 535676
rect 246604 535674 247204 535676
rect 282604 535674 283204 535676
rect 318604 535674 319204 535676
rect 354604 535674 355204 535676
rect 390604 535674 391204 535676
rect 426604 535674 427204 535676
rect 462604 535674 463204 535676
rect 498604 535674 499204 535676
rect 534604 535674 535204 535676
rect 570604 535674 571204 535676
rect 591900 535674 592500 535676
rect -6696 532676 -6096 532678
rect 27004 532676 27604 532678
rect 63004 532676 63604 532678
rect 99004 532676 99604 532678
rect 135004 532676 135604 532678
rect 171004 532676 171604 532678
rect 207004 532676 207604 532678
rect 243004 532676 243604 532678
rect 279004 532676 279604 532678
rect 315004 532676 315604 532678
rect 351004 532676 351604 532678
rect 387004 532676 387604 532678
rect 423004 532676 423604 532678
rect 459004 532676 459604 532678
rect 495004 532676 495604 532678
rect 531004 532676 531604 532678
rect 567004 532676 567604 532678
rect 590020 532676 590620 532678
rect -6696 532654 590620 532676
rect -6696 532418 -6514 532654
rect -6278 532418 27186 532654
rect 27422 532418 63186 532654
rect 63422 532418 99186 532654
rect 99422 532418 135186 532654
rect 135422 532418 171186 532654
rect 171422 532418 207186 532654
rect 207422 532418 243186 532654
rect 243422 532418 279186 532654
rect 279422 532418 315186 532654
rect 315422 532418 351186 532654
rect 351422 532418 387186 532654
rect 387422 532418 423186 532654
rect 423422 532418 459186 532654
rect 459422 532418 495186 532654
rect 495422 532418 531186 532654
rect 531422 532418 567186 532654
rect 567422 532418 590202 532654
rect 590438 532418 590620 532654
rect -6696 532334 590620 532418
rect -6696 532098 -6514 532334
rect -6278 532098 27186 532334
rect 27422 532098 63186 532334
rect 63422 532098 99186 532334
rect 99422 532098 135186 532334
rect 135422 532098 171186 532334
rect 171422 532098 207186 532334
rect 207422 532098 243186 532334
rect 243422 532098 279186 532334
rect 279422 532098 315186 532334
rect 315422 532098 351186 532334
rect 351422 532098 387186 532334
rect 387422 532098 423186 532334
rect 423422 532098 459186 532334
rect 459422 532098 495186 532334
rect 495422 532098 531186 532334
rect 531422 532098 567186 532334
rect 567422 532098 590202 532334
rect 590438 532098 590620 532334
rect -6696 532076 590620 532098
rect -6696 532074 -6096 532076
rect 27004 532074 27604 532076
rect 63004 532074 63604 532076
rect 99004 532074 99604 532076
rect 135004 532074 135604 532076
rect 171004 532074 171604 532076
rect 207004 532074 207604 532076
rect 243004 532074 243604 532076
rect 279004 532074 279604 532076
rect 315004 532074 315604 532076
rect 351004 532074 351604 532076
rect 387004 532074 387604 532076
rect 423004 532074 423604 532076
rect 459004 532074 459604 532076
rect 495004 532074 495604 532076
rect 531004 532074 531604 532076
rect 567004 532074 567604 532076
rect 590020 532074 590620 532076
rect -4816 529076 -4216 529078
rect 23404 529076 24004 529078
rect 59404 529076 60004 529078
rect 95404 529076 96004 529078
rect 131404 529076 132004 529078
rect 167404 529076 168004 529078
rect 203404 529076 204004 529078
rect 239404 529076 240004 529078
rect 275404 529076 276004 529078
rect 311404 529076 312004 529078
rect 347404 529076 348004 529078
rect 383404 529076 384004 529078
rect 419404 529076 420004 529078
rect 455404 529076 456004 529078
rect 491404 529076 492004 529078
rect 527404 529076 528004 529078
rect 563404 529076 564004 529078
rect 588140 529076 588740 529078
rect -4816 529054 588740 529076
rect -4816 528818 -4634 529054
rect -4398 528818 23586 529054
rect 23822 528818 59586 529054
rect 59822 528818 95586 529054
rect 95822 528818 131586 529054
rect 131822 528818 167586 529054
rect 167822 528818 203586 529054
rect 203822 528818 239586 529054
rect 239822 528818 275586 529054
rect 275822 528818 311586 529054
rect 311822 528818 347586 529054
rect 347822 528818 383586 529054
rect 383822 528818 419586 529054
rect 419822 528818 455586 529054
rect 455822 528818 491586 529054
rect 491822 528818 527586 529054
rect 527822 528818 563586 529054
rect 563822 528818 588322 529054
rect 588558 528818 588740 529054
rect -4816 528734 588740 528818
rect -4816 528498 -4634 528734
rect -4398 528498 23586 528734
rect 23822 528498 59586 528734
rect 59822 528498 95586 528734
rect 95822 528498 131586 528734
rect 131822 528498 167586 528734
rect 167822 528498 203586 528734
rect 203822 528498 239586 528734
rect 239822 528498 275586 528734
rect 275822 528498 311586 528734
rect 311822 528498 347586 528734
rect 347822 528498 383586 528734
rect 383822 528498 419586 528734
rect 419822 528498 455586 528734
rect 455822 528498 491586 528734
rect 491822 528498 527586 528734
rect 527822 528498 563586 528734
rect 563822 528498 588322 528734
rect 588558 528498 588740 528734
rect -4816 528476 588740 528498
rect -4816 528474 -4216 528476
rect 23404 528474 24004 528476
rect 59404 528474 60004 528476
rect 95404 528474 96004 528476
rect 131404 528474 132004 528476
rect 167404 528474 168004 528476
rect 203404 528474 204004 528476
rect 239404 528474 240004 528476
rect 275404 528474 276004 528476
rect 311404 528474 312004 528476
rect 347404 528474 348004 528476
rect 383404 528474 384004 528476
rect 419404 528474 420004 528476
rect 455404 528474 456004 528476
rect 491404 528474 492004 528476
rect 527404 528474 528004 528476
rect 563404 528474 564004 528476
rect 588140 528474 588740 528476
rect -2936 525476 -2336 525478
rect 19804 525476 20404 525478
rect 55804 525476 56404 525478
rect 91804 525476 92404 525478
rect 127804 525476 128404 525478
rect 163804 525476 164404 525478
rect 199804 525476 200404 525478
rect 235804 525476 236404 525478
rect 271804 525476 272404 525478
rect 307804 525476 308404 525478
rect 343804 525476 344404 525478
rect 379804 525476 380404 525478
rect 415804 525476 416404 525478
rect 451804 525476 452404 525478
rect 487804 525476 488404 525478
rect 523804 525476 524404 525478
rect 559804 525476 560404 525478
rect 586260 525476 586860 525478
rect -2936 525454 586860 525476
rect -2936 525218 -2754 525454
rect -2518 525218 19986 525454
rect 20222 525218 55986 525454
rect 56222 525218 91986 525454
rect 92222 525218 127986 525454
rect 128222 525218 163986 525454
rect 164222 525218 199986 525454
rect 200222 525218 235986 525454
rect 236222 525218 271986 525454
rect 272222 525218 307986 525454
rect 308222 525218 343986 525454
rect 344222 525218 379986 525454
rect 380222 525218 415986 525454
rect 416222 525218 451986 525454
rect 452222 525218 487986 525454
rect 488222 525218 523986 525454
rect 524222 525218 559986 525454
rect 560222 525218 586442 525454
rect 586678 525218 586860 525454
rect -2936 525134 586860 525218
rect -2936 524898 -2754 525134
rect -2518 524898 19986 525134
rect 20222 524898 55986 525134
rect 56222 524898 91986 525134
rect 92222 524898 127986 525134
rect 128222 524898 163986 525134
rect 164222 524898 199986 525134
rect 200222 524898 235986 525134
rect 236222 524898 271986 525134
rect 272222 524898 307986 525134
rect 308222 524898 343986 525134
rect 344222 524898 379986 525134
rect 380222 524898 415986 525134
rect 416222 524898 451986 525134
rect 452222 524898 487986 525134
rect 488222 524898 523986 525134
rect 524222 524898 559986 525134
rect 560222 524898 586442 525134
rect 586678 524898 586860 525134
rect -2936 524876 586860 524898
rect -2936 524874 -2336 524876
rect 19804 524874 20404 524876
rect 55804 524874 56404 524876
rect 91804 524874 92404 524876
rect 127804 524874 128404 524876
rect 163804 524874 164404 524876
rect 199804 524874 200404 524876
rect 235804 524874 236404 524876
rect 271804 524874 272404 524876
rect 307804 524874 308404 524876
rect 343804 524874 344404 524876
rect 379804 524874 380404 524876
rect 415804 524874 416404 524876
rect 451804 524874 452404 524876
rect 487804 524874 488404 524876
rect 523804 524874 524404 524876
rect 559804 524874 560404 524876
rect 586260 524874 586860 524876
rect -7636 518276 -7036 518278
rect 12604 518276 13204 518278
rect 48604 518276 49204 518278
rect 84604 518276 85204 518278
rect 120604 518276 121204 518278
rect 156604 518276 157204 518278
rect 192604 518276 193204 518278
rect 228604 518276 229204 518278
rect 264604 518276 265204 518278
rect 300604 518276 301204 518278
rect 336604 518276 337204 518278
rect 372604 518276 373204 518278
rect 408604 518276 409204 518278
rect 444604 518276 445204 518278
rect 480604 518276 481204 518278
rect 516604 518276 517204 518278
rect 552604 518276 553204 518278
rect 590960 518276 591560 518278
rect -8576 518254 592500 518276
rect -8576 518018 -7454 518254
rect -7218 518018 12786 518254
rect 13022 518018 48786 518254
rect 49022 518018 84786 518254
rect 85022 518018 120786 518254
rect 121022 518018 156786 518254
rect 157022 518018 192786 518254
rect 193022 518018 228786 518254
rect 229022 518018 264786 518254
rect 265022 518018 300786 518254
rect 301022 518018 336786 518254
rect 337022 518018 372786 518254
rect 373022 518018 408786 518254
rect 409022 518018 444786 518254
rect 445022 518018 480786 518254
rect 481022 518018 516786 518254
rect 517022 518018 552786 518254
rect 553022 518018 591142 518254
rect 591378 518018 592500 518254
rect -8576 517934 592500 518018
rect -8576 517698 -7454 517934
rect -7218 517698 12786 517934
rect 13022 517698 48786 517934
rect 49022 517698 84786 517934
rect 85022 517698 120786 517934
rect 121022 517698 156786 517934
rect 157022 517698 192786 517934
rect 193022 517698 228786 517934
rect 229022 517698 264786 517934
rect 265022 517698 300786 517934
rect 301022 517698 336786 517934
rect 337022 517698 372786 517934
rect 373022 517698 408786 517934
rect 409022 517698 444786 517934
rect 445022 517698 480786 517934
rect 481022 517698 516786 517934
rect 517022 517698 552786 517934
rect 553022 517698 591142 517934
rect 591378 517698 592500 517934
rect -8576 517676 592500 517698
rect -7636 517674 -7036 517676
rect 12604 517674 13204 517676
rect 48604 517674 49204 517676
rect 84604 517674 85204 517676
rect 120604 517674 121204 517676
rect 156604 517674 157204 517676
rect 192604 517674 193204 517676
rect 228604 517674 229204 517676
rect 264604 517674 265204 517676
rect 300604 517674 301204 517676
rect 336604 517674 337204 517676
rect 372604 517674 373204 517676
rect 408604 517674 409204 517676
rect 444604 517674 445204 517676
rect 480604 517674 481204 517676
rect 516604 517674 517204 517676
rect 552604 517674 553204 517676
rect 590960 517674 591560 517676
rect -5756 514676 -5156 514678
rect 9004 514676 9604 514678
rect 45004 514676 45604 514678
rect 81004 514676 81604 514678
rect 117004 514676 117604 514678
rect 153004 514676 153604 514678
rect 189004 514676 189604 514678
rect 225004 514676 225604 514678
rect 261004 514676 261604 514678
rect 297004 514676 297604 514678
rect 333004 514676 333604 514678
rect 369004 514676 369604 514678
rect 405004 514676 405604 514678
rect 441004 514676 441604 514678
rect 477004 514676 477604 514678
rect 513004 514676 513604 514678
rect 549004 514676 549604 514678
rect 589080 514676 589680 514678
rect -6696 514654 590620 514676
rect -6696 514418 -5574 514654
rect -5338 514418 9186 514654
rect 9422 514418 45186 514654
rect 45422 514418 81186 514654
rect 81422 514418 117186 514654
rect 117422 514418 153186 514654
rect 153422 514418 189186 514654
rect 189422 514418 225186 514654
rect 225422 514418 261186 514654
rect 261422 514418 297186 514654
rect 297422 514418 333186 514654
rect 333422 514418 369186 514654
rect 369422 514418 405186 514654
rect 405422 514418 441186 514654
rect 441422 514418 477186 514654
rect 477422 514418 513186 514654
rect 513422 514418 549186 514654
rect 549422 514418 589262 514654
rect 589498 514418 590620 514654
rect -6696 514334 590620 514418
rect -6696 514098 -5574 514334
rect -5338 514098 9186 514334
rect 9422 514098 45186 514334
rect 45422 514098 81186 514334
rect 81422 514098 117186 514334
rect 117422 514098 153186 514334
rect 153422 514098 189186 514334
rect 189422 514098 225186 514334
rect 225422 514098 261186 514334
rect 261422 514098 297186 514334
rect 297422 514098 333186 514334
rect 333422 514098 369186 514334
rect 369422 514098 405186 514334
rect 405422 514098 441186 514334
rect 441422 514098 477186 514334
rect 477422 514098 513186 514334
rect 513422 514098 549186 514334
rect 549422 514098 589262 514334
rect 589498 514098 590620 514334
rect -6696 514076 590620 514098
rect -5756 514074 -5156 514076
rect 9004 514074 9604 514076
rect 45004 514074 45604 514076
rect 81004 514074 81604 514076
rect 117004 514074 117604 514076
rect 153004 514074 153604 514076
rect 189004 514074 189604 514076
rect 225004 514074 225604 514076
rect 261004 514074 261604 514076
rect 297004 514074 297604 514076
rect 333004 514074 333604 514076
rect 369004 514074 369604 514076
rect 405004 514074 405604 514076
rect 441004 514074 441604 514076
rect 477004 514074 477604 514076
rect 513004 514074 513604 514076
rect 549004 514074 549604 514076
rect 589080 514074 589680 514076
rect -3876 511076 -3276 511078
rect 5404 511076 6004 511078
rect 41404 511076 42004 511078
rect 77404 511076 78004 511078
rect 113404 511076 114004 511078
rect 149404 511076 150004 511078
rect 185404 511076 186004 511078
rect 221404 511076 222004 511078
rect 257404 511076 258004 511078
rect 293404 511076 294004 511078
rect 329404 511076 330004 511078
rect 365404 511076 366004 511078
rect 401404 511076 402004 511078
rect 437404 511076 438004 511078
rect 473404 511076 474004 511078
rect 509404 511076 510004 511078
rect 545404 511076 546004 511078
rect 581404 511076 582004 511078
rect 587200 511076 587800 511078
rect -4816 511054 588740 511076
rect -4816 510818 -3694 511054
rect -3458 510818 5586 511054
rect 5822 510818 41586 511054
rect 41822 510818 77586 511054
rect 77822 510818 113586 511054
rect 113822 510818 149586 511054
rect 149822 510818 185586 511054
rect 185822 510818 221586 511054
rect 221822 510818 257586 511054
rect 257822 510818 293586 511054
rect 293822 510818 329586 511054
rect 329822 510818 365586 511054
rect 365822 510818 401586 511054
rect 401822 510818 437586 511054
rect 437822 510818 473586 511054
rect 473822 510818 509586 511054
rect 509822 510818 545586 511054
rect 545822 510818 581586 511054
rect 581822 510818 587382 511054
rect 587618 510818 588740 511054
rect -4816 510734 588740 510818
rect -4816 510498 -3694 510734
rect -3458 510498 5586 510734
rect 5822 510498 41586 510734
rect 41822 510498 77586 510734
rect 77822 510498 113586 510734
rect 113822 510498 149586 510734
rect 149822 510498 185586 510734
rect 185822 510498 221586 510734
rect 221822 510498 257586 510734
rect 257822 510498 293586 510734
rect 293822 510498 329586 510734
rect 329822 510498 365586 510734
rect 365822 510498 401586 510734
rect 401822 510498 437586 510734
rect 437822 510498 473586 510734
rect 473822 510498 509586 510734
rect 509822 510498 545586 510734
rect 545822 510498 581586 510734
rect 581822 510498 587382 510734
rect 587618 510498 588740 510734
rect -4816 510476 588740 510498
rect -3876 510474 -3276 510476
rect 5404 510474 6004 510476
rect 41404 510474 42004 510476
rect 77404 510474 78004 510476
rect 113404 510474 114004 510476
rect 149404 510474 150004 510476
rect 185404 510474 186004 510476
rect 221404 510474 222004 510476
rect 257404 510474 258004 510476
rect 293404 510474 294004 510476
rect 329404 510474 330004 510476
rect 365404 510474 366004 510476
rect 401404 510474 402004 510476
rect 437404 510474 438004 510476
rect 473404 510474 474004 510476
rect 509404 510474 510004 510476
rect 545404 510474 546004 510476
rect 581404 510474 582004 510476
rect 587200 510474 587800 510476
rect -1996 507476 -1396 507478
rect 1804 507476 2404 507478
rect 37804 507476 38404 507478
rect 73804 507476 74404 507478
rect 109804 507476 110404 507478
rect 145804 507476 146404 507478
rect 181804 507476 182404 507478
rect 217804 507476 218404 507478
rect 253804 507476 254404 507478
rect 289804 507476 290404 507478
rect 325804 507476 326404 507478
rect 361804 507476 362404 507478
rect 397804 507476 398404 507478
rect 433804 507476 434404 507478
rect 469804 507476 470404 507478
rect 505804 507476 506404 507478
rect 541804 507476 542404 507478
rect 577804 507476 578404 507478
rect 585320 507476 585920 507478
rect -2936 507454 586860 507476
rect -2936 507218 -1814 507454
rect -1578 507218 1986 507454
rect 2222 507218 37986 507454
rect 38222 507218 73986 507454
rect 74222 507218 109986 507454
rect 110222 507218 145986 507454
rect 146222 507218 181986 507454
rect 182222 507218 217986 507454
rect 218222 507218 253986 507454
rect 254222 507218 289986 507454
rect 290222 507218 325986 507454
rect 326222 507218 361986 507454
rect 362222 507218 397986 507454
rect 398222 507218 433986 507454
rect 434222 507218 469986 507454
rect 470222 507218 505986 507454
rect 506222 507218 541986 507454
rect 542222 507218 577986 507454
rect 578222 507218 585502 507454
rect 585738 507218 586860 507454
rect -2936 507134 586860 507218
rect -2936 506898 -1814 507134
rect -1578 506898 1986 507134
rect 2222 506898 37986 507134
rect 38222 506898 73986 507134
rect 74222 506898 109986 507134
rect 110222 506898 145986 507134
rect 146222 506898 181986 507134
rect 182222 506898 217986 507134
rect 218222 506898 253986 507134
rect 254222 506898 289986 507134
rect 290222 506898 325986 507134
rect 326222 506898 361986 507134
rect 362222 506898 397986 507134
rect 398222 506898 433986 507134
rect 434222 506898 469986 507134
rect 470222 506898 505986 507134
rect 506222 506898 541986 507134
rect 542222 506898 577986 507134
rect 578222 506898 585502 507134
rect 585738 506898 586860 507134
rect -2936 506876 586860 506898
rect -1996 506874 -1396 506876
rect 1804 506874 2404 506876
rect 37804 506874 38404 506876
rect 73804 506874 74404 506876
rect 109804 506874 110404 506876
rect 145804 506874 146404 506876
rect 181804 506874 182404 506876
rect 217804 506874 218404 506876
rect 253804 506874 254404 506876
rect 289804 506874 290404 506876
rect 325804 506874 326404 506876
rect 361804 506874 362404 506876
rect 397804 506874 398404 506876
rect 433804 506874 434404 506876
rect 469804 506874 470404 506876
rect 505804 506874 506404 506876
rect 541804 506874 542404 506876
rect 577804 506874 578404 506876
rect 585320 506874 585920 506876
rect -8576 500276 -7976 500278
rect 30604 500276 31204 500278
rect 66604 500276 67204 500278
rect 102604 500276 103204 500278
rect 138604 500276 139204 500278
rect 174604 500276 175204 500278
rect 210604 500276 211204 500278
rect 246604 500276 247204 500278
rect 282604 500276 283204 500278
rect 318604 500276 319204 500278
rect 354604 500276 355204 500278
rect 390604 500276 391204 500278
rect 426604 500276 427204 500278
rect 462604 500276 463204 500278
rect 498604 500276 499204 500278
rect 534604 500276 535204 500278
rect 570604 500276 571204 500278
rect 591900 500276 592500 500278
rect -8576 500254 592500 500276
rect -8576 500018 -8394 500254
rect -8158 500018 30786 500254
rect 31022 500018 66786 500254
rect 67022 500018 102786 500254
rect 103022 500018 138786 500254
rect 139022 500018 174786 500254
rect 175022 500018 210786 500254
rect 211022 500018 246786 500254
rect 247022 500018 282786 500254
rect 283022 500018 318786 500254
rect 319022 500018 354786 500254
rect 355022 500018 390786 500254
rect 391022 500018 426786 500254
rect 427022 500018 462786 500254
rect 463022 500018 498786 500254
rect 499022 500018 534786 500254
rect 535022 500018 570786 500254
rect 571022 500018 592082 500254
rect 592318 500018 592500 500254
rect -8576 499934 592500 500018
rect -8576 499698 -8394 499934
rect -8158 499698 30786 499934
rect 31022 499698 66786 499934
rect 67022 499698 102786 499934
rect 103022 499698 138786 499934
rect 139022 499698 174786 499934
rect 175022 499698 210786 499934
rect 211022 499698 246786 499934
rect 247022 499698 282786 499934
rect 283022 499698 318786 499934
rect 319022 499698 354786 499934
rect 355022 499698 390786 499934
rect 391022 499698 426786 499934
rect 427022 499698 462786 499934
rect 463022 499698 498786 499934
rect 499022 499698 534786 499934
rect 535022 499698 570786 499934
rect 571022 499698 592082 499934
rect 592318 499698 592500 499934
rect -8576 499676 592500 499698
rect -8576 499674 -7976 499676
rect 30604 499674 31204 499676
rect 66604 499674 67204 499676
rect 102604 499674 103204 499676
rect 138604 499674 139204 499676
rect 174604 499674 175204 499676
rect 210604 499674 211204 499676
rect 246604 499674 247204 499676
rect 282604 499674 283204 499676
rect 318604 499674 319204 499676
rect 354604 499674 355204 499676
rect 390604 499674 391204 499676
rect 426604 499674 427204 499676
rect 462604 499674 463204 499676
rect 498604 499674 499204 499676
rect 534604 499674 535204 499676
rect 570604 499674 571204 499676
rect 591900 499674 592500 499676
rect -6696 496676 -6096 496678
rect 27004 496676 27604 496678
rect 63004 496676 63604 496678
rect 99004 496676 99604 496678
rect 135004 496676 135604 496678
rect 171004 496676 171604 496678
rect 207004 496676 207604 496678
rect 243004 496676 243604 496678
rect 279004 496676 279604 496678
rect 315004 496676 315604 496678
rect 351004 496676 351604 496678
rect 387004 496676 387604 496678
rect 423004 496676 423604 496678
rect 459004 496676 459604 496678
rect 495004 496676 495604 496678
rect 531004 496676 531604 496678
rect 567004 496676 567604 496678
rect 590020 496676 590620 496678
rect -6696 496654 590620 496676
rect -6696 496418 -6514 496654
rect -6278 496418 27186 496654
rect 27422 496418 63186 496654
rect 63422 496418 99186 496654
rect 99422 496418 135186 496654
rect 135422 496418 171186 496654
rect 171422 496418 207186 496654
rect 207422 496418 243186 496654
rect 243422 496418 279186 496654
rect 279422 496418 315186 496654
rect 315422 496418 351186 496654
rect 351422 496418 387186 496654
rect 387422 496418 423186 496654
rect 423422 496418 459186 496654
rect 459422 496418 495186 496654
rect 495422 496418 531186 496654
rect 531422 496418 567186 496654
rect 567422 496418 590202 496654
rect 590438 496418 590620 496654
rect -6696 496334 590620 496418
rect -6696 496098 -6514 496334
rect -6278 496098 27186 496334
rect 27422 496098 63186 496334
rect 63422 496098 99186 496334
rect 99422 496098 135186 496334
rect 135422 496098 171186 496334
rect 171422 496098 207186 496334
rect 207422 496098 243186 496334
rect 243422 496098 279186 496334
rect 279422 496098 315186 496334
rect 315422 496098 351186 496334
rect 351422 496098 387186 496334
rect 387422 496098 423186 496334
rect 423422 496098 459186 496334
rect 459422 496098 495186 496334
rect 495422 496098 531186 496334
rect 531422 496098 567186 496334
rect 567422 496098 590202 496334
rect 590438 496098 590620 496334
rect -6696 496076 590620 496098
rect -6696 496074 -6096 496076
rect 27004 496074 27604 496076
rect 63004 496074 63604 496076
rect 99004 496074 99604 496076
rect 135004 496074 135604 496076
rect 171004 496074 171604 496076
rect 207004 496074 207604 496076
rect 243004 496074 243604 496076
rect 279004 496074 279604 496076
rect 315004 496074 315604 496076
rect 351004 496074 351604 496076
rect 387004 496074 387604 496076
rect 423004 496074 423604 496076
rect 459004 496074 459604 496076
rect 495004 496074 495604 496076
rect 531004 496074 531604 496076
rect 567004 496074 567604 496076
rect 590020 496074 590620 496076
rect -4816 493076 -4216 493078
rect 23404 493076 24004 493078
rect 59404 493076 60004 493078
rect 95404 493076 96004 493078
rect 131404 493076 132004 493078
rect 167404 493076 168004 493078
rect 203404 493076 204004 493078
rect 239404 493076 240004 493078
rect 275404 493076 276004 493078
rect 311404 493076 312004 493078
rect 347404 493076 348004 493078
rect 383404 493076 384004 493078
rect 419404 493076 420004 493078
rect 455404 493076 456004 493078
rect 491404 493076 492004 493078
rect 527404 493076 528004 493078
rect 563404 493076 564004 493078
rect 588140 493076 588740 493078
rect -4816 493054 588740 493076
rect -4816 492818 -4634 493054
rect -4398 492818 23586 493054
rect 23822 492818 59586 493054
rect 59822 492818 95586 493054
rect 95822 492818 131586 493054
rect 131822 492818 167586 493054
rect 167822 492818 203586 493054
rect 203822 492818 239586 493054
rect 239822 492818 275586 493054
rect 275822 492818 311586 493054
rect 311822 492818 347586 493054
rect 347822 492818 383586 493054
rect 383822 492818 419586 493054
rect 419822 492818 455586 493054
rect 455822 492818 491586 493054
rect 491822 492818 527586 493054
rect 527822 492818 563586 493054
rect 563822 492818 588322 493054
rect 588558 492818 588740 493054
rect -4816 492734 588740 492818
rect -4816 492498 -4634 492734
rect -4398 492498 23586 492734
rect 23822 492498 59586 492734
rect 59822 492498 95586 492734
rect 95822 492498 131586 492734
rect 131822 492498 167586 492734
rect 167822 492498 203586 492734
rect 203822 492498 239586 492734
rect 239822 492498 275586 492734
rect 275822 492498 311586 492734
rect 311822 492498 347586 492734
rect 347822 492498 383586 492734
rect 383822 492498 419586 492734
rect 419822 492498 455586 492734
rect 455822 492498 491586 492734
rect 491822 492498 527586 492734
rect 527822 492498 563586 492734
rect 563822 492498 588322 492734
rect 588558 492498 588740 492734
rect -4816 492476 588740 492498
rect -4816 492474 -4216 492476
rect 23404 492474 24004 492476
rect 59404 492474 60004 492476
rect 95404 492474 96004 492476
rect 131404 492474 132004 492476
rect 167404 492474 168004 492476
rect 203404 492474 204004 492476
rect 239404 492474 240004 492476
rect 275404 492474 276004 492476
rect 311404 492474 312004 492476
rect 347404 492474 348004 492476
rect 383404 492474 384004 492476
rect 419404 492474 420004 492476
rect 455404 492474 456004 492476
rect 491404 492474 492004 492476
rect 527404 492474 528004 492476
rect 563404 492474 564004 492476
rect 588140 492474 588740 492476
rect -2936 489476 -2336 489478
rect 19804 489476 20404 489478
rect 55804 489476 56404 489478
rect 91804 489476 92404 489478
rect 127804 489476 128404 489478
rect 163804 489476 164404 489478
rect 199804 489476 200404 489478
rect 235804 489476 236404 489478
rect 271804 489476 272404 489478
rect 307804 489476 308404 489478
rect 343804 489476 344404 489478
rect 379804 489476 380404 489478
rect 415804 489476 416404 489478
rect 451804 489476 452404 489478
rect 487804 489476 488404 489478
rect 523804 489476 524404 489478
rect 559804 489476 560404 489478
rect 586260 489476 586860 489478
rect -2936 489454 586860 489476
rect -2936 489218 -2754 489454
rect -2518 489218 19986 489454
rect 20222 489218 55986 489454
rect 56222 489218 91986 489454
rect 92222 489218 127986 489454
rect 128222 489218 163986 489454
rect 164222 489218 199986 489454
rect 200222 489218 235986 489454
rect 236222 489218 271986 489454
rect 272222 489218 307986 489454
rect 308222 489218 343986 489454
rect 344222 489218 379986 489454
rect 380222 489218 415986 489454
rect 416222 489218 451986 489454
rect 452222 489218 487986 489454
rect 488222 489218 523986 489454
rect 524222 489218 559986 489454
rect 560222 489218 586442 489454
rect 586678 489218 586860 489454
rect -2936 489134 586860 489218
rect -2936 488898 -2754 489134
rect -2518 488898 19986 489134
rect 20222 488898 55986 489134
rect 56222 488898 91986 489134
rect 92222 488898 127986 489134
rect 128222 488898 163986 489134
rect 164222 488898 199986 489134
rect 200222 488898 235986 489134
rect 236222 488898 271986 489134
rect 272222 488898 307986 489134
rect 308222 488898 343986 489134
rect 344222 488898 379986 489134
rect 380222 488898 415986 489134
rect 416222 488898 451986 489134
rect 452222 488898 487986 489134
rect 488222 488898 523986 489134
rect 524222 488898 559986 489134
rect 560222 488898 586442 489134
rect 586678 488898 586860 489134
rect -2936 488876 586860 488898
rect -2936 488874 -2336 488876
rect 19804 488874 20404 488876
rect 55804 488874 56404 488876
rect 91804 488874 92404 488876
rect 127804 488874 128404 488876
rect 163804 488874 164404 488876
rect 199804 488874 200404 488876
rect 235804 488874 236404 488876
rect 271804 488874 272404 488876
rect 307804 488874 308404 488876
rect 343804 488874 344404 488876
rect 379804 488874 380404 488876
rect 415804 488874 416404 488876
rect 451804 488874 452404 488876
rect 487804 488874 488404 488876
rect 523804 488874 524404 488876
rect 559804 488874 560404 488876
rect 586260 488874 586860 488876
rect -7636 482276 -7036 482278
rect 12604 482276 13204 482278
rect 48604 482276 49204 482278
rect 84604 482276 85204 482278
rect 120604 482276 121204 482278
rect 156604 482276 157204 482278
rect 192604 482276 193204 482278
rect 228604 482276 229204 482278
rect 264604 482276 265204 482278
rect 300604 482276 301204 482278
rect 336604 482276 337204 482278
rect 372604 482276 373204 482278
rect 408604 482276 409204 482278
rect 444604 482276 445204 482278
rect 480604 482276 481204 482278
rect 516604 482276 517204 482278
rect 552604 482276 553204 482278
rect 590960 482276 591560 482278
rect -8576 482254 592500 482276
rect -8576 482018 -7454 482254
rect -7218 482018 12786 482254
rect 13022 482018 48786 482254
rect 49022 482018 84786 482254
rect 85022 482018 120786 482254
rect 121022 482018 156786 482254
rect 157022 482018 192786 482254
rect 193022 482018 228786 482254
rect 229022 482018 264786 482254
rect 265022 482018 300786 482254
rect 301022 482018 336786 482254
rect 337022 482018 372786 482254
rect 373022 482018 408786 482254
rect 409022 482018 444786 482254
rect 445022 482018 480786 482254
rect 481022 482018 516786 482254
rect 517022 482018 552786 482254
rect 553022 482018 591142 482254
rect 591378 482018 592500 482254
rect -8576 481934 592500 482018
rect -8576 481698 -7454 481934
rect -7218 481698 12786 481934
rect 13022 481698 48786 481934
rect 49022 481698 84786 481934
rect 85022 481698 120786 481934
rect 121022 481698 156786 481934
rect 157022 481698 192786 481934
rect 193022 481698 228786 481934
rect 229022 481698 264786 481934
rect 265022 481698 300786 481934
rect 301022 481698 336786 481934
rect 337022 481698 372786 481934
rect 373022 481698 408786 481934
rect 409022 481698 444786 481934
rect 445022 481698 480786 481934
rect 481022 481698 516786 481934
rect 517022 481698 552786 481934
rect 553022 481698 591142 481934
rect 591378 481698 592500 481934
rect -8576 481676 592500 481698
rect -7636 481674 -7036 481676
rect 12604 481674 13204 481676
rect 48604 481674 49204 481676
rect 84604 481674 85204 481676
rect 120604 481674 121204 481676
rect 156604 481674 157204 481676
rect 192604 481674 193204 481676
rect 228604 481674 229204 481676
rect 264604 481674 265204 481676
rect 300604 481674 301204 481676
rect 336604 481674 337204 481676
rect 372604 481674 373204 481676
rect 408604 481674 409204 481676
rect 444604 481674 445204 481676
rect 480604 481674 481204 481676
rect 516604 481674 517204 481676
rect 552604 481674 553204 481676
rect 590960 481674 591560 481676
rect -5756 478676 -5156 478678
rect 9004 478676 9604 478678
rect 45004 478676 45604 478678
rect 81004 478676 81604 478678
rect 117004 478676 117604 478678
rect 153004 478676 153604 478678
rect 189004 478676 189604 478678
rect 225004 478676 225604 478678
rect 261004 478676 261604 478678
rect 297004 478676 297604 478678
rect 333004 478676 333604 478678
rect 369004 478676 369604 478678
rect 405004 478676 405604 478678
rect 441004 478676 441604 478678
rect 477004 478676 477604 478678
rect 513004 478676 513604 478678
rect 549004 478676 549604 478678
rect 589080 478676 589680 478678
rect -6696 478654 590620 478676
rect -6696 478418 -5574 478654
rect -5338 478418 9186 478654
rect 9422 478418 45186 478654
rect 45422 478418 81186 478654
rect 81422 478418 117186 478654
rect 117422 478418 153186 478654
rect 153422 478418 189186 478654
rect 189422 478418 225186 478654
rect 225422 478418 261186 478654
rect 261422 478418 297186 478654
rect 297422 478418 333186 478654
rect 333422 478418 369186 478654
rect 369422 478418 405186 478654
rect 405422 478418 441186 478654
rect 441422 478418 477186 478654
rect 477422 478418 513186 478654
rect 513422 478418 549186 478654
rect 549422 478418 589262 478654
rect 589498 478418 590620 478654
rect -6696 478334 590620 478418
rect -6696 478098 -5574 478334
rect -5338 478098 9186 478334
rect 9422 478098 45186 478334
rect 45422 478098 81186 478334
rect 81422 478098 117186 478334
rect 117422 478098 153186 478334
rect 153422 478098 189186 478334
rect 189422 478098 225186 478334
rect 225422 478098 261186 478334
rect 261422 478098 297186 478334
rect 297422 478098 333186 478334
rect 333422 478098 369186 478334
rect 369422 478098 405186 478334
rect 405422 478098 441186 478334
rect 441422 478098 477186 478334
rect 477422 478098 513186 478334
rect 513422 478098 549186 478334
rect 549422 478098 589262 478334
rect 589498 478098 590620 478334
rect -6696 478076 590620 478098
rect -5756 478074 -5156 478076
rect 9004 478074 9604 478076
rect 45004 478074 45604 478076
rect 81004 478074 81604 478076
rect 117004 478074 117604 478076
rect 153004 478074 153604 478076
rect 189004 478074 189604 478076
rect 225004 478074 225604 478076
rect 261004 478074 261604 478076
rect 297004 478074 297604 478076
rect 333004 478074 333604 478076
rect 369004 478074 369604 478076
rect 405004 478074 405604 478076
rect 441004 478074 441604 478076
rect 477004 478074 477604 478076
rect 513004 478074 513604 478076
rect 549004 478074 549604 478076
rect 589080 478074 589680 478076
rect -3876 475076 -3276 475078
rect 5404 475076 6004 475078
rect 41404 475076 42004 475078
rect 77404 475076 78004 475078
rect 113404 475076 114004 475078
rect 149404 475076 150004 475078
rect 185404 475076 186004 475078
rect 221404 475076 222004 475078
rect 257404 475076 258004 475078
rect 293404 475076 294004 475078
rect 329404 475076 330004 475078
rect 365404 475076 366004 475078
rect 401404 475076 402004 475078
rect 437404 475076 438004 475078
rect 473404 475076 474004 475078
rect 509404 475076 510004 475078
rect 545404 475076 546004 475078
rect 581404 475076 582004 475078
rect 587200 475076 587800 475078
rect -4816 475054 588740 475076
rect -4816 474818 -3694 475054
rect -3458 474818 5586 475054
rect 5822 474818 41586 475054
rect 41822 474818 77586 475054
rect 77822 474818 113586 475054
rect 113822 474818 149586 475054
rect 149822 474818 185586 475054
rect 185822 474818 221586 475054
rect 221822 474818 257586 475054
rect 257822 474818 293586 475054
rect 293822 474818 329586 475054
rect 329822 474818 365586 475054
rect 365822 474818 401586 475054
rect 401822 474818 437586 475054
rect 437822 474818 473586 475054
rect 473822 474818 509586 475054
rect 509822 474818 545586 475054
rect 545822 474818 581586 475054
rect 581822 474818 587382 475054
rect 587618 474818 588740 475054
rect -4816 474734 588740 474818
rect -4816 474498 -3694 474734
rect -3458 474498 5586 474734
rect 5822 474498 41586 474734
rect 41822 474498 77586 474734
rect 77822 474498 113586 474734
rect 113822 474498 149586 474734
rect 149822 474498 185586 474734
rect 185822 474498 221586 474734
rect 221822 474498 257586 474734
rect 257822 474498 293586 474734
rect 293822 474498 329586 474734
rect 329822 474498 365586 474734
rect 365822 474498 401586 474734
rect 401822 474498 437586 474734
rect 437822 474498 473586 474734
rect 473822 474498 509586 474734
rect 509822 474498 545586 474734
rect 545822 474498 581586 474734
rect 581822 474498 587382 474734
rect 587618 474498 588740 474734
rect -4816 474476 588740 474498
rect -3876 474474 -3276 474476
rect 5404 474474 6004 474476
rect 41404 474474 42004 474476
rect 77404 474474 78004 474476
rect 113404 474474 114004 474476
rect 149404 474474 150004 474476
rect 185404 474474 186004 474476
rect 221404 474474 222004 474476
rect 257404 474474 258004 474476
rect 293404 474474 294004 474476
rect 329404 474474 330004 474476
rect 365404 474474 366004 474476
rect 401404 474474 402004 474476
rect 437404 474474 438004 474476
rect 473404 474474 474004 474476
rect 509404 474474 510004 474476
rect 545404 474474 546004 474476
rect 581404 474474 582004 474476
rect 587200 474474 587800 474476
rect -1996 471476 -1396 471478
rect 1804 471476 2404 471478
rect 37804 471476 38404 471478
rect 73804 471476 74404 471478
rect 109804 471476 110404 471478
rect 145804 471476 146404 471478
rect 181804 471476 182404 471478
rect 217804 471476 218404 471478
rect 253804 471476 254404 471478
rect 289804 471476 290404 471478
rect 325804 471476 326404 471478
rect 361804 471476 362404 471478
rect 397804 471476 398404 471478
rect 433804 471476 434404 471478
rect 469804 471476 470404 471478
rect 505804 471476 506404 471478
rect 541804 471476 542404 471478
rect 577804 471476 578404 471478
rect 585320 471476 585920 471478
rect -2936 471454 586860 471476
rect -2936 471218 -1814 471454
rect -1578 471218 1986 471454
rect 2222 471218 37986 471454
rect 38222 471218 73986 471454
rect 74222 471218 109986 471454
rect 110222 471218 145986 471454
rect 146222 471218 181986 471454
rect 182222 471218 217986 471454
rect 218222 471218 253986 471454
rect 254222 471218 289986 471454
rect 290222 471218 325986 471454
rect 326222 471218 361986 471454
rect 362222 471218 397986 471454
rect 398222 471218 433986 471454
rect 434222 471218 469986 471454
rect 470222 471218 505986 471454
rect 506222 471218 541986 471454
rect 542222 471218 577986 471454
rect 578222 471218 585502 471454
rect 585738 471218 586860 471454
rect -2936 471134 586860 471218
rect -2936 470898 -1814 471134
rect -1578 470898 1986 471134
rect 2222 470898 37986 471134
rect 38222 470898 73986 471134
rect 74222 470898 109986 471134
rect 110222 470898 145986 471134
rect 146222 470898 181986 471134
rect 182222 470898 217986 471134
rect 218222 470898 253986 471134
rect 254222 470898 289986 471134
rect 290222 470898 325986 471134
rect 326222 470898 361986 471134
rect 362222 470898 397986 471134
rect 398222 470898 433986 471134
rect 434222 470898 469986 471134
rect 470222 470898 505986 471134
rect 506222 470898 541986 471134
rect 542222 470898 577986 471134
rect 578222 470898 585502 471134
rect 585738 470898 586860 471134
rect -2936 470876 586860 470898
rect -1996 470874 -1396 470876
rect 1804 470874 2404 470876
rect 37804 470874 38404 470876
rect 73804 470874 74404 470876
rect 109804 470874 110404 470876
rect 145804 470874 146404 470876
rect 181804 470874 182404 470876
rect 217804 470874 218404 470876
rect 253804 470874 254404 470876
rect 289804 470874 290404 470876
rect 325804 470874 326404 470876
rect 361804 470874 362404 470876
rect 397804 470874 398404 470876
rect 433804 470874 434404 470876
rect 469804 470874 470404 470876
rect 505804 470874 506404 470876
rect 541804 470874 542404 470876
rect 577804 470874 578404 470876
rect 585320 470874 585920 470876
rect -8576 464276 -7976 464278
rect 30604 464276 31204 464278
rect 66604 464276 67204 464278
rect 102604 464276 103204 464278
rect 138604 464276 139204 464278
rect 174604 464276 175204 464278
rect 210604 464276 211204 464278
rect 246604 464276 247204 464278
rect 282604 464276 283204 464278
rect 318604 464276 319204 464278
rect 354604 464276 355204 464278
rect 390604 464276 391204 464278
rect 426604 464276 427204 464278
rect 462604 464276 463204 464278
rect 498604 464276 499204 464278
rect 534604 464276 535204 464278
rect 570604 464276 571204 464278
rect 591900 464276 592500 464278
rect -8576 464254 592500 464276
rect -8576 464018 -8394 464254
rect -8158 464018 30786 464254
rect 31022 464018 66786 464254
rect 67022 464018 102786 464254
rect 103022 464018 138786 464254
rect 139022 464018 174786 464254
rect 175022 464018 210786 464254
rect 211022 464018 246786 464254
rect 247022 464018 282786 464254
rect 283022 464018 318786 464254
rect 319022 464018 354786 464254
rect 355022 464018 390786 464254
rect 391022 464018 426786 464254
rect 427022 464018 462786 464254
rect 463022 464018 498786 464254
rect 499022 464018 534786 464254
rect 535022 464018 570786 464254
rect 571022 464018 592082 464254
rect 592318 464018 592500 464254
rect -8576 463934 592500 464018
rect -8576 463698 -8394 463934
rect -8158 463698 30786 463934
rect 31022 463698 66786 463934
rect 67022 463698 102786 463934
rect 103022 463698 138786 463934
rect 139022 463698 174786 463934
rect 175022 463698 210786 463934
rect 211022 463698 246786 463934
rect 247022 463698 282786 463934
rect 283022 463698 318786 463934
rect 319022 463698 354786 463934
rect 355022 463698 390786 463934
rect 391022 463698 426786 463934
rect 427022 463698 462786 463934
rect 463022 463698 498786 463934
rect 499022 463698 534786 463934
rect 535022 463698 570786 463934
rect 571022 463698 592082 463934
rect 592318 463698 592500 463934
rect -8576 463676 592500 463698
rect -8576 463674 -7976 463676
rect 30604 463674 31204 463676
rect 66604 463674 67204 463676
rect 102604 463674 103204 463676
rect 138604 463674 139204 463676
rect 174604 463674 175204 463676
rect 210604 463674 211204 463676
rect 246604 463674 247204 463676
rect 282604 463674 283204 463676
rect 318604 463674 319204 463676
rect 354604 463674 355204 463676
rect 390604 463674 391204 463676
rect 426604 463674 427204 463676
rect 462604 463674 463204 463676
rect 498604 463674 499204 463676
rect 534604 463674 535204 463676
rect 570604 463674 571204 463676
rect 591900 463674 592500 463676
rect -6696 460676 -6096 460678
rect 27004 460676 27604 460678
rect 63004 460676 63604 460678
rect 99004 460676 99604 460678
rect 135004 460676 135604 460678
rect 171004 460676 171604 460678
rect 207004 460676 207604 460678
rect 243004 460676 243604 460678
rect 279004 460676 279604 460678
rect 315004 460676 315604 460678
rect 351004 460676 351604 460678
rect 387004 460676 387604 460678
rect 423004 460676 423604 460678
rect 459004 460676 459604 460678
rect 495004 460676 495604 460678
rect 531004 460676 531604 460678
rect 567004 460676 567604 460678
rect 590020 460676 590620 460678
rect -6696 460654 590620 460676
rect -6696 460418 -6514 460654
rect -6278 460418 27186 460654
rect 27422 460418 63186 460654
rect 63422 460418 99186 460654
rect 99422 460418 135186 460654
rect 135422 460418 171186 460654
rect 171422 460418 207186 460654
rect 207422 460418 243186 460654
rect 243422 460418 279186 460654
rect 279422 460418 315186 460654
rect 315422 460418 351186 460654
rect 351422 460418 387186 460654
rect 387422 460418 423186 460654
rect 423422 460418 459186 460654
rect 459422 460418 495186 460654
rect 495422 460418 531186 460654
rect 531422 460418 567186 460654
rect 567422 460418 590202 460654
rect 590438 460418 590620 460654
rect -6696 460334 590620 460418
rect -6696 460098 -6514 460334
rect -6278 460098 27186 460334
rect 27422 460098 63186 460334
rect 63422 460098 99186 460334
rect 99422 460098 135186 460334
rect 135422 460098 171186 460334
rect 171422 460098 207186 460334
rect 207422 460098 243186 460334
rect 243422 460098 279186 460334
rect 279422 460098 315186 460334
rect 315422 460098 351186 460334
rect 351422 460098 387186 460334
rect 387422 460098 423186 460334
rect 423422 460098 459186 460334
rect 459422 460098 495186 460334
rect 495422 460098 531186 460334
rect 531422 460098 567186 460334
rect 567422 460098 590202 460334
rect 590438 460098 590620 460334
rect -6696 460076 590620 460098
rect -6696 460074 -6096 460076
rect 27004 460074 27604 460076
rect 63004 460074 63604 460076
rect 99004 460074 99604 460076
rect 135004 460074 135604 460076
rect 171004 460074 171604 460076
rect 207004 460074 207604 460076
rect 243004 460074 243604 460076
rect 279004 460074 279604 460076
rect 315004 460074 315604 460076
rect 351004 460074 351604 460076
rect 387004 460074 387604 460076
rect 423004 460074 423604 460076
rect 459004 460074 459604 460076
rect 495004 460074 495604 460076
rect 531004 460074 531604 460076
rect 567004 460074 567604 460076
rect 590020 460074 590620 460076
rect -4816 457076 -4216 457078
rect 23404 457076 24004 457078
rect 59404 457076 60004 457078
rect 95404 457076 96004 457078
rect 131404 457076 132004 457078
rect 167404 457076 168004 457078
rect 203404 457076 204004 457078
rect 239404 457076 240004 457078
rect 275404 457076 276004 457078
rect 311404 457076 312004 457078
rect 347404 457076 348004 457078
rect 383404 457076 384004 457078
rect 419404 457076 420004 457078
rect 455404 457076 456004 457078
rect 491404 457076 492004 457078
rect 527404 457076 528004 457078
rect 563404 457076 564004 457078
rect 588140 457076 588740 457078
rect -4816 457054 588740 457076
rect -4816 456818 -4634 457054
rect -4398 456818 23586 457054
rect 23822 456818 59586 457054
rect 59822 456818 95586 457054
rect 95822 456818 131586 457054
rect 131822 456818 167586 457054
rect 167822 456818 203586 457054
rect 203822 456818 239586 457054
rect 239822 456818 275586 457054
rect 275822 456818 311586 457054
rect 311822 456818 347586 457054
rect 347822 456818 383586 457054
rect 383822 456818 419586 457054
rect 419822 456818 455586 457054
rect 455822 456818 491586 457054
rect 491822 456818 527586 457054
rect 527822 456818 563586 457054
rect 563822 456818 588322 457054
rect 588558 456818 588740 457054
rect -4816 456734 588740 456818
rect -4816 456498 -4634 456734
rect -4398 456498 23586 456734
rect 23822 456498 59586 456734
rect 59822 456498 95586 456734
rect 95822 456498 131586 456734
rect 131822 456498 167586 456734
rect 167822 456498 203586 456734
rect 203822 456498 239586 456734
rect 239822 456498 275586 456734
rect 275822 456498 311586 456734
rect 311822 456498 347586 456734
rect 347822 456498 383586 456734
rect 383822 456498 419586 456734
rect 419822 456498 455586 456734
rect 455822 456498 491586 456734
rect 491822 456498 527586 456734
rect 527822 456498 563586 456734
rect 563822 456498 588322 456734
rect 588558 456498 588740 456734
rect -4816 456476 588740 456498
rect -4816 456474 -4216 456476
rect 23404 456474 24004 456476
rect 59404 456474 60004 456476
rect 95404 456474 96004 456476
rect 131404 456474 132004 456476
rect 167404 456474 168004 456476
rect 203404 456474 204004 456476
rect 239404 456474 240004 456476
rect 275404 456474 276004 456476
rect 311404 456474 312004 456476
rect 347404 456474 348004 456476
rect 383404 456474 384004 456476
rect 419404 456474 420004 456476
rect 455404 456474 456004 456476
rect 491404 456474 492004 456476
rect 527404 456474 528004 456476
rect 563404 456474 564004 456476
rect 588140 456474 588740 456476
rect -2936 453476 -2336 453478
rect 19804 453476 20404 453478
rect 55804 453476 56404 453478
rect 91804 453476 92404 453478
rect 127804 453476 128404 453478
rect 163804 453476 164404 453478
rect 199804 453476 200404 453478
rect 235804 453476 236404 453478
rect 271804 453476 272404 453478
rect 307804 453476 308404 453478
rect 343804 453476 344404 453478
rect 379804 453476 380404 453478
rect 415804 453476 416404 453478
rect 451804 453476 452404 453478
rect 487804 453476 488404 453478
rect 523804 453476 524404 453478
rect 559804 453476 560404 453478
rect 586260 453476 586860 453478
rect -2936 453454 586860 453476
rect -2936 453218 -2754 453454
rect -2518 453218 19986 453454
rect 20222 453218 55986 453454
rect 56222 453218 91986 453454
rect 92222 453218 127986 453454
rect 128222 453218 163986 453454
rect 164222 453218 199986 453454
rect 200222 453218 235986 453454
rect 236222 453218 271986 453454
rect 272222 453218 307986 453454
rect 308222 453218 343986 453454
rect 344222 453218 379986 453454
rect 380222 453218 415986 453454
rect 416222 453218 451986 453454
rect 452222 453218 487986 453454
rect 488222 453218 523986 453454
rect 524222 453218 559986 453454
rect 560222 453218 586442 453454
rect 586678 453218 586860 453454
rect -2936 453134 586860 453218
rect -2936 452898 -2754 453134
rect -2518 452898 19986 453134
rect 20222 452898 55986 453134
rect 56222 452898 91986 453134
rect 92222 452898 127986 453134
rect 128222 452898 163986 453134
rect 164222 452898 199986 453134
rect 200222 452898 235986 453134
rect 236222 452898 271986 453134
rect 272222 452898 307986 453134
rect 308222 452898 343986 453134
rect 344222 452898 379986 453134
rect 380222 452898 415986 453134
rect 416222 452898 451986 453134
rect 452222 452898 487986 453134
rect 488222 452898 523986 453134
rect 524222 452898 559986 453134
rect 560222 452898 586442 453134
rect 586678 452898 586860 453134
rect -2936 452876 586860 452898
rect -2936 452874 -2336 452876
rect 19804 452874 20404 452876
rect 55804 452874 56404 452876
rect 91804 452874 92404 452876
rect 127804 452874 128404 452876
rect 163804 452874 164404 452876
rect 199804 452874 200404 452876
rect 235804 452874 236404 452876
rect 271804 452874 272404 452876
rect 307804 452874 308404 452876
rect 343804 452874 344404 452876
rect 379804 452874 380404 452876
rect 415804 452874 416404 452876
rect 451804 452874 452404 452876
rect 487804 452874 488404 452876
rect 523804 452874 524404 452876
rect 559804 452874 560404 452876
rect 586260 452874 586860 452876
rect -7636 446276 -7036 446278
rect 12604 446276 13204 446278
rect 48604 446276 49204 446278
rect 84604 446276 85204 446278
rect 120604 446276 121204 446278
rect 156604 446276 157204 446278
rect 192604 446276 193204 446278
rect 228604 446276 229204 446278
rect 264604 446276 265204 446278
rect 300604 446276 301204 446278
rect 336604 446276 337204 446278
rect 372604 446276 373204 446278
rect 408604 446276 409204 446278
rect 444604 446276 445204 446278
rect 480604 446276 481204 446278
rect 516604 446276 517204 446278
rect 552604 446276 553204 446278
rect 590960 446276 591560 446278
rect -8576 446254 592500 446276
rect -8576 446018 -7454 446254
rect -7218 446018 12786 446254
rect 13022 446018 48786 446254
rect 49022 446018 84786 446254
rect 85022 446018 120786 446254
rect 121022 446018 156786 446254
rect 157022 446018 192786 446254
rect 193022 446018 228786 446254
rect 229022 446018 264786 446254
rect 265022 446018 300786 446254
rect 301022 446018 336786 446254
rect 337022 446018 372786 446254
rect 373022 446018 408786 446254
rect 409022 446018 444786 446254
rect 445022 446018 480786 446254
rect 481022 446018 516786 446254
rect 517022 446018 552786 446254
rect 553022 446018 591142 446254
rect 591378 446018 592500 446254
rect -8576 445934 592500 446018
rect -8576 445698 -7454 445934
rect -7218 445698 12786 445934
rect 13022 445698 48786 445934
rect 49022 445698 84786 445934
rect 85022 445698 120786 445934
rect 121022 445698 156786 445934
rect 157022 445698 192786 445934
rect 193022 445698 228786 445934
rect 229022 445698 264786 445934
rect 265022 445698 300786 445934
rect 301022 445698 336786 445934
rect 337022 445698 372786 445934
rect 373022 445698 408786 445934
rect 409022 445698 444786 445934
rect 445022 445698 480786 445934
rect 481022 445698 516786 445934
rect 517022 445698 552786 445934
rect 553022 445698 591142 445934
rect 591378 445698 592500 445934
rect -8576 445676 592500 445698
rect -7636 445674 -7036 445676
rect 12604 445674 13204 445676
rect 48604 445674 49204 445676
rect 84604 445674 85204 445676
rect 120604 445674 121204 445676
rect 156604 445674 157204 445676
rect 192604 445674 193204 445676
rect 228604 445674 229204 445676
rect 264604 445674 265204 445676
rect 300604 445674 301204 445676
rect 336604 445674 337204 445676
rect 372604 445674 373204 445676
rect 408604 445674 409204 445676
rect 444604 445674 445204 445676
rect 480604 445674 481204 445676
rect 516604 445674 517204 445676
rect 552604 445674 553204 445676
rect 590960 445674 591560 445676
rect -5756 442676 -5156 442678
rect 9004 442676 9604 442678
rect 45004 442676 45604 442678
rect 81004 442676 81604 442678
rect 117004 442676 117604 442678
rect 153004 442676 153604 442678
rect 189004 442676 189604 442678
rect 225004 442676 225604 442678
rect 261004 442676 261604 442678
rect 297004 442676 297604 442678
rect 333004 442676 333604 442678
rect 369004 442676 369604 442678
rect 405004 442676 405604 442678
rect 441004 442676 441604 442678
rect 477004 442676 477604 442678
rect 513004 442676 513604 442678
rect 549004 442676 549604 442678
rect 589080 442676 589680 442678
rect -6696 442654 590620 442676
rect -6696 442418 -5574 442654
rect -5338 442418 9186 442654
rect 9422 442418 45186 442654
rect 45422 442418 81186 442654
rect 81422 442418 117186 442654
rect 117422 442418 153186 442654
rect 153422 442418 189186 442654
rect 189422 442418 225186 442654
rect 225422 442418 261186 442654
rect 261422 442418 297186 442654
rect 297422 442418 333186 442654
rect 333422 442418 369186 442654
rect 369422 442418 405186 442654
rect 405422 442418 441186 442654
rect 441422 442418 477186 442654
rect 477422 442418 513186 442654
rect 513422 442418 549186 442654
rect 549422 442418 589262 442654
rect 589498 442418 590620 442654
rect -6696 442334 590620 442418
rect -6696 442098 -5574 442334
rect -5338 442098 9186 442334
rect 9422 442098 45186 442334
rect 45422 442098 81186 442334
rect 81422 442098 117186 442334
rect 117422 442098 153186 442334
rect 153422 442098 189186 442334
rect 189422 442098 225186 442334
rect 225422 442098 261186 442334
rect 261422 442098 297186 442334
rect 297422 442098 333186 442334
rect 333422 442098 369186 442334
rect 369422 442098 405186 442334
rect 405422 442098 441186 442334
rect 441422 442098 477186 442334
rect 477422 442098 513186 442334
rect 513422 442098 549186 442334
rect 549422 442098 589262 442334
rect 589498 442098 590620 442334
rect -6696 442076 590620 442098
rect -5756 442074 -5156 442076
rect 9004 442074 9604 442076
rect 45004 442074 45604 442076
rect 81004 442074 81604 442076
rect 117004 442074 117604 442076
rect 153004 442074 153604 442076
rect 189004 442074 189604 442076
rect 225004 442074 225604 442076
rect 261004 442074 261604 442076
rect 297004 442074 297604 442076
rect 333004 442074 333604 442076
rect 369004 442074 369604 442076
rect 405004 442074 405604 442076
rect 441004 442074 441604 442076
rect 477004 442074 477604 442076
rect 513004 442074 513604 442076
rect 549004 442074 549604 442076
rect 589080 442074 589680 442076
rect -3876 439076 -3276 439078
rect 5404 439076 6004 439078
rect 41404 439076 42004 439078
rect 77404 439076 78004 439078
rect 113404 439076 114004 439078
rect 149404 439076 150004 439078
rect 185404 439076 186004 439078
rect 221404 439076 222004 439078
rect 257404 439076 258004 439078
rect 293404 439076 294004 439078
rect 329404 439076 330004 439078
rect 365404 439076 366004 439078
rect 401404 439076 402004 439078
rect 437404 439076 438004 439078
rect 473404 439076 474004 439078
rect 509404 439076 510004 439078
rect 545404 439076 546004 439078
rect 581404 439076 582004 439078
rect 587200 439076 587800 439078
rect -4816 439054 588740 439076
rect -4816 438818 -3694 439054
rect -3458 438818 5586 439054
rect 5822 438818 41586 439054
rect 41822 438818 77586 439054
rect 77822 438818 113586 439054
rect 113822 438818 149586 439054
rect 149822 438818 185586 439054
rect 185822 438818 221586 439054
rect 221822 438818 257586 439054
rect 257822 438818 293586 439054
rect 293822 438818 329586 439054
rect 329822 438818 365586 439054
rect 365822 438818 401586 439054
rect 401822 438818 437586 439054
rect 437822 438818 473586 439054
rect 473822 438818 509586 439054
rect 509822 438818 545586 439054
rect 545822 438818 581586 439054
rect 581822 438818 587382 439054
rect 587618 438818 588740 439054
rect -4816 438734 588740 438818
rect -4816 438498 -3694 438734
rect -3458 438498 5586 438734
rect 5822 438498 41586 438734
rect 41822 438498 77586 438734
rect 77822 438498 113586 438734
rect 113822 438498 149586 438734
rect 149822 438498 185586 438734
rect 185822 438498 221586 438734
rect 221822 438498 257586 438734
rect 257822 438498 293586 438734
rect 293822 438498 329586 438734
rect 329822 438498 365586 438734
rect 365822 438498 401586 438734
rect 401822 438498 437586 438734
rect 437822 438498 473586 438734
rect 473822 438498 509586 438734
rect 509822 438498 545586 438734
rect 545822 438498 581586 438734
rect 581822 438498 587382 438734
rect 587618 438498 588740 438734
rect -4816 438476 588740 438498
rect -3876 438474 -3276 438476
rect 5404 438474 6004 438476
rect 41404 438474 42004 438476
rect 77404 438474 78004 438476
rect 113404 438474 114004 438476
rect 149404 438474 150004 438476
rect 185404 438474 186004 438476
rect 221404 438474 222004 438476
rect 257404 438474 258004 438476
rect 293404 438474 294004 438476
rect 329404 438474 330004 438476
rect 365404 438474 366004 438476
rect 401404 438474 402004 438476
rect 437404 438474 438004 438476
rect 473404 438474 474004 438476
rect 509404 438474 510004 438476
rect 545404 438474 546004 438476
rect 581404 438474 582004 438476
rect 587200 438474 587800 438476
rect -1996 435476 -1396 435478
rect 1804 435476 2404 435478
rect 37804 435476 38404 435478
rect 73804 435476 74404 435478
rect 109804 435476 110404 435478
rect 145804 435476 146404 435478
rect 181804 435476 182404 435478
rect 217804 435476 218404 435478
rect 253804 435476 254404 435478
rect 289804 435476 290404 435478
rect 325804 435476 326404 435478
rect 361804 435476 362404 435478
rect 397804 435476 398404 435478
rect 433804 435476 434404 435478
rect 469804 435476 470404 435478
rect 505804 435476 506404 435478
rect 541804 435476 542404 435478
rect 577804 435476 578404 435478
rect 585320 435476 585920 435478
rect -2936 435454 586860 435476
rect -2936 435218 -1814 435454
rect -1578 435218 1986 435454
rect 2222 435218 37986 435454
rect 38222 435218 73986 435454
rect 74222 435218 109986 435454
rect 110222 435218 145986 435454
rect 146222 435218 181986 435454
rect 182222 435218 217986 435454
rect 218222 435218 253986 435454
rect 254222 435218 289986 435454
rect 290222 435218 325986 435454
rect 326222 435218 361986 435454
rect 362222 435218 397986 435454
rect 398222 435218 433986 435454
rect 434222 435218 469986 435454
rect 470222 435218 505986 435454
rect 506222 435218 541986 435454
rect 542222 435218 577986 435454
rect 578222 435218 585502 435454
rect 585738 435218 586860 435454
rect -2936 435134 586860 435218
rect -2936 434898 -1814 435134
rect -1578 434898 1986 435134
rect 2222 434898 37986 435134
rect 38222 434898 73986 435134
rect 74222 434898 109986 435134
rect 110222 434898 145986 435134
rect 146222 434898 181986 435134
rect 182222 434898 217986 435134
rect 218222 434898 253986 435134
rect 254222 434898 289986 435134
rect 290222 434898 325986 435134
rect 326222 434898 361986 435134
rect 362222 434898 397986 435134
rect 398222 434898 433986 435134
rect 434222 434898 469986 435134
rect 470222 434898 505986 435134
rect 506222 434898 541986 435134
rect 542222 434898 577986 435134
rect 578222 434898 585502 435134
rect 585738 434898 586860 435134
rect -2936 434876 586860 434898
rect -1996 434874 -1396 434876
rect 1804 434874 2404 434876
rect 37804 434874 38404 434876
rect 73804 434874 74404 434876
rect 109804 434874 110404 434876
rect 145804 434874 146404 434876
rect 181804 434874 182404 434876
rect 217804 434874 218404 434876
rect 253804 434874 254404 434876
rect 289804 434874 290404 434876
rect 325804 434874 326404 434876
rect 361804 434874 362404 434876
rect 397804 434874 398404 434876
rect 433804 434874 434404 434876
rect 469804 434874 470404 434876
rect 505804 434874 506404 434876
rect 541804 434874 542404 434876
rect 577804 434874 578404 434876
rect 585320 434874 585920 434876
rect -8576 428276 -7976 428278
rect 30604 428276 31204 428278
rect 66604 428276 67204 428278
rect 102604 428276 103204 428278
rect 138604 428276 139204 428278
rect 174604 428276 175204 428278
rect 210604 428276 211204 428278
rect 246604 428276 247204 428278
rect 282604 428276 283204 428278
rect 318604 428276 319204 428278
rect 354604 428276 355204 428278
rect 390604 428276 391204 428278
rect 426604 428276 427204 428278
rect 462604 428276 463204 428278
rect 498604 428276 499204 428278
rect 534604 428276 535204 428278
rect 570604 428276 571204 428278
rect 591900 428276 592500 428278
rect -8576 428254 592500 428276
rect -8576 428018 -8394 428254
rect -8158 428018 30786 428254
rect 31022 428018 66786 428254
rect 67022 428018 102786 428254
rect 103022 428018 138786 428254
rect 139022 428018 174786 428254
rect 175022 428018 210786 428254
rect 211022 428018 246786 428254
rect 247022 428018 282786 428254
rect 283022 428018 318786 428254
rect 319022 428018 354786 428254
rect 355022 428018 390786 428254
rect 391022 428018 426786 428254
rect 427022 428018 462786 428254
rect 463022 428018 498786 428254
rect 499022 428018 534786 428254
rect 535022 428018 570786 428254
rect 571022 428018 592082 428254
rect 592318 428018 592500 428254
rect -8576 427934 592500 428018
rect -8576 427698 -8394 427934
rect -8158 427698 30786 427934
rect 31022 427698 66786 427934
rect 67022 427698 102786 427934
rect 103022 427698 138786 427934
rect 139022 427698 174786 427934
rect 175022 427698 210786 427934
rect 211022 427698 246786 427934
rect 247022 427698 282786 427934
rect 283022 427698 318786 427934
rect 319022 427698 354786 427934
rect 355022 427698 390786 427934
rect 391022 427698 426786 427934
rect 427022 427698 462786 427934
rect 463022 427698 498786 427934
rect 499022 427698 534786 427934
rect 535022 427698 570786 427934
rect 571022 427698 592082 427934
rect 592318 427698 592500 427934
rect -8576 427676 592500 427698
rect -8576 427674 -7976 427676
rect 30604 427674 31204 427676
rect 66604 427674 67204 427676
rect 102604 427674 103204 427676
rect 138604 427674 139204 427676
rect 174604 427674 175204 427676
rect 210604 427674 211204 427676
rect 246604 427674 247204 427676
rect 282604 427674 283204 427676
rect 318604 427674 319204 427676
rect 354604 427674 355204 427676
rect 390604 427674 391204 427676
rect 426604 427674 427204 427676
rect 462604 427674 463204 427676
rect 498604 427674 499204 427676
rect 534604 427674 535204 427676
rect 570604 427674 571204 427676
rect 591900 427674 592500 427676
rect -6696 424676 -6096 424678
rect 27004 424676 27604 424678
rect 63004 424676 63604 424678
rect 99004 424676 99604 424678
rect 135004 424676 135604 424678
rect 171004 424676 171604 424678
rect 207004 424676 207604 424678
rect 243004 424676 243604 424678
rect 279004 424676 279604 424678
rect 315004 424676 315604 424678
rect 351004 424676 351604 424678
rect 387004 424676 387604 424678
rect 423004 424676 423604 424678
rect 459004 424676 459604 424678
rect 495004 424676 495604 424678
rect 531004 424676 531604 424678
rect 567004 424676 567604 424678
rect 590020 424676 590620 424678
rect -6696 424654 590620 424676
rect -6696 424418 -6514 424654
rect -6278 424418 27186 424654
rect 27422 424418 63186 424654
rect 63422 424418 99186 424654
rect 99422 424418 135186 424654
rect 135422 424418 171186 424654
rect 171422 424418 207186 424654
rect 207422 424418 243186 424654
rect 243422 424418 279186 424654
rect 279422 424418 315186 424654
rect 315422 424418 351186 424654
rect 351422 424418 387186 424654
rect 387422 424418 423186 424654
rect 423422 424418 459186 424654
rect 459422 424418 495186 424654
rect 495422 424418 531186 424654
rect 531422 424418 567186 424654
rect 567422 424418 590202 424654
rect 590438 424418 590620 424654
rect -6696 424334 590620 424418
rect -6696 424098 -6514 424334
rect -6278 424098 27186 424334
rect 27422 424098 63186 424334
rect 63422 424098 99186 424334
rect 99422 424098 135186 424334
rect 135422 424098 171186 424334
rect 171422 424098 207186 424334
rect 207422 424098 243186 424334
rect 243422 424098 279186 424334
rect 279422 424098 315186 424334
rect 315422 424098 351186 424334
rect 351422 424098 387186 424334
rect 387422 424098 423186 424334
rect 423422 424098 459186 424334
rect 459422 424098 495186 424334
rect 495422 424098 531186 424334
rect 531422 424098 567186 424334
rect 567422 424098 590202 424334
rect 590438 424098 590620 424334
rect -6696 424076 590620 424098
rect -6696 424074 -6096 424076
rect 27004 424074 27604 424076
rect 63004 424074 63604 424076
rect 99004 424074 99604 424076
rect 135004 424074 135604 424076
rect 171004 424074 171604 424076
rect 207004 424074 207604 424076
rect 243004 424074 243604 424076
rect 279004 424074 279604 424076
rect 315004 424074 315604 424076
rect 351004 424074 351604 424076
rect 387004 424074 387604 424076
rect 423004 424074 423604 424076
rect 459004 424074 459604 424076
rect 495004 424074 495604 424076
rect 531004 424074 531604 424076
rect 567004 424074 567604 424076
rect 590020 424074 590620 424076
rect -4816 421076 -4216 421078
rect 23404 421076 24004 421078
rect 59404 421076 60004 421078
rect 95404 421076 96004 421078
rect 131404 421076 132004 421078
rect 167404 421076 168004 421078
rect 203404 421076 204004 421078
rect 239404 421076 240004 421078
rect 275404 421076 276004 421078
rect 311404 421076 312004 421078
rect 347404 421076 348004 421078
rect 383404 421076 384004 421078
rect 419404 421076 420004 421078
rect 455404 421076 456004 421078
rect 491404 421076 492004 421078
rect 527404 421076 528004 421078
rect 563404 421076 564004 421078
rect 588140 421076 588740 421078
rect -4816 421054 588740 421076
rect -4816 420818 -4634 421054
rect -4398 420818 23586 421054
rect 23822 420818 59586 421054
rect 59822 420818 95586 421054
rect 95822 420818 131586 421054
rect 131822 420818 167586 421054
rect 167822 420818 203586 421054
rect 203822 420818 239586 421054
rect 239822 420818 275586 421054
rect 275822 420818 311586 421054
rect 311822 420818 347586 421054
rect 347822 420818 383586 421054
rect 383822 420818 419586 421054
rect 419822 420818 455586 421054
rect 455822 420818 491586 421054
rect 491822 420818 527586 421054
rect 527822 420818 563586 421054
rect 563822 420818 588322 421054
rect 588558 420818 588740 421054
rect -4816 420734 588740 420818
rect -4816 420498 -4634 420734
rect -4398 420498 23586 420734
rect 23822 420498 59586 420734
rect 59822 420498 95586 420734
rect 95822 420498 131586 420734
rect 131822 420498 167586 420734
rect 167822 420498 203586 420734
rect 203822 420498 239586 420734
rect 239822 420498 275586 420734
rect 275822 420498 311586 420734
rect 311822 420498 347586 420734
rect 347822 420498 383586 420734
rect 383822 420498 419586 420734
rect 419822 420498 455586 420734
rect 455822 420498 491586 420734
rect 491822 420498 527586 420734
rect 527822 420498 563586 420734
rect 563822 420498 588322 420734
rect 588558 420498 588740 420734
rect -4816 420476 588740 420498
rect -4816 420474 -4216 420476
rect 23404 420474 24004 420476
rect 59404 420474 60004 420476
rect 95404 420474 96004 420476
rect 131404 420474 132004 420476
rect 167404 420474 168004 420476
rect 203404 420474 204004 420476
rect 239404 420474 240004 420476
rect 275404 420474 276004 420476
rect 311404 420474 312004 420476
rect 347404 420474 348004 420476
rect 383404 420474 384004 420476
rect 419404 420474 420004 420476
rect 455404 420474 456004 420476
rect 491404 420474 492004 420476
rect 527404 420474 528004 420476
rect 563404 420474 564004 420476
rect 588140 420474 588740 420476
rect -2936 417476 -2336 417478
rect 19804 417476 20404 417478
rect 55804 417476 56404 417478
rect 91804 417476 92404 417478
rect 127804 417476 128404 417478
rect 163804 417476 164404 417478
rect 199804 417476 200404 417478
rect 235804 417476 236404 417478
rect 271804 417476 272404 417478
rect 307804 417476 308404 417478
rect 343804 417476 344404 417478
rect 379804 417476 380404 417478
rect 415804 417476 416404 417478
rect 451804 417476 452404 417478
rect 487804 417476 488404 417478
rect 523804 417476 524404 417478
rect 559804 417476 560404 417478
rect 586260 417476 586860 417478
rect -2936 417454 586860 417476
rect -2936 417218 -2754 417454
rect -2518 417218 19986 417454
rect 20222 417218 55986 417454
rect 56222 417218 91986 417454
rect 92222 417218 127986 417454
rect 128222 417218 163986 417454
rect 164222 417218 199986 417454
rect 200222 417218 235986 417454
rect 236222 417218 271986 417454
rect 272222 417218 307986 417454
rect 308222 417218 343986 417454
rect 344222 417218 379986 417454
rect 380222 417218 415986 417454
rect 416222 417218 451986 417454
rect 452222 417218 487986 417454
rect 488222 417218 523986 417454
rect 524222 417218 559986 417454
rect 560222 417218 586442 417454
rect 586678 417218 586860 417454
rect -2936 417134 586860 417218
rect -2936 416898 -2754 417134
rect -2518 416898 19986 417134
rect 20222 416898 55986 417134
rect 56222 416898 91986 417134
rect 92222 416898 127986 417134
rect 128222 416898 163986 417134
rect 164222 416898 199986 417134
rect 200222 416898 235986 417134
rect 236222 416898 271986 417134
rect 272222 416898 307986 417134
rect 308222 416898 343986 417134
rect 344222 416898 379986 417134
rect 380222 416898 415986 417134
rect 416222 416898 451986 417134
rect 452222 416898 487986 417134
rect 488222 416898 523986 417134
rect 524222 416898 559986 417134
rect 560222 416898 586442 417134
rect 586678 416898 586860 417134
rect -2936 416876 586860 416898
rect -2936 416874 -2336 416876
rect 19804 416874 20404 416876
rect 55804 416874 56404 416876
rect 91804 416874 92404 416876
rect 127804 416874 128404 416876
rect 163804 416874 164404 416876
rect 199804 416874 200404 416876
rect 235804 416874 236404 416876
rect 271804 416874 272404 416876
rect 307804 416874 308404 416876
rect 343804 416874 344404 416876
rect 379804 416874 380404 416876
rect 415804 416874 416404 416876
rect 451804 416874 452404 416876
rect 487804 416874 488404 416876
rect 523804 416874 524404 416876
rect 559804 416874 560404 416876
rect 586260 416874 586860 416876
rect -7636 410276 -7036 410278
rect 12604 410276 13204 410278
rect 48604 410276 49204 410278
rect 84604 410276 85204 410278
rect 120604 410276 121204 410278
rect 156604 410276 157204 410278
rect 192604 410276 193204 410278
rect 228604 410276 229204 410278
rect 336604 410276 337204 410278
rect 372604 410276 373204 410278
rect 408604 410276 409204 410278
rect 444604 410276 445204 410278
rect 480604 410276 481204 410278
rect 516604 410276 517204 410278
rect 552604 410276 553204 410278
rect 590960 410276 591560 410278
rect -8576 410254 592500 410276
rect -8576 410018 -7454 410254
rect -7218 410018 12786 410254
rect 13022 410018 48786 410254
rect 49022 410018 84786 410254
rect 85022 410018 120786 410254
rect 121022 410018 156786 410254
rect 157022 410018 192786 410254
rect 193022 410018 228786 410254
rect 229022 410018 336786 410254
rect 337022 410018 372786 410254
rect 373022 410018 408786 410254
rect 409022 410018 444786 410254
rect 445022 410018 480786 410254
rect 481022 410018 516786 410254
rect 517022 410018 552786 410254
rect 553022 410018 591142 410254
rect 591378 410018 592500 410254
rect -8576 409934 592500 410018
rect -8576 409698 -7454 409934
rect -7218 409698 12786 409934
rect 13022 409698 48786 409934
rect 49022 409698 84786 409934
rect 85022 409698 120786 409934
rect 121022 409698 156786 409934
rect 157022 409698 192786 409934
rect 193022 409698 228786 409934
rect 229022 409698 336786 409934
rect 337022 409698 372786 409934
rect 373022 409698 408786 409934
rect 409022 409698 444786 409934
rect 445022 409698 480786 409934
rect 481022 409698 516786 409934
rect 517022 409698 552786 409934
rect 553022 409698 591142 409934
rect 591378 409698 592500 409934
rect -8576 409676 592500 409698
rect -7636 409674 -7036 409676
rect 12604 409674 13204 409676
rect 48604 409674 49204 409676
rect 84604 409674 85204 409676
rect 120604 409674 121204 409676
rect 156604 409674 157204 409676
rect 192604 409674 193204 409676
rect 228604 409674 229204 409676
rect 336604 409674 337204 409676
rect 372604 409674 373204 409676
rect 408604 409674 409204 409676
rect 444604 409674 445204 409676
rect 480604 409674 481204 409676
rect 516604 409674 517204 409676
rect 552604 409674 553204 409676
rect 590960 409674 591560 409676
rect -5756 406676 -5156 406678
rect 9004 406676 9604 406678
rect 45004 406676 45604 406678
rect 81004 406676 81604 406678
rect 117004 406676 117604 406678
rect 153004 406676 153604 406678
rect 189004 406676 189604 406678
rect 225004 406676 225604 406678
rect 333004 406676 333604 406678
rect 369004 406676 369604 406678
rect 405004 406676 405604 406678
rect 441004 406676 441604 406678
rect 477004 406676 477604 406678
rect 513004 406676 513604 406678
rect 549004 406676 549604 406678
rect 589080 406676 589680 406678
rect -6696 406654 590620 406676
rect -6696 406418 -5574 406654
rect -5338 406418 9186 406654
rect 9422 406418 45186 406654
rect 45422 406418 81186 406654
rect 81422 406418 117186 406654
rect 117422 406418 153186 406654
rect 153422 406418 189186 406654
rect 189422 406418 225186 406654
rect 225422 406418 333186 406654
rect 333422 406418 369186 406654
rect 369422 406418 405186 406654
rect 405422 406418 441186 406654
rect 441422 406418 477186 406654
rect 477422 406418 513186 406654
rect 513422 406418 549186 406654
rect 549422 406418 589262 406654
rect 589498 406418 590620 406654
rect -6696 406334 590620 406418
rect -6696 406098 -5574 406334
rect -5338 406098 9186 406334
rect 9422 406098 45186 406334
rect 45422 406098 81186 406334
rect 81422 406098 117186 406334
rect 117422 406098 153186 406334
rect 153422 406098 189186 406334
rect 189422 406098 225186 406334
rect 225422 406098 333186 406334
rect 333422 406098 369186 406334
rect 369422 406098 405186 406334
rect 405422 406098 441186 406334
rect 441422 406098 477186 406334
rect 477422 406098 513186 406334
rect 513422 406098 549186 406334
rect 549422 406098 589262 406334
rect 589498 406098 590620 406334
rect -6696 406076 590620 406098
rect -5756 406074 -5156 406076
rect 9004 406074 9604 406076
rect 45004 406074 45604 406076
rect 81004 406074 81604 406076
rect 117004 406074 117604 406076
rect 153004 406074 153604 406076
rect 189004 406074 189604 406076
rect 225004 406074 225604 406076
rect 333004 406074 333604 406076
rect 369004 406074 369604 406076
rect 405004 406074 405604 406076
rect 441004 406074 441604 406076
rect 477004 406074 477604 406076
rect 513004 406074 513604 406076
rect 549004 406074 549604 406076
rect 589080 406074 589680 406076
rect -3876 403076 -3276 403078
rect 5404 403076 6004 403078
rect 41404 403076 42004 403078
rect 77404 403076 78004 403078
rect 113404 403076 114004 403078
rect 149404 403076 150004 403078
rect 185404 403076 186004 403078
rect 221404 403076 222004 403078
rect 329404 403076 330004 403078
rect 365404 403076 366004 403078
rect 401404 403076 402004 403078
rect 437404 403076 438004 403078
rect 473404 403076 474004 403078
rect 509404 403076 510004 403078
rect 545404 403076 546004 403078
rect 581404 403076 582004 403078
rect 587200 403076 587800 403078
rect -4816 403054 588740 403076
rect -4816 402818 -3694 403054
rect -3458 402818 5586 403054
rect 5822 402818 41586 403054
rect 41822 402818 77586 403054
rect 77822 402818 113586 403054
rect 113822 402818 149586 403054
rect 149822 402818 185586 403054
rect 185822 402818 221586 403054
rect 221822 402818 329586 403054
rect 329822 402818 365586 403054
rect 365822 402818 401586 403054
rect 401822 402818 437586 403054
rect 437822 402818 473586 403054
rect 473822 402818 509586 403054
rect 509822 402818 545586 403054
rect 545822 402818 581586 403054
rect 581822 402818 587382 403054
rect 587618 402818 588740 403054
rect -4816 402734 588740 402818
rect -4816 402498 -3694 402734
rect -3458 402498 5586 402734
rect 5822 402498 41586 402734
rect 41822 402498 77586 402734
rect 77822 402498 113586 402734
rect 113822 402498 149586 402734
rect 149822 402498 185586 402734
rect 185822 402498 221586 402734
rect 221822 402498 329586 402734
rect 329822 402498 365586 402734
rect 365822 402498 401586 402734
rect 401822 402498 437586 402734
rect 437822 402498 473586 402734
rect 473822 402498 509586 402734
rect 509822 402498 545586 402734
rect 545822 402498 581586 402734
rect 581822 402498 587382 402734
rect 587618 402498 588740 402734
rect -4816 402476 588740 402498
rect -3876 402474 -3276 402476
rect 5404 402474 6004 402476
rect 41404 402474 42004 402476
rect 77404 402474 78004 402476
rect 113404 402474 114004 402476
rect 149404 402474 150004 402476
rect 185404 402474 186004 402476
rect 221404 402474 222004 402476
rect 329404 402474 330004 402476
rect 365404 402474 366004 402476
rect 401404 402474 402004 402476
rect 437404 402474 438004 402476
rect 473404 402474 474004 402476
rect 509404 402474 510004 402476
rect 545404 402474 546004 402476
rect 581404 402474 582004 402476
rect 587200 402474 587800 402476
rect -1996 399476 -1396 399478
rect 1804 399476 2404 399478
rect 37804 399476 38404 399478
rect 73804 399476 74404 399478
rect 109804 399476 110404 399478
rect 145804 399476 146404 399478
rect 181804 399476 182404 399478
rect 217804 399476 218404 399478
rect 325804 399476 326404 399478
rect 361804 399476 362404 399478
rect 397804 399476 398404 399478
rect 433804 399476 434404 399478
rect 469804 399476 470404 399478
rect 505804 399476 506404 399478
rect 541804 399476 542404 399478
rect 577804 399476 578404 399478
rect 585320 399476 585920 399478
rect -2936 399454 586860 399476
rect -2936 399218 -1814 399454
rect -1578 399218 1986 399454
rect 2222 399218 37986 399454
rect 38222 399218 73986 399454
rect 74222 399218 109986 399454
rect 110222 399218 145986 399454
rect 146222 399218 181986 399454
rect 182222 399218 217986 399454
rect 218222 399218 325986 399454
rect 326222 399218 361986 399454
rect 362222 399218 397986 399454
rect 398222 399218 433986 399454
rect 434222 399218 469986 399454
rect 470222 399218 505986 399454
rect 506222 399218 541986 399454
rect 542222 399218 577986 399454
rect 578222 399218 585502 399454
rect 585738 399218 586860 399454
rect -2936 399134 586860 399218
rect -2936 398898 -1814 399134
rect -1578 398898 1986 399134
rect 2222 398898 37986 399134
rect 38222 398898 73986 399134
rect 74222 398898 109986 399134
rect 110222 398898 145986 399134
rect 146222 398898 181986 399134
rect 182222 398898 217986 399134
rect 218222 398898 325986 399134
rect 326222 398898 361986 399134
rect 362222 398898 397986 399134
rect 398222 398898 433986 399134
rect 434222 398898 469986 399134
rect 470222 398898 505986 399134
rect 506222 398898 541986 399134
rect 542222 398898 577986 399134
rect 578222 398898 585502 399134
rect 585738 398898 586860 399134
rect -2936 398876 586860 398898
rect -1996 398874 -1396 398876
rect 1804 398874 2404 398876
rect 37804 398874 38404 398876
rect 73804 398874 74404 398876
rect 109804 398874 110404 398876
rect 145804 398874 146404 398876
rect 181804 398874 182404 398876
rect 217804 398874 218404 398876
rect 325804 398874 326404 398876
rect 361804 398874 362404 398876
rect 397804 398874 398404 398876
rect 433804 398874 434404 398876
rect 469804 398874 470404 398876
rect 505804 398874 506404 398876
rect 541804 398874 542404 398876
rect 577804 398874 578404 398876
rect 585320 398874 585920 398876
rect -8576 392276 -7976 392278
rect 30604 392276 31204 392278
rect 66604 392276 67204 392278
rect 102604 392276 103204 392278
rect 138604 392276 139204 392278
rect 174604 392276 175204 392278
rect 210604 392276 211204 392278
rect 318604 392276 319204 392278
rect 354604 392276 355204 392278
rect 390604 392276 391204 392278
rect 426604 392276 427204 392278
rect 462604 392276 463204 392278
rect 498604 392276 499204 392278
rect 534604 392276 535204 392278
rect 570604 392276 571204 392278
rect 591900 392276 592500 392278
rect -8576 392254 592500 392276
rect -8576 392018 -8394 392254
rect -8158 392018 30786 392254
rect 31022 392018 66786 392254
rect 67022 392018 102786 392254
rect 103022 392018 138786 392254
rect 139022 392018 174786 392254
rect 175022 392018 210786 392254
rect 211022 392018 318786 392254
rect 319022 392018 354786 392254
rect 355022 392018 390786 392254
rect 391022 392018 426786 392254
rect 427022 392018 462786 392254
rect 463022 392018 498786 392254
rect 499022 392018 534786 392254
rect 535022 392018 570786 392254
rect 571022 392018 592082 392254
rect 592318 392018 592500 392254
rect -8576 391934 592500 392018
rect -8576 391698 -8394 391934
rect -8158 391698 30786 391934
rect 31022 391698 66786 391934
rect 67022 391698 102786 391934
rect 103022 391698 138786 391934
rect 139022 391698 174786 391934
rect 175022 391698 210786 391934
rect 211022 391698 318786 391934
rect 319022 391698 354786 391934
rect 355022 391698 390786 391934
rect 391022 391698 426786 391934
rect 427022 391698 462786 391934
rect 463022 391698 498786 391934
rect 499022 391698 534786 391934
rect 535022 391698 570786 391934
rect 571022 391698 592082 391934
rect 592318 391698 592500 391934
rect -8576 391676 592500 391698
rect -8576 391674 -7976 391676
rect 30604 391674 31204 391676
rect 66604 391674 67204 391676
rect 102604 391674 103204 391676
rect 138604 391674 139204 391676
rect 174604 391674 175204 391676
rect 210604 391674 211204 391676
rect 318604 391674 319204 391676
rect 354604 391674 355204 391676
rect 390604 391674 391204 391676
rect 426604 391674 427204 391676
rect 462604 391674 463204 391676
rect 498604 391674 499204 391676
rect 534604 391674 535204 391676
rect 570604 391674 571204 391676
rect 591900 391674 592500 391676
rect -6696 388676 -6096 388678
rect 27004 388676 27604 388678
rect 63004 388676 63604 388678
rect 99004 388676 99604 388678
rect 135004 388676 135604 388678
rect 171004 388676 171604 388678
rect 207004 388676 207604 388678
rect 315004 388676 315604 388678
rect 351004 388676 351604 388678
rect 387004 388676 387604 388678
rect 423004 388676 423604 388678
rect 459004 388676 459604 388678
rect 495004 388676 495604 388678
rect 531004 388676 531604 388678
rect 567004 388676 567604 388678
rect 590020 388676 590620 388678
rect -6696 388654 590620 388676
rect -6696 388418 -6514 388654
rect -6278 388418 27186 388654
rect 27422 388418 63186 388654
rect 63422 388418 99186 388654
rect 99422 388418 135186 388654
rect 135422 388418 171186 388654
rect 171422 388418 207186 388654
rect 207422 388418 315186 388654
rect 315422 388418 351186 388654
rect 351422 388418 387186 388654
rect 387422 388418 423186 388654
rect 423422 388418 459186 388654
rect 459422 388418 495186 388654
rect 495422 388418 531186 388654
rect 531422 388418 567186 388654
rect 567422 388418 590202 388654
rect 590438 388418 590620 388654
rect -6696 388334 590620 388418
rect -6696 388098 -6514 388334
rect -6278 388098 27186 388334
rect 27422 388098 63186 388334
rect 63422 388098 99186 388334
rect 99422 388098 135186 388334
rect 135422 388098 171186 388334
rect 171422 388098 207186 388334
rect 207422 388098 315186 388334
rect 315422 388098 351186 388334
rect 351422 388098 387186 388334
rect 387422 388098 423186 388334
rect 423422 388098 459186 388334
rect 459422 388098 495186 388334
rect 495422 388098 531186 388334
rect 531422 388098 567186 388334
rect 567422 388098 590202 388334
rect 590438 388098 590620 388334
rect -6696 388076 590620 388098
rect -6696 388074 -6096 388076
rect 27004 388074 27604 388076
rect 63004 388074 63604 388076
rect 99004 388074 99604 388076
rect 135004 388074 135604 388076
rect 171004 388074 171604 388076
rect 207004 388074 207604 388076
rect 315004 388074 315604 388076
rect 351004 388074 351604 388076
rect 387004 388074 387604 388076
rect 423004 388074 423604 388076
rect 459004 388074 459604 388076
rect 495004 388074 495604 388076
rect 531004 388074 531604 388076
rect 567004 388074 567604 388076
rect 590020 388074 590620 388076
rect -4816 385076 -4216 385078
rect 23404 385076 24004 385078
rect 59404 385076 60004 385078
rect 95404 385076 96004 385078
rect 131404 385076 132004 385078
rect 167404 385076 168004 385078
rect 203404 385076 204004 385078
rect 311404 385076 312004 385078
rect 347404 385076 348004 385078
rect 383404 385076 384004 385078
rect 419404 385076 420004 385078
rect 455404 385076 456004 385078
rect 491404 385076 492004 385078
rect 527404 385076 528004 385078
rect 563404 385076 564004 385078
rect 588140 385076 588740 385078
rect -4816 385054 588740 385076
rect -4816 384818 -4634 385054
rect -4398 384818 23586 385054
rect 23822 384818 59586 385054
rect 59822 384818 95586 385054
rect 95822 384818 131586 385054
rect 131822 384818 167586 385054
rect 167822 384818 203586 385054
rect 203822 384818 311586 385054
rect 311822 384818 347586 385054
rect 347822 384818 383586 385054
rect 383822 384818 419586 385054
rect 419822 384818 455586 385054
rect 455822 384818 491586 385054
rect 491822 384818 527586 385054
rect 527822 384818 563586 385054
rect 563822 384818 588322 385054
rect 588558 384818 588740 385054
rect -4816 384734 588740 384818
rect -4816 384498 -4634 384734
rect -4398 384498 23586 384734
rect 23822 384498 59586 384734
rect 59822 384498 95586 384734
rect 95822 384498 131586 384734
rect 131822 384498 167586 384734
rect 167822 384498 203586 384734
rect 203822 384498 311586 384734
rect 311822 384498 347586 384734
rect 347822 384498 383586 384734
rect 383822 384498 419586 384734
rect 419822 384498 455586 384734
rect 455822 384498 491586 384734
rect 491822 384498 527586 384734
rect 527822 384498 563586 384734
rect 563822 384498 588322 384734
rect 588558 384498 588740 384734
rect -4816 384476 588740 384498
rect -4816 384474 -4216 384476
rect 23404 384474 24004 384476
rect 59404 384474 60004 384476
rect 95404 384474 96004 384476
rect 131404 384474 132004 384476
rect 167404 384474 168004 384476
rect 203404 384474 204004 384476
rect 311404 384474 312004 384476
rect 347404 384474 348004 384476
rect 383404 384474 384004 384476
rect 419404 384474 420004 384476
rect 455404 384474 456004 384476
rect 491404 384474 492004 384476
rect 527404 384474 528004 384476
rect 563404 384474 564004 384476
rect 588140 384474 588740 384476
rect -2936 381476 -2336 381478
rect 19804 381476 20404 381478
rect 55804 381476 56404 381478
rect 91804 381476 92404 381478
rect 127804 381476 128404 381478
rect 163804 381476 164404 381478
rect 199804 381476 200404 381478
rect 307804 381476 308404 381478
rect 343804 381476 344404 381478
rect 379804 381476 380404 381478
rect 415804 381476 416404 381478
rect 451804 381476 452404 381478
rect 487804 381476 488404 381478
rect 523804 381476 524404 381478
rect 559804 381476 560404 381478
rect 586260 381476 586860 381478
rect -2936 381454 586860 381476
rect -2936 381218 -2754 381454
rect -2518 381218 19986 381454
rect 20222 381218 55986 381454
rect 56222 381218 91986 381454
rect 92222 381218 127986 381454
rect 128222 381218 163986 381454
rect 164222 381218 199986 381454
rect 200222 381218 307986 381454
rect 308222 381218 343986 381454
rect 344222 381218 379986 381454
rect 380222 381218 415986 381454
rect 416222 381218 451986 381454
rect 452222 381218 487986 381454
rect 488222 381218 523986 381454
rect 524222 381218 559986 381454
rect 560222 381218 586442 381454
rect 586678 381218 586860 381454
rect -2936 381134 586860 381218
rect -2936 380898 -2754 381134
rect -2518 380898 19986 381134
rect 20222 380898 55986 381134
rect 56222 380898 91986 381134
rect 92222 380898 127986 381134
rect 128222 380898 163986 381134
rect 164222 380898 199986 381134
rect 200222 380898 307986 381134
rect 308222 380898 343986 381134
rect 344222 380898 379986 381134
rect 380222 380898 415986 381134
rect 416222 380898 451986 381134
rect 452222 380898 487986 381134
rect 488222 380898 523986 381134
rect 524222 380898 559986 381134
rect 560222 380898 586442 381134
rect 586678 380898 586860 381134
rect -2936 380876 586860 380898
rect -2936 380874 -2336 380876
rect 19804 380874 20404 380876
rect 55804 380874 56404 380876
rect 91804 380874 92404 380876
rect 127804 380874 128404 380876
rect 163804 380874 164404 380876
rect 199804 380874 200404 380876
rect 307804 380874 308404 380876
rect 343804 380874 344404 380876
rect 379804 380874 380404 380876
rect 415804 380874 416404 380876
rect 451804 380874 452404 380876
rect 487804 380874 488404 380876
rect 523804 380874 524404 380876
rect 559804 380874 560404 380876
rect 586260 380874 586860 380876
rect -7636 374276 -7036 374278
rect 12604 374276 13204 374278
rect 48604 374276 49204 374278
rect 84604 374276 85204 374278
rect 120604 374276 121204 374278
rect 156604 374276 157204 374278
rect 192604 374276 193204 374278
rect 228604 374276 229204 374278
rect 336604 374276 337204 374278
rect 372604 374276 373204 374278
rect 408604 374276 409204 374278
rect 444604 374276 445204 374278
rect 480604 374276 481204 374278
rect 516604 374276 517204 374278
rect 552604 374276 553204 374278
rect 590960 374276 591560 374278
rect -8576 374254 592500 374276
rect -8576 374018 -7454 374254
rect -7218 374018 12786 374254
rect 13022 374018 48786 374254
rect 49022 374018 84786 374254
rect 85022 374018 120786 374254
rect 121022 374018 156786 374254
rect 157022 374018 192786 374254
rect 193022 374018 228786 374254
rect 229022 374018 336786 374254
rect 337022 374018 372786 374254
rect 373022 374018 408786 374254
rect 409022 374018 444786 374254
rect 445022 374018 480786 374254
rect 481022 374018 516786 374254
rect 517022 374018 552786 374254
rect 553022 374018 591142 374254
rect 591378 374018 592500 374254
rect -8576 373934 592500 374018
rect -8576 373698 -7454 373934
rect -7218 373698 12786 373934
rect 13022 373698 48786 373934
rect 49022 373698 84786 373934
rect 85022 373698 120786 373934
rect 121022 373698 156786 373934
rect 157022 373698 192786 373934
rect 193022 373698 228786 373934
rect 229022 373698 336786 373934
rect 337022 373698 372786 373934
rect 373022 373698 408786 373934
rect 409022 373698 444786 373934
rect 445022 373698 480786 373934
rect 481022 373698 516786 373934
rect 517022 373698 552786 373934
rect 553022 373698 591142 373934
rect 591378 373698 592500 373934
rect -8576 373676 592500 373698
rect -7636 373674 -7036 373676
rect 12604 373674 13204 373676
rect 48604 373674 49204 373676
rect 84604 373674 85204 373676
rect 120604 373674 121204 373676
rect 156604 373674 157204 373676
rect 192604 373674 193204 373676
rect 228604 373674 229204 373676
rect 336604 373674 337204 373676
rect 372604 373674 373204 373676
rect 408604 373674 409204 373676
rect 444604 373674 445204 373676
rect 480604 373674 481204 373676
rect 516604 373674 517204 373676
rect 552604 373674 553204 373676
rect 590960 373674 591560 373676
rect -5756 370676 -5156 370678
rect 9004 370676 9604 370678
rect 45004 370676 45604 370678
rect 81004 370676 81604 370678
rect 117004 370676 117604 370678
rect 153004 370676 153604 370678
rect 189004 370676 189604 370678
rect 225004 370676 225604 370678
rect 333004 370676 333604 370678
rect 369004 370676 369604 370678
rect 405004 370676 405604 370678
rect 441004 370676 441604 370678
rect 477004 370676 477604 370678
rect 513004 370676 513604 370678
rect 549004 370676 549604 370678
rect 589080 370676 589680 370678
rect -6696 370654 590620 370676
rect -6696 370418 -5574 370654
rect -5338 370418 9186 370654
rect 9422 370418 45186 370654
rect 45422 370418 81186 370654
rect 81422 370418 117186 370654
rect 117422 370418 153186 370654
rect 153422 370418 189186 370654
rect 189422 370418 225186 370654
rect 225422 370418 333186 370654
rect 333422 370418 369186 370654
rect 369422 370418 405186 370654
rect 405422 370418 441186 370654
rect 441422 370418 477186 370654
rect 477422 370418 513186 370654
rect 513422 370418 549186 370654
rect 549422 370418 589262 370654
rect 589498 370418 590620 370654
rect -6696 370334 590620 370418
rect -6696 370098 -5574 370334
rect -5338 370098 9186 370334
rect 9422 370098 45186 370334
rect 45422 370098 81186 370334
rect 81422 370098 117186 370334
rect 117422 370098 153186 370334
rect 153422 370098 189186 370334
rect 189422 370098 225186 370334
rect 225422 370098 333186 370334
rect 333422 370098 369186 370334
rect 369422 370098 405186 370334
rect 405422 370098 441186 370334
rect 441422 370098 477186 370334
rect 477422 370098 513186 370334
rect 513422 370098 549186 370334
rect 549422 370098 589262 370334
rect 589498 370098 590620 370334
rect -6696 370076 590620 370098
rect -5756 370074 -5156 370076
rect 9004 370074 9604 370076
rect 45004 370074 45604 370076
rect 81004 370074 81604 370076
rect 117004 370074 117604 370076
rect 153004 370074 153604 370076
rect 189004 370074 189604 370076
rect 225004 370074 225604 370076
rect 333004 370074 333604 370076
rect 369004 370074 369604 370076
rect 405004 370074 405604 370076
rect 441004 370074 441604 370076
rect 477004 370074 477604 370076
rect 513004 370074 513604 370076
rect 549004 370074 549604 370076
rect 589080 370074 589680 370076
rect -3876 367076 -3276 367078
rect 5404 367076 6004 367078
rect 41404 367076 42004 367078
rect 77404 367076 78004 367078
rect 113404 367076 114004 367078
rect 149404 367076 150004 367078
rect 185404 367076 186004 367078
rect 221404 367076 222004 367078
rect 329404 367076 330004 367078
rect 365404 367076 366004 367078
rect 401404 367076 402004 367078
rect 437404 367076 438004 367078
rect 473404 367076 474004 367078
rect 509404 367076 510004 367078
rect 545404 367076 546004 367078
rect 581404 367076 582004 367078
rect 587200 367076 587800 367078
rect -4816 367054 588740 367076
rect -4816 366818 -3694 367054
rect -3458 366818 5586 367054
rect 5822 366818 41586 367054
rect 41822 366818 77586 367054
rect 77822 366818 113586 367054
rect 113822 366818 149586 367054
rect 149822 366818 185586 367054
rect 185822 366818 221586 367054
rect 221822 366818 329586 367054
rect 329822 366818 365586 367054
rect 365822 366818 401586 367054
rect 401822 366818 437586 367054
rect 437822 366818 473586 367054
rect 473822 366818 509586 367054
rect 509822 366818 545586 367054
rect 545822 366818 581586 367054
rect 581822 366818 587382 367054
rect 587618 366818 588740 367054
rect -4816 366734 588740 366818
rect -4816 366498 -3694 366734
rect -3458 366498 5586 366734
rect 5822 366498 41586 366734
rect 41822 366498 77586 366734
rect 77822 366498 113586 366734
rect 113822 366498 149586 366734
rect 149822 366498 185586 366734
rect 185822 366498 221586 366734
rect 221822 366498 329586 366734
rect 329822 366498 365586 366734
rect 365822 366498 401586 366734
rect 401822 366498 437586 366734
rect 437822 366498 473586 366734
rect 473822 366498 509586 366734
rect 509822 366498 545586 366734
rect 545822 366498 581586 366734
rect 581822 366498 587382 366734
rect 587618 366498 588740 366734
rect -4816 366476 588740 366498
rect -3876 366474 -3276 366476
rect 5404 366474 6004 366476
rect 41404 366474 42004 366476
rect 77404 366474 78004 366476
rect 113404 366474 114004 366476
rect 149404 366474 150004 366476
rect 185404 366474 186004 366476
rect 221404 366474 222004 366476
rect 329404 366474 330004 366476
rect 365404 366474 366004 366476
rect 401404 366474 402004 366476
rect 437404 366474 438004 366476
rect 473404 366474 474004 366476
rect 509404 366474 510004 366476
rect 545404 366474 546004 366476
rect 581404 366474 582004 366476
rect 587200 366474 587800 366476
rect -1996 363476 -1396 363478
rect 1804 363476 2404 363478
rect 37804 363476 38404 363478
rect 73804 363476 74404 363478
rect 109804 363476 110404 363478
rect 145804 363476 146404 363478
rect 181804 363476 182404 363478
rect 217804 363476 218404 363478
rect 325804 363476 326404 363478
rect 361804 363476 362404 363478
rect 397804 363476 398404 363478
rect 433804 363476 434404 363478
rect 469804 363476 470404 363478
rect 505804 363476 506404 363478
rect 541804 363476 542404 363478
rect 577804 363476 578404 363478
rect 585320 363476 585920 363478
rect -2936 363454 586860 363476
rect -2936 363218 -1814 363454
rect -1578 363218 1986 363454
rect 2222 363218 37986 363454
rect 38222 363218 73986 363454
rect 74222 363218 109986 363454
rect 110222 363218 145986 363454
rect 146222 363218 181986 363454
rect 182222 363218 217986 363454
rect 218222 363218 325986 363454
rect 326222 363218 361986 363454
rect 362222 363218 397986 363454
rect 398222 363218 433986 363454
rect 434222 363218 469986 363454
rect 470222 363218 505986 363454
rect 506222 363218 541986 363454
rect 542222 363218 577986 363454
rect 578222 363218 585502 363454
rect 585738 363218 586860 363454
rect -2936 363134 586860 363218
rect -2936 362898 -1814 363134
rect -1578 362898 1986 363134
rect 2222 362898 37986 363134
rect 38222 362898 73986 363134
rect 74222 362898 109986 363134
rect 110222 362898 145986 363134
rect 146222 362898 181986 363134
rect 182222 362898 217986 363134
rect 218222 362898 325986 363134
rect 326222 362898 361986 363134
rect 362222 362898 397986 363134
rect 398222 362898 433986 363134
rect 434222 362898 469986 363134
rect 470222 362898 505986 363134
rect 506222 362898 541986 363134
rect 542222 362898 577986 363134
rect 578222 362898 585502 363134
rect 585738 362898 586860 363134
rect -2936 362876 586860 362898
rect -1996 362874 -1396 362876
rect 1804 362874 2404 362876
rect 37804 362874 38404 362876
rect 73804 362874 74404 362876
rect 109804 362874 110404 362876
rect 145804 362874 146404 362876
rect 181804 362874 182404 362876
rect 217804 362874 218404 362876
rect 325804 362874 326404 362876
rect 361804 362874 362404 362876
rect 397804 362874 398404 362876
rect 433804 362874 434404 362876
rect 469804 362874 470404 362876
rect 505804 362874 506404 362876
rect 541804 362874 542404 362876
rect 577804 362874 578404 362876
rect 585320 362874 585920 362876
rect -8576 356276 -7976 356278
rect 30604 356276 31204 356278
rect 66604 356276 67204 356278
rect 102604 356276 103204 356278
rect 138604 356276 139204 356278
rect 174604 356276 175204 356278
rect 210604 356276 211204 356278
rect 318604 356276 319204 356278
rect 354604 356276 355204 356278
rect 390604 356276 391204 356278
rect 426604 356276 427204 356278
rect 462604 356276 463204 356278
rect 498604 356276 499204 356278
rect 534604 356276 535204 356278
rect 570604 356276 571204 356278
rect 591900 356276 592500 356278
rect -8576 356254 592500 356276
rect -8576 356018 -8394 356254
rect -8158 356018 30786 356254
rect 31022 356018 66786 356254
rect 67022 356018 102786 356254
rect 103022 356018 138786 356254
rect 139022 356018 174786 356254
rect 175022 356018 210786 356254
rect 211022 356018 318786 356254
rect 319022 356018 354786 356254
rect 355022 356018 390786 356254
rect 391022 356018 426786 356254
rect 427022 356018 462786 356254
rect 463022 356018 498786 356254
rect 499022 356018 534786 356254
rect 535022 356018 570786 356254
rect 571022 356018 592082 356254
rect 592318 356018 592500 356254
rect -8576 355934 592500 356018
rect -8576 355698 -8394 355934
rect -8158 355698 30786 355934
rect 31022 355698 66786 355934
rect 67022 355698 102786 355934
rect 103022 355698 138786 355934
rect 139022 355698 174786 355934
rect 175022 355698 210786 355934
rect 211022 355698 318786 355934
rect 319022 355698 354786 355934
rect 355022 355698 390786 355934
rect 391022 355698 426786 355934
rect 427022 355698 462786 355934
rect 463022 355698 498786 355934
rect 499022 355698 534786 355934
rect 535022 355698 570786 355934
rect 571022 355698 592082 355934
rect 592318 355698 592500 355934
rect -8576 355676 592500 355698
rect -8576 355674 -7976 355676
rect 30604 355674 31204 355676
rect 66604 355674 67204 355676
rect 102604 355674 103204 355676
rect 138604 355674 139204 355676
rect 174604 355674 175204 355676
rect 210604 355674 211204 355676
rect 318604 355674 319204 355676
rect 354604 355674 355204 355676
rect 390604 355674 391204 355676
rect 426604 355674 427204 355676
rect 462604 355674 463204 355676
rect 498604 355674 499204 355676
rect 534604 355674 535204 355676
rect 570604 355674 571204 355676
rect 591900 355674 592500 355676
rect -6696 352676 -6096 352678
rect 27004 352676 27604 352678
rect 63004 352676 63604 352678
rect 99004 352676 99604 352678
rect 135004 352676 135604 352678
rect 171004 352676 171604 352678
rect 207004 352676 207604 352678
rect 315004 352676 315604 352678
rect 351004 352676 351604 352678
rect 387004 352676 387604 352678
rect 423004 352676 423604 352678
rect 459004 352676 459604 352678
rect 495004 352676 495604 352678
rect 531004 352676 531604 352678
rect 567004 352676 567604 352678
rect 590020 352676 590620 352678
rect -6696 352654 590620 352676
rect -6696 352418 -6514 352654
rect -6278 352418 27186 352654
rect 27422 352418 63186 352654
rect 63422 352418 99186 352654
rect 99422 352418 135186 352654
rect 135422 352418 171186 352654
rect 171422 352418 207186 352654
rect 207422 352418 315186 352654
rect 315422 352418 351186 352654
rect 351422 352418 387186 352654
rect 387422 352418 423186 352654
rect 423422 352418 459186 352654
rect 459422 352418 495186 352654
rect 495422 352418 531186 352654
rect 531422 352418 567186 352654
rect 567422 352418 590202 352654
rect 590438 352418 590620 352654
rect -6696 352334 590620 352418
rect -6696 352098 -6514 352334
rect -6278 352098 27186 352334
rect 27422 352098 63186 352334
rect 63422 352098 99186 352334
rect 99422 352098 135186 352334
rect 135422 352098 171186 352334
rect 171422 352098 207186 352334
rect 207422 352098 315186 352334
rect 315422 352098 351186 352334
rect 351422 352098 387186 352334
rect 387422 352098 423186 352334
rect 423422 352098 459186 352334
rect 459422 352098 495186 352334
rect 495422 352098 531186 352334
rect 531422 352098 567186 352334
rect 567422 352098 590202 352334
rect 590438 352098 590620 352334
rect -6696 352076 590620 352098
rect -6696 352074 -6096 352076
rect 27004 352074 27604 352076
rect 63004 352074 63604 352076
rect 99004 352074 99604 352076
rect 135004 352074 135604 352076
rect 171004 352074 171604 352076
rect 207004 352074 207604 352076
rect 315004 352074 315604 352076
rect 351004 352074 351604 352076
rect 387004 352074 387604 352076
rect 423004 352074 423604 352076
rect 459004 352074 459604 352076
rect 495004 352074 495604 352076
rect 531004 352074 531604 352076
rect 567004 352074 567604 352076
rect 590020 352074 590620 352076
rect -4816 349076 -4216 349078
rect 23404 349076 24004 349078
rect 59404 349076 60004 349078
rect 95404 349076 96004 349078
rect 131404 349076 132004 349078
rect 167404 349076 168004 349078
rect 203404 349076 204004 349078
rect 311404 349076 312004 349078
rect 347404 349076 348004 349078
rect 383404 349076 384004 349078
rect 419404 349076 420004 349078
rect 455404 349076 456004 349078
rect 491404 349076 492004 349078
rect 527404 349076 528004 349078
rect 563404 349076 564004 349078
rect 588140 349076 588740 349078
rect -4816 349054 588740 349076
rect -4816 348818 -4634 349054
rect -4398 348818 23586 349054
rect 23822 348818 59586 349054
rect 59822 348818 95586 349054
rect 95822 348818 131586 349054
rect 131822 348818 167586 349054
rect 167822 348818 203586 349054
rect 203822 348818 311586 349054
rect 311822 348818 347586 349054
rect 347822 348818 383586 349054
rect 383822 348818 419586 349054
rect 419822 348818 455586 349054
rect 455822 348818 491586 349054
rect 491822 348818 527586 349054
rect 527822 348818 563586 349054
rect 563822 348818 588322 349054
rect 588558 348818 588740 349054
rect -4816 348734 588740 348818
rect -4816 348498 -4634 348734
rect -4398 348498 23586 348734
rect 23822 348498 59586 348734
rect 59822 348498 95586 348734
rect 95822 348498 131586 348734
rect 131822 348498 167586 348734
rect 167822 348498 203586 348734
rect 203822 348498 311586 348734
rect 311822 348498 347586 348734
rect 347822 348498 383586 348734
rect 383822 348498 419586 348734
rect 419822 348498 455586 348734
rect 455822 348498 491586 348734
rect 491822 348498 527586 348734
rect 527822 348498 563586 348734
rect 563822 348498 588322 348734
rect 588558 348498 588740 348734
rect -4816 348476 588740 348498
rect -4816 348474 -4216 348476
rect 23404 348474 24004 348476
rect 59404 348474 60004 348476
rect 95404 348474 96004 348476
rect 131404 348474 132004 348476
rect 167404 348474 168004 348476
rect 203404 348474 204004 348476
rect 311404 348474 312004 348476
rect 347404 348474 348004 348476
rect 383404 348474 384004 348476
rect 419404 348474 420004 348476
rect 455404 348474 456004 348476
rect 491404 348474 492004 348476
rect 527404 348474 528004 348476
rect 563404 348474 564004 348476
rect 588140 348474 588740 348476
rect -2936 345476 -2336 345478
rect 19804 345476 20404 345478
rect 55804 345476 56404 345478
rect 91804 345476 92404 345478
rect 127804 345476 128404 345478
rect 163804 345476 164404 345478
rect 199804 345476 200404 345478
rect 307804 345476 308404 345478
rect 343804 345476 344404 345478
rect 379804 345476 380404 345478
rect 415804 345476 416404 345478
rect 451804 345476 452404 345478
rect 487804 345476 488404 345478
rect 523804 345476 524404 345478
rect 559804 345476 560404 345478
rect 586260 345476 586860 345478
rect -2936 345454 586860 345476
rect -2936 345218 -2754 345454
rect -2518 345218 19986 345454
rect 20222 345218 55986 345454
rect 56222 345218 91986 345454
rect 92222 345218 127986 345454
rect 128222 345218 163986 345454
rect 164222 345218 199986 345454
rect 200222 345218 307986 345454
rect 308222 345218 343986 345454
rect 344222 345218 379986 345454
rect 380222 345218 415986 345454
rect 416222 345218 451986 345454
rect 452222 345218 487986 345454
rect 488222 345218 523986 345454
rect 524222 345218 559986 345454
rect 560222 345218 586442 345454
rect 586678 345218 586860 345454
rect -2936 345134 586860 345218
rect -2936 344898 -2754 345134
rect -2518 344898 19986 345134
rect 20222 344898 55986 345134
rect 56222 344898 91986 345134
rect 92222 344898 127986 345134
rect 128222 344898 163986 345134
rect 164222 344898 199986 345134
rect 200222 344898 307986 345134
rect 308222 344898 343986 345134
rect 344222 344898 379986 345134
rect 380222 344898 415986 345134
rect 416222 344898 451986 345134
rect 452222 344898 487986 345134
rect 488222 344898 523986 345134
rect 524222 344898 559986 345134
rect 560222 344898 586442 345134
rect 586678 344898 586860 345134
rect -2936 344876 586860 344898
rect -2936 344874 -2336 344876
rect 19804 344874 20404 344876
rect 55804 344874 56404 344876
rect 91804 344874 92404 344876
rect 127804 344874 128404 344876
rect 163804 344874 164404 344876
rect 199804 344874 200404 344876
rect 307804 344874 308404 344876
rect 343804 344874 344404 344876
rect 379804 344874 380404 344876
rect 415804 344874 416404 344876
rect 451804 344874 452404 344876
rect 487804 344874 488404 344876
rect 523804 344874 524404 344876
rect 559804 344874 560404 344876
rect 586260 344874 586860 344876
rect -7636 338276 -7036 338278
rect 12604 338276 13204 338278
rect 48604 338276 49204 338278
rect 84604 338276 85204 338278
rect 120604 338276 121204 338278
rect 156604 338276 157204 338278
rect 192604 338276 193204 338278
rect 228604 338276 229204 338278
rect 336604 338276 337204 338278
rect 372604 338276 373204 338278
rect 408604 338276 409204 338278
rect 444604 338276 445204 338278
rect 480604 338276 481204 338278
rect 516604 338276 517204 338278
rect 552604 338276 553204 338278
rect 590960 338276 591560 338278
rect -8576 338254 592500 338276
rect -8576 338018 -7454 338254
rect -7218 338018 12786 338254
rect 13022 338018 48786 338254
rect 49022 338018 84786 338254
rect 85022 338018 120786 338254
rect 121022 338018 156786 338254
rect 157022 338018 192786 338254
rect 193022 338018 228786 338254
rect 229022 338018 336786 338254
rect 337022 338018 372786 338254
rect 373022 338018 408786 338254
rect 409022 338018 444786 338254
rect 445022 338018 480786 338254
rect 481022 338018 516786 338254
rect 517022 338018 552786 338254
rect 553022 338018 591142 338254
rect 591378 338018 592500 338254
rect -8576 337934 592500 338018
rect -8576 337698 -7454 337934
rect -7218 337698 12786 337934
rect 13022 337698 48786 337934
rect 49022 337698 84786 337934
rect 85022 337698 120786 337934
rect 121022 337698 156786 337934
rect 157022 337698 192786 337934
rect 193022 337698 228786 337934
rect 229022 337698 336786 337934
rect 337022 337698 372786 337934
rect 373022 337698 408786 337934
rect 409022 337698 444786 337934
rect 445022 337698 480786 337934
rect 481022 337698 516786 337934
rect 517022 337698 552786 337934
rect 553022 337698 591142 337934
rect 591378 337698 592500 337934
rect -8576 337676 592500 337698
rect -7636 337674 -7036 337676
rect 12604 337674 13204 337676
rect 48604 337674 49204 337676
rect 84604 337674 85204 337676
rect 120604 337674 121204 337676
rect 156604 337674 157204 337676
rect 192604 337674 193204 337676
rect 228604 337674 229204 337676
rect 336604 337674 337204 337676
rect 372604 337674 373204 337676
rect 408604 337674 409204 337676
rect 444604 337674 445204 337676
rect 480604 337674 481204 337676
rect 516604 337674 517204 337676
rect 552604 337674 553204 337676
rect 590960 337674 591560 337676
rect -5756 334676 -5156 334678
rect 9004 334676 9604 334678
rect 45004 334676 45604 334678
rect 81004 334676 81604 334678
rect 117004 334676 117604 334678
rect 153004 334676 153604 334678
rect 189004 334676 189604 334678
rect 225004 334676 225604 334678
rect 261004 334676 261604 334678
rect 297004 334676 297604 334678
rect 333004 334676 333604 334678
rect 369004 334676 369604 334678
rect 405004 334676 405604 334678
rect 441004 334676 441604 334678
rect 477004 334676 477604 334678
rect 513004 334676 513604 334678
rect 549004 334676 549604 334678
rect 589080 334676 589680 334678
rect -6696 334654 590620 334676
rect -6696 334418 -5574 334654
rect -5338 334418 9186 334654
rect 9422 334418 45186 334654
rect 45422 334418 81186 334654
rect 81422 334418 117186 334654
rect 117422 334418 153186 334654
rect 153422 334418 189186 334654
rect 189422 334418 225186 334654
rect 225422 334418 261186 334654
rect 261422 334418 297186 334654
rect 297422 334418 333186 334654
rect 333422 334418 369186 334654
rect 369422 334418 405186 334654
rect 405422 334418 441186 334654
rect 441422 334418 477186 334654
rect 477422 334418 513186 334654
rect 513422 334418 549186 334654
rect 549422 334418 589262 334654
rect 589498 334418 590620 334654
rect -6696 334334 590620 334418
rect -6696 334098 -5574 334334
rect -5338 334098 9186 334334
rect 9422 334098 45186 334334
rect 45422 334098 81186 334334
rect 81422 334098 117186 334334
rect 117422 334098 153186 334334
rect 153422 334098 189186 334334
rect 189422 334098 225186 334334
rect 225422 334098 261186 334334
rect 261422 334098 297186 334334
rect 297422 334098 333186 334334
rect 333422 334098 369186 334334
rect 369422 334098 405186 334334
rect 405422 334098 441186 334334
rect 441422 334098 477186 334334
rect 477422 334098 513186 334334
rect 513422 334098 549186 334334
rect 549422 334098 589262 334334
rect 589498 334098 590620 334334
rect -6696 334076 590620 334098
rect -5756 334074 -5156 334076
rect 9004 334074 9604 334076
rect 45004 334074 45604 334076
rect 81004 334074 81604 334076
rect 117004 334074 117604 334076
rect 153004 334074 153604 334076
rect 189004 334074 189604 334076
rect 225004 334074 225604 334076
rect 261004 334074 261604 334076
rect 297004 334074 297604 334076
rect 333004 334074 333604 334076
rect 369004 334074 369604 334076
rect 405004 334074 405604 334076
rect 441004 334074 441604 334076
rect 477004 334074 477604 334076
rect 513004 334074 513604 334076
rect 549004 334074 549604 334076
rect 589080 334074 589680 334076
rect -3876 331076 -3276 331078
rect 5404 331076 6004 331078
rect 41404 331076 42004 331078
rect 77404 331076 78004 331078
rect 113404 331076 114004 331078
rect 149404 331076 150004 331078
rect 185404 331076 186004 331078
rect 221404 331076 222004 331078
rect 257404 331076 258004 331078
rect 293404 331076 294004 331078
rect 329404 331076 330004 331078
rect 365404 331076 366004 331078
rect 401404 331076 402004 331078
rect 437404 331076 438004 331078
rect 473404 331076 474004 331078
rect 509404 331076 510004 331078
rect 545404 331076 546004 331078
rect 581404 331076 582004 331078
rect 587200 331076 587800 331078
rect -4816 331054 588740 331076
rect -4816 330818 -3694 331054
rect -3458 330818 5586 331054
rect 5822 330818 41586 331054
rect 41822 330818 77586 331054
rect 77822 330818 113586 331054
rect 113822 330818 149586 331054
rect 149822 330818 185586 331054
rect 185822 330818 221586 331054
rect 221822 330818 257586 331054
rect 257822 330818 293586 331054
rect 293822 330818 329586 331054
rect 329822 330818 365586 331054
rect 365822 330818 401586 331054
rect 401822 330818 437586 331054
rect 437822 330818 473586 331054
rect 473822 330818 509586 331054
rect 509822 330818 545586 331054
rect 545822 330818 581586 331054
rect 581822 330818 587382 331054
rect 587618 330818 588740 331054
rect -4816 330734 588740 330818
rect -4816 330498 -3694 330734
rect -3458 330498 5586 330734
rect 5822 330498 41586 330734
rect 41822 330498 77586 330734
rect 77822 330498 113586 330734
rect 113822 330498 149586 330734
rect 149822 330498 185586 330734
rect 185822 330498 221586 330734
rect 221822 330498 257586 330734
rect 257822 330498 293586 330734
rect 293822 330498 329586 330734
rect 329822 330498 365586 330734
rect 365822 330498 401586 330734
rect 401822 330498 437586 330734
rect 437822 330498 473586 330734
rect 473822 330498 509586 330734
rect 509822 330498 545586 330734
rect 545822 330498 581586 330734
rect 581822 330498 587382 330734
rect 587618 330498 588740 330734
rect -4816 330476 588740 330498
rect -3876 330474 -3276 330476
rect 5404 330474 6004 330476
rect 41404 330474 42004 330476
rect 77404 330474 78004 330476
rect 113404 330474 114004 330476
rect 149404 330474 150004 330476
rect 185404 330474 186004 330476
rect 221404 330474 222004 330476
rect 257404 330474 258004 330476
rect 293404 330474 294004 330476
rect 329404 330474 330004 330476
rect 365404 330474 366004 330476
rect 401404 330474 402004 330476
rect 437404 330474 438004 330476
rect 473404 330474 474004 330476
rect 509404 330474 510004 330476
rect 545404 330474 546004 330476
rect 581404 330474 582004 330476
rect 587200 330474 587800 330476
rect -1996 327476 -1396 327478
rect 1804 327476 2404 327478
rect 37804 327476 38404 327478
rect 73804 327476 74404 327478
rect 109804 327476 110404 327478
rect 145804 327476 146404 327478
rect 181804 327476 182404 327478
rect 217804 327476 218404 327478
rect 253804 327476 254404 327478
rect 289804 327476 290404 327478
rect 325804 327476 326404 327478
rect 361804 327476 362404 327478
rect 397804 327476 398404 327478
rect 433804 327476 434404 327478
rect 469804 327476 470404 327478
rect 505804 327476 506404 327478
rect 541804 327476 542404 327478
rect 577804 327476 578404 327478
rect 585320 327476 585920 327478
rect -2936 327454 586860 327476
rect -2936 327218 -1814 327454
rect -1578 327218 1986 327454
rect 2222 327218 37986 327454
rect 38222 327218 73986 327454
rect 74222 327218 109986 327454
rect 110222 327218 145986 327454
rect 146222 327218 181986 327454
rect 182222 327218 217986 327454
rect 218222 327218 253986 327454
rect 254222 327218 289986 327454
rect 290222 327218 325986 327454
rect 326222 327218 361986 327454
rect 362222 327218 397986 327454
rect 398222 327218 433986 327454
rect 434222 327218 469986 327454
rect 470222 327218 505986 327454
rect 506222 327218 541986 327454
rect 542222 327218 577986 327454
rect 578222 327218 585502 327454
rect 585738 327218 586860 327454
rect -2936 327134 586860 327218
rect -2936 326898 -1814 327134
rect -1578 326898 1986 327134
rect 2222 326898 37986 327134
rect 38222 326898 73986 327134
rect 74222 326898 109986 327134
rect 110222 326898 145986 327134
rect 146222 326898 181986 327134
rect 182222 326898 217986 327134
rect 218222 326898 253986 327134
rect 254222 326898 289986 327134
rect 290222 326898 325986 327134
rect 326222 326898 361986 327134
rect 362222 326898 397986 327134
rect 398222 326898 433986 327134
rect 434222 326898 469986 327134
rect 470222 326898 505986 327134
rect 506222 326898 541986 327134
rect 542222 326898 577986 327134
rect 578222 326898 585502 327134
rect 585738 326898 586860 327134
rect -2936 326876 586860 326898
rect -1996 326874 -1396 326876
rect 1804 326874 2404 326876
rect 37804 326874 38404 326876
rect 73804 326874 74404 326876
rect 109804 326874 110404 326876
rect 145804 326874 146404 326876
rect 181804 326874 182404 326876
rect 217804 326874 218404 326876
rect 253804 326874 254404 326876
rect 289804 326874 290404 326876
rect 325804 326874 326404 326876
rect 361804 326874 362404 326876
rect 397804 326874 398404 326876
rect 433804 326874 434404 326876
rect 469804 326874 470404 326876
rect 505804 326874 506404 326876
rect 541804 326874 542404 326876
rect 577804 326874 578404 326876
rect 585320 326874 585920 326876
rect -8576 320276 -7976 320278
rect 30604 320276 31204 320278
rect 66604 320276 67204 320278
rect 102604 320276 103204 320278
rect 138604 320276 139204 320278
rect 174604 320276 175204 320278
rect 210604 320276 211204 320278
rect 246604 320276 247204 320278
rect 282604 320276 283204 320278
rect 318604 320276 319204 320278
rect 354604 320276 355204 320278
rect 390604 320276 391204 320278
rect 426604 320276 427204 320278
rect 462604 320276 463204 320278
rect 498604 320276 499204 320278
rect 534604 320276 535204 320278
rect 570604 320276 571204 320278
rect 591900 320276 592500 320278
rect -8576 320254 592500 320276
rect -8576 320018 -8394 320254
rect -8158 320018 30786 320254
rect 31022 320018 66786 320254
rect 67022 320018 102786 320254
rect 103022 320018 138786 320254
rect 139022 320018 174786 320254
rect 175022 320018 210786 320254
rect 211022 320018 246786 320254
rect 247022 320018 282786 320254
rect 283022 320018 318786 320254
rect 319022 320018 354786 320254
rect 355022 320018 390786 320254
rect 391022 320018 426786 320254
rect 427022 320018 462786 320254
rect 463022 320018 498786 320254
rect 499022 320018 534786 320254
rect 535022 320018 570786 320254
rect 571022 320018 592082 320254
rect 592318 320018 592500 320254
rect -8576 319934 592500 320018
rect -8576 319698 -8394 319934
rect -8158 319698 30786 319934
rect 31022 319698 66786 319934
rect 67022 319698 102786 319934
rect 103022 319698 138786 319934
rect 139022 319698 174786 319934
rect 175022 319698 210786 319934
rect 211022 319698 246786 319934
rect 247022 319698 282786 319934
rect 283022 319698 318786 319934
rect 319022 319698 354786 319934
rect 355022 319698 390786 319934
rect 391022 319698 426786 319934
rect 427022 319698 462786 319934
rect 463022 319698 498786 319934
rect 499022 319698 534786 319934
rect 535022 319698 570786 319934
rect 571022 319698 592082 319934
rect 592318 319698 592500 319934
rect -8576 319676 592500 319698
rect -8576 319674 -7976 319676
rect 30604 319674 31204 319676
rect 66604 319674 67204 319676
rect 102604 319674 103204 319676
rect 138604 319674 139204 319676
rect 174604 319674 175204 319676
rect 210604 319674 211204 319676
rect 246604 319674 247204 319676
rect 282604 319674 283204 319676
rect 318604 319674 319204 319676
rect 354604 319674 355204 319676
rect 390604 319674 391204 319676
rect 426604 319674 427204 319676
rect 462604 319674 463204 319676
rect 498604 319674 499204 319676
rect 534604 319674 535204 319676
rect 570604 319674 571204 319676
rect 591900 319674 592500 319676
rect -6696 316676 -6096 316678
rect 27004 316676 27604 316678
rect 63004 316676 63604 316678
rect 99004 316676 99604 316678
rect 135004 316676 135604 316678
rect 171004 316676 171604 316678
rect 207004 316676 207604 316678
rect 243004 316676 243604 316678
rect 279004 316676 279604 316678
rect 315004 316676 315604 316678
rect 351004 316676 351604 316678
rect 387004 316676 387604 316678
rect 423004 316676 423604 316678
rect 459004 316676 459604 316678
rect 495004 316676 495604 316678
rect 531004 316676 531604 316678
rect 567004 316676 567604 316678
rect 590020 316676 590620 316678
rect -6696 316654 590620 316676
rect -6696 316418 -6514 316654
rect -6278 316418 27186 316654
rect 27422 316418 63186 316654
rect 63422 316418 99186 316654
rect 99422 316418 135186 316654
rect 135422 316418 171186 316654
rect 171422 316418 207186 316654
rect 207422 316418 243186 316654
rect 243422 316418 279186 316654
rect 279422 316418 315186 316654
rect 315422 316418 351186 316654
rect 351422 316418 387186 316654
rect 387422 316418 423186 316654
rect 423422 316418 459186 316654
rect 459422 316418 495186 316654
rect 495422 316418 531186 316654
rect 531422 316418 567186 316654
rect 567422 316418 590202 316654
rect 590438 316418 590620 316654
rect -6696 316334 590620 316418
rect -6696 316098 -6514 316334
rect -6278 316098 27186 316334
rect 27422 316098 63186 316334
rect 63422 316098 99186 316334
rect 99422 316098 135186 316334
rect 135422 316098 171186 316334
rect 171422 316098 207186 316334
rect 207422 316098 243186 316334
rect 243422 316098 279186 316334
rect 279422 316098 315186 316334
rect 315422 316098 351186 316334
rect 351422 316098 387186 316334
rect 387422 316098 423186 316334
rect 423422 316098 459186 316334
rect 459422 316098 495186 316334
rect 495422 316098 531186 316334
rect 531422 316098 567186 316334
rect 567422 316098 590202 316334
rect 590438 316098 590620 316334
rect -6696 316076 590620 316098
rect -6696 316074 -6096 316076
rect 27004 316074 27604 316076
rect 63004 316074 63604 316076
rect 99004 316074 99604 316076
rect 135004 316074 135604 316076
rect 171004 316074 171604 316076
rect 207004 316074 207604 316076
rect 243004 316074 243604 316076
rect 279004 316074 279604 316076
rect 315004 316074 315604 316076
rect 351004 316074 351604 316076
rect 387004 316074 387604 316076
rect 423004 316074 423604 316076
rect 459004 316074 459604 316076
rect 495004 316074 495604 316076
rect 531004 316074 531604 316076
rect 567004 316074 567604 316076
rect 590020 316074 590620 316076
rect -4816 313076 -4216 313078
rect 23404 313076 24004 313078
rect 59404 313076 60004 313078
rect 95404 313076 96004 313078
rect 131404 313076 132004 313078
rect 167404 313076 168004 313078
rect 203404 313076 204004 313078
rect 239404 313076 240004 313078
rect 275404 313076 276004 313078
rect 311404 313076 312004 313078
rect 347404 313076 348004 313078
rect 383404 313076 384004 313078
rect 419404 313076 420004 313078
rect 455404 313076 456004 313078
rect 491404 313076 492004 313078
rect 527404 313076 528004 313078
rect 563404 313076 564004 313078
rect 588140 313076 588740 313078
rect -4816 313054 588740 313076
rect -4816 312818 -4634 313054
rect -4398 312818 23586 313054
rect 23822 312818 59586 313054
rect 59822 312818 95586 313054
rect 95822 312818 131586 313054
rect 131822 312818 167586 313054
rect 167822 312818 203586 313054
rect 203822 312818 239586 313054
rect 239822 312818 275586 313054
rect 275822 312818 311586 313054
rect 311822 312818 347586 313054
rect 347822 312818 383586 313054
rect 383822 312818 419586 313054
rect 419822 312818 455586 313054
rect 455822 312818 491586 313054
rect 491822 312818 527586 313054
rect 527822 312818 563586 313054
rect 563822 312818 588322 313054
rect 588558 312818 588740 313054
rect -4816 312734 588740 312818
rect -4816 312498 -4634 312734
rect -4398 312498 23586 312734
rect 23822 312498 59586 312734
rect 59822 312498 95586 312734
rect 95822 312498 131586 312734
rect 131822 312498 167586 312734
rect 167822 312498 203586 312734
rect 203822 312498 239586 312734
rect 239822 312498 275586 312734
rect 275822 312498 311586 312734
rect 311822 312498 347586 312734
rect 347822 312498 383586 312734
rect 383822 312498 419586 312734
rect 419822 312498 455586 312734
rect 455822 312498 491586 312734
rect 491822 312498 527586 312734
rect 527822 312498 563586 312734
rect 563822 312498 588322 312734
rect 588558 312498 588740 312734
rect -4816 312476 588740 312498
rect -4816 312474 -4216 312476
rect 23404 312474 24004 312476
rect 59404 312474 60004 312476
rect 95404 312474 96004 312476
rect 131404 312474 132004 312476
rect 167404 312474 168004 312476
rect 203404 312474 204004 312476
rect 239404 312474 240004 312476
rect 275404 312474 276004 312476
rect 311404 312474 312004 312476
rect 347404 312474 348004 312476
rect 383404 312474 384004 312476
rect 419404 312474 420004 312476
rect 455404 312474 456004 312476
rect 491404 312474 492004 312476
rect 527404 312474 528004 312476
rect 563404 312474 564004 312476
rect 588140 312474 588740 312476
rect -2936 309476 -2336 309478
rect 19804 309476 20404 309478
rect 55804 309476 56404 309478
rect 91804 309476 92404 309478
rect 127804 309476 128404 309478
rect 163804 309476 164404 309478
rect 199804 309476 200404 309478
rect 235804 309476 236404 309478
rect 271804 309476 272404 309478
rect 307804 309476 308404 309478
rect 343804 309476 344404 309478
rect 379804 309476 380404 309478
rect 415804 309476 416404 309478
rect 451804 309476 452404 309478
rect 487804 309476 488404 309478
rect 523804 309476 524404 309478
rect 559804 309476 560404 309478
rect 586260 309476 586860 309478
rect -2936 309454 586860 309476
rect -2936 309218 -2754 309454
rect -2518 309218 19986 309454
rect 20222 309218 55986 309454
rect 56222 309218 91986 309454
rect 92222 309218 127986 309454
rect 128222 309218 163986 309454
rect 164222 309218 199986 309454
rect 200222 309218 235986 309454
rect 236222 309218 271986 309454
rect 272222 309218 307986 309454
rect 308222 309218 343986 309454
rect 344222 309218 379986 309454
rect 380222 309218 415986 309454
rect 416222 309218 451986 309454
rect 452222 309218 487986 309454
rect 488222 309218 523986 309454
rect 524222 309218 559986 309454
rect 560222 309218 586442 309454
rect 586678 309218 586860 309454
rect -2936 309134 586860 309218
rect -2936 308898 -2754 309134
rect -2518 308898 19986 309134
rect 20222 308898 55986 309134
rect 56222 308898 91986 309134
rect 92222 308898 127986 309134
rect 128222 308898 163986 309134
rect 164222 308898 199986 309134
rect 200222 308898 235986 309134
rect 236222 308898 271986 309134
rect 272222 308898 307986 309134
rect 308222 308898 343986 309134
rect 344222 308898 379986 309134
rect 380222 308898 415986 309134
rect 416222 308898 451986 309134
rect 452222 308898 487986 309134
rect 488222 308898 523986 309134
rect 524222 308898 559986 309134
rect 560222 308898 586442 309134
rect 586678 308898 586860 309134
rect -2936 308876 586860 308898
rect -2936 308874 -2336 308876
rect 19804 308874 20404 308876
rect 55804 308874 56404 308876
rect 91804 308874 92404 308876
rect 127804 308874 128404 308876
rect 163804 308874 164404 308876
rect 199804 308874 200404 308876
rect 235804 308874 236404 308876
rect 271804 308874 272404 308876
rect 307804 308874 308404 308876
rect 343804 308874 344404 308876
rect 379804 308874 380404 308876
rect 415804 308874 416404 308876
rect 451804 308874 452404 308876
rect 487804 308874 488404 308876
rect 523804 308874 524404 308876
rect 559804 308874 560404 308876
rect 586260 308874 586860 308876
rect -7636 302276 -7036 302278
rect 12604 302276 13204 302278
rect 48604 302276 49204 302278
rect 84604 302276 85204 302278
rect 120604 302276 121204 302278
rect 156604 302276 157204 302278
rect 192604 302276 193204 302278
rect 228604 302276 229204 302278
rect 264604 302276 265204 302278
rect 300604 302276 301204 302278
rect 336604 302276 337204 302278
rect 372604 302276 373204 302278
rect 408604 302276 409204 302278
rect 444604 302276 445204 302278
rect 480604 302276 481204 302278
rect 516604 302276 517204 302278
rect 552604 302276 553204 302278
rect 590960 302276 591560 302278
rect -8576 302254 592500 302276
rect -8576 302018 -7454 302254
rect -7218 302018 12786 302254
rect 13022 302018 48786 302254
rect 49022 302018 84786 302254
rect 85022 302018 120786 302254
rect 121022 302018 156786 302254
rect 157022 302018 192786 302254
rect 193022 302018 228786 302254
rect 229022 302018 264786 302254
rect 265022 302018 300786 302254
rect 301022 302018 336786 302254
rect 337022 302018 372786 302254
rect 373022 302018 408786 302254
rect 409022 302018 444786 302254
rect 445022 302018 480786 302254
rect 481022 302018 516786 302254
rect 517022 302018 552786 302254
rect 553022 302018 591142 302254
rect 591378 302018 592500 302254
rect -8576 301934 592500 302018
rect -8576 301698 -7454 301934
rect -7218 301698 12786 301934
rect 13022 301698 48786 301934
rect 49022 301698 84786 301934
rect 85022 301698 120786 301934
rect 121022 301698 156786 301934
rect 157022 301698 192786 301934
rect 193022 301698 228786 301934
rect 229022 301698 264786 301934
rect 265022 301698 300786 301934
rect 301022 301698 336786 301934
rect 337022 301698 372786 301934
rect 373022 301698 408786 301934
rect 409022 301698 444786 301934
rect 445022 301698 480786 301934
rect 481022 301698 516786 301934
rect 517022 301698 552786 301934
rect 553022 301698 591142 301934
rect 591378 301698 592500 301934
rect -8576 301676 592500 301698
rect -7636 301674 -7036 301676
rect 12604 301674 13204 301676
rect 48604 301674 49204 301676
rect 84604 301674 85204 301676
rect 120604 301674 121204 301676
rect 156604 301674 157204 301676
rect 192604 301674 193204 301676
rect 228604 301674 229204 301676
rect 264604 301674 265204 301676
rect 300604 301674 301204 301676
rect 336604 301674 337204 301676
rect 372604 301674 373204 301676
rect 408604 301674 409204 301676
rect 444604 301674 445204 301676
rect 480604 301674 481204 301676
rect 516604 301674 517204 301676
rect 552604 301674 553204 301676
rect 590960 301674 591560 301676
rect -5756 298676 -5156 298678
rect 9004 298676 9604 298678
rect 45004 298676 45604 298678
rect 81004 298676 81604 298678
rect 117004 298676 117604 298678
rect 153004 298676 153604 298678
rect 189004 298676 189604 298678
rect 225004 298676 225604 298678
rect 261004 298676 261604 298678
rect 297004 298676 297604 298678
rect 333004 298676 333604 298678
rect 369004 298676 369604 298678
rect 405004 298676 405604 298678
rect 441004 298676 441604 298678
rect 477004 298676 477604 298678
rect 513004 298676 513604 298678
rect 549004 298676 549604 298678
rect 589080 298676 589680 298678
rect -6696 298654 590620 298676
rect -6696 298418 -5574 298654
rect -5338 298418 9186 298654
rect 9422 298418 45186 298654
rect 45422 298418 81186 298654
rect 81422 298418 117186 298654
rect 117422 298418 153186 298654
rect 153422 298418 189186 298654
rect 189422 298418 225186 298654
rect 225422 298418 261186 298654
rect 261422 298418 297186 298654
rect 297422 298418 333186 298654
rect 333422 298418 369186 298654
rect 369422 298418 405186 298654
rect 405422 298418 441186 298654
rect 441422 298418 477186 298654
rect 477422 298418 513186 298654
rect 513422 298418 549186 298654
rect 549422 298418 589262 298654
rect 589498 298418 590620 298654
rect -6696 298334 590620 298418
rect -6696 298098 -5574 298334
rect -5338 298098 9186 298334
rect 9422 298098 45186 298334
rect 45422 298098 81186 298334
rect 81422 298098 117186 298334
rect 117422 298098 153186 298334
rect 153422 298098 189186 298334
rect 189422 298098 225186 298334
rect 225422 298098 261186 298334
rect 261422 298098 297186 298334
rect 297422 298098 333186 298334
rect 333422 298098 369186 298334
rect 369422 298098 405186 298334
rect 405422 298098 441186 298334
rect 441422 298098 477186 298334
rect 477422 298098 513186 298334
rect 513422 298098 549186 298334
rect 549422 298098 589262 298334
rect 589498 298098 590620 298334
rect -6696 298076 590620 298098
rect -5756 298074 -5156 298076
rect 9004 298074 9604 298076
rect 45004 298074 45604 298076
rect 81004 298074 81604 298076
rect 117004 298074 117604 298076
rect 153004 298074 153604 298076
rect 189004 298074 189604 298076
rect 225004 298074 225604 298076
rect 261004 298074 261604 298076
rect 297004 298074 297604 298076
rect 333004 298074 333604 298076
rect 369004 298074 369604 298076
rect 405004 298074 405604 298076
rect 441004 298074 441604 298076
rect 477004 298074 477604 298076
rect 513004 298074 513604 298076
rect 549004 298074 549604 298076
rect 589080 298074 589680 298076
rect -3876 295076 -3276 295078
rect 5404 295076 6004 295078
rect 41404 295076 42004 295078
rect 77404 295076 78004 295078
rect 113404 295076 114004 295078
rect 149404 295076 150004 295078
rect 185404 295076 186004 295078
rect 221404 295076 222004 295078
rect 257404 295076 258004 295078
rect 293404 295076 294004 295078
rect 329404 295076 330004 295078
rect 365404 295076 366004 295078
rect 401404 295076 402004 295078
rect 437404 295076 438004 295078
rect 473404 295076 474004 295078
rect 509404 295076 510004 295078
rect 545404 295076 546004 295078
rect 581404 295076 582004 295078
rect 587200 295076 587800 295078
rect -4816 295054 588740 295076
rect -4816 294818 -3694 295054
rect -3458 294818 5586 295054
rect 5822 294818 41586 295054
rect 41822 294818 77586 295054
rect 77822 294818 113586 295054
rect 113822 294818 149586 295054
rect 149822 294818 185586 295054
rect 185822 294818 221586 295054
rect 221822 294818 257586 295054
rect 257822 294818 293586 295054
rect 293822 294818 329586 295054
rect 329822 294818 365586 295054
rect 365822 294818 401586 295054
rect 401822 294818 437586 295054
rect 437822 294818 473586 295054
rect 473822 294818 509586 295054
rect 509822 294818 545586 295054
rect 545822 294818 581586 295054
rect 581822 294818 587382 295054
rect 587618 294818 588740 295054
rect -4816 294734 588740 294818
rect -4816 294498 -3694 294734
rect -3458 294498 5586 294734
rect 5822 294498 41586 294734
rect 41822 294498 77586 294734
rect 77822 294498 113586 294734
rect 113822 294498 149586 294734
rect 149822 294498 185586 294734
rect 185822 294498 221586 294734
rect 221822 294498 257586 294734
rect 257822 294498 293586 294734
rect 293822 294498 329586 294734
rect 329822 294498 365586 294734
rect 365822 294498 401586 294734
rect 401822 294498 437586 294734
rect 437822 294498 473586 294734
rect 473822 294498 509586 294734
rect 509822 294498 545586 294734
rect 545822 294498 581586 294734
rect 581822 294498 587382 294734
rect 587618 294498 588740 294734
rect -4816 294476 588740 294498
rect -3876 294474 -3276 294476
rect 5404 294474 6004 294476
rect 41404 294474 42004 294476
rect 77404 294474 78004 294476
rect 113404 294474 114004 294476
rect 149404 294474 150004 294476
rect 185404 294474 186004 294476
rect 221404 294474 222004 294476
rect 257404 294474 258004 294476
rect 293404 294474 294004 294476
rect 329404 294474 330004 294476
rect 365404 294474 366004 294476
rect 401404 294474 402004 294476
rect 437404 294474 438004 294476
rect 473404 294474 474004 294476
rect 509404 294474 510004 294476
rect 545404 294474 546004 294476
rect 581404 294474 582004 294476
rect 587200 294474 587800 294476
rect -1996 291476 -1396 291478
rect 1804 291476 2404 291478
rect 37804 291476 38404 291478
rect 73804 291476 74404 291478
rect 109804 291476 110404 291478
rect 145804 291476 146404 291478
rect 181804 291476 182404 291478
rect 217804 291476 218404 291478
rect 253804 291476 254404 291478
rect 289804 291476 290404 291478
rect 325804 291476 326404 291478
rect 361804 291476 362404 291478
rect 397804 291476 398404 291478
rect 433804 291476 434404 291478
rect 469804 291476 470404 291478
rect 505804 291476 506404 291478
rect 541804 291476 542404 291478
rect 577804 291476 578404 291478
rect 585320 291476 585920 291478
rect -2936 291454 586860 291476
rect -2936 291218 -1814 291454
rect -1578 291218 1986 291454
rect 2222 291218 37986 291454
rect 38222 291218 73986 291454
rect 74222 291218 109986 291454
rect 110222 291218 145986 291454
rect 146222 291218 181986 291454
rect 182222 291218 217986 291454
rect 218222 291218 253986 291454
rect 254222 291218 289986 291454
rect 290222 291218 325986 291454
rect 326222 291218 361986 291454
rect 362222 291218 397986 291454
rect 398222 291218 433986 291454
rect 434222 291218 469986 291454
rect 470222 291218 505986 291454
rect 506222 291218 541986 291454
rect 542222 291218 577986 291454
rect 578222 291218 585502 291454
rect 585738 291218 586860 291454
rect -2936 291134 586860 291218
rect -2936 290898 -1814 291134
rect -1578 290898 1986 291134
rect 2222 290898 37986 291134
rect 38222 290898 73986 291134
rect 74222 290898 109986 291134
rect 110222 290898 145986 291134
rect 146222 290898 181986 291134
rect 182222 290898 217986 291134
rect 218222 290898 253986 291134
rect 254222 290898 289986 291134
rect 290222 290898 325986 291134
rect 326222 290898 361986 291134
rect 362222 290898 397986 291134
rect 398222 290898 433986 291134
rect 434222 290898 469986 291134
rect 470222 290898 505986 291134
rect 506222 290898 541986 291134
rect 542222 290898 577986 291134
rect 578222 290898 585502 291134
rect 585738 290898 586860 291134
rect -2936 290876 586860 290898
rect -1996 290874 -1396 290876
rect 1804 290874 2404 290876
rect 37804 290874 38404 290876
rect 73804 290874 74404 290876
rect 109804 290874 110404 290876
rect 145804 290874 146404 290876
rect 181804 290874 182404 290876
rect 217804 290874 218404 290876
rect 253804 290874 254404 290876
rect 289804 290874 290404 290876
rect 325804 290874 326404 290876
rect 361804 290874 362404 290876
rect 397804 290874 398404 290876
rect 433804 290874 434404 290876
rect 469804 290874 470404 290876
rect 505804 290874 506404 290876
rect 541804 290874 542404 290876
rect 577804 290874 578404 290876
rect 585320 290874 585920 290876
rect -8576 284276 -7976 284278
rect 30604 284276 31204 284278
rect 66604 284276 67204 284278
rect 102604 284276 103204 284278
rect 138604 284276 139204 284278
rect 174604 284276 175204 284278
rect 210604 284276 211204 284278
rect 246604 284276 247204 284278
rect 282604 284276 283204 284278
rect 318604 284276 319204 284278
rect 354604 284276 355204 284278
rect 390604 284276 391204 284278
rect 426604 284276 427204 284278
rect 462604 284276 463204 284278
rect 498604 284276 499204 284278
rect 534604 284276 535204 284278
rect 570604 284276 571204 284278
rect 591900 284276 592500 284278
rect -8576 284254 592500 284276
rect -8576 284018 -8394 284254
rect -8158 284018 30786 284254
rect 31022 284018 66786 284254
rect 67022 284018 102786 284254
rect 103022 284018 138786 284254
rect 139022 284018 174786 284254
rect 175022 284018 210786 284254
rect 211022 284018 246786 284254
rect 247022 284018 282786 284254
rect 283022 284018 318786 284254
rect 319022 284018 354786 284254
rect 355022 284018 390786 284254
rect 391022 284018 426786 284254
rect 427022 284018 462786 284254
rect 463022 284018 498786 284254
rect 499022 284018 534786 284254
rect 535022 284018 570786 284254
rect 571022 284018 592082 284254
rect 592318 284018 592500 284254
rect -8576 283934 592500 284018
rect -8576 283698 -8394 283934
rect -8158 283698 30786 283934
rect 31022 283698 66786 283934
rect 67022 283698 102786 283934
rect 103022 283698 138786 283934
rect 139022 283698 174786 283934
rect 175022 283698 210786 283934
rect 211022 283698 246786 283934
rect 247022 283698 282786 283934
rect 283022 283698 318786 283934
rect 319022 283698 354786 283934
rect 355022 283698 390786 283934
rect 391022 283698 426786 283934
rect 427022 283698 462786 283934
rect 463022 283698 498786 283934
rect 499022 283698 534786 283934
rect 535022 283698 570786 283934
rect 571022 283698 592082 283934
rect 592318 283698 592500 283934
rect -8576 283676 592500 283698
rect -8576 283674 -7976 283676
rect 30604 283674 31204 283676
rect 66604 283674 67204 283676
rect 102604 283674 103204 283676
rect 138604 283674 139204 283676
rect 174604 283674 175204 283676
rect 210604 283674 211204 283676
rect 246604 283674 247204 283676
rect 282604 283674 283204 283676
rect 318604 283674 319204 283676
rect 354604 283674 355204 283676
rect 390604 283674 391204 283676
rect 426604 283674 427204 283676
rect 462604 283674 463204 283676
rect 498604 283674 499204 283676
rect 534604 283674 535204 283676
rect 570604 283674 571204 283676
rect 591900 283674 592500 283676
rect -6696 280676 -6096 280678
rect 27004 280676 27604 280678
rect 63004 280676 63604 280678
rect 99004 280676 99604 280678
rect 135004 280676 135604 280678
rect 171004 280676 171604 280678
rect 207004 280676 207604 280678
rect 243004 280676 243604 280678
rect 279004 280676 279604 280678
rect 315004 280676 315604 280678
rect 351004 280676 351604 280678
rect 387004 280676 387604 280678
rect 423004 280676 423604 280678
rect 459004 280676 459604 280678
rect 495004 280676 495604 280678
rect 531004 280676 531604 280678
rect 567004 280676 567604 280678
rect 590020 280676 590620 280678
rect -6696 280654 590620 280676
rect -6696 280418 -6514 280654
rect -6278 280418 27186 280654
rect 27422 280418 63186 280654
rect 63422 280418 99186 280654
rect 99422 280418 135186 280654
rect 135422 280418 171186 280654
rect 171422 280418 207186 280654
rect 207422 280418 243186 280654
rect 243422 280418 279186 280654
rect 279422 280418 315186 280654
rect 315422 280418 351186 280654
rect 351422 280418 387186 280654
rect 387422 280418 423186 280654
rect 423422 280418 459186 280654
rect 459422 280418 495186 280654
rect 495422 280418 531186 280654
rect 531422 280418 567186 280654
rect 567422 280418 590202 280654
rect 590438 280418 590620 280654
rect -6696 280334 590620 280418
rect -6696 280098 -6514 280334
rect -6278 280098 27186 280334
rect 27422 280098 63186 280334
rect 63422 280098 99186 280334
rect 99422 280098 135186 280334
rect 135422 280098 171186 280334
rect 171422 280098 207186 280334
rect 207422 280098 243186 280334
rect 243422 280098 279186 280334
rect 279422 280098 315186 280334
rect 315422 280098 351186 280334
rect 351422 280098 387186 280334
rect 387422 280098 423186 280334
rect 423422 280098 459186 280334
rect 459422 280098 495186 280334
rect 495422 280098 531186 280334
rect 531422 280098 567186 280334
rect 567422 280098 590202 280334
rect 590438 280098 590620 280334
rect -6696 280076 590620 280098
rect -6696 280074 -6096 280076
rect 27004 280074 27604 280076
rect 63004 280074 63604 280076
rect 99004 280074 99604 280076
rect 135004 280074 135604 280076
rect 171004 280074 171604 280076
rect 207004 280074 207604 280076
rect 243004 280074 243604 280076
rect 279004 280074 279604 280076
rect 315004 280074 315604 280076
rect 351004 280074 351604 280076
rect 387004 280074 387604 280076
rect 423004 280074 423604 280076
rect 459004 280074 459604 280076
rect 495004 280074 495604 280076
rect 531004 280074 531604 280076
rect 567004 280074 567604 280076
rect 590020 280074 590620 280076
rect -4816 277076 -4216 277078
rect 23404 277076 24004 277078
rect 59404 277076 60004 277078
rect 95404 277076 96004 277078
rect 131404 277076 132004 277078
rect 167404 277076 168004 277078
rect 203404 277076 204004 277078
rect 239404 277076 240004 277078
rect 275404 277076 276004 277078
rect 311404 277076 312004 277078
rect 347404 277076 348004 277078
rect 383404 277076 384004 277078
rect 419404 277076 420004 277078
rect 455404 277076 456004 277078
rect 491404 277076 492004 277078
rect 527404 277076 528004 277078
rect 563404 277076 564004 277078
rect 588140 277076 588740 277078
rect -4816 277054 588740 277076
rect -4816 276818 -4634 277054
rect -4398 276818 23586 277054
rect 23822 276818 59586 277054
rect 59822 276818 95586 277054
rect 95822 276818 131586 277054
rect 131822 276818 167586 277054
rect 167822 276818 203586 277054
rect 203822 276818 239586 277054
rect 239822 276818 275586 277054
rect 275822 276818 311586 277054
rect 311822 276818 347586 277054
rect 347822 276818 383586 277054
rect 383822 276818 419586 277054
rect 419822 276818 455586 277054
rect 455822 276818 491586 277054
rect 491822 276818 527586 277054
rect 527822 276818 563586 277054
rect 563822 276818 588322 277054
rect 588558 276818 588740 277054
rect -4816 276734 588740 276818
rect -4816 276498 -4634 276734
rect -4398 276498 23586 276734
rect 23822 276498 59586 276734
rect 59822 276498 95586 276734
rect 95822 276498 131586 276734
rect 131822 276498 167586 276734
rect 167822 276498 203586 276734
rect 203822 276498 239586 276734
rect 239822 276498 275586 276734
rect 275822 276498 311586 276734
rect 311822 276498 347586 276734
rect 347822 276498 383586 276734
rect 383822 276498 419586 276734
rect 419822 276498 455586 276734
rect 455822 276498 491586 276734
rect 491822 276498 527586 276734
rect 527822 276498 563586 276734
rect 563822 276498 588322 276734
rect 588558 276498 588740 276734
rect -4816 276476 588740 276498
rect -4816 276474 -4216 276476
rect 23404 276474 24004 276476
rect 59404 276474 60004 276476
rect 95404 276474 96004 276476
rect 131404 276474 132004 276476
rect 167404 276474 168004 276476
rect 203404 276474 204004 276476
rect 239404 276474 240004 276476
rect 275404 276474 276004 276476
rect 311404 276474 312004 276476
rect 347404 276474 348004 276476
rect 383404 276474 384004 276476
rect 419404 276474 420004 276476
rect 455404 276474 456004 276476
rect 491404 276474 492004 276476
rect 527404 276474 528004 276476
rect 563404 276474 564004 276476
rect 588140 276474 588740 276476
rect -2936 273476 -2336 273478
rect 19804 273476 20404 273478
rect 55804 273476 56404 273478
rect 91804 273476 92404 273478
rect 127804 273476 128404 273478
rect 163804 273476 164404 273478
rect 199804 273476 200404 273478
rect 235804 273476 236404 273478
rect 271804 273476 272404 273478
rect 307804 273476 308404 273478
rect 343804 273476 344404 273478
rect 379804 273476 380404 273478
rect 415804 273476 416404 273478
rect 451804 273476 452404 273478
rect 487804 273476 488404 273478
rect 523804 273476 524404 273478
rect 559804 273476 560404 273478
rect 586260 273476 586860 273478
rect -2936 273454 586860 273476
rect -2936 273218 -2754 273454
rect -2518 273218 19986 273454
rect 20222 273218 55986 273454
rect 56222 273218 91986 273454
rect 92222 273218 127986 273454
rect 128222 273218 163986 273454
rect 164222 273218 199986 273454
rect 200222 273218 235986 273454
rect 236222 273218 271986 273454
rect 272222 273218 307986 273454
rect 308222 273218 343986 273454
rect 344222 273218 379986 273454
rect 380222 273218 415986 273454
rect 416222 273218 451986 273454
rect 452222 273218 487986 273454
rect 488222 273218 523986 273454
rect 524222 273218 559986 273454
rect 560222 273218 586442 273454
rect 586678 273218 586860 273454
rect -2936 273134 586860 273218
rect -2936 272898 -2754 273134
rect -2518 272898 19986 273134
rect 20222 272898 55986 273134
rect 56222 272898 91986 273134
rect 92222 272898 127986 273134
rect 128222 272898 163986 273134
rect 164222 272898 199986 273134
rect 200222 272898 235986 273134
rect 236222 272898 271986 273134
rect 272222 272898 307986 273134
rect 308222 272898 343986 273134
rect 344222 272898 379986 273134
rect 380222 272898 415986 273134
rect 416222 272898 451986 273134
rect 452222 272898 487986 273134
rect 488222 272898 523986 273134
rect 524222 272898 559986 273134
rect 560222 272898 586442 273134
rect 586678 272898 586860 273134
rect -2936 272876 586860 272898
rect -2936 272874 -2336 272876
rect 19804 272874 20404 272876
rect 55804 272874 56404 272876
rect 91804 272874 92404 272876
rect 127804 272874 128404 272876
rect 163804 272874 164404 272876
rect 199804 272874 200404 272876
rect 235804 272874 236404 272876
rect 271804 272874 272404 272876
rect 307804 272874 308404 272876
rect 343804 272874 344404 272876
rect 379804 272874 380404 272876
rect 415804 272874 416404 272876
rect 451804 272874 452404 272876
rect 487804 272874 488404 272876
rect 523804 272874 524404 272876
rect 559804 272874 560404 272876
rect 586260 272874 586860 272876
rect -7636 266276 -7036 266278
rect 12604 266276 13204 266278
rect 48604 266276 49204 266278
rect 84604 266276 85204 266278
rect 120604 266276 121204 266278
rect 156604 266276 157204 266278
rect 192604 266276 193204 266278
rect 228604 266276 229204 266278
rect 264604 266276 265204 266278
rect 300604 266276 301204 266278
rect 336604 266276 337204 266278
rect 372604 266276 373204 266278
rect 408604 266276 409204 266278
rect 444604 266276 445204 266278
rect 480604 266276 481204 266278
rect 516604 266276 517204 266278
rect 552604 266276 553204 266278
rect 590960 266276 591560 266278
rect -8576 266254 592500 266276
rect -8576 266018 -7454 266254
rect -7218 266018 12786 266254
rect 13022 266018 48786 266254
rect 49022 266018 84786 266254
rect 85022 266018 120786 266254
rect 121022 266018 156786 266254
rect 157022 266018 192786 266254
rect 193022 266018 228786 266254
rect 229022 266018 264786 266254
rect 265022 266018 300786 266254
rect 301022 266018 336786 266254
rect 337022 266018 372786 266254
rect 373022 266018 408786 266254
rect 409022 266018 444786 266254
rect 445022 266018 480786 266254
rect 481022 266018 516786 266254
rect 517022 266018 552786 266254
rect 553022 266018 591142 266254
rect 591378 266018 592500 266254
rect -8576 265934 592500 266018
rect -8576 265698 -7454 265934
rect -7218 265698 12786 265934
rect 13022 265698 48786 265934
rect 49022 265698 84786 265934
rect 85022 265698 120786 265934
rect 121022 265698 156786 265934
rect 157022 265698 192786 265934
rect 193022 265698 228786 265934
rect 229022 265698 264786 265934
rect 265022 265698 300786 265934
rect 301022 265698 336786 265934
rect 337022 265698 372786 265934
rect 373022 265698 408786 265934
rect 409022 265698 444786 265934
rect 445022 265698 480786 265934
rect 481022 265698 516786 265934
rect 517022 265698 552786 265934
rect 553022 265698 591142 265934
rect 591378 265698 592500 265934
rect -8576 265676 592500 265698
rect -7636 265674 -7036 265676
rect 12604 265674 13204 265676
rect 48604 265674 49204 265676
rect 84604 265674 85204 265676
rect 120604 265674 121204 265676
rect 156604 265674 157204 265676
rect 192604 265674 193204 265676
rect 228604 265674 229204 265676
rect 264604 265674 265204 265676
rect 300604 265674 301204 265676
rect 336604 265674 337204 265676
rect 372604 265674 373204 265676
rect 408604 265674 409204 265676
rect 444604 265674 445204 265676
rect 480604 265674 481204 265676
rect 516604 265674 517204 265676
rect 552604 265674 553204 265676
rect 590960 265674 591560 265676
rect -5756 262676 -5156 262678
rect 9004 262676 9604 262678
rect 45004 262676 45604 262678
rect 81004 262676 81604 262678
rect 117004 262676 117604 262678
rect 153004 262676 153604 262678
rect 189004 262676 189604 262678
rect 225004 262676 225604 262678
rect 261004 262676 261604 262678
rect 297004 262676 297604 262678
rect 333004 262676 333604 262678
rect 369004 262676 369604 262678
rect 405004 262676 405604 262678
rect 441004 262676 441604 262678
rect 477004 262676 477604 262678
rect 513004 262676 513604 262678
rect 549004 262676 549604 262678
rect 589080 262676 589680 262678
rect -6696 262654 590620 262676
rect -6696 262418 -5574 262654
rect -5338 262418 9186 262654
rect 9422 262418 45186 262654
rect 45422 262418 81186 262654
rect 81422 262418 117186 262654
rect 117422 262418 153186 262654
rect 153422 262418 189186 262654
rect 189422 262418 225186 262654
rect 225422 262418 261186 262654
rect 261422 262418 297186 262654
rect 297422 262418 333186 262654
rect 333422 262418 369186 262654
rect 369422 262418 405186 262654
rect 405422 262418 441186 262654
rect 441422 262418 477186 262654
rect 477422 262418 513186 262654
rect 513422 262418 549186 262654
rect 549422 262418 589262 262654
rect 589498 262418 590620 262654
rect -6696 262334 590620 262418
rect -6696 262098 -5574 262334
rect -5338 262098 9186 262334
rect 9422 262098 45186 262334
rect 45422 262098 81186 262334
rect 81422 262098 117186 262334
rect 117422 262098 153186 262334
rect 153422 262098 189186 262334
rect 189422 262098 225186 262334
rect 225422 262098 261186 262334
rect 261422 262098 297186 262334
rect 297422 262098 333186 262334
rect 333422 262098 369186 262334
rect 369422 262098 405186 262334
rect 405422 262098 441186 262334
rect 441422 262098 477186 262334
rect 477422 262098 513186 262334
rect 513422 262098 549186 262334
rect 549422 262098 589262 262334
rect 589498 262098 590620 262334
rect -6696 262076 590620 262098
rect -5756 262074 -5156 262076
rect 9004 262074 9604 262076
rect 45004 262074 45604 262076
rect 81004 262074 81604 262076
rect 117004 262074 117604 262076
rect 153004 262074 153604 262076
rect 189004 262074 189604 262076
rect 225004 262074 225604 262076
rect 261004 262074 261604 262076
rect 297004 262074 297604 262076
rect 333004 262074 333604 262076
rect 369004 262074 369604 262076
rect 405004 262074 405604 262076
rect 441004 262074 441604 262076
rect 477004 262074 477604 262076
rect 513004 262074 513604 262076
rect 549004 262074 549604 262076
rect 589080 262074 589680 262076
rect -3876 259076 -3276 259078
rect 5404 259076 6004 259078
rect 41404 259076 42004 259078
rect 77404 259076 78004 259078
rect 113404 259076 114004 259078
rect 149404 259076 150004 259078
rect 185404 259076 186004 259078
rect 221404 259076 222004 259078
rect 257404 259076 258004 259078
rect 293404 259076 294004 259078
rect 329404 259076 330004 259078
rect 365404 259076 366004 259078
rect 401404 259076 402004 259078
rect 437404 259076 438004 259078
rect 473404 259076 474004 259078
rect 509404 259076 510004 259078
rect 545404 259076 546004 259078
rect 581404 259076 582004 259078
rect 587200 259076 587800 259078
rect -4816 259054 588740 259076
rect -4816 258818 -3694 259054
rect -3458 258818 5586 259054
rect 5822 258818 41586 259054
rect 41822 258818 77586 259054
rect 77822 258818 113586 259054
rect 113822 258818 149586 259054
rect 149822 258818 185586 259054
rect 185822 258818 221586 259054
rect 221822 258818 257586 259054
rect 257822 258818 293586 259054
rect 293822 258818 329586 259054
rect 329822 258818 365586 259054
rect 365822 258818 401586 259054
rect 401822 258818 437586 259054
rect 437822 258818 473586 259054
rect 473822 258818 509586 259054
rect 509822 258818 545586 259054
rect 545822 258818 581586 259054
rect 581822 258818 587382 259054
rect 587618 258818 588740 259054
rect -4816 258734 588740 258818
rect -4816 258498 -3694 258734
rect -3458 258498 5586 258734
rect 5822 258498 41586 258734
rect 41822 258498 77586 258734
rect 77822 258498 113586 258734
rect 113822 258498 149586 258734
rect 149822 258498 185586 258734
rect 185822 258498 221586 258734
rect 221822 258498 257586 258734
rect 257822 258498 293586 258734
rect 293822 258498 329586 258734
rect 329822 258498 365586 258734
rect 365822 258498 401586 258734
rect 401822 258498 437586 258734
rect 437822 258498 473586 258734
rect 473822 258498 509586 258734
rect 509822 258498 545586 258734
rect 545822 258498 581586 258734
rect 581822 258498 587382 258734
rect 587618 258498 588740 258734
rect -4816 258476 588740 258498
rect -3876 258474 -3276 258476
rect 5404 258474 6004 258476
rect 41404 258474 42004 258476
rect 77404 258474 78004 258476
rect 113404 258474 114004 258476
rect 149404 258474 150004 258476
rect 185404 258474 186004 258476
rect 221404 258474 222004 258476
rect 257404 258474 258004 258476
rect 293404 258474 294004 258476
rect 329404 258474 330004 258476
rect 365404 258474 366004 258476
rect 401404 258474 402004 258476
rect 437404 258474 438004 258476
rect 473404 258474 474004 258476
rect 509404 258474 510004 258476
rect 545404 258474 546004 258476
rect 581404 258474 582004 258476
rect 587200 258474 587800 258476
rect -1996 255476 -1396 255478
rect 1804 255476 2404 255478
rect 37804 255476 38404 255478
rect 73804 255476 74404 255478
rect 109804 255476 110404 255478
rect 145804 255476 146404 255478
rect 181804 255476 182404 255478
rect 217804 255476 218404 255478
rect 253804 255476 254404 255478
rect 289804 255476 290404 255478
rect 325804 255476 326404 255478
rect 361804 255476 362404 255478
rect 397804 255476 398404 255478
rect 433804 255476 434404 255478
rect 469804 255476 470404 255478
rect 505804 255476 506404 255478
rect 541804 255476 542404 255478
rect 577804 255476 578404 255478
rect 585320 255476 585920 255478
rect -2936 255454 586860 255476
rect -2936 255218 -1814 255454
rect -1578 255218 1986 255454
rect 2222 255218 37986 255454
rect 38222 255218 73986 255454
rect 74222 255218 109986 255454
rect 110222 255218 145986 255454
rect 146222 255218 181986 255454
rect 182222 255218 217986 255454
rect 218222 255218 253986 255454
rect 254222 255218 289986 255454
rect 290222 255218 325986 255454
rect 326222 255218 361986 255454
rect 362222 255218 397986 255454
rect 398222 255218 433986 255454
rect 434222 255218 469986 255454
rect 470222 255218 505986 255454
rect 506222 255218 541986 255454
rect 542222 255218 577986 255454
rect 578222 255218 585502 255454
rect 585738 255218 586860 255454
rect -2936 255134 586860 255218
rect -2936 254898 -1814 255134
rect -1578 254898 1986 255134
rect 2222 254898 37986 255134
rect 38222 254898 73986 255134
rect 74222 254898 109986 255134
rect 110222 254898 145986 255134
rect 146222 254898 181986 255134
rect 182222 254898 217986 255134
rect 218222 254898 253986 255134
rect 254222 254898 289986 255134
rect 290222 254898 325986 255134
rect 326222 254898 361986 255134
rect 362222 254898 397986 255134
rect 398222 254898 433986 255134
rect 434222 254898 469986 255134
rect 470222 254898 505986 255134
rect 506222 254898 541986 255134
rect 542222 254898 577986 255134
rect 578222 254898 585502 255134
rect 585738 254898 586860 255134
rect -2936 254876 586860 254898
rect -1996 254874 -1396 254876
rect 1804 254874 2404 254876
rect 37804 254874 38404 254876
rect 73804 254874 74404 254876
rect 109804 254874 110404 254876
rect 145804 254874 146404 254876
rect 181804 254874 182404 254876
rect 217804 254874 218404 254876
rect 253804 254874 254404 254876
rect 289804 254874 290404 254876
rect 325804 254874 326404 254876
rect 361804 254874 362404 254876
rect 397804 254874 398404 254876
rect 433804 254874 434404 254876
rect 469804 254874 470404 254876
rect 505804 254874 506404 254876
rect 541804 254874 542404 254876
rect 577804 254874 578404 254876
rect 585320 254874 585920 254876
rect -8576 248276 -7976 248278
rect 30604 248276 31204 248278
rect 66604 248276 67204 248278
rect 102604 248276 103204 248278
rect 138604 248276 139204 248278
rect 174604 248276 175204 248278
rect 210604 248276 211204 248278
rect 246604 248276 247204 248278
rect 282604 248276 283204 248278
rect 318604 248276 319204 248278
rect 354604 248276 355204 248278
rect 390604 248276 391204 248278
rect 426604 248276 427204 248278
rect 462604 248276 463204 248278
rect 498604 248276 499204 248278
rect 534604 248276 535204 248278
rect 570604 248276 571204 248278
rect 591900 248276 592500 248278
rect -8576 248254 592500 248276
rect -8576 248018 -8394 248254
rect -8158 248018 30786 248254
rect 31022 248018 66786 248254
rect 67022 248018 102786 248254
rect 103022 248018 138786 248254
rect 139022 248018 174786 248254
rect 175022 248018 210786 248254
rect 211022 248018 246786 248254
rect 247022 248018 282786 248254
rect 283022 248018 318786 248254
rect 319022 248018 354786 248254
rect 355022 248018 390786 248254
rect 391022 248018 426786 248254
rect 427022 248018 462786 248254
rect 463022 248018 498786 248254
rect 499022 248018 534786 248254
rect 535022 248018 570786 248254
rect 571022 248018 592082 248254
rect 592318 248018 592500 248254
rect -8576 247934 592500 248018
rect -8576 247698 -8394 247934
rect -8158 247698 30786 247934
rect 31022 247698 66786 247934
rect 67022 247698 102786 247934
rect 103022 247698 138786 247934
rect 139022 247698 174786 247934
rect 175022 247698 210786 247934
rect 211022 247698 246786 247934
rect 247022 247698 282786 247934
rect 283022 247698 318786 247934
rect 319022 247698 354786 247934
rect 355022 247698 390786 247934
rect 391022 247698 426786 247934
rect 427022 247698 462786 247934
rect 463022 247698 498786 247934
rect 499022 247698 534786 247934
rect 535022 247698 570786 247934
rect 571022 247698 592082 247934
rect 592318 247698 592500 247934
rect -8576 247676 592500 247698
rect -8576 247674 -7976 247676
rect 30604 247674 31204 247676
rect 66604 247674 67204 247676
rect 102604 247674 103204 247676
rect 138604 247674 139204 247676
rect 174604 247674 175204 247676
rect 210604 247674 211204 247676
rect 246604 247674 247204 247676
rect 282604 247674 283204 247676
rect 318604 247674 319204 247676
rect 354604 247674 355204 247676
rect 390604 247674 391204 247676
rect 426604 247674 427204 247676
rect 462604 247674 463204 247676
rect 498604 247674 499204 247676
rect 534604 247674 535204 247676
rect 570604 247674 571204 247676
rect 591900 247674 592500 247676
rect -6696 244676 -6096 244678
rect 27004 244676 27604 244678
rect 63004 244676 63604 244678
rect 99004 244676 99604 244678
rect 135004 244676 135604 244678
rect 171004 244676 171604 244678
rect 207004 244676 207604 244678
rect 243004 244676 243604 244678
rect 279004 244676 279604 244678
rect 315004 244676 315604 244678
rect 351004 244676 351604 244678
rect 387004 244676 387604 244678
rect 423004 244676 423604 244678
rect 459004 244676 459604 244678
rect 495004 244676 495604 244678
rect 531004 244676 531604 244678
rect 567004 244676 567604 244678
rect 590020 244676 590620 244678
rect -6696 244654 590620 244676
rect -6696 244418 -6514 244654
rect -6278 244418 27186 244654
rect 27422 244418 63186 244654
rect 63422 244418 99186 244654
rect 99422 244418 135186 244654
rect 135422 244418 171186 244654
rect 171422 244418 207186 244654
rect 207422 244418 243186 244654
rect 243422 244418 279186 244654
rect 279422 244418 315186 244654
rect 315422 244418 351186 244654
rect 351422 244418 387186 244654
rect 387422 244418 423186 244654
rect 423422 244418 459186 244654
rect 459422 244418 495186 244654
rect 495422 244418 531186 244654
rect 531422 244418 567186 244654
rect 567422 244418 590202 244654
rect 590438 244418 590620 244654
rect -6696 244334 590620 244418
rect -6696 244098 -6514 244334
rect -6278 244098 27186 244334
rect 27422 244098 63186 244334
rect 63422 244098 99186 244334
rect 99422 244098 135186 244334
rect 135422 244098 171186 244334
rect 171422 244098 207186 244334
rect 207422 244098 243186 244334
rect 243422 244098 279186 244334
rect 279422 244098 315186 244334
rect 315422 244098 351186 244334
rect 351422 244098 387186 244334
rect 387422 244098 423186 244334
rect 423422 244098 459186 244334
rect 459422 244098 495186 244334
rect 495422 244098 531186 244334
rect 531422 244098 567186 244334
rect 567422 244098 590202 244334
rect 590438 244098 590620 244334
rect -6696 244076 590620 244098
rect -6696 244074 -6096 244076
rect 27004 244074 27604 244076
rect 63004 244074 63604 244076
rect 99004 244074 99604 244076
rect 135004 244074 135604 244076
rect 171004 244074 171604 244076
rect 207004 244074 207604 244076
rect 243004 244074 243604 244076
rect 279004 244074 279604 244076
rect 315004 244074 315604 244076
rect 351004 244074 351604 244076
rect 387004 244074 387604 244076
rect 423004 244074 423604 244076
rect 459004 244074 459604 244076
rect 495004 244074 495604 244076
rect 531004 244074 531604 244076
rect 567004 244074 567604 244076
rect 590020 244074 590620 244076
rect -4816 241076 -4216 241078
rect 23404 241076 24004 241078
rect 59404 241076 60004 241078
rect 95404 241076 96004 241078
rect 131404 241076 132004 241078
rect 167404 241076 168004 241078
rect 203404 241076 204004 241078
rect 239404 241076 240004 241078
rect 275404 241076 276004 241078
rect 311404 241076 312004 241078
rect 347404 241076 348004 241078
rect 383404 241076 384004 241078
rect 419404 241076 420004 241078
rect 455404 241076 456004 241078
rect 491404 241076 492004 241078
rect 527404 241076 528004 241078
rect 563404 241076 564004 241078
rect 588140 241076 588740 241078
rect -4816 241054 588740 241076
rect -4816 240818 -4634 241054
rect -4398 240818 23586 241054
rect 23822 240818 59586 241054
rect 59822 240818 95586 241054
rect 95822 240818 131586 241054
rect 131822 240818 167586 241054
rect 167822 240818 203586 241054
rect 203822 240818 239586 241054
rect 239822 240818 275586 241054
rect 275822 240818 311586 241054
rect 311822 240818 347586 241054
rect 347822 240818 383586 241054
rect 383822 240818 419586 241054
rect 419822 240818 455586 241054
rect 455822 240818 491586 241054
rect 491822 240818 527586 241054
rect 527822 240818 563586 241054
rect 563822 240818 588322 241054
rect 588558 240818 588740 241054
rect -4816 240734 588740 240818
rect -4816 240498 -4634 240734
rect -4398 240498 23586 240734
rect 23822 240498 59586 240734
rect 59822 240498 95586 240734
rect 95822 240498 131586 240734
rect 131822 240498 167586 240734
rect 167822 240498 203586 240734
rect 203822 240498 239586 240734
rect 239822 240498 275586 240734
rect 275822 240498 311586 240734
rect 311822 240498 347586 240734
rect 347822 240498 383586 240734
rect 383822 240498 419586 240734
rect 419822 240498 455586 240734
rect 455822 240498 491586 240734
rect 491822 240498 527586 240734
rect 527822 240498 563586 240734
rect 563822 240498 588322 240734
rect 588558 240498 588740 240734
rect -4816 240476 588740 240498
rect -4816 240474 -4216 240476
rect 23404 240474 24004 240476
rect 59404 240474 60004 240476
rect 95404 240474 96004 240476
rect 131404 240474 132004 240476
rect 167404 240474 168004 240476
rect 203404 240474 204004 240476
rect 239404 240474 240004 240476
rect 275404 240474 276004 240476
rect 311404 240474 312004 240476
rect 347404 240474 348004 240476
rect 383404 240474 384004 240476
rect 419404 240474 420004 240476
rect 455404 240474 456004 240476
rect 491404 240474 492004 240476
rect 527404 240474 528004 240476
rect 563404 240474 564004 240476
rect 588140 240474 588740 240476
rect -2936 237476 -2336 237478
rect 19804 237476 20404 237478
rect 55804 237476 56404 237478
rect 91804 237476 92404 237478
rect 127804 237476 128404 237478
rect 163804 237476 164404 237478
rect 199804 237476 200404 237478
rect 235804 237476 236404 237478
rect 271804 237476 272404 237478
rect 307804 237476 308404 237478
rect 343804 237476 344404 237478
rect 379804 237476 380404 237478
rect 415804 237476 416404 237478
rect 451804 237476 452404 237478
rect 487804 237476 488404 237478
rect 523804 237476 524404 237478
rect 559804 237476 560404 237478
rect 586260 237476 586860 237478
rect -2936 237454 586860 237476
rect -2936 237218 -2754 237454
rect -2518 237218 19986 237454
rect 20222 237218 55986 237454
rect 56222 237218 91986 237454
rect 92222 237218 127986 237454
rect 128222 237218 163986 237454
rect 164222 237218 199986 237454
rect 200222 237218 235986 237454
rect 236222 237218 271986 237454
rect 272222 237218 307986 237454
rect 308222 237218 343986 237454
rect 344222 237218 379986 237454
rect 380222 237218 415986 237454
rect 416222 237218 451986 237454
rect 452222 237218 487986 237454
rect 488222 237218 523986 237454
rect 524222 237218 559986 237454
rect 560222 237218 586442 237454
rect 586678 237218 586860 237454
rect -2936 237134 586860 237218
rect -2936 236898 -2754 237134
rect -2518 236898 19986 237134
rect 20222 236898 55986 237134
rect 56222 236898 91986 237134
rect 92222 236898 127986 237134
rect 128222 236898 163986 237134
rect 164222 236898 199986 237134
rect 200222 236898 235986 237134
rect 236222 236898 271986 237134
rect 272222 236898 307986 237134
rect 308222 236898 343986 237134
rect 344222 236898 379986 237134
rect 380222 236898 415986 237134
rect 416222 236898 451986 237134
rect 452222 236898 487986 237134
rect 488222 236898 523986 237134
rect 524222 236898 559986 237134
rect 560222 236898 586442 237134
rect 586678 236898 586860 237134
rect -2936 236876 586860 236898
rect -2936 236874 -2336 236876
rect 19804 236874 20404 236876
rect 55804 236874 56404 236876
rect 91804 236874 92404 236876
rect 127804 236874 128404 236876
rect 163804 236874 164404 236876
rect 199804 236874 200404 236876
rect 235804 236874 236404 236876
rect 271804 236874 272404 236876
rect 307804 236874 308404 236876
rect 343804 236874 344404 236876
rect 379804 236874 380404 236876
rect 415804 236874 416404 236876
rect 451804 236874 452404 236876
rect 487804 236874 488404 236876
rect 523804 236874 524404 236876
rect 559804 236874 560404 236876
rect 586260 236874 586860 236876
rect -7636 230276 -7036 230278
rect 12604 230276 13204 230278
rect 48604 230276 49204 230278
rect 84604 230276 85204 230278
rect 120604 230276 121204 230278
rect 156604 230276 157204 230278
rect 192604 230276 193204 230278
rect 228604 230276 229204 230278
rect 264604 230276 265204 230278
rect 300604 230276 301204 230278
rect 336604 230276 337204 230278
rect 372604 230276 373204 230278
rect 408604 230276 409204 230278
rect 444604 230276 445204 230278
rect 480604 230276 481204 230278
rect 516604 230276 517204 230278
rect 552604 230276 553204 230278
rect 590960 230276 591560 230278
rect -8576 230254 592500 230276
rect -8576 230018 -7454 230254
rect -7218 230018 12786 230254
rect 13022 230018 48786 230254
rect 49022 230018 84786 230254
rect 85022 230018 120786 230254
rect 121022 230018 156786 230254
rect 157022 230018 192786 230254
rect 193022 230018 228786 230254
rect 229022 230018 264786 230254
rect 265022 230018 300786 230254
rect 301022 230018 336786 230254
rect 337022 230018 372786 230254
rect 373022 230018 408786 230254
rect 409022 230018 444786 230254
rect 445022 230018 480786 230254
rect 481022 230018 516786 230254
rect 517022 230018 552786 230254
rect 553022 230018 591142 230254
rect 591378 230018 592500 230254
rect -8576 229934 592500 230018
rect -8576 229698 -7454 229934
rect -7218 229698 12786 229934
rect 13022 229698 48786 229934
rect 49022 229698 84786 229934
rect 85022 229698 120786 229934
rect 121022 229698 156786 229934
rect 157022 229698 192786 229934
rect 193022 229698 228786 229934
rect 229022 229698 264786 229934
rect 265022 229698 300786 229934
rect 301022 229698 336786 229934
rect 337022 229698 372786 229934
rect 373022 229698 408786 229934
rect 409022 229698 444786 229934
rect 445022 229698 480786 229934
rect 481022 229698 516786 229934
rect 517022 229698 552786 229934
rect 553022 229698 591142 229934
rect 591378 229698 592500 229934
rect -8576 229676 592500 229698
rect -7636 229674 -7036 229676
rect 12604 229674 13204 229676
rect 48604 229674 49204 229676
rect 84604 229674 85204 229676
rect 120604 229674 121204 229676
rect 156604 229674 157204 229676
rect 192604 229674 193204 229676
rect 228604 229674 229204 229676
rect 264604 229674 265204 229676
rect 300604 229674 301204 229676
rect 336604 229674 337204 229676
rect 372604 229674 373204 229676
rect 408604 229674 409204 229676
rect 444604 229674 445204 229676
rect 480604 229674 481204 229676
rect 516604 229674 517204 229676
rect 552604 229674 553204 229676
rect 590960 229674 591560 229676
rect -5756 226676 -5156 226678
rect 9004 226676 9604 226678
rect 45004 226676 45604 226678
rect 81004 226676 81604 226678
rect 117004 226676 117604 226678
rect 153004 226676 153604 226678
rect 189004 226676 189604 226678
rect 225004 226676 225604 226678
rect 261004 226676 261604 226678
rect 297004 226676 297604 226678
rect 333004 226676 333604 226678
rect 369004 226676 369604 226678
rect 405004 226676 405604 226678
rect 441004 226676 441604 226678
rect 477004 226676 477604 226678
rect 513004 226676 513604 226678
rect 549004 226676 549604 226678
rect 589080 226676 589680 226678
rect -6696 226654 590620 226676
rect -6696 226418 -5574 226654
rect -5338 226418 9186 226654
rect 9422 226418 45186 226654
rect 45422 226418 81186 226654
rect 81422 226418 117186 226654
rect 117422 226418 153186 226654
rect 153422 226418 189186 226654
rect 189422 226418 225186 226654
rect 225422 226418 261186 226654
rect 261422 226418 297186 226654
rect 297422 226418 333186 226654
rect 333422 226418 369186 226654
rect 369422 226418 405186 226654
rect 405422 226418 441186 226654
rect 441422 226418 477186 226654
rect 477422 226418 513186 226654
rect 513422 226418 549186 226654
rect 549422 226418 589262 226654
rect 589498 226418 590620 226654
rect -6696 226334 590620 226418
rect -6696 226098 -5574 226334
rect -5338 226098 9186 226334
rect 9422 226098 45186 226334
rect 45422 226098 81186 226334
rect 81422 226098 117186 226334
rect 117422 226098 153186 226334
rect 153422 226098 189186 226334
rect 189422 226098 225186 226334
rect 225422 226098 261186 226334
rect 261422 226098 297186 226334
rect 297422 226098 333186 226334
rect 333422 226098 369186 226334
rect 369422 226098 405186 226334
rect 405422 226098 441186 226334
rect 441422 226098 477186 226334
rect 477422 226098 513186 226334
rect 513422 226098 549186 226334
rect 549422 226098 589262 226334
rect 589498 226098 590620 226334
rect -6696 226076 590620 226098
rect -5756 226074 -5156 226076
rect 9004 226074 9604 226076
rect 45004 226074 45604 226076
rect 81004 226074 81604 226076
rect 117004 226074 117604 226076
rect 153004 226074 153604 226076
rect 189004 226074 189604 226076
rect 225004 226074 225604 226076
rect 261004 226074 261604 226076
rect 297004 226074 297604 226076
rect 333004 226074 333604 226076
rect 369004 226074 369604 226076
rect 405004 226074 405604 226076
rect 441004 226074 441604 226076
rect 477004 226074 477604 226076
rect 513004 226074 513604 226076
rect 549004 226074 549604 226076
rect 589080 226074 589680 226076
rect -3876 223076 -3276 223078
rect 5404 223076 6004 223078
rect 41404 223076 42004 223078
rect 77404 223076 78004 223078
rect 113404 223076 114004 223078
rect 149404 223076 150004 223078
rect 185404 223076 186004 223078
rect 221404 223076 222004 223078
rect 257404 223076 258004 223078
rect 293404 223076 294004 223078
rect 329404 223076 330004 223078
rect 365404 223076 366004 223078
rect 401404 223076 402004 223078
rect 437404 223076 438004 223078
rect 473404 223076 474004 223078
rect 509404 223076 510004 223078
rect 545404 223076 546004 223078
rect 581404 223076 582004 223078
rect 587200 223076 587800 223078
rect -4816 223054 588740 223076
rect -4816 222818 -3694 223054
rect -3458 222818 5586 223054
rect 5822 222818 41586 223054
rect 41822 222818 77586 223054
rect 77822 222818 113586 223054
rect 113822 222818 149586 223054
rect 149822 222818 185586 223054
rect 185822 222818 221586 223054
rect 221822 222818 257586 223054
rect 257822 222818 293586 223054
rect 293822 222818 329586 223054
rect 329822 222818 365586 223054
rect 365822 222818 401586 223054
rect 401822 222818 437586 223054
rect 437822 222818 473586 223054
rect 473822 222818 509586 223054
rect 509822 222818 545586 223054
rect 545822 222818 581586 223054
rect 581822 222818 587382 223054
rect 587618 222818 588740 223054
rect -4816 222734 588740 222818
rect -4816 222498 -3694 222734
rect -3458 222498 5586 222734
rect 5822 222498 41586 222734
rect 41822 222498 77586 222734
rect 77822 222498 113586 222734
rect 113822 222498 149586 222734
rect 149822 222498 185586 222734
rect 185822 222498 221586 222734
rect 221822 222498 257586 222734
rect 257822 222498 293586 222734
rect 293822 222498 329586 222734
rect 329822 222498 365586 222734
rect 365822 222498 401586 222734
rect 401822 222498 437586 222734
rect 437822 222498 473586 222734
rect 473822 222498 509586 222734
rect 509822 222498 545586 222734
rect 545822 222498 581586 222734
rect 581822 222498 587382 222734
rect 587618 222498 588740 222734
rect -4816 222476 588740 222498
rect -3876 222474 -3276 222476
rect 5404 222474 6004 222476
rect 41404 222474 42004 222476
rect 77404 222474 78004 222476
rect 113404 222474 114004 222476
rect 149404 222474 150004 222476
rect 185404 222474 186004 222476
rect 221404 222474 222004 222476
rect 257404 222474 258004 222476
rect 293404 222474 294004 222476
rect 329404 222474 330004 222476
rect 365404 222474 366004 222476
rect 401404 222474 402004 222476
rect 437404 222474 438004 222476
rect 473404 222474 474004 222476
rect 509404 222474 510004 222476
rect 545404 222474 546004 222476
rect 581404 222474 582004 222476
rect 587200 222474 587800 222476
rect -1996 219476 -1396 219478
rect 1804 219476 2404 219478
rect 37804 219476 38404 219478
rect 73804 219476 74404 219478
rect 109804 219476 110404 219478
rect 145804 219476 146404 219478
rect 181804 219476 182404 219478
rect 217804 219476 218404 219478
rect 253804 219476 254404 219478
rect 289804 219476 290404 219478
rect 325804 219476 326404 219478
rect 361804 219476 362404 219478
rect 397804 219476 398404 219478
rect 433804 219476 434404 219478
rect 469804 219476 470404 219478
rect 505804 219476 506404 219478
rect 541804 219476 542404 219478
rect 577804 219476 578404 219478
rect 585320 219476 585920 219478
rect -2936 219454 586860 219476
rect -2936 219218 -1814 219454
rect -1578 219218 1986 219454
rect 2222 219218 37986 219454
rect 38222 219218 73986 219454
rect 74222 219218 109986 219454
rect 110222 219218 145986 219454
rect 146222 219218 181986 219454
rect 182222 219218 217986 219454
rect 218222 219218 253986 219454
rect 254222 219218 289986 219454
rect 290222 219218 325986 219454
rect 326222 219218 361986 219454
rect 362222 219218 397986 219454
rect 398222 219218 433986 219454
rect 434222 219218 469986 219454
rect 470222 219218 505986 219454
rect 506222 219218 541986 219454
rect 542222 219218 577986 219454
rect 578222 219218 585502 219454
rect 585738 219218 586860 219454
rect -2936 219134 586860 219218
rect -2936 218898 -1814 219134
rect -1578 218898 1986 219134
rect 2222 218898 37986 219134
rect 38222 218898 73986 219134
rect 74222 218898 109986 219134
rect 110222 218898 145986 219134
rect 146222 218898 181986 219134
rect 182222 218898 217986 219134
rect 218222 218898 253986 219134
rect 254222 218898 289986 219134
rect 290222 218898 325986 219134
rect 326222 218898 361986 219134
rect 362222 218898 397986 219134
rect 398222 218898 433986 219134
rect 434222 218898 469986 219134
rect 470222 218898 505986 219134
rect 506222 218898 541986 219134
rect 542222 218898 577986 219134
rect 578222 218898 585502 219134
rect 585738 218898 586860 219134
rect -2936 218876 586860 218898
rect -1996 218874 -1396 218876
rect 1804 218874 2404 218876
rect 37804 218874 38404 218876
rect 73804 218874 74404 218876
rect 109804 218874 110404 218876
rect 145804 218874 146404 218876
rect 181804 218874 182404 218876
rect 217804 218874 218404 218876
rect 253804 218874 254404 218876
rect 289804 218874 290404 218876
rect 325804 218874 326404 218876
rect 361804 218874 362404 218876
rect 397804 218874 398404 218876
rect 433804 218874 434404 218876
rect 469804 218874 470404 218876
rect 505804 218874 506404 218876
rect 541804 218874 542404 218876
rect 577804 218874 578404 218876
rect 585320 218874 585920 218876
rect -8576 212276 -7976 212278
rect 30604 212276 31204 212278
rect 66604 212276 67204 212278
rect 102604 212276 103204 212278
rect 138604 212276 139204 212278
rect 174604 212276 175204 212278
rect 210604 212276 211204 212278
rect 246604 212276 247204 212278
rect 282604 212276 283204 212278
rect 318604 212276 319204 212278
rect 354604 212276 355204 212278
rect 390604 212276 391204 212278
rect 426604 212276 427204 212278
rect 462604 212276 463204 212278
rect 498604 212276 499204 212278
rect 534604 212276 535204 212278
rect 570604 212276 571204 212278
rect 591900 212276 592500 212278
rect -8576 212254 592500 212276
rect -8576 212018 -8394 212254
rect -8158 212018 30786 212254
rect 31022 212018 66786 212254
rect 67022 212018 102786 212254
rect 103022 212018 138786 212254
rect 139022 212018 174786 212254
rect 175022 212018 210786 212254
rect 211022 212018 246786 212254
rect 247022 212018 282786 212254
rect 283022 212018 318786 212254
rect 319022 212018 354786 212254
rect 355022 212018 390786 212254
rect 391022 212018 426786 212254
rect 427022 212018 462786 212254
rect 463022 212018 498786 212254
rect 499022 212018 534786 212254
rect 535022 212018 570786 212254
rect 571022 212018 592082 212254
rect 592318 212018 592500 212254
rect -8576 211934 592500 212018
rect -8576 211698 -8394 211934
rect -8158 211698 30786 211934
rect 31022 211698 66786 211934
rect 67022 211698 102786 211934
rect 103022 211698 138786 211934
rect 139022 211698 174786 211934
rect 175022 211698 210786 211934
rect 211022 211698 246786 211934
rect 247022 211698 282786 211934
rect 283022 211698 318786 211934
rect 319022 211698 354786 211934
rect 355022 211698 390786 211934
rect 391022 211698 426786 211934
rect 427022 211698 462786 211934
rect 463022 211698 498786 211934
rect 499022 211698 534786 211934
rect 535022 211698 570786 211934
rect 571022 211698 592082 211934
rect 592318 211698 592500 211934
rect -8576 211676 592500 211698
rect -8576 211674 -7976 211676
rect 30604 211674 31204 211676
rect 66604 211674 67204 211676
rect 102604 211674 103204 211676
rect 138604 211674 139204 211676
rect 174604 211674 175204 211676
rect 210604 211674 211204 211676
rect 246604 211674 247204 211676
rect 282604 211674 283204 211676
rect 318604 211674 319204 211676
rect 354604 211674 355204 211676
rect 390604 211674 391204 211676
rect 426604 211674 427204 211676
rect 462604 211674 463204 211676
rect 498604 211674 499204 211676
rect 534604 211674 535204 211676
rect 570604 211674 571204 211676
rect 591900 211674 592500 211676
rect -6696 208676 -6096 208678
rect 27004 208676 27604 208678
rect 63004 208676 63604 208678
rect 99004 208676 99604 208678
rect 135004 208676 135604 208678
rect 171004 208676 171604 208678
rect 207004 208676 207604 208678
rect 243004 208676 243604 208678
rect 279004 208676 279604 208678
rect 315004 208676 315604 208678
rect 351004 208676 351604 208678
rect 387004 208676 387604 208678
rect 423004 208676 423604 208678
rect 459004 208676 459604 208678
rect 495004 208676 495604 208678
rect 531004 208676 531604 208678
rect 567004 208676 567604 208678
rect 590020 208676 590620 208678
rect -6696 208654 590620 208676
rect -6696 208418 -6514 208654
rect -6278 208418 27186 208654
rect 27422 208418 63186 208654
rect 63422 208418 99186 208654
rect 99422 208418 135186 208654
rect 135422 208418 171186 208654
rect 171422 208418 207186 208654
rect 207422 208418 243186 208654
rect 243422 208418 279186 208654
rect 279422 208418 315186 208654
rect 315422 208418 351186 208654
rect 351422 208418 387186 208654
rect 387422 208418 423186 208654
rect 423422 208418 459186 208654
rect 459422 208418 495186 208654
rect 495422 208418 531186 208654
rect 531422 208418 567186 208654
rect 567422 208418 590202 208654
rect 590438 208418 590620 208654
rect -6696 208334 590620 208418
rect -6696 208098 -6514 208334
rect -6278 208098 27186 208334
rect 27422 208098 63186 208334
rect 63422 208098 99186 208334
rect 99422 208098 135186 208334
rect 135422 208098 171186 208334
rect 171422 208098 207186 208334
rect 207422 208098 243186 208334
rect 243422 208098 279186 208334
rect 279422 208098 315186 208334
rect 315422 208098 351186 208334
rect 351422 208098 387186 208334
rect 387422 208098 423186 208334
rect 423422 208098 459186 208334
rect 459422 208098 495186 208334
rect 495422 208098 531186 208334
rect 531422 208098 567186 208334
rect 567422 208098 590202 208334
rect 590438 208098 590620 208334
rect -6696 208076 590620 208098
rect -6696 208074 -6096 208076
rect 27004 208074 27604 208076
rect 63004 208074 63604 208076
rect 99004 208074 99604 208076
rect 135004 208074 135604 208076
rect 171004 208074 171604 208076
rect 207004 208074 207604 208076
rect 243004 208074 243604 208076
rect 279004 208074 279604 208076
rect 315004 208074 315604 208076
rect 351004 208074 351604 208076
rect 387004 208074 387604 208076
rect 423004 208074 423604 208076
rect 459004 208074 459604 208076
rect 495004 208074 495604 208076
rect 531004 208074 531604 208076
rect 567004 208074 567604 208076
rect 590020 208074 590620 208076
rect -4816 205076 -4216 205078
rect 23404 205076 24004 205078
rect 59404 205076 60004 205078
rect 95404 205076 96004 205078
rect 131404 205076 132004 205078
rect 167404 205076 168004 205078
rect 203404 205076 204004 205078
rect 239404 205076 240004 205078
rect 275404 205076 276004 205078
rect 311404 205076 312004 205078
rect 347404 205076 348004 205078
rect 383404 205076 384004 205078
rect 419404 205076 420004 205078
rect 455404 205076 456004 205078
rect 491404 205076 492004 205078
rect 527404 205076 528004 205078
rect 563404 205076 564004 205078
rect 588140 205076 588740 205078
rect -4816 205054 588740 205076
rect -4816 204818 -4634 205054
rect -4398 204818 23586 205054
rect 23822 204818 59586 205054
rect 59822 204818 95586 205054
rect 95822 204818 131586 205054
rect 131822 204818 167586 205054
rect 167822 204818 203586 205054
rect 203822 204818 239586 205054
rect 239822 204818 275586 205054
rect 275822 204818 311586 205054
rect 311822 204818 347586 205054
rect 347822 204818 383586 205054
rect 383822 204818 419586 205054
rect 419822 204818 455586 205054
rect 455822 204818 491586 205054
rect 491822 204818 527586 205054
rect 527822 204818 563586 205054
rect 563822 204818 588322 205054
rect 588558 204818 588740 205054
rect -4816 204734 588740 204818
rect -4816 204498 -4634 204734
rect -4398 204498 23586 204734
rect 23822 204498 59586 204734
rect 59822 204498 95586 204734
rect 95822 204498 131586 204734
rect 131822 204498 167586 204734
rect 167822 204498 203586 204734
rect 203822 204498 239586 204734
rect 239822 204498 275586 204734
rect 275822 204498 311586 204734
rect 311822 204498 347586 204734
rect 347822 204498 383586 204734
rect 383822 204498 419586 204734
rect 419822 204498 455586 204734
rect 455822 204498 491586 204734
rect 491822 204498 527586 204734
rect 527822 204498 563586 204734
rect 563822 204498 588322 204734
rect 588558 204498 588740 204734
rect -4816 204476 588740 204498
rect -4816 204474 -4216 204476
rect 23404 204474 24004 204476
rect 59404 204474 60004 204476
rect 95404 204474 96004 204476
rect 131404 204474 132004 204476
rect 167404 204474 168004 204476
rect 203404 204474 204004 204476
rect 239404 204474 240004 204476
rect 275404 204474 276004 204476
rect 311404 204474 312004 204476
rect 347404 204474 348004 204476
rect 383404 204474 384004 204476
rect 419404 204474 420004 204476
rect 455404 204474 456004 204476
rect 491404 204474 492004 204476
rect 527404 204474 528004 204476
rect 563404 204474 564004 204476
rect 588140 204474 588740 204476
rect -2936 201476 -2336 201478
rect 19804 201476 20404 201478
rect 55804 201476 56404 201478
rect 91804 201476 92404 201478
rect 127804 201476 128404 201478
rect 163804 201476 164404 201478
rect 199804 201476 200404 201478
rect 235804 201476 236404 201478
rect 271804 201476 272404 201478
rect 307804 201476 308404 201478
rect 343804 201476 344404 201478
rect 379804 201476 380404 201478
rect 415804 201476 416404 201478
rect 451804 201476 452404 201478
rect 487804 201476 488404 201478
rect 523804 201476 524404 201478
rect 559804 201476 560404 201478
rect 586260 201476 586860 201478
rect -2936 201454 586860 201476
rect -2936 201218 -2754 201454
rect -2518 201218 19986 201454
rect 20222 201218 55986 201454
rect 56222 201218 91986 201454
rect 92222 201218 127986 201454
rect 128222 201218 163986 201454
rect 164222 201218 199986 201454
rect 200222 201218 235986 201454
rect 236222 201218 271986 201454
rect 272222 201218 307986 201454
rect 308222 201218 343986 201454
rect 344222 201218 379986 201454
rect 380222 201218 415986 201454
rect 416222 201218 451986 201454
rect 452222 201218 487986 201454
rect 488222 201218 523986 201454
rect 524222 201218 559986 201454
rect 560222 201218 586442 201454
rect 586678 201218 586860 201454
rect -2936 201134 586860 201218
rect -2936 200898 -2754 201134
rect -2518 200898 19986 201134
rect 20222 200898 55986 201134
rect 56222 200898 91986 201134
rect 92222 200898 127986 201134
rect 128222 200898 163986 201134
rect 164222 200898 199986 201134
rect 200222 200898 235986 201134
rect 236222 200898 271986 201134
rect 272222 200898 307986 201134
rect 308222 200898 343986 201134
rect 344222 200898 379986 201134
rect 380222 200898 415986 201134
rect 416222 200898 451986 201134
rect 452222 200898 487986 201134
rect 488222 200898 523986 201134
rect 524222 200898 559986 201134
rect 560222 200898 586442 201134
rect 586678 200898 586860 201134
rect -2936 200876 586860 200898
rect -2936 200874 -2336 200876
rect 19804 200874 20404 200876
rect 55804 200874 56404 200876
rect 91804 200874 92404 200876
rect 127804 200874 128404 200876
rect 163804 200874 164404 200876
rect 199804 200874 200404 200876
rect 235804 200874 236404 200876
rect 271804 200874 272404 200876
rect 307804 200874 308404 200876
rect 343804 200874 344404 200876
rect 379804 200874 380404 200876
rect 415804 200874 416404 200876
rect 451804 200874 452404 200876
rect 487804 200874 488404 200876
rect 523804 200874 524404 200876
rect 559804 200874 560404 200876
rect 586260 200874 586860 200876
rect -7636 194276 -7036 194278
rect 12604 194276 13204 194278
rect 48604 194276 49204 194278
rect 84604 194276 85204 194278
rect 120604 194276 121204 194278
rect 156604 194276 157204 194278
rect 192604 194276 193204 194278
rect 228604 194276 229204 194278
rect 264604 194276 265204 194278
rect 300604 194276 301204 194278
rect 336604 194276 337204 194278
rect 372604 194276 373204 194278
rect 408604 194276 409204 194278
rect 444604 194276 445204 194278
rect 480604 194276 481204 194278
rect 516604 194276 517204 194278
rect 552604 194276 553204 194278
rect 590960 194276 591560 194278
rect -8576 194254 592500 194276
rect -8576 194018 -7454 194254
rect -7218 194018 12786 194254
rect 13022 194018 48786 194254
rect 49022 194018 84786 194254
rect 85022 194018 120786 194254
rect 121022 194018 156786 194254
rect 157022 194018 192786 194254
rect 193022 194018 228786 194254
rect 229022 194018 264786 194254
rect 265022 194018 300786 194254
rect 301022 194018 336786 194254
rect 337022 194018 372786 194254
rect 373022 194018 408786 194254
rect 409022 194018 444786 194254
rect 445022 194018 480786 194254
rect 481022 194018 516786 194254
rect 517022 194018 552786 194254
rect 553022 194018 591142 194254
rect 591378 194018 592500 194254
rect -8576 193934 592500 194018
rect -8576 193698 -7454 193934
rect -7218 193698 12786 193934
rect 13022 193698 48786 193934
rect 49022 193698 84786 193934
rect 85022 193698 120786 193934
rect 121022 193698 156786 193934
rect 157022 193698 192786 193934
rect 193022 193698 228786 193934
rect 229022 193698 264786 193934
rect 265022 193698 300786 193934
rect 301022 193698 336786 193934
rect 337022 193698 372786 193934
rect 373022 193698 408786 193934
rect 409022 193698 444786 193934
rect 445022 193698 480786 193934
rect 481022 193698 516786 193934
rect 517022 193698 552786 193934
rect 553022 193698 591142 193934
rect 591378 193698 592500 193934
rect -8576 193676 592500 193698
rect -7636 193674 -7036 193676
rect 12604 193674 13204 193676
rect 48604 193674 49204 193676
rect 84604 193674 85204 193676
rect 120604 193674 121204 193676
rect 156604 193674 157204 193676
rect 192604 193674 193204 193676
rect 228604 193674 229204 193676
rect 264604 193674 265204 193676
rect 300604 193674 301204 193676
rect 336604 193674 337204 193676
rect 372604 193674 373204 193676
rect 408604 193674 409204 193676
rect 444604 193674 445204 193676
rect 480604 193674 481204 193676
rect 516604 193674 517204 193676
rect 552604 193674 553204 193676
rect 590960 193674 591560 193676
rect -5756 190676 -5156 190678
rect 9004 190676 9604 190678
rect 45004 190676 45604 190678
rect 81004 190676 81604 190678
rect 117004 190676 117604 190678
rect 153004 190676 153604 190678
rect 189004 190676 189604 190678
rect 225004 190676 225604 190678
rect 261004 190676 261604 190678
rect 297004 190676 297604 190678
rect 333004 190676 333604 190678
rect 369004 190676 369604 190678
rect 405004 190676 405604 190678
rect 441004 190676 441604 190678
rect 477004 190676 477604 190678
rect 513004 190676 513604 190678
rect 549004 190676 549604 190678
rect 589080 190676 589680 190678
rect -6696 190654 590620 190676
rect -6696 190418 -5574 190654
rect -5338 190418 9186 190654
rect 9422 190418 45186 190654
rect 45422 190418 81186 190654
rect 81422 190418 117186 190654
rect 117422 190418 153186 190654
rect 153422 190418 189186 190654
rect 189422 190418 225186 190654
rect 225422 190418 261186 190654
rect 261422 190418 297186 190654
rect 297422 190418 333186 190654
rect 333422 190418 369186 190654
rect 369422 190418 405186 190654
rect 405422 190418 441186 190654
rect 441422 190418 477186 190654
rect 477422 190418 513186 190654
rect 513422 190418 549186 190654
rect 549422 190418 589262 190654
rect 589498 190418 590620 190654
rect -6696 190334 590620 190418
rect -6696 190098 -5574 190334
rect -5338 190098 9186 190334
rect 9422 190098 45186 190334
rect 45422 190098 81186 190334
rect 81422 190098 117186 190334
rect 117422 190098 153186 190334
rect 153422 190098 189186 190334
rect 189422 190098 225186 190334
rect 225422 190098 261186 190334
rect 261422 190098 297186 190334
rect 297422 190098 333186 190334
rect 333422 190098 369186 190334
rect 369422 190098 405186 190334
rect 405422 190098 441186 190334
rect 441422 190098 477186 190334
rect 477422 190098 513186 190334
rect 513422 190098 549186 190334
rect 549422 190098 589262 190334
rect 589498 190098 590620 190334
rect -6696 190076 590620 190098
rect -5756 190074 -5156 190076
rect 9004 190074 9604 190076
rect 45004 190074 45604 190076
rect 81004 190074 81604 190076
rect 117004 190074 117604 190076
rect 153004 190074 153604 190076
rect 189004 190074 189604 190076
rect 225004 190074 225604 190076
rect 261004 190074 261604 190076
rect 297004 190074 297604 190076
rect 333004 190074 333604 190076
rect 369004 190074 369604 190076
rect 405004 190074 405604 190076
rect 441004 190074 441604 190076
rect 477004 190074 477604 190076
rect 513004 190074 513604 190076
rect 549004 190074 549604 190076
rect 589080 190074 589680 190076
rect -3876 187076 -3276 187078
rect 5404 187076 6004 187078
rect 41404 187076 42004 187078
rect 77404 187076 78004 187078
rect 113404 187076 114004 187078
rect 149404 187076 150004 187078
rect 185404 187076 186004 187078
rect 221404 187076 222004 187078
rect 257404 187076 258004 187078
rect 293404 187076 294004 187078
rect 329404 187076 330004 187078
rect 365404 187076 366004 187078
rect 401404 187076 402004 187078
rect 437404 187076 438004 187078
rect 473404 187076 474004 187078
rect 509404 187076 510004 187078
rect 545404 187076 546004 187078
rect 581404 187076 582004 187078
rect 587200 187076 587800 187078
rect -4816 187054 588740 187076
rect -4816 186818 -3694 187054
rect -3458 186818 5586 187054
rect 5822 186818 41586 187054
rect 41822 186818 77586 187054
rect 77822 186818 113586 187054
rect 113822 186818 149586 187054
rect 149822 186818 185586 187054
rect 185822 186818 221586 187054
rect 221822 186818 257586 187054
rect 257822 186818 293586 187054
rect 293822 186818 329586 187054
rect 329822 186818 365586 187054
rect 365822 186818 401586 187054
rect 401822 186818 437586 187054
rect 437822 186818 473586 187054
rect 473822 186818 509586 187054
rect 509822 186818 545586 187054
rect 545822 186818 581586 187054
rect 581822 186818 587382 187054
rect 587618 186818 588740 187054
rect -4816 186734 588740 186818
rect -4816 186498 -3694 186734
rect -3458 186498 5586 186734
rect 5822 186498 41586 186734
rect 41822 186498 77586 186734
rect 77822 186498 113586 186734
rect 113822 186498 149586 186734
rect 149822 186498 185586 186734
rect 185822 186498 221586 186734
rect 221822 186498 257586 186734
rect 257822 186498 293586 186734
rect 293822 186498 329586 186734
rect 329822 186498 365586 186734
rect 365822 186498 401586 186734
rect 401822 186498 437586 186734
rect 437822 186498 473586 186734
rect 473822 186498 509586 186734
rect 509822 186498 545586 186734
rect 545822 186498 581586 186734
rect 581822 186498 587382 186734
rect 587618 186498 588740 186734
rect -4816 186476 588740 186498
rect -3876 186474 -3276 186476
rect 5404 186474 6004 186476
rect 41404 186474 42004 186476
rect 77404 186474 78004 186476
rect 113404 186474 114004 186476
rect 149404 186474 150004 186476
rect 185404 186474 186004 186476
rect 221404 186474 222004 186476
rect 257404 186474 258004 186476
rect 293404 186474 294004 186476
rect 329404 186474 330004 186476
rect 365404 186474 366004 186476
rect 401404 186474 402004 186476
rect 437404 186474 438004 186476
rect 473404 186474 474004 186476
rect 509404 186474 510004 186476
rect 545404 186474 546004 186476
rect 581404 186474 582004 186476
rect 587200 186474 587800 186476
rect -1996 183476 -1396 183478
rect 1804 183476 2404 183478
rect 37804 183476 38404 183478
rect 73804 183476 74404 183478
rect 109804 183476 110404 183478
rect 145804 183476 146404 183478
rect 181804 183476 182404 183478
rect 217804 183476 218404 183478
rect 253804 183476 254404 183478
rect 289804 183476 290404 183478
rect 325804 183476 326404 183478
rect 361804 183476 362404 183478
rect 397804 183476 398404 183478
rect 433804 183476 434404 183478
rect 469804 183476 470404 183478
rect 505804 183476 506404 183478
rect 541804 183476 542404 183478
rect 577804 183476 578404 183478
rect 585320 183476 585920 183478
rect -2936 183454 586860 183476
rect -2936 183218 -1814 183454
rect -1578 183218 1986 183454
rect 2222 183218 37986 183454
rect 38222 183218 73986 183454
rect 74222 183218 109986 183454
rect 110222 183218 145986 183454
rect 146222 183218 181986 183454
rect 182222 183218 217986 183454
rect 218222 183218 253986 183454
rect 254222 183218 289986 183454
rect 290222 183218 325986 183454
rect 326222 183218 361986 183454
rect 362222 183218 397986 183454
rect 398222 183218 433986 183454
rect 434222 183218 469986 183454
rect 470222 183218 505986 183454
rect 506222 183218 541986 183454
rect 542222 183218 577986 183454
rect 578222 183218 585502 183454
rect 585738 183218 586860 183454
rect -2936 183134 586860 183218
rect -2936 182898 -1814 183134
rect -1578 182898 1986 183134
rect 2222 182898 37986 183134
rect 38222 182898 73986 183134
rect 74222 182898 109986 183134
rect 110222 182898 145986 183134
rect 146222 182898 181986 183134
rect 182222 182898 217986 183134
rect 218222 182898 253986 183134
rect 254222 182898 289986 183134
rect 290222 182898 325986 183134
rect 326222 182898 361986 183134
rect 362222 182898 397986 183134
rect 398222 182898 433986 183134
rect 434222 182898 469986 183134
rect 470222 182898 505986 183134
rect 506222 182898 541986 183134
rect 542222 182898 577986 183134
rect 578222 182898 585502 183134
rect 585738 182898 586860 183134
rect -2936 182876 586860 182898
rect -1996 182874 -1396 182876
rect 1804 182874 2404 182876
rect 37804 182874 38404 182876
rect 73804 182874 74404 182876
rect 109804 182874 110404 182876
rect 145804 182874 146404 182876
rect 181804 182874 182404 182876
rect 217804 182874 218404 182876
rect 253804 182874 254404 182876
rect 289804 182874 290404 182876
rect 325804 182874 326404 182876
rect 361804 182874 362404 182876
rect 397804 182874 398404 182876
rect 433804 182874 434404 182876
rect 469804 182874 470404 182876
rect 505804 182874 506404 182876
rect 541804 182874 542404 182876
rect 577804 182874 578404 182876
rect 585320 182874 585920 182876
rect -8576 176276 -7976 176278
rect 30604 176276 31204 176278
rect 66604 176276 67204 176278
rect 102604 176276 103204 176278
rect 138604 176276 139204 176278
rect 174604 176276 175204 176278
rect 210604 176276 211204 176278
rect 246604 176276 247204 176278
rect 282604 176276 283204 176278
rect 318604 176276 319204 176278
rect 354604 176276 355204 176278
rect 390604 176276 391204 176278
rect 426604 176276 427204 176278
rect 462604 176276 463204 176278
rect 498604 176276 499204 176278
rect 534604 176276 535204 176278
rect 570604 176276 571204 176278
rect 591900 176276 592500 176278
rect -8576 176254 592500 176276
rect -8576 176018 -8394 176254
rect -8158 176018 30786 176254
rect 31022 176018 66786 176254
rect 67022 176018 102786 176254
rect 103022 176018 138786 176254
rect 139022 176018 174786 176254
rect 175022 176018 210786 176254
rect 211022 176018 246786 176254
rect 247022 176018 282786 176254
rect 283022 176018 318786 176254
rect 319022 176018 354786 176254
rect 355022 176018 390786 176254
rect 391022 176018 426786 176254
rect 427022 176018 462786 176254
rect 463022 176018 498786 176254
rect 499022 176018 534786 176254
rect 535022 176018 570786 176254
rect 571022 176018 592082 176254
rect 592318 176018 592500 176254
rect -8576 175934 592500 176018
rect -8576 175698 -8394 175934
rect -8158 175698 30786 175934
rect 31022 175698 66786 175934
rect 67022 175698 102786 175934
rect 103022 175698 138786 175934
rect 139022 175698 174786 175934
rect 175022 175698 210786 175934
rect 211022 175698 246786 175934
rect 247022 175698 282786 175934
rect 283022 175698 318786 175934
rect 319022 175698 354786 175934
rect 355022 175698 390786 175934
rect 391022 175698 426786 175934
rect 427022 175698 462786 175934
rect 463022 175698 498786 175934
rect 499022 175698 534786 175934
rect 535022 175698 570786 175934
rect 571022 175698 592082 175934
rect 592318 175698 592500 175934
rect -8576 175676 592500 175698
rect -8576 175674 -7976 175676
rect 30604 175674 31204 175676
rect 66604 175674 67204 175676
rect 102604 175674 103204 175676
rect 138604 175674 139204 175676
rect 174604 175674 175204 175676
rect 210604 175674 211204 175676
rect 246604 175674 247204 175676
rect 282604 175674 283204 175676
rect 318604 175674 319204 175676
rect 354604 175674 355204 175676
rect 390604 175674 391204 175676
rect 426604 175674 427204 175676
rect 462604 175674 463204 175676
rect 498604 175674 499204 175676
rect 534604 175674 535204 175676
rect 570604 175674 571204 175676
rect 591900 175674 592500 175676
rect -6696 172676 -6096 172678
rect 27004 172676 27604 172678
rect 63004 172676 63604 172678
rect 99004 172676 99604 172678
rect 135004 172676 135604 172678
rect 171004 172676 171604 172678
rect 207004 172676 207604 172678
rect 243004 172676 243604 172678
rect 279004 172676 279604 172678
rect 315004 172676 315604 172678
rect 351004 172676 351604 172678
rect 387004 172676 387604 172678
rect 423004 172676 423604 172678
rect 459004 172676 459604 172678
rect 495004 172676 495604 172678
rect 531004 172676 531604 172678
rect 567004 172676 567604 172678
rect 590020 172676 590620 172678
rect -6696 172654 590620 172676
rect -6696 172418 -6514 172654
rect -6278 172418 27186 172654
rect 27422 172418 63186 172654
rect 63422 172418 99186 172654
rect 99422 172418 135186 172654
rect 135422 172418 171186 172654
rect 171422 172418 207186 172654
rect 207422 172418 243186 172654
rect 243422 172418 279186 172654
rect 279422 172418 315186 172654
rect 315422 172418 351186 172654
rect 351422 172418 387186 172654
rect 387422 172418 423186 172654
rect 423422 172418 459186 172654
rect 459422 172418 495186 172654
rect 495422 172418 531186 172654
rect 531422 172418 567186 172654
rect 567422 172418 590202 172654
rect 590438 172418 590620 172654
rect -6696 172334 590620 172418
rect -6696 172098 -6514 172334
rect -6278 172098 27186 172334
rect 27422 172098 63186 172334
rect 63422 172098 99186 172334
rect 99422 172098 135186 172334
rect 135422 172098 171186 172334
rect 171422 172098 207186 172334
rect 207422 172098 243186 172334
rect 243422 172098 279186 172334
rect 279422 172098 315186 172334
rect 315422 172098 351186 172334
rect 351422 172098 387186 172334
rect 387422 172098 423186 172334
rect 423422 172098 459186 172334
rect 459422 172098 495186 172334
rect 495422 172098 531186 172334
rect 531422 172098 567186 172334
rect 567422 172098 590202 172334
rect 590438 172098 590620 172334
rect -6696 172076 590620 172098
rect -6696 172074 -6096 172076
rect 27004 172074 27604 172076
rect 63004 172074 63604 172076
rect 99004 172074 99604 172076
rect 135004 172074 135604 172076
rect 171004 172074 171604 172076
rect 207004 172074 207604 172076
rect 243004 172074 243604 172076
rect 279004 172074 279604 172076
rect 315004 172074 315604 172076
rect 351004 172074 351604 172076
rect 387004 172074 387604 172076
rect 423004 172074 423604 172076
rect 459004 172074 459604 172076
rect 495004 172074 495604 172076
rect 531004 172074 531604 172076
rect 567004 172074 567604 172076
rect 590020 172074 590620 172076
rect -4816 169076 -4216 169078
rect 23404 169076 24004 169078
rect 59404 169076 60004 169078
rect 95404 169076 96004 169078
rect 131404 169076 132004 169078
rect 167404 169076 168004 169078
rect 203404 169076 204004 169078
rect 239404 169076 240004 169078
rect 275404 169076 276004 169078
rect 311404 169076 312004 169078
rect 347404 169076 348004 169078
rect 383404 169076 384004 169078
rect 419404 169076 420004 169078
rect 455404 169076 456004 169078
rect 491404 169076 492004 169078
rect 527404 169076 528004 169078
rect 563404 169076 564004 169078
rect 588140 169076 588740 169078
rect -4816 169054 588740 169076
rect -4816 168818 -4634 169054
rect -4398 168818 23586 169054
rect 23822 168818 59586 169054
rect 59822 168818 95586 169054
rect 95822 168818 131586 169054
rect 131822 168818 167586 169054
rect 167822 168818 203586 169054
rect 203822 168818 239586 169054
rect 239822 168818 275586 169054
rect 275822 168818 311586 169054
rect 311822 168818 347586 169054
rect 347822 168818 383586 169054
rect 383822 168818 419586 169054
rect 419822 168818 455586 169054
rect 455822 168818 491586 169054
rect 491822 168818 527586 169054
rect 527822 168818 563586 169054
rect 563822 168818 588322 169054
rect 588558 168818 588740 169054
rect -4816 168734 588740 168818
rect -4816 168498 -4634 168734
rect -4398 168498 23586 168734
rect 23822 168498 59586 168734
rect 59822 168498 95586 168734
rect 95822 168498 131586 168734
rect 131822 168498 167586 168734
rect 167822 168498 203586 168734
rect 203822 168498 239586 168734
rect 239822 168498 275586 168734
rect 275822 168498 311586 168734
rect 311822 168498 347586 168734
rect 347822 168498 383586 168734
rect 383822 168498 419586 168734
rect 419822 168498 455586 168734
rect 455822 168498 491586 168734
rect 491822 168498 527586 168734
rect 527822 168498 563586 168734
rect 563822 168498 588322 168734
rect 588558 168498 588740 168734
rect -4816 168476 588740 168498
rect -4816 168474 -4216 168476
rect 23404 168474 24004 168476
rect 59404 168474 60004 168476
rect 95404 168474 96004 168476
rect 131404 168474 132004 168476
rect 167404 168474 168004 168476
rect 203404 168474 204004 168476
rect 239404 168474 240004 168476
rect 275404 168474 276004 168476
rect 311404 168474 312004 168476
rect 347404 168474 348004 168476
rect 383404 168474 384004 168476
rect 419404 168474 420004 168476
rect 455404 168474 456004 168476
rect 491404 168474 492004 168476
rect 527404 168474 528004 168476
rect 563404 168474 564004 168476
rect 588140 168474 588740 168476
rect -2936 165476 -2336 165478
rect 19804 165476 20404 165478
rect 55804 165476 56404 165478
rect 91804 165476 92404 165478
rect 127804 165476 128404 165478
rect 163804 165476 164404 165478
rect 199804 165476 200404 165478
rect 235804 165476 236404 165478
rect 271804 165476 272404 165478
rect 307804 165476 308404 165478
rect 343804 165476 344404 165478
rect 379804 165476 380404 165478
rect 415804 165476 416404 165478
rect 451804 165476 452404 165478
rect 487804 165476 488404 165478
rect 523804 165476 524404 165478
rect 559804 165476 560404 165478
rect 586260 165476 586860 165478
rect -2936 165454 586860 165476
rect -2936 165218 -2754 165454
rect -2518 165218 19986 165454
rect 20222 165218 55986 165454
rect 56222 165218 91986 165454
rect 92222 165218 127986 165454
rect 128222 165218 163986 165454
rect 164222 165218 199986 165454
rect 200222 165218 235986 165454
rect 236222 165218 271986 165454
rect 272222 165218 307986 165454
rect 308222 165218 343986 165454
rect 344222 165218 379986 165454
rect 380222 165218 415986 165454
rect 416222 165218 451986 165454
rect 452222 165218 487986 165454
rect 488222 165218 523986 165454
rect 524222 165218 559986 165454
rect 560222 165218 586442 165454
rect 586678 165218 586860 165454
rect -2936 165134 586860 165218
rect -2936 164898 -2754 165134
rect -2518 164898 19986 165134
rect 20222 164898 55986 165134
rect 56222 164898 91986 165134
rect 92222 164898 127986 165134
rect 128222 164898 163986 165134
rect 164222 164898 199986 165134
rect 200222 164898 235986 165134
rect 236222 164898 271986 165134
rect 272222 164898 307986 165134
rect 308222 164898 343986 165134
rect 344222 164898 379986 165134
rect 380222 164898 415986 165134
rect 416222 164898 451986 165134
rect 452222 164898 487986 165134
rect 488222 164898 523986 165134
rect 524222 164898 559986 165134
rect 560222 164898 586442 165134
rect 586678 164898 586860 165134
rect -2936 164876 586860 164898
rect -2936 164874 -2336 164876
rect 19804 164874 20404 164876
rect 55804 164874 56404 164876
rect 91804 164874 92404 164876
rect 127804 164874 128404 164876
rect 163804 164874 164404 164876
rect 199804 164874 200404 164876
rect 235804 164874 236404 164876
rect 271804 164874 272404 164876
rect 307804 164874 308404 164876
rect 343804 164874 344404 164876
rect 379804 164874 380404 164876
rect 415804 164874 416404 164876
rect 451804 164874 452404 164876
rect 487804 164874 488404 164876
rect 523804 164874 524404 164876
rect 559804 164874 560404 164876
rect 586260 164874 586860 164876
rect -7636 158276 -7036 158278
rect 12604 158276 13204 158278
rect 48604 158276 49204 158278
rect 84604 158276 85204 158278
rect 120604 158276 121204 158278
rect 156604 158276 157204 158278
rect 192604 158276 193204 158278
rect 228604 158276 229204 158278
rect 264604 158276 265204 158278
rect 300604 158276 301204 158278
rect 336604 158276 337204 158278
rect 372604 158276 373204 158278
rect 408604 158276 409204 158278
rect 444604 158276 445204 158278
rect 480604 158276 481204 158278
rect 516604 158276 517204 158278
rect 552604 158276 553204 158278
rect 590960 158276 591560 158278
rect -8576 158254 592500 158276
rect -8576 158018 -7454 158254
rect -7218 158018 12786 158254
rect 13022 158018 48786 158254
rect 49022 158018 84786 158254
rect 85022 158018 120786 158254
rect 121022 158018 156786 158254
rect 157022 158018 192786 158254
rect 193022 158018 228786 158254
rect 229022 158018 264786 158254
rect 265022 158018 300786 158254
rect 301022 158018 336786 158254
rect 337022 158018 372786 158254
rect 373022 158018 408786 158254
rect 409022 158018 444786 158254
rect 445022 158018 480786 158254
rect 481022 158018 516786 158254
rect 517022 158018 552786 158254
rect 553022 158018 591142 158254
rect 591378 158018 592500 158254
rect -8576 157934 592500 158018
rect -8576 157698 -7454 157934
rect -7218 157698 12786 157934
rect 13022 157698 48786 157934
rect 49022 157698 84786 157934
rect 85022 157698 120786 157934
rect 121022 157698 156786 157934
rect 157022 157698 192786 157934
rect 193022 157698 228786 157934
rect 229022 157698 264786 157934
rect 265022 157698 300786 157934
rect 301022 157698 336786 157934
rect 337022 157698 372786 157934
rect 373022 157698 408786 157934
rect 409022 157698 444786 157934
rect 445022 157698 480786 157934
rect 481022 157698 516786 157934
rect 517022 157698 552786 157934
rect 553022 157698 591142 157934
rect 591378 157698 592500 157934
rect -8576 157676 592500 157698
rect -7636 157674 -7036 157676
rect 12604 157674 13204 157676
rect 48604 157674 49204 157676
rect 84604 157674 85204 157676
rect 120604 157674 121204 157676
rect 156604 157674 157204 157676
rect 192604 157674 193204 157676
rect 228604 157674 229204 157676
rect 264604 157674 265204 157676
rect 300604 157674 301204 157676
rect 336604 157674 337204 157676
rect 372604 157674 373204 157676
rect 408604 157674 409204 157676
rect 444604 157674 445204 157676
rect 480604 157674 481204 157676
rect 516604 157674 517204 157676
rect 552604 157674 553204 157676
rect 590960 157674 591560 157676
rect -5756 154676 -5156 154678
rect 9004 154676 9604 154678
rect 45004 154676 45604 154678
rect 81004 154676 81604 154678
rect 117004 154676 117604 154678
rect 153004 154676 153604 154678
rect 189004 154676 189604 154678
rect 225004 154676 225604 154678
rect 261004 154676 261604 154678
rect 297004 154676 297604 154678
rect 333004 154676 333604 154678
rect 369004 154676 369604 154678
rect 405004 154676 405604 154678
rect 441004 154676 441604 154678
rect 477004 154676 477604 154678
rect 513004 154676 513604 154678
rect 549004 154676 549604 154678
rect 589080 154676 589680 154678
rect -6696 154654 590620 154676
rect -6696 154418 -5574 154654
rect -5338 154418 9186 154654
rect 9422 154418 45186 154654
rect 45422 154418 81186 154654
rect 81422 154418 117186 154654
rect 117422 154418 153186 154654
rect 153422 154418 189186 154654
rect 189422 154418 225186 154654
rect 225422 154418 261186 154654
rect 261422 154418 297186 154654
rect 297422 154418 333186 154654
rect 333422 154418 369186 154654
rect 369422 154418 405186 154654
rect 405422 154418 441186 154654
rect 441422 154418 477186 154654
rect 477422 154418 513186 154654
rect 513422 154418 549186 154654
rect 549422 154418 589262 154654
rect 589498 154418 590620 154654
rect -6696 154334 590620 154418
rect -6696 154098 -5574 154334
rect -5338 154098 9186 154334
rect 9422 154098 45186 154334
rect 45422 154098 81186 154334
rect 81422 154098 117186 154334
rect 117422 154098 153186 154334
rect 153422 154098 189186 154334
rect 189422 154098 225186 154334
rect 225422 154098 261186 154334
rect 261422 154098 297186 154334
rect 297422 154098 333186 154334
rect 333422 154098 369186 154334
rect 369422 154098 405186 154334
rect 405422 154098 441186 154334
rect 441422 154098 477186 154334
rect 477422 154098 513186 154334
rect 513422 154098 549186 154334
rect 549422 154098 589262 154334
rect 589498 154098 590620 154334
rect -6696 154076 590620 154098
rect -5756 154074 -5156 154076
rect 9004 154074 9604 154076
rect 45004 154074 45604 154076
rect 81004 154074 81604 154076
rect 117004 154074 117604 154076
rect 153004 154074 153604 154076
rect 189004 154074 189604 154076
rect 225004 154074 225604 154076
rect 261004 154074 261604 154076
rect 297004 154074 297604 154076
rect 333004 154074 333604 154076
rect 369004 154074 369604 154076
rect 405004 154074 405604 154076
rect 441004 154074 441604 154076
rect 477004 154074 477604 154076
rect 513004 154074 513604 154076
rect 549004 154074 549604 154076
rect 589080 154074 589680 154076
rect -3876 151076 -3276 151078
rect 5404 151076 6004 151078
rect 41404 151076 42004 151078
rect 77404 151076 78004 151078
rect 113404 151076 114004 151078
rect 149404 151076 150004 151078
rect 185404 151076 186004 151078
rect 221404 151076 222004 151078
rect 257404 151076 258004 151078
rect 293404 151076 294004 151078
rect 329404 151076 330004 151078
rect 365404 151076 366004 151078
rect 401404 151076 402004 151078
rect 437404 151076 438004 151078
rect 473404 151076 474004 151078
rect 509404 151076 510004 151078
rect 545404 151076 546004 151078
rect 581404 151076 582004 151078
rect 587200 151076 587800 151078
rect -4816 151054 588740 151076
rect -4816 150818 -3694 151054
rect -3458 150818 5586 151054
rect 5822 150818 41586 151054
rect 41822 150818 77586 151054
rect 77822 150818 113586 151054
rect 113822 150818 149586 151054
rect 149822 150818 185586 151054
rect 185822 150818 221586 151054
rect 221822 150818 257586 151054
rect 257822 150818 293586 151054
rect 293822 150818 329586 151054
rect 329822 150818 365586 151054
rect 365822 150818 401586 151054
rect 401822 150818 437586 151054
rect 437822 150818 473586 151054
rect 473822 150818 509586 151054
rect 509822 150818 545586 151054
rect 545822 150818 581586 151054
rect 581822 150818 587382 151054
rect 587618 150818 588740 151054
rect -4816 150734 588740 150818
rect -4816 150498 -3694 150734
rect -3458 150498 5586 150734
rect 5822 150498 41586 150734
rect 41822 150498 77586 150734
rect 77822 150498 113586 150734
rect 113822 150498 149586 150734
rect 149822 150498 185586 150734
rect 185822 150498 221586 150734
rect 221822 150498 257586 150734
rect 257822 150498 293586 150734
rect 293822 150498 329586 150734
rect 329822 150498 365586 150734
rect 365822 150498 401586 150734
rect 401822 150498 437586 150734
rect 437822 150498 473586 150734
rect 473822 150498 509586 150734
rect 509822 150498 545586 150734
rect 545822 150498 581586 150734
rect 581822 150498 587382 150734
rect 587618 150498 588740 150734
rect -4816 150476 588740 150498
rect -3876 150474 -3276 150476
rect 5404 150474 6004 150476
rect 41404 150474 42004 150476
rect 77404 150474 78004 150476
rect 113404 150474 114004 150476
rect 149404 150474 150004 150476
rect 185404 150474 186004 150476
rect 221404 150474 222004 150476
rect 257404 150474 258004 150476
rect 293404 150474 294004 150476
rect 329404 150474 330004 150476
rect 365404 150474 366004 150476
rect 401404 150474 402004 150476
rect 437404 150474 438004 150476
rect 473404 150474 474004 150476
rect 509404 150474 510004 150476
rect 545404 150474 546004 150476
rect 581404 150474 582004 150476
rect 587200 150474 587800 150476
rect -1996 147476 -1396 147478
rect 1804 147476 2404 147478
rect 37804 147476 38404 147478
rect 73804 147476 74404 147478
rect 109804 147476 110404 147478
rect 145804 147476 146404 147478
rect 181804 147476 182404 147478
rect 217804 147476 218404 147478
rect 253804 147476 254404 147478
rect 289804 147476 290404 147478
rect 325804 147476 326404 147478
rect 361804 147476 362404 147478
rect 397804 147476 398404 147478
rect 433804 147476 434404 147478
rect 469804 147476 470404 147478
rect 505804 147476 506404 147478
rect 541804 147476 542404 147478
rect 577804 147476 578404 147478
rect 585320 147476 585920 147478
rect -2936 147454 586860 147476
rect -2936 147218 -1814 147454
rect -1578 147218 1986 147454
rect 2222 147218 37986 147454
rect 38222 147218 73986 147454
rect 74222 147218 109986 147454
rect 110222 147218 145986 147454
rect 146222 147218 181986 147454
rect 182222 147218 217986 147454
rect 218222 147218 253986 147454
rect 254222 147218 289986 147454
rect 290222 147218 325986 147454
rect 326222 147218 361986 147454
rect 362222 147218 397986 147454
rect 398222 147218 433986 147454
rect 434222 147218 469986 147454
rect 470222 147218 505986 147454
rect 506222 147218 541986 147454
rect 542222 147218 577986 147454
rect 578222 147218 585502 147454
rect 585738 147218 586860 147454
rect -2936 147134 586860 147218
rect -2936 146898 -1814 147134
rect -1578 146898 1986 147134
rect 2222 146898 37986 147134
rect 38222 146898 73986 147134
rect 74222 146898 109986 147134
rect 110222 146898 145986 147134
rect 146222 146898 181986 147134
rect 182222 146898 217986 147134
rect 218222 146898 253986 147134
rect 254222 146898 289986 147134
rect 290222 146898 325986 147134
rect 326222 146898 361986 147134
rect 362222 146898 397986 147134
rect 398222 146898 433986 147134
rect 434222 146898 469986 147134
rect 470222 146898 505986 147134
rect 506222 146898 541986 147134
rect 542222 146898 577986 147134
rect 578222 146898 585502 147134
rect 585738 146898 586860 147134
rect -2936 146876 586860 146898
rect -1996 146874 -1396 146876
rect 1804 146874 2404 146876
rect 37804 146874 38404 146876
rect 73804 146874 74404 146876
rect 109804 146874 110404 146876
rect 145804 146874 146404 146876
rect 181804 146874 182404 146876
rect 217804 146874 218404 146876
rect 253804 146874 254404 146876
rect 289804 146874 290404 146876
rect 325804 146874 326404 146876
rect 361804 146874 362404 146876
rect 397804 146874 398404 146876
rect 433804 146874 434404 146876
rect 469804 146874 470404 146876
rect 505804 146874 506404 146876
rect 541804 146874 542404 146876
rect 577804 146874 578404 146876
rect 585320 146874 585920 146876
rect -8576 140276 -7976 140278
rect 30604 140276 31204 140278
rect 66604 140276 67204 140278
rect 102604 140276 103204 140278
rect 138604 140276 139204 140278
rect 174604 140276 175204 140278
rect 210604 140276 211204 140278
rect 246604 140276 247204 140278
rect 282604 140276 283204 140278
rect 318604 140276 319204 140278
rect 354604 140276 355204 140278
rect 390604 140276 391204 140278
rect 426604 140276 427204 140278
rect 462604 140276 463204 140278
rect 498604 140276 499204 140278
rect 534604 140276 535204 140278
rect 570604 140276 571204 140278
rect 591900 140276 592500 140278
rect -8576 140254 592500 140276
rect -8576 140018 -8394 140254
rect -8158 140018 30786 140254
rect 31022 140018 66786 140254
rect 67022 140018 102786 140254
rect 103022 140018 138786 140254
rect 139022 140018 174786 140254
rect 175022 140018 210786 140254
rect 211022 140018 246786 140254
rect 247022 140018 282786 140254
rect 283022 140018 318786 140254
rect 319022 140018 354786 140254
rect 355022 140018 390786 140254
rect 391022 140018 426786 140254
rect 427022 140018 462786 140254
rect 463022 140018 498786 140254
rect 499022 140018 534786 140254
rect 535022 140018 570786 140254
rect 571022 140018 592082 140254
rect 592318 140018 592500 140254
rect -8576 139934 592500 140018
rect -8576 139698 -8394 139934
rect -8158 139698 30786 139934
rect 31022 139698 66786 139934
rect 67022 139698 102786 139934
rect 103022 139698 138786 139934
rect 139022 139698 174786 139934
rect 175022 139698 210786 139934
rect 211022 139698 246786 139934
rect 247022 139698 282786 139934
rect 283022 139698 318786 139934
rect 319022 139698 354786 139934
rect 355022 139698 390786 139934
rect 391022 139698 426786 139934
rect 427022 139698 462786 139934
rect 463022 139698 498786 139934
rect 499022 139698 534786 139934
rect 535022 139698 570786 139934
rect 571022 139698 592082 139934
rect 592318 139698 592500 139934
rect -8576 139676 592500 139698
rect -8576 139674 -7976 139676
rect 30604 139674 31204 139676
rect 66604 139674 67204 139676
rect 102604 139674 103204 139676
rect 138604 139674 139204 139676
rect 174604 139674 175204 139676
rect 210604 139674 211204 139676
rect 246604 139674 247204 139676
rect 282604 139674 283204 139676
rect 318604 139674 319204 139676
rect 354604 139674 355204 139676
rect 390604 139674 391204 139676
rect 426604 139674 427204 139676
rect 462604 139674 463204 139676
rect 498604 139674 499204 139676
rect 534604 139674 535204 139676
rect 570604 139674 571204 139676
rect 591900 139674 592500 139676
rect -6696 136676 -6096 136678
rect 27004 136676 27604 136678
rect 63004 136676 63604 136678
rect 99004 136676 99604 136678
rect 135004 136676 135604 136678
rect 171004 136676 171604 136678
rect 207004 136676 207604 136678
rect 243004 136676 243604 136678
rect 279004 136676 279604 136678
rect 315004 136676 315604 136678
rect 351004 136676 351604 136678
rect 387004 136676 387604 136678
rect 423004 136676 423604 136678
rect 459004 136676 459604 136678
rect 495004 136676 495604 136678
rect 531004 136676 531604 136678
rect 567004 136676 567604 136678
rect 590020 136676 590620 136678
rect -6696 136654 590620 136676
rect -6696 136418 -6514 136654
rect -6278 136418 27186 136654
rect 27422 136418 63186 136654
rect 63422 136418 99186 136654
rect 99422 136418 135186 136654
rect 135422 136418 171186 136654
rect 171422 136418 207186 136654
rect 207422 136418 243186 136654
rect 243422 136418 279186 136654
rect 279422 136418 315186 136654
rect 315422 136418 351186 136654
rect 351422 136418 387186 136654
rect 387422 136418 423186 136654
rect 423422 136418 459186 136654
rect 459422 136418 495186 136654
rect 495422 136418 531186 136654
rect 531422 136418 567186 136654
rect 567422 136418 590202 136654
rect 590438 136418 590620 136654
rect -6696 136334 590620 136418
rect -6696 136098 -6514 136334
rect -6278 136098 27186 136334
rect 27422 136098 63186 136334
rect 63422 136098 99186 136334
rect 99422 136098 135186 136334
rect 135422 136098 171186 136334
rect 171422 136098 207186 136334
rect 207422 136098 243186 136334
rect 243422 136098 279186 136334
rect 279422 136098 315186 136334
rect 315422 136098 351186 136334
rect 351422 136098 387186 136334
rect 387422 136098 423186 136334
rect 423422 136098 459186 136334
rect 459422 136098 495186 136334
rect 495422 136098 531186 136334
rect 531422 136098 567186 136334
rect 567422 136098 590202 136334
rect 590438 136098 590620 136334
rect -6696 136076 590620 136098
rect -6696 136074 -6096 136076
rect 27004 136074 27604 136076
rect 63004 136074 63604 136076
rect 99004 136074 99604 136076
rect 135004 136074 135604 136076
rect 171004 136074 171604 136076
rect 207004 136074 207604 136076
rect 243004 136074 243604 136076
rect 279004 136074 279604 136076
rect 315004 136074 315604 136076
rect 351004 136074 351604 136076
rect 387004 136074 387604 136076
rect 423004 136074 423604 136076
rect 459004 136074 459604 136076
rect 495004 136074 495604 136076
rect 531004 136074 531604 136076
rect 567004 136074 567604 136076
rect 590020 136074 590620 136076
rect -4816 133076 -4216 133078
rect 23404 133076 24004 133078
rect 59404 133076 60004 133078
rect 95404 133076 96004 133078
rect 131404 133076 132004 133078
rect 167404 133076 168004 133078
rect 203404 133076 204004 133078
rect 239404 133076 240004 133078
rect 275404 133076 276004 133078
rect 311404 133076 312004 133078
rect 347404 133076 348004 133078
rect 383404 133076 384004 133078
rect 419404 133076 420004 133078
rect 455404 133076 456004 133078
rect 491404 133076 492004 133078
rect 527404 133076 528004 133078
rect 563404 133076 564004 133078
rect 588140 133076 588740 133078
rect -4816 133054 588740 133076
rect -4816 132818 -4634 133054
rect -4398 132818 23586 133054
rect 23822 132818 59586 133054
rect 59822 132818 95586 133054
rect 95822 132818 131586 133054
rect 131822 132818 167586 133054
rect 167822 132818 203586 133054
rect 203822 132818 239586 133054
rect 239822 132818 275586 133054
rect 275822 132818 311586 133054
rect 311822 132818 347586 133054
rect 347822 132818 383586 133054
rect 383822 132818 419586 133054
rect 419822 132818 455586 133054
rect 455822 132818 491586 133054
rect 491822 132818 527586 133054
rect 527822 132818 563586 133054
rect 563822 132818 588322 133054
rect 588558 132818 588740 133054
rect -4816 132734 588740 132818
rect -4816 132498 -4634 132734
rect -4398 132498 23586 132734
rect 23822 132498 59586 132734
rect 59822 132498 95586 132734
rect 95822 132498 131586 132734
rect 131822 132498 167586 132734
rect 167822 132498 203586 132734
rect 203822 132498 239586 132734
rect 239822 132498 275586 132734
rect 275822 132498 311586 132734
rect 311822 132498 347586 132734
rect 347822 132498 383586 132734
rect 383822 132498 419586 132734
rect 419822 132498 455586 132734
rect 455822 132498 491586 132734
rect 491822 132498 527586 132734
rect 527822 132498 563586 132734
rect 563822 132498 588322 132734
rect 588558 132498 588740 132734
rect -4816 132476 588740 132498
rect -4816 132474 -4216 132476
rect 23404 132474 24004 132476
rect 59404 132474 60004 132476
rect 95404 132474 96004 132476
rect 131404 132474 132004 132476
rect 167404 132474 168004 132476
rect 203404 132474 204004 132476
rect 239404 132474 240004 132476
rect 275404 132474 276004 132476
rect 311404 132474 312004 132476
rect 347404 132474 348004 132476
rect 383404 132474 384004 132476
rect 419404 132474 420004 132476
rect 455404 132474 456004 132476
rect 491404 132474 492004 132476
rect 527404 132474 528004 132476
rect 563404 132474 564004 132476
rect 588140 132474 588740 132476
rect -2936 129476 -2336 129478
rect 19804 129476 20404 129478
rect 55804 129476 56404 129478
rect 91804 129476 92404 129478
rect 127804 129476 128404 129478
rect 163804 129476 164404 129478
rect 199804 129476 200404 129478
rect 235804 129476 236404 129478
rect 271804 129476 272404 129478
rect 307804 129476 308404 129478
rect 343804 129476 344404 129478
rect 379804 129476 380404 129478
rect 415804 129476 416404 129478
rect 451804 129476 452404 129478
rect 487804 129476 488404 129478
rect 523804 129476 524404 129478
rect 559804 129476 560404 129478
rect 586260 129476 586860 129478
rect -2936 129454 586860 129476
rect -2936 129218 -2754 129454
rect -2518 129218 19986 129454
rect 20222 129218 55986 129454
rect 56222 129218 91986 129454
rect 92222 129218 127986 129454
rect 128222 129218 163986 129454
rect 164222 129218 199986 129454
rect 200222 129218 235986 129454
rect 236222 129218 271986 129454
rect 272222 129218 307986 129454
rect 308222 129218 343986 129454
rect 344222 129218 379986 129454
rect 380222 129218 415986 129454
rect 416222 129218 451986 129454
rect 452222 129218 487986 129454
rect 488222 129218 523986 129454
rect 524222 129218 559986 129454
rect 560222 129218 586442 129454
rect 586678 129218 586860 129454
rect -2936 129134 586860 129218
rect -2936 128898 -2754 129134
rect -2518 128898 19986 129134
rect 20222 128898 55986 129134
rect 56222 128898 91986 129134
rect 92222 128898 127986 129134
rect 128222 128898 163986 129134
rect 164222 128898 199986 129134
rect 200222 128898 235986 129134
rect 236222 128898 271986 129134
rect 272222 128898 307986 129134
rect 308222 128898 343986 129134
rect 344222 128898 379986 129134
rect 380222 128898 415986 129134
rect 416222 128898 451986 129134
rect 452222 128898 487986 129134
rect 488222 128898 523986 129134
rect 524222 128898 559986 129134
rect 560222 128898 586442 129134
rect 586678 128898 586860 129134
rect -2936 128876 586860 128898
rect -2936 128874 -2336 128876
rect 19804 128874 20404 128876
rect 55804 128874 56404 128876
rect 91804 128874 92404 128876
rect 127804 128874 128404 128876
rect 163804 128874 164404 128876
rect 199804 128874 200404 128876
rect 235804 128874 236404 128876
rect 271804 128874 272404 128876
rect 307804 128874 308404 128876
rect 343804 128874 344404 128876
rect 379804 128874 380404 128876
rect 415804 128874 416404 128876
rect 451804 128874 452404 128876
rect 487804 128874 488404 128876
rect 523804 128874 524404 128876
rect 559804 128874 560404 128876
rect 586260 128874 586860 128876
rect -7636 122276 -7036 122278
rect 12604 122276 13204 122278
rect 48604 122276 49204 122278
rect 84604 122276 85204 122278
rect 120604 122276 121204 122278
rect 156604 122276 157204 122278
rect 192604 122276 193204 122278
rect 228604 122276 229204 122278
rect 264604 122276 265204 122278
rect 300604 122276 301204 122278
rect 336604 122276 337204 122278
rect 372604 122276 373204 122278
rect 408604 122276 409204 122278
rect 444604 122276 445204 122278
rect 480604 122276 481204 122278
rect 516604 122276 517204 122278
rect 552604 122276 553204 122278
rect 590960 122276 591560 122278
rect -8576 122254 592500 122276
rect -8576 122018 -7454 122254
rect -7218 122018 12786 122254
rect 13022 122018 48786 122254
rect 49022 122018 84786 122254
rect 85022 122018 120786 122254
rect 121022 122018 156786 122254
rect 157022 122018 192786 122254
rect 193022 122018 228786 122254
rect 229022 122018 264786 122254
rect 265022 122018 300786 122254
rect 301022 122018 336786 122254
rect 337022 122018 372786 122254
rect 373022 122018 408786 122254
rect 409022 122018 444786 122254
rect 445022 122018 480786 122254
rect 481022 122018 516786 122254
rect 517022 122018 552786 122254
rect 553022 122018 591142 122254
rect 591378 122018 592500 122254
rect -8576 121934 592500 122018
rect -8576 121698 -7454 121934
rect -7218 121698 12786 121934
rect 13022 121698 48786 121934
rect 49022 121698 84786 121934
rect 85022 121698 120786 121934
rect 121022 121698 156786 121934
rect 157022 121698 192786 121934
rect 193022 121698 228786 121934
rect 229022 121698 264786 121934
rect 265022 121698 300786 121934
rect 301022 121698 336786 121934
rect 337022 121698 372786 121934
rect 373022 121698 408786 121934
rect 409022 121698 444786 121934
rect 445022 121698 480786 121934
rect 481022 121698 516786 121934
rect 517022 121698 552786 121934
rect 553022 121698 591142 121934
rect 591378 121698 592500 121934
rect -8576 121676 592500 121698
rect -7636 121674 -7036 121676
rect 12604 121674 13204 121676
rect 48604 121674 49204 121676
rect 84604 121674 85204 121676
rect 120604 121674 121204 121676
rect 156604 121674 157204 121676
rect 192604 121674 193204 121676
rect 228604 121674 229204 121676
rect 264604 121674 265204 121676
rect 300604 121674 301204 121676
rect 336604 121674 337204 121676
rect 372604 121674 373204 121676
rect 408604 121674 409204 121676
rect 444604 121674 445204 121676
rect 480604 121674 481204 121676
rect 516604 121674 517204 121676
rect 552604 121674 553204 121676
rect 590960 121674 591560 121676
rect -5756 118676 -5156 118678
rect 9004 118676 9604 118678
rect 45004 118676 45604 118678
rect 81004 118676 81604 118678
rect 117004 118676 117604 118678
rect 153004 118676 153604 118678
rect 189004 118676 189604 118678
rect 225004 118676 225604 118678
rect 261004 118676 261604 118678
rect 297004 118676 297604 118678
rect 333004 118676 333604 118678
rect 369004 118676 369604 118678
rect 405004 118676 405604 118678
rect 441004 118676 441604 118678
rect 477004 118676 477604 118678
rect 513004 118676 513604 118678
rect 549004 118676 549604 118678
rect 589080 118676 589680 118678
rect -6696 118654 590620 118676
rect -6696 118418 -5574 118654
rect -5338 118418 9186 118654
rect 9422 118418 45186 118654
rect 45422 118418 81186 118654
rect 81422 118418 117186 118654
rect 117422 118418 153186 118654
rect 153422 118418 189186 118654
rect 189422 118418 225186 118654
rect 225422 118418 261186 118654
rect 261422 118418 297186 118654
rect 297422 118418 333186 118654
rect 333422 118418 369186 118654
rect 369422 118418 405186 118654
rect 405422 118418 441186 118654
rect 441422 118418 477186 118654
rect 477422 118418 513186 118654
rect 513422 118418 549186 118654
rect 549422 118418 589262 118654
rect 589498 118418 590620 118654
rect -6696 118334 590620 118418
rect -6696 118098 -5574 118334
rect -5338 118098 9186 118334
rect 9422 118098 45186 118334
rect 45422 118098 81186 118334
rect 81422 118098 117186 118334
rect 117422 118098 153186 118334
rect 153422 118098 189186 118334
rect 189422 118098 225186 118334
rect 225422 118098 261186 118334
rect 261422 118098 297186 118334
rect 297422 118098 333186 118334
rect 333422 118098 369186 118334
rect 369422 118098 405186 118334
rect 405422 118098 441186 118334
rect 441422 118098 477186 118334
rect 477422 118098 513186 118334
rect 513422 118098 549186 118334
rect 549422 118098 589262 118334
rect 589498 118098 590620 118334
rect -6696 118076 590620 118098
rect -5756 118074 -5156 118076
rect 9004 118074 9604 118076
rect 45004 118074 45604 118076
rect 81004 118074 81604 118076
rect 117004 118074 117604 118076
rect 153004 118074 153604 118076
rect 189004 118074 189604 118076
rect 225004 118074 225604 118076
rect 261004 118074 261604 118076
rect 297004 118074 297604 118076
rect 333004 118074 333604 118076
rect 369004 118074 369604 118076
rect 405004 118074 405604 118076
rect 441004 118074 441604 118076
rect 477004 118074 477604 118076
rect 513004 118074 513604 118076
rect 549004 118074 549604 118076
rect 589080 118074 589680 118076
rect -3876 115076 -3276 115078
rect 5404 115076 6004 115078
rect 41404 115076 42004 115078
rect 77404 115076 78004 115078
rect 113404 115076 114004 115078
rect 149404 115076 150004 115078
rect 185404 115076 186004 115078
rect 221404 115076 222004 115078
rect 257404 115076 258004 115078
rect 293404 115076 294004 115078
rect 329404 115076 330004 115078
rect 365404 115076 366004 115078
rect 401404 115076 402004 115078
rect 437404 115076 438004 115078
rect 473404 115076 474004 115078
rect 509404 115076 510004 115078
rect 545404 115076 546004 115078
rect 581404 115076 582004 115078
rect 587200 115076 587800 115078
rect -4816 115054 588740 115076
rect -4816 114818 -3694 115054
rect -3458 114818 5586 115054
rect 5822 114818 41586 115054
rect 41822 114818 77586 115054
rect 77822 114818 113586 115054
rect 113822 114818 149586 115054
rect 149822 114818 185586 115054
rect 185822 114818 221586 115054
rect 221822 114818 257586 115054
rect 257822 114818 293586 115054
rect 293822 114818 329586 115054
rect 329822 114818 365586 115054
rect 365822 114818 401586 115054
rect 401822 114818 437586 115054
rect 437822 114818 473586 115054
rect 473822 114818 509586 115054
rect 509822 114818 545586 115054
rect 545822 114818 581586 115054
rect 581822 114818 587382 115054
rect 587618 114818 588740 115054
rect -4816 114734 588740 114818
rect -4816 114498 -3694 114734
rect -3458 114498 5586 114734
rect 5822 114498 41586 114734
rect 41822 114498 77586 114734
rect 77822 114498 113586 114734
rect 113822 114498 149586 114734
rect 149822 114498 185586 114734
rect 185822 114498 221586 114734
rect 221822 114498 257586 114734
rect 257822 114498 293586 114734
rect 293822 114498 329586 114734
rect 329822 114498 365586 114734
rect 365822 114498 401586 114734
rect 401822 114498 437586 114734
rect 437822 114498 473586 114734
rect 473822 114498 509586 114734
rect 509822 114498 545586 114734
rect 545822 114498 581586 114734
rect 581822 114498 587382 114734
rect 587618 114498 588740 114734
rect -4816 114476 588740 114498
rect -3876 114474 -3276 114476
rect 5404 114474 6004 114476
rect 41404 114474 42004 114476
rect 77404 114474 78004 114476
rect 113404 114474 114004 114476
rect 149404 114474 150004 114476
rect 185404 114474 186004 114476
rect 221404 114474 222004 114476
rect 257404 114474 258004 114476
rect 293404 114474 294004 114476
rect 329404 114474 330004 114476
rect 365404 114474 366004 114476
rect 401404 114474 402004 114476
rect 437404 114474 438004 114476
rect 473404 114474 474004 114476
rect 509404 114474 510004 114476
rect 545404 114474 546004 114476
rect 581404 114474 582004 114476
rect 587200 114474 587800 114476
rect -1996 111476 -1396 111478
rect 1804 111476 2404 111478
rect 37804 111476 38404 111478
rect 73804 111476 74404 111478
rect 109804 111476 110404 111478
rect 145804 111476 146404 111478
rect 181804 111476 182404 111478
rect 217804 111476 218404 111478
rect 253804 111476 254404 111478
rect 289804 111476 290404 111478
rect 325804 111476 326404 111478
rect 361804 111476 362404 111478
rect 397804 111476 398404 111478
rect 433804 111476 434404 111478
rect 469804 111476 470404 111478
rect 505804 111476 506404 111478
rect 541804 111476 542404 111478
rect 577804 111476 578404 111478
rect 585320 111476 585920 111478
rect -2936 111454 586860 111476
rect -2936 111218 -1814 111454
rect -1578 111218 1986 111454
rect 2222 111218 37986 111454
rect 38222 111218 73986 111454
rect 74222 111218 109986 111454
rect 110222 111218 145986 111454
rect 146222 111218 181986 111454
rect 182222 111218 217986 111454
rect 218222 111218 253986 111454
rect 254222 111218 289986 111454
rect 290222 111218 325986 111454
rect 326222 111218 361986 111454
rect 362222 111218 397986 111454
rect 398222 111218 433986 111454
rect 434222 111218 469986 111454
rect 470222 111218 505986 111454
rect 506222 111218 541986 111454
rect 542222 111218 577986 111454
rect 578222 111218 585502 111454
rect 585738 111218 586860 111454
rect -2936 111134 586860 111218
rect -2936 110898 -1814 111134
rect -1578 110898 1986 111134
rect 2222 110898 37986 111134
rect 38222 110898 73986 111134
rect 74222 110898 109986 111134
rect 110222 110898 145986 111134
rect 146222 110898 181986 111134
rect 182222 110898 217986 111134
rect 218222 110898 253986 111134
rect 254222 110898 289986 111134
rect 290222 110898 325986 111134
rect 326222 110898 361986 111134
rect 362222 110898 397986 111134
rect 398222 110898 433986 111134
rect 434222 110898 469986 111134
rect 470222 110898 505986 111134
rect 506222 110898 541986 111134
rect 542222 110898 577986 111134
rect 578222 110898 585502 111134
rect 585738 110898 586860 111134
rect -2936 110876 586860 110898
rect -1996 110874 -1396 110876
rect 1804 110874 2404 110876
rect 37804 110874 38404 110876
rect 73804 110874 74404 110876
rect 109804 110874 110404 110876
rect 145804 110874 146404 110876
rect 181804 110874 182404 110876
rect 217804 110874 218404 110876
rect 253804 110874 254404 110876
rect 289804 110874 290404 110876
rect 325804 110874 326404 110876
rect 361804 110874 362404 110876
rect 397804 110874 398404 110876
rect 433804 110874 434404 110876
rect 469804 110874 470404 110876
rect 505804 110874 506404 110876
rect 541804 110874 542404 110876
rect 577804 110874 578404 110876
rect 585320 110874 585920 110876
rect -8576 104276 -7976 104278
rect 30604 104276 31204 104278
rect 66604 104276 67204 104278
rect 102604 104276 103204 104278
rect 138604 104276 139204 104278
rect 174604 104276 175204 104278
rect 210604 104276 211204 104278
rect 246604 104276 247204 104278
rect 282604 104276 283204 104278
rect 318604 104276 319204 104278
rect 354604 104276 355204 104278
rect 390604 104276 391204 104278
rect 426604 104276 427204 104278
rect 462604 104276 463204 104278
rect 498604 104276 499204 104278
rect 534604 104276 535204 104278
rect 570604 104276 571204 104278
rect 591900 104276 592500 104278
rect -8576 104254 592500 104276
rect -8576 104018 -8394 104254
rect -8158 104018 30786 104254
rect 31022 104018 66786 104254
rect 67022 104018 102786 104254
rect 103022 104018 138786 104254
rect 139022 104018 174786 104254
rect 175022 104018 210786 104254
rect 211022 104018 246786 104254
rect 247022 104018 282786 104254
rect 283022 104018 318786 104254
rect 319022 104018 354786 104254
rect 355022 104018 390786 104254
rect 391022 104018 426786 104254
rect 427022 104018 462786 104254
rect 463022 104018 498786 104254
rect 499022 104018 534786 104254
rect 535022 104018 570786 104254
rect 571022 104018 592082 104254
rect 592318 104018 592500 104254
rect -8576 103934 592500 104018
rect -8576 103698 -8394 103934
rect -8158 103698 30786 103934
rect 31022 103698 66786 103934
rect 67022 103698 102786 103934
rect 103022 103698 138786 103934
rect 139022 103698 174786 103934
rect 175022 103698 210786 103934
rect 211022 103698 246786 103934
rect 247022 103698 282786 103934
rect 283022 103698 318786 103934
rect 319022 103698 354786 103934
rect 355022 103698 390786 103934
rect 391022 103698 426786 103934
rect 427022 103698 462786 103934
rect 463022 103698 498786 103934
rect 499022 103698 534786 103934
rect 535022 103698 570786 103934
rect 571022 103698 592082 103934
rect 592318 103698 592500 103934
rect -8576 103676 592500 103698
rect -8576 103674 -7976 103676
rect 30604 103674 31204 103676
rect 66604 103674 67204 103676
rect 102604 103674 103204 103676
rect 138604 103674 139204 103676
rect 174604 103674 175204 103676
rect 210604 103674 211204 103676
rect 246604 103674 247204 103676
rect 282604 103674 283204 103676
rect 318604 103674 319204 103676
rect 354604 103674 355204 103676
rect 390604 103674 391204 103676
rect 426604 103674 427204 103676
rect 462604 103674 463204 103676
rect 498604 103674 499204 103676
rect 534604 103674 535204 103676
rect 570604 103674 571204 103676
rect 591900 103674 592500 103676
rect -6696 100676 -6096 100678
rect 27004 100676 27604 100678
rect 63004 100676 63604 100678
rect 99004 100676 99604 100678
rect 135004 100676 135604 100678
rect 171004 100676 171604 100678
rect 207004 100676 207604 100678
rect 243004 100676 243604 100678
rect 279004 100676 279604 100678
rect 315004 100676 315604 100678
rect 351004 100676 351604 100678
rect 387004 100676 387604 100678
rect 423004 100676 423604 100678
rect 459004 100676 459604 100678
rect 495004 100676 495604 100678
rect 531004 100676 531604 100678
rect 567004 100676 567604 100678
rect 590020 100676 590620 100678
rect -6696 100654 590620 100676
rect -6696 100418 -6514 100654
rect -6278 100418 27186 100654
rect 27422 100418 63186 100654
rect 63422 100418 99186 100654
rect 99422 100418 135186 100654
rect 135422 100418 171186 100654
rect 171422 100418 207186 100654
rect 207422 100418 243186 100654
rect 243422 100418 279186 100654
rect 279422 100418 315186 100654
rect 315422 100418 351186 100654
rect 351422 100418 387186 100654
rect 387422 100418 423186 100654
rect 423422 100418 459186 100654
rect 459422 100418 495186 100654
rect 495422 100418 531186 100654
rect 531422 100418 567186 100654
rect 567422 100418 590202 100654
rect 590438 100418 590620 100654
rect -6696 100334 590620 100418
rect -6696 100098 -6514 100334
rect -6278 100098 27186 100334
rect 27422 100098 63186 100334
rect 63422 100098 99186 100334
rect 99422 100098 135186 100334
rect 135422 100098 171186 100334
rect 171422 100098 207186 100334
rect 207422 100098 243186 100334
rect 243422 100098 279186 100334
rect 279422 100098 315186 100334
rect 315422 100098 351186 100334
rect 351422 100098 387186 100334
rect 387422 100098 423186 100334
rect 423422 100098 459186 100334
rect 459422 100098 495186 100334
rect 495422 100098 531186 100334
rect 531422 100098 567186 100334
rect 567422 100098 590202 100334
rect 590438 100098 590620 100334
rect -6696 100076 590620 100098
rect -6696 100074 -6096 100076
rect 27004 100074 27604 100076
rect 63004 100074 63604 100076
rect 99004 100074 99604 100076
rect 135004 100074 135604 100076
rect 171004 100074 171604 100076
rect 207004 100074 207604 100076
rect 243004 100074 243604 100076
rect 279004 100074 279604 100076
rect 315004 100074 315604 100076
rect 351004 100074 351604 100076
rect 387004 100074 387604 100076
rect 423004 100074 423604 100076
rect 459004 100074 459604 100076
rect 495004 100074 495604 100076
rect 531004 100074 531604 100076
rect 567004 100074 567604 100076
rect 590020 100074 590620 100076
rect -4816 97076 -4216 97078
rect 23404 97076 24004 97078
rect 59404 97076 60004 97078
rect 95404 97076 96004 97078
rect 131404 97076 132004 97078
rect 167404 97076 168004 97078
rect 203404 97076 204004 97078
rect 239404 97076 240004 97078
rect 275404 97076 276004 97078
rect 311404 97076 312004 97078
rect 347404 97076 348004 97078
rect 383404 97076 384004 97078
rect 419404 97076 420004 97078
rect 455404 97076 456004 97078
rect 491404 97076 492004 97078
rect 527404 97076 528004 97078
rect 563404 97076 564004 97078
rect 588140 97076 588740 97078
rect -4816 97054 588740 97076
rect -4816 96818 -4634 97054
rect -4398 96818 23586 97054
rect 23822 96818 59586 97054
rect 59822 96818 95586 97054
rect 95822 96818 131586 97054
rect 131822 96818 167586 97054
rect 167822 96818 203586 97054
rect 203822 96818 239586 97054
rect 239822 96818 275586 97054
rect 275822 96818 311586 97054
rect 311822 96818 347586 97054
rect 347822 96818 383586 97054
rect 383822 96818 419586 97054
rect 419822 96818 455586 97054
rect 455822 96818 491586 97054
rect 491822 96818 527586 97054
rect 527822 96818 563586 97054
rect 563822 96818 588322 97054
rect 588558 96818 588740 97054
rect -4816 96734 588740 96818
rect -4816 96498 -4634 96734
rect -4398 96498 23586 96734
rect 23822 96498 59586 96734
rect 59822 96498 95586 96734
rect 95822 96498 131586 96734
rect 131822 96498 167586 96734
rect 167822 96498 203586 96734
rect 203822 96498 239586 96734
rect 239822 96498 275586 96734
rect 275822 96498 311586 96734
rect 311822 96498 347586 96734
rect 347822 96498 383586 96734
rect 383822 96498 419586 96734
rect 419822 96498 455586 96734
rect 455822 96498 491586 96734
rect 491822 96498 527586 96734
rect 527822 96498 563586 96734
rect 563822 96498 588322 96734
rect 588558 96498 588740 96734
rect -4816 96476 588740 96498
rect -4816 96474 -4216 96476
rect 23404 96474 24004 96476
rect 59404 96474 60004 96476
rect 95404 96474 96004 96476
rect 131404 96474 132004 96476
rect 167404 96474 168004 96476
rect 203404 96474 204004 96476
rect 239404 96474 240004 96476
rect 275404 96474 276004 96476
rect 311404 96474 312004 96476
rect 347404 96474 348004 96476
rect 383404 96474 384004 96476
rect 419404 96474 420004 96476
rect 455404 96474 456004 96476
rect 491404 96474 492004 96476
rect 527404 96474 528004 96476
rect 563404 96474 564004 96476
rect 588140 96474 588740 96476
rect -2936 93476 -2336 93478
rect 19804 93476 20404 93478
rect 55804 93476 56404 93478
rect 91804 93476 92404 93478
rect 127804 93476 128404 93478
rect 163804 93476 164404 93478
rect 199804 93476 200404 93478
rect 235804 93476 236404 93478
rect 271804 93476 272404 93478
rect 307804 93476 308404 93478
rect 343804 93476 344404 93478
rect 379804 93476 380404 93478
rect 415804 93476 416404 93478
rect 451804 93476 452404 93478
rect 487804 93476 488404 93478
rect 523804 93476 524404 93478
rect 559804 93476 560404 93478
rect 586260 93476 586860 93478
rect -2936 93454 586860 93476
rect -2936 93218 -2754 93454
rect -2518 93218 19986 93454
rect 20222 93218 55986 93454
rect 56222 93218 91986 93454
rect 92222 93218 127986 93454
rect 128222 93218 163986 93454
rect 164222 93218 199986 93454
rect 200222 93218 235986 93454
rect 236222 93218 271986 93454
rect 272222 93218 307986 93454
rect 308222 93218 343986 93454
rect 344222 93218 379986 93454
rect 380222 93218 415986 93454
rect 416222 93218 451986 93454
rect 452222 93218 487986 93454
rect 488222 93218 523986 93454
rect 524222 93218 559986 93454
rect 560222 93218 586442 93454
rect 586678 93218 586860 93454
rect -2936 93134 586860 93218
rect -2936 92898 -2754 93134
rect -2518 92898 19986 93134
rect 20222 92898 55986 93134
rect 56222 92898 91986 93134
rect 92222 92898 127986 93134
rect 128222 92898 163986 93134
rect 164222 92898 199986 93134
rect 200222 92898 235986 93134
rect 236222 92898 271986 93134
rect 272222 92898 307986 93134
rect 308222 92898 343986 93134
rect 344222 92898 379986 93134
rect 380222 92898 415986 93134
rect 416222 92898 451986 93134
rect 452222 92898 487986 93134
rect 488222 92898 523986 93134
rect 524222 92898 559986 93134
rect 560222 92898 586442 93134
rect 586678 92898 586860 93134
rect -2936 92876 586860 92898
rect -2936 92874 -2336 92876
rect 19804 92874 20404 92876
rect 55804 92874 56404 92876
rect 91804 92874 92404 92876
rect 127804 92874 128404 92876
rect 163804 92874 164404 92876
rect 199804 92874 200404 92876
rect 235804 92874 236404 92876
rect 271804 92874 272404 92876
rect 307804 92874 308404 92876
rect 343804 92874 344404 92876
rect 379804 92874 380404 92876
rect 415804 92874 416404 92876
rect 451804 92874 452404 92876
rect 487804 92874 488404 92876
rect 523804 92874 524404 92876
rect 559804 92874 560404 92876
rect 586260 92874 586860 92876
rect -7636 86276 -7036 86278
rect 12604 86276 13204 86278
rect 48604 86276 49204 86278
rect 84604 86276 85204 86278
rect 120604 86276 121204 86278
rect 156604 86276 157204 86278
rect 192604 86276 193204 86278
rect 228604 86276 229204 86278
rect 264604 86276 265204 86278
rect 300604 86276 301204 86278
rect 336604 86276 337204 86278
rect 372604 86276 373204 86278
rect 408604 86276 409204 86278
rect 444604 86276 445204 86278
rect 480604 86276 481204 86278
rect 516604 86276 517204 86278
rect 552604 86276 553204 86278
rect 590960 86276 591560 86278
rect -8576 86254 592500 86276
rect -8576 86018 -7454 86254
rect -7218 86018 12786 86254
rect 13022 86018 48786 86254
rect 49022 86018 84786 86254
rect 85022 86018 120786 86254
rect 121022 86018 156786 86254
rect 157022 86018 192786 86254
rect 193022 86018 228786 86254
rect 229022 86018 264786 86254
rect 265022 86018 300786 86254
rect 301022 86018 336786 86254
rect 337022 86018 372786 86254
rect 373022 86018 408786 86254
rect 409022 86018 444786 86254
rect 445022 86018 480786 86254
rect 481022 86018 516786 86254
rect 517022 86018 552786 86254
rect 553022 86018 591142 86254
rect 591378 86018 592500 86254
rect -8576 85934 592500 86018
rect -8576 85698 -7454 85934
rect -7218 85698 12786 85934
rect 13022 85698 48786 85934
rect 49022 85698 84786 85934
rect 85022 85698 120786 85934
rect 121022 85698 156786 85934
rect 157022 85698 192786 85934
rect 193022 85698 228786 85934
rect 229022 85698 264786 85934
rect 265022 85698 300786 85934
rect 301022 85698 336786 85934
rect 337022 85698 372786 85934
rect 373022 85698 408786 85934
rect 409022 85698 444786 85934
rect 445022 85698 480786 85934
rect 481022 85698 516786 85934
rect 517022 85698 552786 85934
rect 553022 85698 591142 85934
rect 591378 85698 592500 85934
rect -8576 85676 592500 85698
rect -7636 85674 -7036 85676
rect 12604 85674 13204 85676
rect 48604 85674 49204 85676
rect 84604 85674 85204 85676
rect 120604 85674 121204 85676
rect 156604 85674 157204 85676
rect 192604 85674 193204 85676
rect 228604 85674 229204 85676
rect 264604 85674 265204 85676
rect 300604 85674 301204 85676
rect 336604 85674 337204 85676
rect 372604 85674 373204 85676
rect 408604 85674 409204 85676
rect 444604 85674 445204 85676
rect 480604 85674 481204 85676
rect 516604 85674 517204 85676
rect 552604 85674 553204 85676
rect 590960 85674 591560 85676
rect -5756 82676 -5156 82678
rect 9004 82676 9604 82678
rect 45004 82676 45604 82678
rect 81004 82676 81604 82678
rect 117004 82676 117604 82678
rect 153004 82676 153604 82678
rect 189004 82676 189604 82678
rect 225004 82676 225604 82678
rect 261004 82676 261604 82678
rect 297004 82676 297604 82678
rect 333004 82676 333604 82678
rect 369004 82676 369604 82678
rect 405004 82676 405604 82678
rect 441004 82676 441604 82678
rect 477004 82676 477604 82678
rect 513004 82676 513604 82678
rect 549004 82676 549604 82678
rect 589080 82676 589680 82678
rect -6696 82654 590620 82676
rect -6696 82418 -5574 82654
rect -5338 82418 9186 82654
rect 9422 82418 45186 82654
rect 45422 82418 81186 82654
rect 81422 82418 117186 82654
rect 117422 82418 153186 82654
rect 153422 82418 189186 82654
rect 189422 82418 225186 82654
rect 225422 82418 261186 82654
rect 261422 82418 297186 82654
rect 297422 82418 333186 82654
rect 333422 82418 369186 82654
rect 369422 82418 405186 82654
rect 405422 82418 441186 82654
rect 441422 82418 477186 82654
rect 477422 82418 513186 82654
rect 513422 82418 549186 82654
rect 549422 82418 589262 82654
rect 589498 82418 590620 82654
rect -6696 82334 590620 82418
rect -6696 82098 -5574 82334
rect -5338 82098 9186 82334
rect 9422 82098 45186 82334
rect 45422 82098 81186 82334
rect 81422 82098 117186 82334
rect 117422 82098 153186 82334
rect 153422 82098 189186 82334
rect 189422 82098 225186 82334
rect 225422 82098 261186 82334
rect 261422 82098 297186 82334
rect 297422 82098 333186 82334
rect 333422 82098 369186 82334
rect 369422 82098 405186 82334
rect 405422 82098 441186 82334
rect 441422 82098 477186 82334
rect 477422 82098 513186 82334
rect 513422 82098 549186 82334
rect 549422 82098 589262 82334
rect 589498 82098 590620 82334
rect -6696 82076 590620 82098
rect -5756 82074 -5156 82076
rect 9004 82074 9604 82076
rect 45004 82074 45604 82076
rect 81004 82074 81604 82076
rect 117004 82074 117604 82076
rect 153004 82074 153604 82076
rect 189004 82074 189604 82076
rect 225004 82074 225604 82076
rect 261004 82074 261604 82076
rect 297004 82074 297604 82076
rect 333004 82074 333604 82076
rect 369004 82074 369604 82076
rect 405004 82074 405604 82076
rect 441004 82074 441604 82076
rect 477004 82074 477604 82076
rect 513004 82074 513604 82076
rect 549004 82074 549604 82076
rect 589080 82074 589680 82076
rect -3876 79076 -3276 79078
rect 5404 79076 6004 79078
rect 41404 79076 42004 79078
rect 77404 79076 78004 79078
rect 113404 79076 114004 79078
rect 149404 79076 150004 79078
rect 185404 79076 186004 79078
rect 221404 79076 222004 79078
rect 257404 79076 258004 79078
rect 293404 79076 294004 79078
rect 329404 79076 330004 79078
rect 365404 79076 366004 79078
rect 401404 79076 402004 79078
rect 437404 79076 438004 79078
rect 473404 79076 474004 79078
rect 509404 79076 510004 79078
rect 545404 79076 546004 79078
rect 581404 79076 582004 79078
rect 587200 79076 587800 79078
rect -4816 79054 588740 79076
rect -4816 78818 -3694 79054
rect -3458 78818 5586 79054
rect 5822 78818 41586 79054
rect 41822 78818 77586 79054
rect 77822 78818 113586 79054
rect 113822 78818 149586 79054
rect 149822 78818 185586 79054
rect 185822 78818 221586 79054
rect 221822 78818 257586 79054
rect 257822 78818 293586 79054
rect 293822 78818 329586 79054
rect 329822 78818 365586 79054
rect 365822 78818 401586 79054
rect 401822 78818 437586 79054
rect 437822 78818 473586 79054
rect 473822 78818 509586 79054
rect 509822 78818 545586 79054
rect 545822 78818 581586 79054
rect 581822 78818 587382 79054
rect 587618 78818 588740 79054
rect -4816 78734 588740 78818
rect -4816 78498 -3694 78734
rect -3458 78498 5586 78734
rect 5822 78498 41586 78734
rect 41822 78498 77586 78734
rect 77822 78498 113586 78734
rect 113822 78498 149586 78734
rect 149822 78498 185586 78734
rect 185822 78498 221586 78734
rect 221822 78498 257586 78734
rect 257822 78498 293586 78734
rect 293822 78498 329586 78734
rect 329822 78498 365586 78734
rect 365822 78498 401586 78734
rect 401822 78498 437586 78734
rect 437822 78498 473586 78734
rect 473822 78498 509586 78734
rect 509822 78498 545586 78734
rect 545822 78498 581586 78734
rect 581822 78498 587382 78734
rect 587618 78498 588740 78734
rect -4816 78476 588740 78498
rect -3876 78474 -3276 78476
rect 5404 78474 6004 78476
rect 41404 78474 42004 78476
rect 77404 78474 78004 78476
rect 113404 78474 114004 78476
rect 149404 78474 150004 78476
rect 185404 78474 186004 78476
rect 221404 78474 222004 78476
rect 257404 78474 258004 78476
rect 293404 78474 294004 78476
rect 329404 78474 330004 78476
rect 365404 78474 366004 78476
rect 401404 78474 402004 78476
rect 437404 78474 438004 78476
rect 473404 78474 474004 78476
rect 509404 78474 510004 78476
rect 545404 78474 546004 78476
rect 581404 78474 582004 78476
rect 587200 78474 587800 78476
rect -1996 75476 -1396 75478
rect 1804 75476 2404 75478
rect 37804 75476 38404 75478
rect 73804 75476 74404 75478
rect 109804 75476 110404 75478
rect 145804 75476 146404 75478
rect 181804 75476 182404 75478
rect 217804 75476 218404 75478
rect 253804 75476 254404 75478
rect 289804 75476 290404 75478
rect 325804 75476 326404 75478
rect 361804 75476 362404 75478
rect 397804 75476 398404 75478
rect 433804 75476 434404 75478
rect 469804 75476 470404 75478
rect 505804 75476 506404 75478
rect 541804 75476 542404 75478
rect 577804 75476 578404 75478
rect 585320 75476 585920 75478
rect -2936 75454 586860 75476
rect -2936 75218 -1814 75454
rect -1578 75218 1986 75454
rect 2222 75218 37986 75454
rect 38222 75218 73986 75454
rect 74222 75218 109986 75454
rect 110222 75218 145986 75454
rect 146222 75218 181986 75454
rect 182222 75218 217986 75454
rect 218222 75218 253986 75454
rect 254222 75218 289986 75454
rect 290222 75218 325986 75454
rect 326222 75218 361986 75454
rect 362222 75218 397986 75454
rect 398222 75218 433986 75454
rect 434222 75218 469986 75454
rect 470222 75218 505986 75454
rect 506222 75218 541986 75454
rect 542222 75218 577986 75454
rect 578222 75218 585502 75454
rect 585738 75218 586860 75454
rect -2936 75134 586860 75218
rect -2936 74898 -1814 75134
rect -1578 74898 1986 75134
rect 2222 74898 37986 75134
rect 38222 74898 73986 75134
rect 74222 74898 109986 75134
rect 110222 74898 145986 75134
rect 146222 74898 181986 75134
rect 182222 74898 217986 75134
rect 218222 74898 253986 75134
rect 254222 74898 289986 75134
rect 290222 74898 325986 75134
rect 326222 74898 361986 75134
rect 362222 74898 397986 75134
rect 398222 74898 433986 75134
rect 434222 74898 469986 75134
rect 470222 74898 505986 75134
rect 506222 74898 541986 75134
rect 542222 74898 577986 75134
rect 578222 74898 585502 75134
rect 585738 74898 586860 75134
rect -2936 74876 586860 74898
rect -1996 74874 -1396 74876
rect 1804 74874 2404 74876
rect 37804 74874 38404 74876
rect 73804 74874 74404 74876
rect 109804 74874 110404 74876
rect 145804 74874 146404 74876
rect 181804 74874 182404 74876
rect 217804 74874 218404 74876
rect 253804 74874 254404 74876
rect 289804 74874 290404 74876
rect 325804 74874 326404 74876
rect 361804 74874 362404 74876
rect 397804 74874 398404 74876
rect 433804 74874 434404 74876
rect 469804 74874 470404 74876
rect 505804 74874 506404 74876
rect 541804 74874 542404 74876
rect 577804 74874 578404 74876
rect 585320 74874 585920 74876
rect -8576 68276 -7976 68278
rect 30604 68276 31204 68278
rect 66604 68276 67204 68278
rect 102604 68276 103204 68278
rect 138604 68276 139204 68278
rect 174604 68276 175204 68278
rect 210604 68276 211204 68278
rect 246604 68276 247204 68278
rect 282604 68276 283204 68278
rect 318604 68276 319204 68278
rect 354604 68276 355204 68278
rect 390604 68276 391204 68278
rect 426604 68276 427204 68278
rect 462604 68276 463204 68278
rect 498604 68276 499204 68278
rect 534604 68276 535204 68278
rect 570604 68276 571204 68278
rect 591900 68276 592500 68278
rect -8576 68254 592500 68276
rect -8576 68018 -8394 68254
rect -8158 68018 30786 68254
rect 31022 68018 66786 68254
rect 67022 68018 102786 68254
rect 103022 68018 138786 68254
rect 139022 68018 174786 68254
rect 175022 68018 210786 68254
rect 211022 68018 246786 68254
rect 247022 68018 282786 68254
rect 283022 68018 318786 68254
rect 319022 68018 354786 68254
rect 355022 68018 390786 68254
rect 391022 68018 426786 68254
rect 427022 68018 462786 68254
rect 463022 68018 498786 68254
rect 499022 68018 534786 68254
rect 535022 68018 570786 68254
rect 571022 68018 592082 68254
rect 592318 68018 592500 68254
rect -8576 67934 592500 68018
rect -8576 67698 -8394 67934
rect -8158 67698 30786 67934
rect 31022 67698 66786 67934
rect 67022 67698 102786 67934
rect 103022 67698 138786 67934
rect 139022 67698 174786 67934
rect 175022 67698 210786 67934
rect 211022 67698 246786 67934
rect 247022 67698 282786 67934
rect 283022 67698 318786 67934
rect 319022 67698 354786 67934
rect 355022 67698 390786 67934
rect 391022 67698 426786 67934
rect 427022 67698 462786 67934
rect 463022 67698 498786 67934
rect 499022 67698 534786 67934
rect 535022 67698 570786 67934
rect 571022 67698 592082 67934
rect 592318 67698 592500 67934
rect -8576 67676 592500 67698
rect -8576 67674 -7976 67676
rect 30604 67674 31204 67676
rect 66604 67674 67204 67676
rect 102604 67674 103204 67676
rect 138604 67674 139204 67676
rect 174604 67674 175204 67676
rect 210604 67674 211204 67676
rect 246604 67674 247204 67676
rect 282604 67674 283204 67676
rect 318604 67674 319204 67676
rect 354604 67674 355204 67676
rect 390604 67674 391204 67676
rect 426604 67674 427204 67676
rect 462604 67674 463204 67676
rect 498604 67674 499204 67676
rect 534604 67674 535204 67676
rect 570604 67674 571204 67676
rect 591900 67674 592500 67676
rect -6696 64676 -6096 64678
rect 27004 64676 27604 64678
rect 63004 64676 63604 64678
rect 99004 64676 99604 64678
rect 135004 64676 135604 64678
rect 171004 64676 171604 64678
rect 207004 64676 207604 64678
rect 243004 64676 243604 64678
rect 279004 64676 279604 64678
rect 315004 64676 315604 64678
rect 351004 64676 351604 64678
rect 387004 64676 387604 64678
rect 423004 64676 423604 64678
rect 459004 64676 459604 64678
rect 495004 64676 495604 64678
rect 531004 64676 531604 64678
rect 567004 64676 567604 64678
rect 590020 64676 590620 64678
rect -6696 64654 590620 64676
rect -6696 64418 -6514 64654
rect -6278 64418 27186 64654
rect 27422 64418 63186 64654
rect 63422 64418 99186 64654
rect 99422 64418 135186 64654
rect 135422 64418 171186 64654
rect 171422 64418 207186 64654
rect 207422 64418 243186 64654
rect 243422 64418 279186 64654
rect 279422 64418 315186 64654
rect 315422 64418 351186 64654
rect 351422 64418 387186 64654
rect 387422 64418 423186 64654
rect 423422 64418 459186 64654
rect 459422 64418 495186 64654
rect 495422 64418 531186 64654
rect 531422 64418 567186 64654
rect 567422 64418 590202 64654
rect 590438 64418 590620 64654
rect -6696 64334 590620 64418
rect -6696 64098 -6514 64334
rect -6278 64098 27186 64334
rect 27422 64098 63186 64334
rect 63422 64098 99186 64334
rect 99422 64098 135186 64334
rect 135422 64098 171186 64334
rect 171422 64098 207186 64334
rect 207422 64098 243186 64334
rect 243422 64098 279186 64334
rect 279422 64098 315186 64334
rect 315422 64098 351186 64334
rect 351422 64098 387186 64334
rect 387422 64098 423186 64334
rect 423422 64098 459186 64334
rect 459422 64098 495186 64334
rect 495422 64098 531186 64334
rect 531422 64098 567186 64334
rect 567422 64098 590202 64334
rect 590438 64098 590620 64334
rect -6696 64076 590620 64098
rect -6696 64074 -6096 64076
rect 27004 64074 27604 64076
rect 63004 64074 63604 64076
rect 99004 64074 99604 64076
rect 135004 64074 135604 64076
rect 171004 64074 171604 64076
rect 207004 64074 207604 64076
rect 243004 64074 243604 64076
rect 279004 64074 279604 64076
rect 315004 64074 315604 64076
rect 351004 64074 351604 64076
rect 387004 64074 387604 64076
rect 423004 64074 423604 64076
rect 459004 64074 459604 64076
rect 495004 64074 495604 64076
rect 531004 64074 531604 64076
rect 567004 64074 567604 64076
rect 590020 64074 590620 64076
rect -4816 61076 -4216 61078
rect 23404 61076 24004 61078
rect 59404 61076 60004 61078
rect 95404 61076 96004 61078
rect 131404 61076 132004 61078
rect 167404 61076 168004 61078
rect 203404 61076 204004 61078
rect 239404 61076 240004 61078
rect 275404 61076 276004 61078
rect 311404 61076 312004 61078
rect 347404 61076 348004 61078
rect 383404 61076 384004 61078
rect 419404 61076 420004 61078
rect 455404 61076 456004 61078
rect 491404 61076 492004 61078
rect 527404 61076 528004 61078
rect 563404 61076 564004 61078
rect 588140 61076 588740 61078
rect -4816 61054 588740 61076
rect -4816 60818 -4634 61054
rect -4398 60818 23586 61054
rect 23822 60818 59586 61054
rect 59822 60818 95586 61054
rect 95822 60818 131586 61054
rect 131822 60818 167586 61054
rect 167822 60818 203586 61054
rect 203822 60818 239586 61054
rect 239822 60818 275586 61054
rect 275822 60818 311586 61054
rect 311822 60818 347586 61054
rect 347822 60818 383586 61054
rect 383822 60818 419586 61054
rect 419822 60818 455586 61054
rect 455822 60818 491586 61054
rect 491822 60818 527586 61054
rect 527822 60818 563586 61054
rect 563822 60818 588322 61054
rect 588558 60818 588740 61054
rect -4816 60734 588740 60818
rect -4816 60498 -4634 60734
rect -4398 60498 23586 60734
rect 23822 60498 59586 60734
rect 59822 60498 95586 60734
rect 95822 60498 131586 60734
rect 131822 60498 167586 60734
rect 167822 60498 203586 60734
rect 203822 60498 239586 60734
rect 239822 60498 275586 60734
rect 275822 60498 311586 60734
rect 311822 60498 347586 60734
rect 347822 60498 383586 60734
rect 383822 60498 419586 60734
rect 419822 60498 455586 60734
rect 455822 60498 491586 60734
rect 491822 60498 527586 60734
rect 527822 60498 563586 60734
rect 563822 60498 588322 60734
rect 588558 60498 588740 60734
rect -4816 60476 588740 60498
rect -4816 60474 -4216 60476
rect 23404 60474 24004 60476
rect 59404 60474 60004 60476
rect 95404 60474 96004 60476
rect 131404 60474 132004 60476
rect 167404 60474 168004 60476
rect 203404 60474 204004 60476
rect 239404 60474 240004 60476
rect 275404 60474 276004 60476
rect 311404 60474 312004 60476
rect 347404 60474 348004 60476
rect 383404 60474 384004 60476
rect 419404 60474 420004 60476
rect 455404 60474 456004 60476
rect 491404 60474 492004 60476
rect 527404 60474 528004 60476
rect 563404 60474 564004 60476
rect 588140 60474 588740 60476
rect -2936 57476 -2336 57478
rect 19804 57476 20404 57478
rect 55804 57476 56404 57478
rect 91804 57476 92404 57478
rect 127804 57476 128404 57478
rect 163804 57476 164404 57478
rect 199804 57476 200404 57478
rect 235804 57476 236404 57478
rect 271804 57476 272404 57478
rect 307804 57476 308404 57478
rect 343804 57476 344404 57478
rect 379804 57476 380404 57478
rect 415804 57476 416404 57478
rect 451804 57476 452404 57478
rect 487804 57476 488404 57478
rect 523804 57476 524404 57478
rect 559804 57476 560404 57478
rect 586260 57476 586860 57478
rect -2936 57454 586860 57476
rect -2936 57218 -2754 57454
rect -2518 57218 19986 57454
rect 20222 57218 55986 57454
rect 56222 57218 91986 57454
rect 92222 57218 127986 57454
rect 128222 57218 163986 57454
rect 164222 57218 199986 57454
rect 200222 57218 235986 57454
rect 236222 57218 271986 57454
rect 272222 57218 307986 57454
rect 308222 57218 343986 57454
rect 344222 57218 379986 57454
rect 380222 57218 415986 57454
rect 416222 57218 451986 57454
rect 452222 57218 487986 57454
rect 488222 57218 523986 57454
rect 524222 57218 559986 57454
rect 560222 57218 586442 57454
rect 586678 57218 586860 57454
rect -2936 57134 586860 57218
rect -2936 56898 -2754 57134
rect -2518 56898 19986 57134
rect 20222 56898 55986 57134
rect 56222 56898 91986 57134
rect 92222 56898 127986 57134
rect 128222 56898 163986 57134
rect 164222 56898 199986 57134
rect 200222 56898 235986 57134
rect 236222 56898 271986 57134
rect 272222 56898 307986 57134
rect 308222 56898 343986 57134
rect 344222 56898 379986 57134
rect 380222 56898 415986 57134
rect 416222 56898 451986 57134
rect 452222 56898 487986 57134
rect 488222 56898 523986 57134
rect 524222 56898 559986 57134
rect 560222 56898 586442 57134
rect 586678 56898 586860 57134
rect -2936 56876 586860 56898
rect -2936 56874 -2336 56876
rect 19804 56874 20404 56876
rect 55804 56874 56404 56876
rect 91804 56874 92404 56876
rect 127804 56874 128404 56876
rect 163804 56874 164404 56876
rect 199804 56874 200404 56876
rect 235804 56874 236404 56876
rect 271804 56874 272404 56876
rect 307804 56874 308404 56876
rect 343804 56874 344404 56876
rect 379804 56874 380404 56876
rect 415804 56874 416404 56876
rect 451804 56874 452404 56876
rect 487804 56874 488404 56876
rect 523804 56874 524404 56876
rect 559804 56874 560404 56876
rect 586260 56874 586860 56876
rect -7636 50276 -7036 50278
rect 12604 50276 13204 50278
rect 48604 50276 49204 50278
rect 84604 50276 85204 50278
rect 120604 50276 121204 50278
rect 156604 50276 157204 50278
rect 192604 50276 193204 50278
rect 228604 50276 229204 50278
rect 264604 50276 265204 50278
rect 300604 50276 301204 50278
rect 336604 50276 337204 50278
rect 372604 50276 373204 50278
rect 408604 50276 409204 50278
rect 444604 50276 445204 50278
rect 480604 50276 481204 50278
rect 516604 50276 517204 50278
rect 552604 50276 553204 50278
rect 590960 50276 591560 50278
rect -8576 50254 592500 50276
rect -8576 50018 -7454 50254
rect -7218 50018 12786 50254
rect 13022 50018 48786 50254
rect 49022 50018 84786 50254
rect 85022 50018 120786 50254
rect 121022 50018 156786 50254
rect 157022 50018 192786 50254
rect 193022 50018 228786 50254
rect 229022 50018 264786 50254
rect 265022 50018 300786 50254
rect 301022 50018 336786 50254
rect 337022 50018 372786 50254
rect 373022 50018 408786 50254
rect 409022 50018 444786 50254
rect 445022 50018 480786 50254
rect 481022 50018 516786 50254
rect 517022 50018 552786 50254
rect 553022 50018 591142 50254
rect 591378 50018 592500 50254
rect -8576 49934 592500 50018
rect -8576 49698 -7454 49934
rect -7218 49698 12786 49934
rect 13022 49698 48786 49934
rect 49022 49698 84786 49934
rect 85022 49698 120786 49934
rect 121022 49698 156786 49934
rect 157022 49698 192786 49934
rect 193022 49698 228786 49934
rect 229022 49698 264786 49934
rect 265022 49698 300786 49934
rect 301022 49698 336786 49934
rect 337022 49698 372786 49934
rect 373022 49698 408786 49934
rect 409022 49698 444786 49934
rect 445022 49698 480786 49934
rect 481022 49698 516786 49934
rect 517022 49698 552786 49934
rect 553022 49698 591142 49934
rect 591378 49698 592500 49934
rect -8576 49676 592500 49698
rect -7636 49674 -7036 49676
rect 12604 49674 13204 49676
rect 48604 49674 49204 49676
rect 84604 49674 85204 49676
rect 120604 49674 121204 49676
rect 156604 49674 157204 49676
rect 192604 49674 193204 49676
rect 228604 49674 229204 49676
rect 264604 49674 265204 49676
rect 300604 49674 301204 49676
rect 336604 49674 337204 49676
rect 372604 49674 373204 49676
rect 408604 49674 409204 49676
rect 444604 49674 445204 49676
rect 480604 49674 481204 49676
rect 516604 49674 517204 49676
rect 552604 49674 553204 49676
rect 590960 49674 591560 49676
rect -5756 46676 -5156 46678
rect 9004 46676 9604 46678
rect 45004 46676 45604 46678
rect 81004 46676 81604 46678
rect 117004 46676 117604 46678
rect 153004 46676 153604 46678
rect 189004 46676 189604 46678
rect 225004 46676 225604 46678
rect 261004 46676 261604 46678
rect 297004 46676 297604 46678
rect 333004 46676 333604 46678
rect 369004 46676 369604 46678
rect 405004 46676 405604 46678
rect 441004 46676 441604 46678
rect 477004 46676 477604 46678
rect 513004 46676 513604 46678
rect 549004 46676 549604 46678
rect 589080 46676 589680 46678
rect -6696 46654 590620 46676
rect -6696 46418 -5574 46654
rect -5338 46418 9186 46654
rect 9422 46418 45186 46654
rect 45422 46418 81186 46654
rect 81422 46418 117186 46654
rect 117422 46418 153186 46654
rect 153422 46418 189186 46654
rect 189422 46418 225186 46654
rect 225422 46418 261186 46654
rect 261422 46418 297186 46654
rect 297422 46418 333186 46654
rect 333422 46418 369186 46654
rect 369422 46418 405186 46654
rect 405422 46418 441186 46654
rect 441422 46418 477186 46654
rect 477422 46418 513186 46654
rect 513422 46418 549186 46654
rect 549422 46418 589262 46654
rect 589498 46418 590620 46654
rect -6696 46334 590620 46418
rect -6696 46098 -5574 46334
rect -5338 46098 9186 46334
rect 9422 46098 45186 46334
rect 45422 46098 81186 46334
rect 81422 46098 117186 46334
rect 117422 46098 153186 46334
rect 153422 46098 189186 46334
rect 189422 46098 225186 46334
rect 225422 46098 261186 46334
rect 261422 46098 297186 46334
rect 297422 46098 333186 46334
rect 333422 46098 369186 46334
rect 369422 46098 405186 46334
rect 405422 46098 441186 46334
rect 441422 46098 477186 46334
rect 477422 46098 513186 46334
rect 513422 46098 549186 46334
rect 549422 46098 589262 46334
rect 589498 46098 590620 46334
rect -6696 46076 590620 46098
rect -5756 46074 -5156 46076
rect 9004 46074 9604 46076
rect 45004 46074 45604 46076
rect 81004 46074 81604 46076
rect 117004 46074 117604 46076
rect 153004 46074 153604 46076
rect 189004 46074 189604 46076
rect 225004 46074 225604 46076
rect 261004 46074 261604 46076
rect 297004 46074 297604 46076
rect 333004 46074 333604 46076
rect 369004 46074 369604 46076
rect 405004 46074 405604 46076
rect 441004 46074 441604 46076
rect 477004 46074 477604 46076
rect 513004 46074 513604 46076
rect 549004 46074 549604 46076
rect 589080 46074 589680 46076
rect -3876 43076 -3276 43078
rect 5404 43076 6004 43078
rect 41404 43076 42004 43078
rect 77404 43076 78004 43078
rect 113404 43076 114004 43078
rect 149404 43076 150004 43078
rect 185404 43076 186004 43078
rect 221404 43076 222004 43078
rect 257404 43076 258004 43078
rect 293404 43076 294004 43078
rect 329404 43076 330004 43078
rect 365404 43076 366004 43078
rect 401404 43076 402004 43078
rect 437404 43076 438004 43078
rect 473404 43076 474004 43078
rect 509404 43076 510004 43078
rect 545404 43076 546004 43078
rect 581404 43076 582004 43078
rect 587200 43076 587800 43078
rect -4816 43054 588740 43076
rect -4816 42818 -3694 43054
rect -3458 42818 5586 43054
rect 5822 42818 41586 43054
rect 41822 42818 77586 43054
rect 77822 42818 113586 43054
rect 113822 42818 149586 43054
rect 149822 42818 185586 43054
rect 185822 42818 221586 43054
rect 221822 42818 257586 43054
rect 257822 42818 293586 43054
rect 293822 42818 329586 43054
rect 329822 42818 365586 43054
rect 365822 42818 401586 43054
rect 401822 42818 437586 43054
rect 437822 42818 473586 43054
rect 473822 42818 509586 43054
rect 509822 42818 545586 43054
rect 545822 42818 581586 43054
rect 581822 42818 587382 43054
rect 587618 42818 588740 43054
rect -4816 42734 588740 42818
rect -4816 42498 -3694 42734
rect -3458 42498 5586 42734
rect 5822 42498 41586 42734
rect 41822 42498 77586 42734
rect 77822 42498 113586 42734
rect 113822 42498 149586 42734
rect 149822 42498 185586 42734
rect 185822 42498 221586 42734
rect 221822 42498 257586 42734
rect 257822 42498 293586 42734
rect 293822 42498 329586 42734
rect 329822 42498 365586 42734
rect 365822 42498 401586 42734
rect 401822 42498 437586 42734
rect 437822 42498 473586 42734
rect 473822 42498 509586 42734
rect 509822 42498 545586 42734
rect 545822 42498 581586 42734
rect 581822 42498 587382 42734
rect 587618 42498 588740 42734
rect -4816 42476 588740 42498
rect -3876 42474 -3276 42476
rect 5404 42474 6004 42476
rect 41404 42474 42004 42476
rect 77404 42474 78004 42476
rect 113404 42474 114004 42476
rect 149404 42474 150004 42476
rect 185404 42474 186004 42476
rect 221404 42474 222004 42476
rect 257404 42474 258004 42476
rect 293404 42474 294004 42476
rect 329404 42474 330004 42476
rect 365404 42474 366004 42476
rect 401404 42474 402004 42476
rect 437404 42474 438004 42476
rect 473404 42474 474004 42476
rect 509404 42474 510004 42476
rect 545404 42474 546004 42476
rect 581404 42474 582004 42476
rect 587200 42474 587800 42476
rect -1996 39476 -1396 39478
rect 1804 39476 2404 39478
rect 37804 39476 38404 39478
rect 73804 39476 74404 39478
rect 109804 39476 110404 39478
rect 145804 39476 146404 39478
rect 181804 39476 182404 39478
rect 217804 39476 218404 39478
rect 253804 39476 254404 39478
rect 289804 39476 290404 39478
rect 325804 39476 326404 39478
rect 361804 39476 362404 39478
rect 397804 39476 398404 39478
rect 433804 39476 434404 39478
rect 469804 39476 470404 39478
rect 505804 39476 506404 39478
rect 541804 39476 542404 39478
rect 577804 39476 578404 39478
rect 585320 39476 585920 39478
rect -2936 39454 586860 39476
rect -2936 39218 -1814 39454
rect -1578 39218 1986 39454
rect 2222 39218 37986 39454
rect 38222 39218 73986 39454
rect 74222 39218 109986 39454
rect 110222 39218 145986 39454
rect 146222 39218 181986 39454
rect 182222 39218 217986 39454
rect 218222 39218 253986 39454
rect 254222 39218 289986 39454
rect 290222 39218 325986 39454
rect 326222 39218 361986 39454
rect 362222 39218 397986 39454
rect 398222 39218 433986 39454
rect 434222 39218 469986 39454
rect 470222 39218 505986 39454
rect 506222 39218 541986 39454
rect 542222 39218 577986 39454
rect 578222 39218 585502 39454
rect 585738 39218 586860 39454
rect -2936 39134 586860 39218
rect -2936 38898 -1814 39134
rect -1578 38898 1986 39134
rect 2222 38898 37986 39134
rect 38222 38898 73986 39134
rect 74222 38898 109986 39134
rect 110222 38898 145986 39134
rect 146222 38898 181986 39134
rect 182222 38898 217986 39134
rect 218222 38898 253986 39134
rect 254222 38898 289986 39134
rect 290222 38898 325986 39134
rect 326222 38898 361986 39134
rect 362222 38898 397986 39134
rect 398222 38898 433986 39134
rect 434222 38898 469986 39134
rect 470222 38898 505986 39134
rect 506222 38898 541986 39134
rect 542222 38898 577986 39134
rect 578222 38898 585502 39134
rect 585738 38898 586860 39134
rect -2936 38876 586860 38898
rect -1996 38874 -1396 38876
rect 1804 38874 2404 38876
rect 37804 38874 38404 38876
rect 73804 38874 74404 38876
rect 109804 38874 110404 38876
rect 145804 38874 146404 38876
rect 181804 38874 182404 38876
rect 217804 38874 218404 38876
rect 253804 38874 254404 38876
rect 289804 38874 290404 38876
rect 325804 38874 326404 38876
rect 361804 38874 362404 38876
rect 397804 38874 398404 38876
rect 433804 38874 434404 38876
rect 469804 38874 470404 38876
rect 505804 38874 506404 38876
rect 541804 38874 542404 38876
rect 577804 38874 578404 38876
rect 585320 38874 585920 38876
rect -8576 32276 -7976 32278
rect 30604 32276 31204 32278
rect 66604 32276 67204 32278
rect 102604 32276 103204 32278
rect 138604 32276 139204 32278
rect 174604 32276 175204 32278
rect 210604 32276 211204 32278
rect 246604 32276 247204 32278
rect 282604 32276 283204 32278
rect 318604 32276 319204 32278
rect 354604 32276 355204 32278
rect 390604 32276 391204 32278
rect 426604 32276 427204 32278
rect 462604 32276 463204 32278
rect 498604 32276 499204 32278
rect 534604 32276 535204 32278
rect 570604 32276 571204 32278
rect 591900 32276 592500 32278
rect -8576 32254 592500 32276
rect -8576 32018 -8394 32254
rect -8158 32018 30786 32254
rect 31022 32018 66786 32254
rect 67022 32018 102786 32254
rect 103022 32018 138786 32254
rect 139022 32018 174786 32254
rect 175022 32018 210786 32254
rect 211022 32018 246786 32254
rect 247022 32018 282786 32254
rect 283022 32018 318786 32254
rect 319022 32018 354786 32254
rect 355022 32018 390786 32254
rect 391022 32018 426786 32254
rect 427022 32018 462786 32254
rect 463022 32018 498786 32254
rect 499022 32018 534786 32254
rect 535022 32018 570786 32254
rect 571022 32018 592082 32254
rect 592318 32018 592500 32254
rect -8576 31934 592500 32018
rect -8576 31698 -8394 31934
rect -8158 31698 30786 31934
rect 31022 31698 66786 31934
rect 67022 31698 102786 31934
rect 103022 31698 138786 31934
rect 139022 31698 174786 31934
rect 175022 31698 210786 31934
rect 211022 31698 246786 31934
rect 247022 31698 282786 31934
rect 283022 31698 318786 31934
rect 319022 31698 354786 31934
rect 355022 31698 390786 31934
rect 391022 31698 426786 31934
rect 427022 31698 462786 31934
rect 463022 31698 498786 31934
rect 499022 31698 534786 31934
rect 535022 31698 570786 31934
rect 571022 31698 592082 31934
rect 592318 31698 592500 31934
rect -8576 31676 592500 31698
rect -8576 31674 -7976 31676
rect 30604 31674 31204 31676
rect 66604 31674 67204 31676
rect 102604 31674 103204 31676
rect 138604 31674 139204 31676
rect 174604 31674 175204 31676
rect 210604 31674 211204 31676
rect 246604 31674 247204 31676
rect 282604 31674 283204 31676
rect 318604 31674 319204 31676
rect 354604 31674 355204 31676
rect 390604 31674 391204 31676
rect 426604 31674 427204 31676
rect 462604 31674 463204 31676
rect 498604 31674 499204 31676
rect 534604 31674 535204 31676
rect 570604 31674 571204 31676
rect 591900 31674 592500 31676
rect -6696 28676 -6096 28678
rect 27004 28676 27604 28678
rect 63004 28676 63604 28678
rect 99004 28676 99604 28678
rect 135004 28676 135604 28678
rect 171004 28676 171604 28678
rect 207004 28676 207604 28678
rect 243004 28676 243604 28678
rect 279004 28676 279604 28678
rect 315004 28676 315604 28678
rect 351004 28676 351604 28678
rect 387004 28676 387604 28678
rect 423004 28676 423604 28678
rect 459004 28676 459604 28678
rect 495004 28676 495604 28678
rect 531004 28676 531604 28678
rect 567004 28676 567604 28678
rect 590020 28676 590620 28678
rect -6696 28654 590620 28676
rect -6696 28418 -6514 28654
rect -6278 28418 27186 28654
rect 27422 28418 63186 28654
rect 63422 28418 99186 28654
rect 99422 28418 135186 28654
rect 135422 28418 171186 28654
rect 171422 28418 207186 28654
rect 207422 28418 243186 28654
rect 243422 28418 279186 28654
rect 279422 28418 315186 28654
rect 315422 28418 351186 28654
rect 351422 28418 387186 28654
rect 387422 28418 423186 28654
rect 423422 28418 459186 28654
rect 459422 28418 495186 28654
rect 495422 28418 531186 28654
rect 531422 28418 567186 28654
rect 567422 28418 590202 28654
rect 590438 28418 590620 28654
rect -6696 28334 590620 28418
rect -6696 28098 -6514 28334
rect -6278 28098 27186 28334
rect 27422 28098 63186 28334
rect 63422 28098 99186 28334
rect 99422 28098 135186 28334
rect 135422 28098 171186 28334
rect 171422 28098 207186 28334
rect 207422 28098 243186 28334
rect 243422 28098 279186 28334
rect 279422 28098 315186 28334
rect 315422 28098 351186 28334
rect 351422 28098 387186 28334
rect 387422 28098 423186 28334
rect 423422 28098 459186 28334
rect 459422 28098 495186 28334
rect 495422 28098 531186 28334
rect 531422 28098 567186 28334
rect 567422 28098 590202 28334
rect 590438 28098 590620 28334
rect -6696 28076 590620 28098
rect -6696 28074 -6096 28076
rect 27004 28074 27604 28076
rect 63004 28074 63604 28076
rect 99004 28074 99604 28076
rect 135004 28074 135604 28076
rect 171004 28074 171604 28076
rect 207004 28074 207604 28076
rect 243004 28074 243604 28076
rect 279004 28074 279604 28076
rect 315004 28074 315604 28076
rect 351004 28074 351604 28076
rect 387004 28074 387604 28076
rect 423004 28074 423604 28076
rect 459004 28074 459604 28076
rect 495004 28074 495604 28076
rect 531004 28074 531604 28076
rect 567004 28074 567604 28076
rect 590020 28074 590620 28076
rect -4816 25076 -4216 25078
rect 23404 25076 24004 25078
rect 59404 25076 60004 25078
rect 95404 25076 96004 25078
rect 131404 25076 132004 25078
rect 167404 25076 168004 25078
rect 203404 25076 204004 25078
rect 239404 25076 240004 25078
rect 275404 25076 276004 25078
rect 311404 25076 312004 25078
rect 347404 25076 348004 25078
rect 383404 25076 384004 25078
rect 419404 25076 420004 25078
rect 455404 25076 456004 25078
rect 491404 25076 492004 25078
rect 527404 25076 528004 25078
rect 563404 25076 564004 25078
rect 588140 25076 588740 25078
rect -4816 25054 588740 25076
rect -4816 24818 -4634 25054
rect -4398 24818 23586 25054
rect 23822 24818 59586 25054
rect 59822 24818 95586 25054
rect 95822 24818 131586 25054
rect 131822 24818 167586 25054
rect 167822 24818 203586 25054
rect 203822 24818 239586 25054
rect 239822 24818 275586 25054
rect 275822 24818 311586 25054
rect 311822 24818 347586 25054
rect 347822 24818 383586 25054
rect 383822 24818 419586 25054
rect 419822 24818 455586 25054
rect 455822 24818 491586 25054
rect 491822 24818 527586 25054
rect 527822 24818 563586 25054
rect 563822 24818 588322 25054
rect 588558 24818 588740 25054
rect -4816 24734 588740 24818
rect -4816 24498 -4634 24734
rect -4398 24498 23586 24734
rect 23822 24498 59586 24734
rect 59822 24498 95586 24734
rect 95822 24498 131586 24734
rect 131822 24498 167586 24734
rect 167822 24498 203586 24734
rect 203822 24498 239586 24734
rect 239822 24498 275586 24734
rect 275822 24498 311586 24734
rect 311822 24498 347586 24734
rect 347822 24498 383586 24734
rect 383822 24498 419586 24734
rect 419822 24498 455586 24734
rect 455822 24498 491586 24734
rect 491822 24498 527586 24734
rect 527822 24498 563586 24734
rect 563822 24498 588322 24734
rect 588558 24498 588740 24734
rect -4816 24476 588740 24498
rect -4816 24474 -4216 24476
rect 23404 24474 24004 24476
rect 59404 24474 60004 24476
rect 95404 24474 96004 24476
rect 131404 24474 132004 24476
rect 167404 24474 168004 24476
rect 203404 24474 204004 24476
rect 239404 24474 240004 24476
rect 275404 24474 276004 24476
rect 311404 24474 312004 24476
rect 347404 24474 348004 24476
rect 383404 24474 384004 24476
rect 419404 24474 420004 24476
rect 455404 24474 456004 24476
rect 491404 24474 492004 24476
rect 527404 24474 528004 24476
rect 563404 24474 564004 24476
rect 588140 24474 588740 24476
rect -2936 21476 -2336 21478
rect 19804 21476 20404 21478
rect 55804 21476 56404 21478
rect 91804 21476 92404 21478
rect 127804 21476 128404 21478
rect 163804 21476 164404 21478
rect 199804 21476 200404 21478
rect 235804 21476 236404 21478
rect 271804 21476 272404 21478
rect 307804 21476 308404 21478
rect 343804 21476 344404 21478
rect 379804 21476 380404 21478
rect 415804 21476 416404 21478
rect 451804 21476 452404 21478
rect 487804 21476 488404 21478
rect 523804 21476 524404 21478
rect 559804 21476 560404 21478
rect 586260 21476 586860 21478
rect -2936 21454 586860 21476
rect -2936 21218 -2754 21454
rect -2518 21218 19986 21454
rect 20222 21218 55986 21454
rect 56222 21218 91986 21454
rect 92222 21218 127986 21454
rect 128222 21218 163986 21454
rect 164222 21218 199986 21454
rect 200222 21218 235986 21454
rect 236222 21218 271986 21454
rect 272222 21218 307986 21454
rect 308222 21218 343986 21454
rect 344222 21218 379986 21454
rect 380222 21218 415986 21454
rect 416222 21218 451986 21454
rect 452222 21218 487986 21454
rect 488222 21218 523986 21454
rect 524222 21218 559986 21454
rect 560222 21218 586442 21454
rect 586678 21218 586860 21454
rect -2936 21134 586860 21218
rect -2936 20898 -2754 21134
rect -2518 20898 19986 21134
rect 20222 20898 55986 21134
rect 56222 20898 91986 21134
rect 92222 20898 127986 21134
rect 128222 20898 163986 21134
rect 164222 20898 199986 21134
rect 200222 20898 235986 21134
rect 236222 20898 271986 21134
rect 272222 20898 307986 21134
rect 308222 20898 343986 21134
rect 344222 20898 379986 21134
rect 380222 20898 415986 21134
rect 416222 20898 451986 21134
rect 452222 20898 487986 21134
rect 488222 20898 523986 21134
rect 524222 20898 559986 21134
rect 560222 20898 586442 21134
rect 586678 20898 586860 21134
rect -2936 20876 586860 20898
rect -2936 20874 -2336 20876
rect 19804 20874 20404 20876
rect 55804 20874 56404 20876
rect 91804 20874 92404 20876
rect 127804 20874 128404 20876
rect 163804 20874 164404 20876
rect 199804 20874 200404 20876
rect 235804 20874 236404 20876
rect 271804 20874 272404 20876
rect 307804 20874 308404 20876
rect 343804 20874 344404 20876
rect 379804 20874 380404 20876
rect 415804 20874 416404 20876
rect 451804 20874 452404 20876
rect 487804 20874 488404 20876
rect 523804 20874 524404 20876
rect 559804 20874 560404 20876
rect 586260 20874 586860 20876
rect -7636 14276 -7036 14278
rect 12604 14276 13204 14278
rect 48604 14276 49204 14278
rect 84604 14276 85204 14278
rect 120604 14276 121204 14278
rect 156604 14276 157204 14278
rect 192604 14276 193204 14278
rect 228604 14276 229204 14278
rect 264604 14276 265204 14278
rect 300604 14276 301204 14278
rect 336604 14276 337204 14278
rect 372604 14276 373204 14278
rect 408604 14276 409204 14278
rect 444604 14276 445204 14278
rect 480604 14276 481204 14278
rect 516604 14276 517204 14278
rect 552604 14276 553204 14278
rect 590960 14276 591560 14278
rect -8576 14254 592500 14276
rect -8576 14018 -7454 14254
rect -7218 14018 12786 14254
rect 13022 14018 48786 14254
rect 49022 14018 84786 14254
rect 85022 14018 120786 14254
rect 121022 14018 156786 14254
rect 157022 14018 192786 14254
rect 193022 14018 228786 14254
rect 229022 14018 264786 14254
rect 265022 14018 300786 14254
rect 301022 14018 336786 14254
rect 337022 14018 372786 14254
rect 373022 14018 408786 14254
rect 409022 14018 444786 14254
rect 445022 14018 480786 14254
rect 481022 14018 516786 14254
rect 517022 14018 552786 14254
rect 553022 14018 591142 14254
rect 591378 14018 592500 14254
rect -8576 13934 592500 14018
rect -8576 13698 -7454 13934
rect -7218 13698 12786 13934
rect 13022 13698 48786 13934
rect 49022 13698 84786 13934
rect 85022 13698 120786 13934
rect 121022 13698 156786 13934
rect 157022 13698 192786 13934
rect 193022 13698 228786 13934
rect 229022 13698 264786 13934
rect 265022 13698 300786 13934
rect 301022 13698 336786 13934
rect 337022 13698 372786 13934
rect 373022 13698 408786 13934
rect 409022 13698 444786 13934
rect 445022 13698 480786 13934
rect 481022 13698 516786 13934
rect 517022 13698 552786 13934
rect 553022 13698 591142 13934
rect 591378 13698 592500 13934
rect -8576 13676 592500 13698
rect -7636 13674 -7036 13676
rect 12604 13674 13204 13676
rect 48604 13674 49204 13676
rect 84604 13674 85204 13676
rect 120604 13674 121204 13676
rect 156604 13674 157204 13676
rect 192604 13674 193204 13676
rect 228604 13674 229204 13676
rect 264604 13674 265204 13676
rect 300604 13674 301204 13676
rect 336604 13674 337204 13676
rect 372604 13674 373204 13676
rect 408604 13674 409204 13676
rect 444604 13674 445204 13676
rect 480604 13674 481204 13676
rect 516604 13674 517204 13676
rect 552604 13674 553204 13676
rect 590960 13674 591560 13676
rect -5756 10676 -5156 10678
rect 9004 10676 9604 10678
rect 45004 10676 45604 10678
rect 81004 10676 81604 10678
rect 117004 10676 117604 10678
rect 153004 10676 153604 10678
rect 189004 10676 189604 10678
rect 225004 10676 225604 10678
rect 261004 10676 261604 10678
rect 297004 10676 297604 10678
rect 333004 10676 333604 10678
rect 369004 10676 369604 10678
rect 405004 10676 405604 10678
rect 441004 10676 441604 10678
rect 477004 10676 477604 10678
rect 513004 10676 513604 10678
rect 549004 10676 549604 10678
rect 589080 10676 589680 10678
rect -6696 10654 590620 10676
rect -6696 10418 -5574 10654
rect -5338 10418 9186 10654
rect 9422 10418 45186 10654
rect 45422 10418 81186 10654
rect 81422 10418 117186 10654
rect 117422 10418 153186 10654
rect 153422 10418 189186 10654
rect 189422 10418 225186 10654
rect 225422 10418 261186 10654
rect 261422 10418 297186 10654
rect 297422 10418 333186 10654
rect 333422 10418 369186 10654
rect 369422 10418 405186 10654
rect 405422 10418 441186 10654
rect 441422 10418 477186 10654
rect 477422 10418 513186 10654
rect 513422 10418 549186 10654
rect 549422 10418 589262 10654
rect 589498 10418 590620 10654
rect -6696 10334 590620 10418
rect -6696 10098 -5574 10334
rect -5338 10098 9186 10334
rect 9422 10098 45186 10334
rect 45422 10098 81186 10334
rect 81422 10098 117186 10334
rect 117422 10098 153186 10334
rect 153422 10098 189186 10334
rect 189422 10098 225186 10334
rect 225422 10098 261186 10334
rect 261422 10098 297186 10334
rect 297422 10098 333186 10334
rect 333422 10098 369186 10334
rect 369422 10098 405186 10334
rect 405422 10098 441186 10334
rect 441422 10098 477186 10334
rect 477422 10098 513186 10334
rect 513422 10098 549186 10334
rect 549422 10098 589262 10334
rect 589498 10098 590620 10334
rect -6696 10076 590620 10098
rect -5756 10074 -5156 10076
rect 9004 10074 9604 10076
rect 45004 10074 45604 10076
rect 81004 10074 81604 10076
rect 117004 10074 117604 10076
rect 153004 10074 153604 10076
rect 189004 10074 189604 10076
rect 225004 10074 225604 10076
rect 261004 10074 261604 10076
rect 297004 10074 297604 10076
rect 333004 10074 333604 10076
rect 369004 10074 369604 10076
rect 405004 10074 405604 10076
rect 441004 10074 441604 10076
rect 477004 10074 477604 10076
rect 513004 10074 513604 10076
rect 549004 10074 549604 10076
rect 589080 10074 589680 10076
rect -3876 7076 -3276 7078
rect 5404 7076 6004 7078
rect 41404 7076 42004 7078
rect 77404 7076 78004 7078
rect 113404 7076 114004 7078
rect 149404 7076 150004 7078
rect 185404 7076 186004 7078
rect 221404 7076 222004 7078
rect 257404 7076 258004 7078
rect 293404 7076 294004 7078
rect 329404 7076 330004 7078
rect 365404 7076 366004 7078
rect 401404 7076 402004 7078
rect 437404 7076 438004 7078
rect 473404 7076 474004 7078
rect 509404 7076 510004 7078
rect 545404 7076 546004 7078
rect 581404 7076 582004 7078
rect 587200 7076 587800 7078
rect -4816 7054 588740 7076
rect -4816 6818 -3694 7054
rect -3458 6818 5586 7054
rect 5822 6818 41586 7054
rect 41822 6818 77586 7054
rect 77822 6818 113586 7054
rect 113822 6818 149586 7054
rect 149822 6818 185586 7054
rect 185822 6818 221586 7054
rect 221822 6818 257586 7054
rect 257822 6818 293586 7054
rect 293822 6818 329586 7054
rect 329822 6818 365586 7054
rect 365822 6818 401586 7054
rect 401822 6818 437586 7054
rect 437822 6818 473586 7054
rect 473822 6818 509586 7054
rect 509822 6818 545586 7054
rect 545822 6818 581586 7054
rect 581822 6818 587382 7054
rect 587618 6818 588740 7054
rect -4816 6734 588740 6818
rect -4816 6498 -3694 6734
rect -3458 6498 5586 6734
rect 5822 6498 41586 6734
rect 41822 6498 77586 6734
rect 77822 6498 113586 6734
rect 113822 6498 149586 6734
rect 149822 6498 185586 6734
rect 185822 6498 221586 6734
rect 221822 6498 257586 6734
rect 257822 6498 293586 6734
rect 293822 6498 329586 6734
rect 329822 6498 365586 6734
rect 365822 6498 401586 6734
rect 401822 6498 437586 6734
rect 437822 6498 473586 6734
rect 473822 6498 509586 6734
rect 509822 6498 545586 6734
rect 545822 6498 581586 6734
rect 581822 6498 587382 6734
rect 587618 6498 588740 6734
rect -4816 6476 588740 6498
rect -3876 6474 -3276 6476
rect 5404 6474 6004 6476
rect 41404 6474 42004 6476
rect 77404 6474 78004 6476
rect 113404 6474 114004 6476
rect 149404 6474 150004 6476
rect 185404 6474 186004 6476
rect 221404 6474 222004 6476
rect 257404 6474 258004 6476
rect 293404 6474 294004 6476
rect 329404 6474 330004 6476
rect 365404 6474 366004 6476
rect 401404 6474 402004 6476
rect 437404 6474 438004 6476
rect 473404 6474 474004 6476
rect 509404 6474 510004 6476
rect 545404 6474 546004 6476
rect 581404 6474 582004 6476
rect 587200 6474 587800 6476
rect -1996 3476 -1396 3478
rect 1804 3476 2404 3478
rect 37804 3476 38404 3478
rect 73804 3476 74404 3478
rect 109804 3476 110404 3478
rect 145804 3476 146404 3478
rect 181804 3476 182404 3478
rect 217804 3476 218404 3478
rect 253804 3476 254404 3478
rect 289804 3476 290404 3478
rect 325804 3476 326404 3478
rect 361804 3476 362404 3478
rect 397804 3476 398404 3478
rect 433804 3476 434404 3478
rect 469804 3476 470404 3478
rect 505804 3476 506404 3478
rect 541804 3476 542404 3478
rect 577804 3476 578404 3478
rect 585320 3476 585920 3478
rect -2936 3454 586860 3476
rect -2936 3218 -1814 3454
rect -1578 3218 1986 3454
rect 2222 3218 37986 3454
rect 38222 3218 73986 3454
rect 74222 3218 109986 3454
rect 110222 3218 145986 3454
rect 146222 3218 181986 3454
rect 182222 3218 217986 3454
rect 218222 3218 253986 3454
rect 254222 3218 289986 3454
rect 290222 3218 325986 3454
rect 326222 3218 361986 3454
rect 362222 3218 397986 3454
rect 398222 3218 433986 3454
rect 434222 3218 469986 3454
rect 470222 3218 505986 3454
rect 506222 3218 541986 3454
rect 542222 3218 577986 3454
rect 578222 3218 585502 3454
rect 585738 3218 586860 3454
rect -2936 3134 586860 3218
rect -2936 2898 -1814 3134
rect -1578 2898 1986 3134
rect 2222 2898 37986 3134
rect 38222 2898 73986 3134
rect 74222 2898 109986 3134
rect 110222 2898 145986 3134
rect 146222 2898 181986 3134
rect 182222 2898 217986 3134
rect 218222 2898 253986 3134
rect 254222 2898 289986 3134
rect 290222 2898 325986 3134
rect 326222 2898 361986 3134
rect 362222 2898 397986 3134
rect 398222 2898 433986 3134
rect 434222 2898 469986 3134
rect 470222 2898 505986 3134
rect 506222 2898 541986 3134
rect 542222 2898 577986 3134
rect 578222 2898 585502 3134
rect 585738 2898 586860 3134
rect -2936 2876 586860 2898
rect -1996 2874 -1396 2876
rect 1804 2874 2404 2876
rect 37804 2874 38404 2876
rect 73804 2874 74404 2876
rect 109804 2874 110404 2876
rect 145804 2874 146404 2876
rect 181804 2874 182404 2876
rect 217804 2874 218404 2876
rect 253804 2874 254404 2876
rect 289804 2874 290404 2876
rect 325804 2874 326404 2876
rect 361804 2874 362404 2876
rect 397804 2874 398404 2876
rect 433804 2874 434404 2876
rect 469804 2874 470404 2876
rect 505804 2874 506404 2876
rect 541804 2874 542404 2876
rect 577804 2874 578404 2876
rect 585320 2874 585920 2876
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 1986 -346
rect 2222 -582 37986 -346
rect 38222 -582 73986 -346
rect 74222 -582 109986 -346
rect 110222 -582 145986 -346
rect 146222 -582 181986 -346
rect 182222 -582 217986 -346
rect 218222 -582 253986 -346
rect 254222 -582 289986 -346
rect 290222 -582 325986 -346
rect 326222 -582 361986 -346
rect 362222 -582 397986 -346
rect 398222 -582 433986 -346
rect 434222 -582 469986 -346
rect 470222 -582 505986 -346
rect 506222 -582 541986 -346
rect 542222 -582 577986 -346
rect 578222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 1986 -666
rect 2222 -902 37986 -666
rect 38222 -902 73986 -666
rect 74222 -902 109986 -666
rect 110222 -902 145986 -666
rect 146222 -902 181986 -666
rect 182222 -902 217986 -666
rect 218222 -902 253986 -666
rect 254222 -902 289986 -666
rect 290222 -902 325986 -666
rect 326222 -902 361986 -666
rect 362222 -902 397986 -666
rect 398222 -902 433986 -666
rect 434222 -902 469986 -666
rect 470222 -902 505986 -666
rect 506222 -902 541986 -666
rect 542222 -902 577986 -666
rect 578222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 19986 -1286
rect 20222 -1522 55986 -1286
rect 56222 -1522 91986 -1286
rect 92222 -1522 127986 -1286
rect 128222 -1522 163986 -1286
rect 164222 -1522 199986 -1286
rect 200222 -1522 235986 -1286
rect 236222 -1522 271986 -1286
rect 272222 -1522 307986 -1286
rect 308222 -1522 343986 -1286
rect 344222 -1522 379986 -1286
rect 380222 -1522 415986 -1286
rect 416222 -1522 451986 -1286
rect 452222 -1522 487986 -1286
rect 488222 -1522 523986 -1286
rect 524222 -1522 559986 -1286
rect 560222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 19986 -1606
rect 20222 -1842 55986 -1606
rect 56222 -1842 91986 -1606
rect 92222 -1842 127986 -1606
rect 128222 -1842 163986 -1606
rect 164222 -1842 199986 -1606
rect 200222 -1842 235986 -1606
rect 236222 -1842 271986 -1606
rect 272222 -1842 307986 -1606
rect 308222 -1842 343986 -1606
rect 344222 -1842 379986 -1606
rect 380222 -1842 415986 -1606
rect 416222 -1842 451986 -1606
rect 452222 -1842 487986 -1606
rect 488222 -1842 523986 -1606
rect 524222 -1842 559986 -1606
rect 560222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 5586 -2226
rect 5822 -2462 41586 -2226
rect 41822 -2462 77586 -2226
rect 77822 -2462 113586 -2226
rect 113822 -2462 149586 -2226
rect 149822 -2462 185586 -2226
rect 185822 -2462 221586 -2226
rect 221822 -2462 257586 -2226
rect 257822 -2462 293586 -2226
rect 293822 -2462 329586 -2226
rect 329822 -2462 365586 -2226
rect 365822 -2462 401586 -2226
rect 401822 -2462 437586 -2226
rect 437822 -2462 473586 -2226
rect 473822 -2462 509586 -2226
rect 509822 -2462 545586 -2226
rect 545822 -2462 581586 -2226
rect 581822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 5586 -2546
rect 5822 -2782 41586 -2546
rect 41822 -2782 77586 -2546
rect 77822 -2782 113586 -2546
rect 113822 -2782 149586 -2546
rect 149822 -2782 185586 -2546
rect 185822 -2782 221586 -2546
rect 221822 -2782 257586 -2546
rect 257822 -2782 293586 -2546
rect 293822 -2782 329586 -2546
rect 329822 -2782 365586 -2546
rect 365822 -2782 401586 -2546
rect 401822 -2782 437586 -2546
rect 437822 -2782 473586 -2546
rect 473822 -2782 509586 -2546
rect 509822 -2782 545586 -2546
rect 545822 -2782 581586 -2546
rect 581822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 23586 -3166
rect 23822 -3402 59586 -3166
rect 59822 -3402 95586 -3166
rect 95822 -3402 131586 -3166
rect 131822 -3402 167586 -3166
rect 167822 -3402 203586 -3166
rect 203822 -3402 239586 -3166
rect 239822 -3402 275586 -3166
rect 275822 -3402 311586 -3166
rect 311822 -3402 347586 -3166
rect 347822 -3402 383586 -3166
rect 383822 -3402 419586 -3166
rect 419822 -3402 455586 -3166
rect 455822 -3402 491586 -3166
rect 491822 -3402 527586 -3166
rect 527822 -3402 563586 -3166
rect 563822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 23586 -3486
rect 23822 -3722 59586 -3486
rect 59822 -3722 95586 -3486
rect 95822 -3722 131586 -3486
rect 131822 -3722 167586 -3486
rect 167822 -3722 203586 -3486
rect 203822 -3722 239586 -3486
rect 239822 -3722 275586 -3486
rect 275822 -3722 311586 -3486
rect 311822 -3722 347586 -3486
rect 347822 -3722 383586 -3486
rect 383822 -3722 419586 -3486
rect 419822 -3722 455586 -3486
rect 455822 -3722 491586 -3486
rect 491822 -3722 527586 -3486
rect 527822 -3722 563586 -3486
rect 563822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 9186 -4106
rect 9422 -4342 45186 -4106
rect 45422 -4342 81186 -4106
rect 81422 -4342 117186 -4106
rect 117422 -4342 153186 -4106
rect 153422 -4342 189186 -4106
rect 189422 -4342 225186 -4106
rect 225422 -4342 261186 -4106
rect 261422 -4342 297186 -4106
rect 297422 -4342 333186 -4106
rect 333422 -4342 369186 -4106
rect 369422 -4342 405186 -4106
rect 405422 -4342 441186 -4106
rect 441422 -4342 477186 -4106
rect 477422 -4342 513186 -4106
rect 513422 -4342 549186 -4106
rect 549422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 9186 -4426
rect 9422 -4662 45186 -4426
rect 45422 -4662 81186 -4426
rect 81422 -4662 117186 -4426
rect 117422 -4662 153186 -4426
rect 153422 -4662 189186 -4426
rect 189422 -4662 225186 -4426
rect 225422 -4662 261186 -4426
rect 261422 -4662 297186 -4426
rect 297422 -4662 333186 -4426
rect 333422 -4662 369186 -4426
rect 369422 -4662 405186 -4426
rect 405422 -4662 441186 -4426
rect 441422 -4662 477186 -4426
rect 477422 -4662 513186 -4426
rect 513422 -4662 549186 -4426
rect 549422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 27186 -5046
rect 27422 -5282 63186 -5046
rect 63422 -5282 99186 -5046
rect 99422 -5282 135186 -5046
rect 135422 -5282 171186 -5046
rect 171422 -5282 207186 -5046
rect 207422 -5282 243186 -5046
rect 243422 -5282 279186 -5046
rect 279422 -5282 315186 -5046
rect 315422 -5282 351186 -5046
rect 351422 -5282 387186 -5046
rect 387422 -5282 423186 -5046
rect 423422 -5282 459186 -5046
rect 459422 -5282 495186 -5046
rect 495422 -5282 531186 -5046
rect 531422 -5282 567186 -5046
rect 567422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 27186 -5366
rect 27422 -5602 63186 -5366
rect 63422 -5602 99186 -5366
rect 99422 -5602 135186 -5366
rect 135422 -5602 171186 -5366
rect 171422 -5602 207186 -5366
rect 207422 -5602 243186 -5366
rect 243422 -5602 279186 -5366
rect 279422 -5602 315186 -5366
rect 315422 -5602 351186 -5366
rect 351422 -5602 387186 -5366
rect 387422 -5602 423186 -5366
rect 423422 -5602 459186 -5366
rect 459422 -5602 495186 -5366
rect 495422 -5602 531186 -5366
rect 531422 -5602 567186 -5366
rect 567422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 12786 -5986
rect 13022 -6222 48786 -5986
rect 49022 -6222 84786 -5986
rect 85022 -6222 120786 -5986
rect 121022 -6222 156786 -5986
rect 157022 -6222 192786 -5986
rect 193022 -6222 228786 -5986
rect 229022 -6222 264786 -5986
rect 265022 -6222 300786 -5986
rect 301022 -6222 336786 -5986
rect 337022 -6222 372786 -5986
rect 373022 -6222 408786 -5986
rect 409022 -6222 444786 -5986
rect 445022 -6222 480786 -5986
rect 481022 -6222 516786 -5986
rect 517022 -6222 552786 -5986
rect 553022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 12786 -6306
rect 13022 -6542 48786 -6306
rect 49022 -6542 84786 -6306
rect 85022 -6542 120786 -6306
rect 121022 -6542 156786 -6306
rect 157022 -6542 192786 -6306
rect 193022 -6542 228786 -6306
rect 229022 -6542 264786 -6306
rect 265022 -6542 300786 -6306
rect 301022 -6542 336786 -6306
rect 337022 -6542 372786 -6306
rect 373022 -6542 408786 -6306
rect 409022 -6542 444786 -6306
rect 445022 -6542 480786 -6306
rect 481022 -6542 516786 -6306
rect 517022 -6542 552786 -6306
rect 553022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 30786 -6926
rect 31022 -7162 66786 -6926
rect 67022 -7162 102786 -6926
rect 103022 -7162 138786 -6926
rect 139022 -7162 174786 -6926
rect 175022 -7162 210786 -6926
rect 211022 -7162 246786 -6926
rect 247022 -7162 282786 -6926
rect 283022 -7162 318786 -6926
rect 319022 -7162 354786 -6926
rect 355022 -7162 390786 -6926
rect 391022 -7162 426786 -6926
rect 427022 -7162 462786 -6926
rect 463022 -7162 498786 -6926
rect 499022 -7162 534786 -6926
rect 535022 -7162 570786 -6926
rect 571022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 30786 -7246
rect 31022 -7482 66786 -7246
rect 67022 -7482 102786 -7246
rect 103022 -7482 138786 -7246
rect 139022 -7482 174786 -7246
rect 175022 -7482 210786 -7246
rect 211022 -7482 246786 -7246
rect 247022 -7482 282786 -7246
rect 283022 -7482 318786 -7246
rect 319022 -7482 354786 -7246
rect 355022 -7482 390786 -7246
rect 391022 -7482 426786 -7246
rect 427022 -7482 462786 -7246
rect 463022 -7482 498786 -7246
rect 499022 -7482 534786 -7246
rect 535022 -7482 570786 -7246
rect 571022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
use adc_wrapper  mprj
timestamp 1626123697
transform 1 0 235000 0 1 338000
box 0 0 70000 70000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 533 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 599 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 600 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 601 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 602 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 603 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 604 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 605 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 606 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 607 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 608 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 609 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 610 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 611 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 612 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 613 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 614 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 615 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 616 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 617 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 618 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 619 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 620 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 621 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 622 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 623 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 624 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 625 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 626 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 627 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 628 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 629 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 630 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 577804 -1864 578404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 541804 -1864 542404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 505804 -1864 506404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 469804 -1864 470404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 433804 -1864 434404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 397804 -1864 398404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 361804 -1864 362404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 325804 -1864 326404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 289804 410000 290404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 253804 410000 254404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 217804 -1864 218404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 181804 -1864 182404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 145804 -1864 146404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 109804 -1864 110404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 73804 -1864 74404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 37804 -1864 38404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 1804 -1864 2404 705800 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 289804 -1864 290404 336000 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 253804 -1864 254404 336000 6 vccd1
port 657 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 658 nsew power bidirectional
rlabel metal5 s -2936 686876 586860 687476 6 vccd1
port 659 nsew power bidirectional
rlabel metal5 s -2936 650876 586860 651476 6 vccd1
port 660 nsew power bidirectional
rlabel metal5 s -2936 614876 586860 615476 6 vccd1
port 661 nsew power bidirectional
rlabel metal5 s -2936 578876 586860 579476 6 vccd1
port 662 nsew power bidirectional
rlabel metal5 s -2936 542876 586860 543476 6 vccd1
port 663 nsew power bidirectional
rlabel metal5 s -2936 506876 586860 507476 6 vccd1
port 664 nsew power bidirectional
rlabel metal5 s -2936 470876 586860 471476 6 vccd1
port 665 nsew power bidirectional
rlabel metal5 s -2936 434876 586860 435476 6 vccd1
port 666 nsew power bidirectional
rlabel metal5 s -2936 398876 586860 399476 6 vccd1
port 667 nsew power bidirectional
rlabel metal5 s -2936 362876 586860 363476 6 vccd1
port 668 nsew power bidirectional
rlabel metal5 s -2936 326876 586860 327476 6 vccd1
port 669 nsew power bidirectional
rlabel metal5 s -2936 290876 586860 291476 6 vccd1
port 670 nsew power bidirectional
rlabel metal5 s -2936 254876 586860 255476 6 vccd1
port 671 nsew power bidirectional
rlabel metal5 s -2936 218876 586860 219476 6 vccd1
port 672 nsew power bidirectional
rlabel metal5 s -2936 182876 586860 183476 6 vccd1
port 673 nsew power bidirectional
rlabel metal5 s -2936 146876 586860 147476 6 vccd1
port 674 nsew power bidirectional
rlabel metal5 s -2936 110876 586860 111476 6 vccd1
port 675 nsew power bidirectional
rlabel metal5 s -2936 74876 586860 75476 6 vccd1
port 676 nsew power bidirectional
rlabel metal5 s -2936 38876 586860 39476 6 vccd1
port 677 nsew power bidirectional
rlabel metal5 s -2936 2876 586860 3476 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 679 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 680 nsew ground bidirectional
rlabel metal4 s 559804 -1864 560404 705800 6 vssd1
port 681 nsew ground bidirectional
rlabel metal4 s 523804 -1864 524404 705800 6 vssd1
port 682 nsew ground bidirectional
rlabel metal4 s 487804 -1864 488404 705800 6 vssd1
port 683 nsew ground bidirectional
rlabel metal4 s 451804 -1864 452404 705800 6 vssd1
port 684 nsew ground bidirectional
rlabel metal4 s 415804 -1864 416404 705800 6 vssd1
port 685 nsew ground bidirectional
rlabel metal4 s 379804 -1864 380404 705800 6 vssd1
port 686 nsew ground bidirectional
rlabel metal4 s 343804 -1864 344404 705800 6 vssd1
port 687 nsew ground bidirectional
rlabel metal4 s 307804 -1864 308404 705800 6 vssd1
port 688 nsew ground bidirectional
rlabel metal4 s 271804 410000 272404 705800 6 vssd1
port 689 nsew ground bidirectional
rlabel metal4 s 235804 410000 236404 705800 6 vssd1
port 690 nsew ground bidirectional
rlabel metal4 s 199804 -1864 200404 705800 6 vssd1
port 691 nsew ground bidirectional
rlabel metal4 s 163804 -1864 164404 705800 6 vssd1
port 692 nsew ground bidirectional
rlabel metal4 s 127804 -1864 128404 705800 6 vssd1
port 693 nsew ground bidirectional
rlabel metal4 s 91804 -1864 92404 705800 6 vssd1
port 694 nsew ground bidirectional
rlabel metal4 s 55804 -1864 56404 705800 6 vssd1
port 695 nsew ground bidirectional
rlabel metal4 s 19804 -1864 20404 705800 6 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 271804 -1864 272404 336000 6 vssd1
port 698 nsew ground bidirectional
rlabel metal4 s 235804 -1864 236404 336000 6 vssd1
port 699 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 700 nsew ground bidirectional
rlabel metal5 s -2936 668876 586860 669476 6 vssd1
port 701 nsew ground bidirectional
rlabel metal5 s -2936 632876 586860 633476 6 vssd1
port 702 nsew ground bidirectional
rlabel metal5 s -2936 596876 586860 597476 6 vssd1
port 703 nsew ground bidirectional
rlabel metal5 s -2936 560876 586860 561476 6 vssd1
port 704 nsew ground bidirectional
rlabel metal5 s -2936 524876 586860 525476 6 vssd1
port 705 nsew ground bidirectional
rlabel metal5 s -2936 488876 586860 489476 6 vssd1
port 706 nsew ground bidirectional
rlabel metal5 s -2936 452876 586860 453476 6 vssd1
port 707 nsew ground bidirectional
rlabel metal5 s -2936 416876 586860 417476 6 vssd1
port 708 nsew ground bidirectional
rlabel metal5 s -2936 380876 586860 381476 6 vssd1
port 709 nsew ground bidirectional
rlabel metal5 s -2936 344876 586860 345476 6 vssd1
port 710 nsew ground bidirectional
rlabel metal5 s -2936 308876 586860 309476 6 vssd1
port 711 nsew ground bidirectional
rlabel metal5 s -2936 272876 586860 273476 6 vssd1
port 712 nsew ground bidirectional
rlabel metal5 s -2936 236876 586860 237476 6 vssd1
port 713 nsew ground bidirectional
rlabel metal5 s -2936 200876 586860 201476 6 vssd1
port 714 nsew ground bidirectional
rlabel metal5 s -2936 164876 586860 165476 6 vssd1
port 715 nsew ground bidirectional
rlabel metal5 s -2936 128876 586860 129476 6 vssd1
port 716 nsew ground bidirectional
rlabel metal5 s -2936 92876 586860 93476 6 vssd1
port 717 nsew ground bidirectional
rlabel metal5 s -2936 56876 586860 57476 6 vssd1
port 718 nsew ground bidirectional
rlabel metal5 s -2936 20876 586860 21476 6 vssd1
port 719 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 721 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 707680 6 vccd2
port 722 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 707680 6 vccd2
port 723 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 707680 6 vccd2
port 724 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 707680 6 vccd2
port 725 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 707680 6 vccd2
port 726 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 707680 6 vccd2
port 727 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 707680 6 vccd2
port 728 nsew power bidirectional
rlabel metal4 s 293404 410000 294004 707680 6 vccd2
port 729 nsew power bidirectional
rlabel metal4 s 257404 410000 258004 707680 6 vccd2
port 730 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 707680 6 vccd2
port 731 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 707680 6 vccd2
port 732 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 707680 6 vccd2
port 733 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 707680 6 vccd2
port 734 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 707680 6 vccd2
port 735 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 707680 6 vccd2
port 736 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2
port 737 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 738 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 739 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 336000 6 vccd2
port 740 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 336000 6 vccd2
port 741 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 742 nsew power bidirectional
rlabel metal5 s -4816 690476 588740 691076 6 vccd2
port 743 nsew power bidirectional
rlabel metal5 s -4816 654476 588740 655076 6 vccd2
port 744 nsew power bidirectional
rlabel metal5 s -4816 618476 588740 619076 6 vccd2
port 745 nsew power bidirectional
rlabel metal5 s -4816 582476 588740 583076 6 vccd2
port 746 nsew power bidirectional
rlabel metal5 s -4816 546476 588740 547076 6 vccd2
port 747 nsew power bidirectional
rlabel metal5 s -4816 510476 588740 511076 6 vccd2
port 748 nsew power bidirectional
rlabel metal5 s -4816 474476 588740 475076 6 vccd2
port 749 nsew power bidirectional
rlabel metal5 s -4816 438476 588740 439076 6 vccd2
port 750 nsew power bidirectional
rlabel metal5 s -4816 402476 588740 403076 6 vccd2
port 751 nsew power bidirectional
rlabel metal5 s -4816 366476 588740 367076 6 vccd2
port 752 nsew power bidirectional
rlabel metal5 s -4816 330476 588740 331076 6 vccd2
port 753 nsew power bidirectional
rlabel metal5 s -4816 294476 588740 295076 6 vccd2
port 754 nsew power bidirectional
rlabel metal5 s -4816 258476 588740 259076 6 vccd2
port 755 nsew power bidirectional
rlabel metal5 s -4816 222476 588740 223076 6 vccd2
port 756 nsew power bidirectional
rlabel metal5 s -4816 186476 588740 187076 6 vccd2
port 757 nsew power bidirectional
rlabel metal5 s -4816 150476 588740 151076 6 vccd2
port 758 nsew power bidirectional
rlabel metal5 s -4816 114476 588740 115076 6 vccd2
port 759 nsew power bidirectional
rlabel metal5 s -4816 78476 588740 79076 6 vccd2
port 760 nsew power bidirectional
rlabel metal5 s -4816 42476 588740 43076 6 vccd2
port 761 nsew power bidirectional
rlabel metal5 s -4816 6476 588740 7076 6 vccd2
port 762 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 764 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 707680 6 vssd2
port 765 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 707680 6 vssd2
port 766 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 707680 6 vssd2
port 767 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 707680 6 vssd2
port 768 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 707680 6 vssd2
port 769 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 707680 6 vssd2
port 770 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 707680 6 vssd2
port 771 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 707680 6 vssd2
port 772 nsew ground bidirectional
rlabel metal4 s 275404 410000 276004 707680 6 vssd2
port 773 nsew ground bidirectional
rlabel metal4 s 239404 410000 240004 707680 6 vssd2
port 774 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 707680 6 vssd2
port 775 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 707680 6 vssd2
port 776 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 707680 6 vssd2
port 777 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 707680 6 vssd2
port 778 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 707680 6 vssd2
port 779 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 707680 6 vssd2
port 780 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 781 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 336000 6 vssd2
port 782 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 336000 6 vssd2
port 783 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 784 nsew ground bidirectional
rlabel metal5 s -4816 672476 588740 673076 6 vssd2
port 785 nsew ground bidirectional
rlabel metal5 s -4816 636476 588740 637076 6 vssd2
port 786 nsew ground bidirectional
rlabel metal5 s -4816 600476 588740 601076 6 vssd2
port 787 nsew ground bidirectional
rlabel metal5 s -4816 564476 588740 565076 6 vssd2
port 788 nsew ground bidirectional
rlabel metal5 s -4816 528476 588740 529076 6 vssd2
port 789 nsew ground bidirectional
rlabel metal5 s -4816 492476 588740 493076 6 vssd2
port 790 nsew ground bidirectional
rlabel metal5 s -4816 456476 588740 457076 6 vssd2
port 791 nsew ground bidirectional
rlabel metal5 s -4816 420476 588740 421076 6 vssd2
port 792 nsew ground bidirectional
rlabel metal5 s -4816 384476 588740 385076 6 vssd2
port 793 nsew ground bidirectional
rlabel metal5 s -4816 348476 588740 349076 6 vssd2
port 794 nsew ground bidirectional
rlabel metal5 s -4816 312476 588740 313076 6 vssd2
port 795 nsew ground bidirectional
rlabel metal5 s -4816 276476 588740 277076 6 vssd2
port 796 nsew ground bidirectional
rlabel metal5 s -4816 240476 588740 241076 6 vssd2
port 797 nsew ground bidirectional
rlabel metal5 s -4816 204476 588740 205076 6 vssd2
port 798 nsew ground bidirectional
rlabel metal5 s -4816 168476 588740 169076 6 vssd2
port 799 nsew ground bidirectional
rlabel metal5 s -4816 132476 588740 133076 6 vssd2
port 800 nsew ground bidirectional
rlabel metal5 s -4816 96476 588740 97076 6 vssd2
port 801 nsew ground bidirectional
rlabel metal5 s -4816 60476 588740 61076 6 vssd2
port 802 nsew ground bidirectional
rlabel metal5 s -4816 24476 588740 25076 6 vssd2
port 803 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 549004 -5624 549604 709560 6 vdda1
port 805 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 709560 6 vdda1
port 806 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 709560 6 vdda1
port 807 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 709560 6 vdda1
port 808 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 709560 6 vdda1
port 809 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 709560 6 vdda1
port 810 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 709560 6 vdda1
port 811 nsew power bidirectional
rlabel metal4 s 297004 410000 297604 709560 6 vdda1
port 812 nsew power bidirectional
rlabel metal4 s 261004 410000 261604 709560 6 vdda1
port 813 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 709560 6 vdda1
port 814 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 709560 6 vdda1
port 815 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 709560 6 vdda1
port 816 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 709560 6 vdda1
port 817 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 709560 6 vdda1
port 818 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 709560 6 vdda1
port 819 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1
port 820 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 821 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 822 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 336000 6 vdda1
port 823 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 336000 6 vdda1
port 824 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 825 nsew power bidirectional
rlabel metal5 s -6696 694076 590620 694676 6 vdda1
port 826 nsew power bidirectional
rlabel metal5 s -6696 658076 590620 658676 6 vdda1
port 827 nsew power bidirectional
rlabel metal5 s -6696 622076 590620 622676 6 vdda1
port 828 nsew power bidirectional
rlabel metal5 s -6696 586076 590620 586676 6 vdda1
port 829 nsew power bidirectional
rlabel metal5 s -6696 550076 590620 550676 6 vdda1
port 830 nsew power bidirectional
rlabel metal5 s -6696 514076 590620 514676 6 vdda1
port 831 nsew power bidirectional
rlabel metal5 s -6696 478076 590620 478676 6 vdda1
port 832 nsew power bidirectional
rlabel metal5 s -6696 442076 590620 442676 6 vdda1
port 833 nsew power bidirectional
rlabel metal5 s -6696 406076 590620 406676 6 vdda1
port 834 nsew power bidirectional
rlabel metal5 s -6696 370076 590620 370676 6 vdda1
port 835 nsew power bidirectional
rlabel metal5 s -6696 334076 590620 334676 6 vdda1
port 836 nsew power bidirectional
rlabel metal5 s -6696 298076 590620 298676 6 vdda1
port 837 nsew power bidirectional
rlabel metal5 s -6696 262076 590620 262676 6 vdda1
port 838 nsew power bidirectional
rlabel metal5 s -6696 226076 590620 226676 6 vdda1
port 839 nsew power bidirectional
rlabel metal5 s -6696 190076 590620 190676 6 vdda1
port 840 nsew power bidirectional
rlabel metal5 s -6696 154076 590620 154676 6 vdda1
port 841 nsew power bidirectional
rlabel metal5 s -6696 118076 590620 118676 6 vdda1
port 842 nsew power bidirectional
rlabel metal5 s -6696 82076 590620 82676 6 vdda1
port 843 nsew power bidirectional
rlabel metal5 s -6696 46076 590620 46676 6 vdda1
port 844 nsew power bidirectional
rlabel metal5 s -6696 10076 590620 10676 6 vdda1
port 845 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 846 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 847 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 709560 6 vssa1
port 848 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 709560 6 vssa1
port 849 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 709560 6 vssa1
port 850 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 709560 6 vssa1
port 851 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 709560 6 vssa1
port 852 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 709560 6 vssa1
port 853 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 709560 6 vssa1
port 854 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 709560 6 vssa1
port 855 nsew ground bidirectional
rlabel metal4 s 279004 410000 279604 709560 6 vssa1
port 856 nsew ground bidirectional
rlabel metal4 s 243004 410000 243604 709560 6 vssa1
port 857 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 709560 6 vssa1
port 858 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 709560 6 vssa1
port 859 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 709560 6 vssa1
port 860 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 709560 6 vssa1
port 861 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 709560 6 vssa1
port 862 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 709560 6 vssa1
port 863 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 864 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 336000 6 vssa1
port 865 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 336000 6 vssa1
port 866 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 867 nsew ground bidirectional
rlabel metal5 s -6696 676076 590620 676676 6 vssa1
port 868 nsew ground bidirectional
rlabel metal5 s -6696 640076 590620 640676 6 vssa1
port 869 nsew ground bidirectional
rlabel metal5 s -6696 604076 590620 604676 6 vssa1
port 870 nsew ground bidirectional
rlabel metal5 s -6696 568076 590620 568676 6 vssa1
port 871 nsew ground bidirectional
rlabel metal5 s -6696 532076 590620 532676 6 vssa1
port 872 nsew ground bidirectional
rlabel metal5 s -6696 496076 590620 496676 6 vssa1
port 873 nsew ground bidirectional
rlabel metal5 s -6696 460076 590620 460676 6 vssa1
port 874 nsew ground bidirectional
rlabel metal5 s -6696 424076 590620 424676 6 vssa1
port 875 nsew ground bidirectional
rlabel metal5 s -6696 388076 590620 388676 6 vssa1
port 876 nsew ground bidirectional
rlabel metal5 s -6696 352076 590620 352676 6 vssa1
port 877 nsew ground bidirectional
rlabel metal5 s -6696 316076 590620 316676 6 vssa1
port 878 nsew ground bidirectional
rlabel metal5 s -6696 280076 590620 280676 6 vssa1
port 879 nsew ground bidirectional
rlabel metal5 s -6696 244076 590620 244676 6 vssa1
port 880 nsew ground bidirectional
rlabel metal5 s -6696 208076 590620 208676 6 vssa1
port 881 nsew ground bidirectional
rlabel metal5 s -6696 172076 590620 172676 6 vssa1
port 882 nsew ground bidirectional
rlabel metal5 s -6696 136076 590620 136676 6 vssa1
port 883 nsew ground bidirectional
rlabel metal5 s -6696 100076 590620 100676 6 vssa1
port 884 nsew ground bidirectional
rlabel metal5 s -6696 64076 590620 64676 6 vssa1
port 885 nsew ground bidirectional
rlabel metal5 s -6696 28076 590620 28676 6 vssa1
port 886 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 887 nsew ground bidirectional
rlabel metal4 s 552604 -7504 553204 711440 6 vdda2
port 888 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 711440 6 vdda2
port 889 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 711440 6 vdda2
port 890 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 711440 6 vdda2
port 891 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 711440 6 vdda2
port 892 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 711440 6 vdda2
port 893 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 711440 6 vdda2
port 894 nsew power bidirectional
rlabel metal4 s 300604 410000 301204 711440 6 vdda2
port 895 nsew power bidirectional
rlabel metal4 s 264604 410000 265204 711440 6 vdda2
port 896 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 711440 6 vdda2
port 897 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 711440 6 vdda2
port 898 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 711440 6 vdda2
port 899 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 711440 6 vdda2
port 900 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 711440 6 vdda2
port 901 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 711440 6 vdda2
port 902 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2
port 903 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 904 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 905 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 336000 6 vdda2
port 906 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 336000 6 vdda2
port 907 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 908 nsew power bidirectional
rlabel metal5 s -8576 697676 592500 698276 6 vdda2
port 909 nsew power bidirectional
rlabel metal5 s -8576 661676 592500 662276 6 vdda2
port 910 nsew power bidirectional
rlabel metal5 s -8576 625676 592500 626276 6 vdda2
port 911 nsew power bidirectional
rlabel metal5 s -8576 589676 592500 590276 6 vdda2
port 912 nsew power bidirectional
rlabel metal5 s -8576 553676 592500 554276 6 vdda2
port 913 nsew power bidirectional
rlabel metal5 s -8576 517676 592500 518276 6 vdda2
port 914 nsew power bidirectional
rlabel metal5 s -8576 481676 592500 482276 6 vdda2
port 915 nsew power bidirectional
rlabel metal5 s -8576 445676 592500 446276 6 vdda2
port 916 nsew power bidirectional
rlabel metal5 s -8576 409676 592500 410276 6 vdda2
port 917 nsew power bidirectional
rlabel metal5 s -8576 373676 592500 374276 6 vdda2
port 918 nsew power bidirectional
rlabel metal5 s -8576 337676 592500 338276 6 vdda2
port 919 nsew power bidirectional
rlabel metal5 s -8576 301676 592500 302276 6 vdda2
port 920 nsew power bidirectional
rlabel metal5 s -8576 265676 592500 266276 6 vdda2
port 921 nsew power bidirectional
rlabel metal5 s -8576 229676 592500 230276 6 vdda2
port 922 nsew power bidirectional
rlabel metal5 s -8576 193676 592500 194276 6 vdda2
port 923 nsew power bidirectional
rlabel metal5 s -8576 157676 592500 158276 6 vdda2
port 924 nsew power bidirectional
rlabel metal5 s -8576 121676 592500 122276 6 vdda2
port 925 nsew power bidirectional
rlabel metal5 s -8576 85676 592500 86276 6 vdda2
port 926 nsew power bidirectional
rlabel metal5 s -8576 49676 592500 50276 6 vdda2
port 927 nsew power bidirectional
rlabel metal5 s -8576 13676 592500 14276 6 vdda2
port 928 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 929 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 930 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 711440 6 vssa2
port 931 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 711440 6 vssa2
port 932 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 711440 6 vssa2
port 933 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 711440 6 vssa2
port 934 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 711440 6 vssa2
port 935 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 711440 6 vssa2
port 936 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 711440 6 vssa2
port 937 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 711440 6 vssa2
port 938 nsew ground bidirectional
rlabel metal4 s 282604 410000 283204 711440 6 vssa2
port 939 nsew ground bidirectional
rlabel metal4 s 246604 410000 247204 711440 6 vssa2
port 940 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 711440 6 vssa2
port 941 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 711440 6 vssa2
port 942 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 711440 6 vssa2
port 943 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 711440 6 vssa2
port 944 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 711440 6 vssa2
port 945 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 711440 6 vssa2
port 946 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 947 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 336000 6 vssa2
port 948 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 336000 6 vssa2
port 949 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 950 nsew ground bidirectional
rlabel metal5 s -8576 679676 592500 680276 6 vssa2
port 951 nsew ground bidirectional
rlabel metal5 s -8576 643676 592500 644276 6 vssa2
port 952 nsew ground bidirectional
rlabel metal5 s -8576 607676 592500 608276 6 vssa2
port 953 nsew ground bidirectional
rlabel metal5 s -8576 571676 592500 572276 6 vssa2
port 954 nsew ground bidirectional
rlabel metal5 s -8576 535676 592500 536276 6 vssa2
port 955 nsew ground bidirectional
rlabel metal5 s -8576 499676 592500 500276 6 vssa2
port 956 nsew ground bidirectional
rlabel metal5 s -8576 463676 592500 464276 6 vssa2
port 957 nsew ground bidirectional
rlabel metal5 s -8576 427676 592500 428276 6 vssa2
port 958 nsew ground bidirectional
rlabel metal5 s -8576 391676 592500 392276 6 vssa2
port 959 nsew ground bidirectional
rlabel metal5 s -8576 355676 592500 356276 6 vssa2
port 960 nsew ground bidirectional
rlabel metal5 s -8576 319676 592500 320276 6 vssa2
port 961 nsew ground bidirectional
rlabel metal5 s -8576 283676 592500 284276 6 vssa2
port 962 nsew ground bidirectional
rlabel metal5 s -8576 247676 592500 248276 6 vssa2
port 963 nsew ground bidirectional
rlabel metal5 s -8576 211676 592500 212276 6 vssa2
port 964 nsew ground bidirectional
rlabel metal5 s -8576 175676 592500 176276 6 vssa2
port 965 nsew ground bidirectional
rlabel metal5 s -8576 139676 592500 140276 6 vssa2
port 966 nsew ground bidirectional
rlabel metal5 s -8576 103676 592500 104276 6 vssa2
port 967 nsew ground bidirectional
rlabel metal5 s -8576 67676 592500 68276 6 vssa2
port 968 nsew ground bidirectional
rlabel metal5 s -8576 31676 592500 32276 6 vssa2
port 969 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 970 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
