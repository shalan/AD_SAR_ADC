magic
tech sky130A
magscale 1 2
timestamp 1626449904
<< obsli1 >>
rect 1104 2159 218868 137649
<< obsm1 >>
rect 198 1776 219774 137828
<< metal2 >>
rect 3054 139200 3110 140000
rect 9126 139200 9182 140000
rect 15198 139200 15254 140000
rect 21362 139200 21418 140000
rect 27434 139200 27490 140000
rect 33598 139200 33654 140000
rect 39670 139200 39726 140000
rect 45742 139200 45798 140000
rect 51906 139200 51962 140000
rect 57978 139200 58034 140000
rect 64142 139200 64198 140000
rect 70214 139200 70270 140000
rect 76378 139200 76434 140000
rect 82450 139200 82506 140000
rect 88522 139200 88578 140000
rect 94686 139200 94742 140000
rect 100758 139200 100814 140000
rect 106922 139200 106978 140000
rect 112994 139200 113050 140000
rect 119066 139200 119122 140000
rect 125230 139200 125286 140000
rect 131302 139200 131358 140000
rect 137466 139200 137522 140000
rect 143538 139200 143594 140000
rect 149702 139200 149758 140000
rect 155774 139200 155830 140000
rect 161846 139200 161902 140000
rect 168010 139200 168066 140000
rect 174082 139200 174138 140000
rect 180246 139200 180302 140000
rect 186318 139200 186374 140000
rect 192390 139200 192446 140000
rect 198554 139200 198610 140000
rect 204626 139200 204682 140000
rect 210790 139200 210846 140000
rect 216862 139200 216918 140000
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23294 0 23350 800
rect 23754 0 23810 800
rect 24214 0 24270 800
rect 24674 0 24730 800
rect 25134 0 25190 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26422 0 26478 800
rect 26882 0 26938 800
rect 27342 0 27398 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28630 0 28686 800
rect 29090 0 29146 800
rect 29550 0 29606 800
rect 30010 0 30066 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34426 0 34482 800
rect 34886 0 34942 800
rect 35346 0 35402 800
rect 35806 0 35862 800
rect 36266 0 36322 800
rect 36634 0 36690 800
rect 37094 0 37150 800
rect 37554 0 37610 800
rect 38014 0 38070 800
rect 38474 0 38530 800
rect 38934 0 38990 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40682 0 40738 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42430 0 42486 800
rect 42890 0 42946 800
rect 43350 0 43406 800
rect 43810 0 43866 800
rect 44270 0 44326 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48226 0 48282 800
rect 48686 0 48742 800
rect 49146 0 49202 800
rect 49606 0 49662 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53562 0 53618 800
rect 54022 0 54078 800
rect 54482 0 54538 800
rect 54942 0 54998 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57150 0 57206 800
rect 57610 0 57666 800
rect 58070 0 58126 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 62026 0 62082 800
rect 62486 0 62542 800
rect 62946 0 63002 800
rect 63406 0 63462 800
rect 63866 0 63922 800
rect 64234 0 64290 800
rect 64694 0 64750 800
rect 65154 0 65210 800
rect 65614 0 65670 800
rect 66074 0 66130 800
rect 66534 0 66590 800
rect 66994 0 67050 800
rect 67362 0 67418 800
rect 67822 0 67878 800
rect 68282 0 68338 800
rect 68742 0 68798 800
rect 69202 0 69258 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70490 0 70546 800
rect 70950 0 71006 800
rect 71410 0 71466 800
rect 71870 0 71926 800
rect 72330 0 72386 800
rect 72698 0 72754 800
rect 73158 0 73214 800
rect 73618 0 73674 800
rect 74078 0 74134 800
rect 74538 0 74594 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75826 0 75882 800
rect 76286 0 76342 800
rect 76746 0 76802 800
rect 77206 0 77262 800
rect 77666 0 77722 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78954 0 79010 800
rect 79414 0 79470 800
rect 79874 0 79930 800
rect 80334 0 80390 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81622 0 81678 800
rect 82082 0 82138 800
rect 82542 0 82598 800
rect 83002 0 83058 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84290 0 84346 800
rect 84750 0 84806 800
rect 85210 0 85266 800
rect 85670 0 85726 800
rect 86130 0 86186 800
rect 86498 0 86554 800
rect 86958 0 87014 800
rect 87418 0 87474 800
rect 87878 0 87934 800
rect 88338 0 88394 800
rect 88798 0 88854 800
rect 89258 0 89314 800
rect 89626 0 89682 800
rect 90086 0 90142 800
rect 90546 0 90602 800
rect 91006 0 91062 800
rect 91466 0 91522 800
rect 91926 0 91982 800
rect 92294 0 92350 800
rect 92754 0 92810 800
rect 93214 0 93270 800
rect 93674 0 93730 800
rect 94134 0 94190 800
rect 94594 0 94650 800
rect 94962 0 95018 800
rect 95422 0 95478 800
rect 95882 0 95938 800
rect 96342 0 96398 800
rect 96802 0 96858 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 98090 0 98146 800
rect 98550 0 98606 800
rect 99010 0 99066 800
rect 99470 0 99526 800
rect 99930 0 99986 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101218 0 101274 800
rect 101678 0 101734 800
rect 102138 0 102194 800
rect 102598 0 102654 800
rect 103058 0 103114 800
rect 103426 0 103482 800
rect 103886 0 103942 800
rect 104346 0 104402 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106554 0 106610 800
rect 107014 0 107070 800
rect 107474 0 107530 800
rect 107934 0 107990 800
rect 108394 0 108450 800
rect 108762 0 108818 800
rect 109222 0 109278 800
rect 109682 0 109738 800
rect 110142 0 110198 800
rect 110602 0 110658 800
rect 111062 0 111118 800
rect 111522 0 111578 800
rect 111890 0 111946 800
rect 112350 0 112406 800
rect 112810 0 112866 800
rect 113270 0 113326 800
rect 113730 0 113786 800
rect 114190 0 114246 800
rect 114558 0 114614 800
rect 115018 0 115074 800
rect 115478 0 115534 800
rect 115938 0 115994 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117686 0 117742 800
rect 118146 0 118202 800
rect 118606 0 118662 800
rect 119066 0 119122 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120354 0 120410 800
rect 120814 0 120870 800
rect 121274 0 121330 800
rect 121734 0 121790 800
rect 122194 0 122250 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123482 0 123538 800
rect 123942 0 123998 800
rect 124402 0 124458 800
rect 124862 0 124918 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126150 0 126206 800
rect 126610 0 126666 800
rect 127070 0 127126 800
rect 127530 0 127586 800
rect 127990 0 128046 800
rect 128358 0 128414 800
rect 128818 0 128874 800
rect 129278 0 129334 800
rect 129738 0 129794 800
rect 130198 0 130254 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131486 0 131542 800
rect 131946 0 132002 800
rect 132406 0 132462 800
rect 132866 0 132922 800
rect 133326 0 133382 800
rect 133786 0 133842 800
rect 134154 0 134210 800
rect 134614 0 134670 800
rect 135074 0 135130 800
rect 135534 0 135590 800
rect 135994 0 136050 800
rect 136454 0 136510 800
rect 136822 0 136878 800
rect 137282 0 137338 800
rect 137742 0 137798 800
rect 138202 0 138258 800
rect 138662 0 138718 800
rect 139122 0 139178 800
rect 139490 0 139546 800
rect 139950 0 140006 800
rect 140410 0 140466 800
rect 140870 0 140926 800
rect 141330 0 141386 800
rect 141790 0 141846 800
rect 142158 0 142214 800
rect 142618 0 142674 800
rect 143078 0 143134 800
rect 143538 0 143594 800
rect 143998 0 144054 800
rect 144458 0 144514 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145746 0 145802 800
rect 146206 0 146262 800
rect 146666 0 146722 800
rect 147126 0 147182 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148414 0 148470 800
rect 148874 0 148930 800
rect 149334 0 149390 800
rect 149794 0 149850 800
rect 150254 0 150310 800
rect 150622 0 150678 800
rect 151082 0 151138 800
rect 151542 0 151598 800
rect 152002 0 152058 800
rect 152462 0 152518 800
rect 152922 0 152978 800
rect 153290 0 153346 800
rect 153750 0 153806 800
rect 154210 0 154266 800
rect 154670 0 154726 800
rect 155130 0 155186 800
rect 155590 0 155646 800
rect 156050 0 156106 800
rect 156418 0 156474 800
rect 156878 0 156934 800
rect 157338 0 157394 800
rect 157798 0 157854 800
rect 158258 0 158314 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159546 0 159602 800
rect 160006 0 160062 800
rect 160466 0 160522 800
rect 160926 0 160982 800
rect 161386 0 161442 800
rect 161754 0 161810 800
rect 162214 0 162270 800
rect 162674 0 162730 800
rect 163134 0 163190 800
rect 163594 0 163650 800
rect 164054 0 164110 800
rect 164422 0 164478 800
rect 164882 0 164938 800
rect 165342 0 165398 800
rect 165802 0 165858 800
rect 166262 0 166318 800
rect 166722 0 166778 800
rect 167182 0 167238 800
rect 167550 0 167606 800
rect 168010 0 168066 800
rect 168470 0 168526 800
rect 168930 0 168986 800
rect 169390 0 169446 800
rect 169850 0 169906 800
rect 170218 0 170274 800
rect 170678 0 170734 800
rect 171138 0 171194 800
rect 171598 0 171654 800
rect 172058 0 172114 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173346 0 173402 800
rect 173806 0 173862 800
rect 174266 0 174322 800
rect 174726 0 174782 800
rect 175186 0 175242 800
rect 175554 0 175610 800
rect 176014 0 176070 800
rect 176474 0 176530 800
rect 176934 0 176990 800
rect 177394 0 177450 800
rect 177854 0 177910 800
rect 178314 0 178370 800
rect 178682 0 178738 800
rect 179142 0 179198 800
rect 179602 0 179658 800
rect 180062 0 180118 800
rect 180522 0 180578 800
rect 180982 0 181038 800
rect 181350 0 181406 800
rect 181810 0 181866 800
rect 182270 0 182326 800
rect 182730 0 182786 800
rect 183190 0 183246 800
rect 183650 0 183706 800
rect 184018 0 184074 800
rect 184478 0 184534 800
rect 184938 0 184994 800
rect 185398 0 185454 800
rect 185858 0 185914 800
rect 186318 0 186374 800
rect 186686 0 186742 800
rect 187146 0 187202 800
rect 187606 0 187662 800
rect 188066 0 188122 800
rect 188526 0 188582 800
rect 188986 0 189042 800
rect 189446 0 189502 800
rect 189814 0 189870 800
rect 190274 0 190330 800
rect 190734 0 190790 800
rect 191194 0 191250 800
rect 191654 0 191710 800
rect 192114 0 192170 800
rect 192482 0 192538 800
rect 192942 0 192998 800
rect 193402 0 193458 800
rect 193862 0 193918 800
rect 194322 0 194378 800
rect 194782 0 194838 800
rect 195150 0 195206 800
rect 195610 0 195666 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 196990 0 197046 800
rect 197450 0 197506 800
rect 197818 0 197874 800
rect 198278 0 198334 800
rect 198738 0 198794 800
rect 199198 0 199254 800
rect 199658 0 199714 800
rect 200118 0 200174 800
rect 200578 0 200634 800
rect 200946 0 201002 800
rect 201406 0 201462 800
rect 201866 0 201922 800
rect 202326 0 202382 800
rect 202786 0 202842 800
rect 203246 0 203302 800
rect 203614 0 203670 800
rect 204074 0 204130 800
rect 204534 0 204590 800
rect 204994 0 205050 800
rect 205454 0 205510 800
rect 205914 0 205970 800
rect 206282 0 206338 800
rect 206742 0 206798 800
rect 207202 0 207258 800
rect 207662 0 207718 800
rect 208122 0 208178 800
rect 208582 0 208638 800
rect 208950 0 209006 800
rect 209410 0 209466 800
rect 209870 0 209926 800
rect 210330 0 210386 800
rect 210790 0 210846 800
rect 211250 0 211306 800
rect 211710 0 211766 800
rect 212078 0 212134 800
rect 212538 0 212594 800
rect 212998 0 213054 800
rect 213458 0 213514 800
rect 213918 0 213974 800
rect 214378 0 214434 800
rect 214746 0 214802 800
rect 215206 0 215262 800
rect 215666 0 215722 800
rect 216126 0 216182 800
rect 216586 0 216642 800
rect 217046 0 217102 800
rect 217414 0 217470 800
rect 217874 0 217930 800
rect 218334 0 218390 800
rect 218794 0 218850 800
rect 219254 0 219310 800
rect 219714 0 219770 800
<< obsm2 >>
rect 204 139144 2998 139200
rect 3166 139144 9070 139200
rect 9238 139144 15142 139200
rect 15310 139144 21306 139200
rect 21474 139144 27378 139200
rect 27546 139144 33542 139200
rect 33710 139144 39614 139200
rect 39782 139144 45686 139200
rect 45854 139144 51850 139200
rect 52018 139144 57922 139200
rect 58090 139144 64086 139200
rect 64254 139144 70158 139200
rect 70326 139144 76322 139200
rect 76490 139144 82394 139200
rect 82562 139144 88466 139200
rect 88634 139144 94630 139200
rect 94798 139144 100702 139200
rect 100870 139144 106866 139200
rect 107034 139144 112938 139200
rect 113106 139144 119010 139200
rect 119178 139144 125174 139200
rect 125342 139144 131246 139200
rect 131414 139144 137410 139200
rect 137578 139144 143482 139200
rect 143650 139144 149646 139200
rect 149814 139144 155718 139200
rect 155886 139144 161790 139200
rect 161958 139144 167954 139200
rect 168122 139144 174026 139200
rect 174194 139144 180190 139200
rect 180358 139144 186262 139200
rect 186430 139144 192334 139200
rect 192502 139144 198498 139200
rect 198666 139144 204570 139200
rect 204738 139144 210734 139200
rect 210902 139144 216806 139200
rect 216974 139144 219768 139200
rect 204 856 219768 139144
rect 314 800 514 856
rect 682 800 974 856
rect 1142 800 1434 856
rect 1602 800 1894 856
rect 2062 800 2354 856
rect 2522 800 2814 856
rect 2982 800 3182 856
rect 3350 800 3642 856
rect 3810 800 4102 856
rect 4270 800 4562 856
rect 4730 800 5022 856
rect 5190 800 5482 856
rect 5650 800 5850 856
rect 6018 800 6310 856
rect 6478 800 6770 856
rect 6938 800 7230 856
rect 7398 800 7690 856
rect 7858 800 8150 856
rect 8318 800 8518 856
rect 8686 800 8978 856
rect 9146 800 9438 856
rect 9606 800 9898 856
rect 10066 800 10358 856
rect 10526 800 10818 856
rect 10986 800 11278 856
rect 11446 800 11646 856
rect 11814 800 12106 856
rect 12274 800 12566 856
rect 12734 800 13026 856
rect 13194 800 13486 856
rect 13654 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14774 856
rect 14942 800 15234 856
rect 15402 800 15694 856
rect 15862 800 16154 856
rect 16322 800 16614 856
rect 16782 800 16982 856
rect 17150 800 17442 856
rect 17610 800 17902 856
rect 18070 800 18362 856
rect 18530 800 18822 856
rect 18990 800 19282 856
rect 19450 800 19650 856
rect 19818 800 20110 856
rect 20278 800 20570 856
rect 20738 800 21030 856
rect 21198 800 21490 856
rect 21658 800 21950 856
rect 22118 800 22410 856
rect 22578 800 22778 856
rect 22946 800 23238 856
rect 23406 800 23698 856
rect 23866 800 24158 856
rect 24326 800 24618 856
rect 24786 800 25078 856
rect 25246 800 25446 856
rect 25614 800 25906 856
rect 26074 800 26366 856
rect 26534 800 26826 856
rect 26994 800 27286 856
rect 27454 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28574 856
rect 28742 800 29034 856
rect 29202 800 29494 856
rect 29662 800 29954 856
rect 30122 800 30414 856
rect 30582 800 30782 856
rect 30950 800 31242 856
rect 31410 800 31702 856
rect 31870 800 32162 856
rect 32330 800 32622 856
rect 32790 800 33082 856
rect 33250 800 33542 856
rect 33710 800 33910 856
rect 34078 800 34370 856
rect 34538 800 34830 856
rect 34998 800 35290 856
rect 35458 800 35750 856
rect 35918 800 36210 856
rect 36378 800 36578 856
rect 36746 800 37038 856
rect 37206 800 37498 856
rect 37666 800 37958 856
rect 38126 800 38418 856
rect 38586 800 38878 856
rect 39046 800 39246 856
rect 39414 800 39706 856
rect 39874 800 40166 856
rect 40334 800 40626 856
rect 40794 800 41086 856
rect 41254 800 41546 856
rect 41714 800 41914 856
rect 42082 800 42374 856
rect 42542 800 42834 856
rect 43002 800 43294 856
rect 43462 800 43754 856
rect 43922 800 44214 856
rect 44382 800 44674 856
rect 44842 800 45042 856
rect 45210 800 45502 856
rect 45670 800 45962 856
rect 46130 800 46422 856
rect 46590 800 46882 856
rect 47050 800 47342 856
rect 47510 800 47710 856
rect 47878 800 48170 856
rect 48338 800 48630 856
rect 48798 800 49090 856
rect 49258 800 49550 856
rect 49718 800 50010 856
rect 50178 800 50378 856
rect 50546 800 50838 856
rect 51006 800 51298 856
rect 51466 800 51758 856
rect 51926 800 52218 856
rect 52386 800 52678 856
rect 52846 800 53046 856
rect 53214 800 53506 856
rect 53674 800 53966 856
rect 54134 800 54426 856
rect 54594 800 54886 856
rect 55054 800 55346 856
rect 55514 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56634 856
rect 56802 800 57094 856
rect 57262 800 57554 856
rect 57722 800 58014 856
rect 58182 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59302 856
rect 59470 800 59762 856
rect 59930 800 60222 856
rect 60390 800 60682 856
rect 60850 800 61142 856
rect 61310 800 61510 856
rect 61678 800 61970 856
rect 62138 800 62430 856
rect 62598 800 62890 856
rect 63058 800 63350 856
rect 63518 800 63810 856
rect 63978 800 64178 856
rect 64346 800 64638 856
rect 64806 800 65098 856
rect 65266 800 65558 856
rect 65726 800 66018 856
rect 66186 800 66478 856
rect 66646 800 66938 856
rect 67106 800 67306 856
rect 67474 800 67766 856
rect 67934 800 68226 856
rect 68394 800 68686 856
rect 68854 800 69146 856
rect 69314 800 69606 856
rect 69774 800 69974 856
rect 70142 800 70434 856
rect 70602 800 70894 856
rect 71062 800 71354 856
rect 71522 800 71814 856
rect 71982 800 72274 856
rect 72442 800 72642 856
rect 72810 800 73102 856
rect 73270 800 73562 856
rect 73730 800 74022 856
rect 74190 800 74482 856
rect 74650 800 74942 856
rect 75110 800 75310 856
rect 75478 800 75770 856
rect 75938 800 76230 856
rect 76398 800 76690 856
rect 76858 800 77150 856
rect 77318 800 77610 856
rect 77778 800 78070 856
rect 78238 800 78438 856
rect 78606 800 78898 856
rect 79066 800 79358 856
rect 79526 800 79818 856
rect 79986 800 80278 856
rect 80446 800 80738 856
rect 80906 800 81106 856
rect 81274 800 81566 856
rect 81734 800 82026 856
rect 82194 800 82486 856
rect 82654 800 82946 856
rect 83114 800 83406 856
rect 83574 800 83774 856
rect 83942 800 84234 856
rect 84402 800 84694 856
rect 84862 800 85154 856
rect 85322 800 85614 856
rect 85782 800 86074 856
rect 86242 800 86442 856
rect 86610 800 86902 856
rect 87070 800 87362 856
rect 87530 800 87822 856
rect 87990 800 88282 856
rect 88450 800 88742 856
rect 88910 800 89202 856
rect 89370 800 89570 856
rect 89738 800 90030 856
rect 90198 800 90490 856
rect 90658 800 90950 856
rect 91118 800 91410 856
rect 91578 800 91870 856
rect 92038 800 92238 856
rect 92406 800 92698 856
rect 92866 800 93158 856
rect 93326 800 93618 856
rect 93786 800 94078 856
rect 94246 800 94538 856
rect 94706 800 94906 856
rect 95074 800 95366 856
rect 95534 800 95826 856
rect 95994 800 96286 856
rect 96454 800 96746 856
rect 96914 800 97206 856
rect 97374 800 97574 856
rect 97742 800 98034 856
rect 98202 800 98494 856
rect 98662 800 98954 856
rect 99122 800 99414 856
rect 99582 800 99874 856
rect 100042 800 100334 856
rect 100502 800 100702 856
rect 100870 800 101162 856
rect 101330 800 101622 856
rect 101790 800 102082 856
rect 102250 800 102542 856
rect 102710 800 103002 856
rect 103170 800 103370 856
rect 103538 800 103830 856
rect 103998 800 104290 856
rect 104458 800 104750 856
rect 104918 800 105210 856
rect 105378 800 105670 856
rect 105838 800 106038 856
rect 106206 800 106498 856
rect 106666 800 106958 856
rect 107126 800 107418 856
rect 107586 800 107878 856
rect 108046 800 108338 856
rect 108506 800 108706 856
rect 108874 800 109166 856
rect 109334 800 109626 856
rect 109794 800 110086 856
rect 110254 800 110546 856
rect 110714 800 111006 856
rect 111174 800 111466 856
rect 111634 800 111834 856
rect 112002 800 112294 856
rect 112462 800 112754 856
rect 112922 800 113214 856
rect 113382 800 113674 856
rect 113842 800 114134 856
rect 114302 800 114502 856
rect 114670 800 114962 856
rect 115130 800 115422 856
rect 115590 800 115882 856
rect 116050 800 116342 856
rect 116510 800 116802 856
rect 116970 800 117170 856
rect 117338 800 117630 856
rect 117798 800 118090 856
rect 118258 800 118550 856
rect 118718 800 119010 856
rect 119178 800 119470 856
rect 119638 800 119838 856
rect 120006 800 120298 856
rect 120466 800 120758 856
rect 120926 800 121218 856
rect 121386 800 121678 856
rect 121846 800 122138 856
rect 122306 800 122598 856
rect 122766 800 122966 856
rect 123134 800 123426 856
rect 123594 800 123886 856
rect 124054 800 124346 856
rect 124514 800 124806 856
rect 124974 800 125266 856
rect 125434 800 125634 856
rect 125802 800 126094 856
rect 126262 800 126554 856
rect 126722 800 127014 856
rect 127182 800 127474 856
rect 127642 800 127934 856
rect 128102 800 128302 856
rect 128470 800 128762 856
rect 128930 800 129222 856
rect 129390 800 129682 856
rect 129850 800 130142 856
rect 130310 800 130602 856
rect 130770 800 130970 856
rect 131138 800 131430 856
rect 131598 800 131890 856
rect 132058 800 132350 856
rect 132518 800 132810 856
rect 132978 800 133270 856
rect 133438 800 133730 856
rect 133898 800 134098 856
rect 134266 800 134558 856
rect 134726 800 135018 856
rect 135186 800 135478 856
rect 135646 800 135938 856
rect 136106 800 136398 856
rect 136566 800 136766 856
rect 136934 800 137226 856
rect 137394 800 137686 856
rect 137854 800 138146 856
rect 138314 800 138606 856
rect 138774 800 139066 856
rect 139234 800 139434 856
rect 139602 800 139894 856
rect 140062 800 140354 856
rect 140522 800 140814 856
rect 140982 800 141274 856
rect 141442 800 141734 856
rect 141902 800 142102 856
rect 142270 800 142562 856
rect 142730 800 143022 856
rect 143190 800 143482 856
rect 143650 800 143942 856
rect 144110 800 144402 856
rect 144570 800 144862 856
rect 145030 800 145230 856
rect 145398 800 145690 856
rect 145858 800 146150 856
rect 146318 800 146610 856
rect 146778 800 147070 856
rect 147238 800 147530 856
rect 147698 800 147898 856
rect 148066 800 148358 856
rect 148526 800 148818 856
rect 148986 800 149278 856
rect 149446 800 149738 856
rect 149906 800 150198 856
rect 150366 800 150566 856
rect 150734 800 151026 856
rect 151194 800 151486 856
rect 151654 800 151946 856
rect 152114 800 152406 856
rect 152574 800 152866 856
rect 153034 800 153234 856
rect 153402 800 153694 856
rect 153862 800 154154 856
rect 154322 800 154614 856
rect 154782 800 155074 856
rect 155242 800 155534 856
rect 155702 800 155994 856
rect 156162 800 156362 856
rect 156530 800 156822 856
rect 156990 800 157282 856
rect 157450 800 157742 856
rect 157910 800 158202 856
rect 158370 800 158662 856
rect 158830 800 159030 856
rect 159198 800 159490 856
rect 159658 800 159950 856
rect 160118 800 160410 856
rect 160578 800 160870 856
rect 161038 800 161330 856
rect 161498 800 161698 856
rect 161866 800 162158 856
rect 162326 800 162618 856
rect 162786 800 163078 856
rect 163246 800 163538 856
rect 163706 800 163998 856
rect 164166 800 164366 856
rect 164534 800 164826 856
rect 164994 800 165286 856
rect 165454 800 165746 856
rect 165914 800 166206 856
rect 166374 800 166666 856
rect 166834 800 167126 856
rect 167294 800 167494 856
rect 167662 800 167954 856
rect 168122 800 168414 856
rect 168582 800 168874 856
rect 169042 800 169334 856
rect 169502 800 169794 856
rect 169962 800 170162 856
rect 170330 800 170622 856
rect 170790 800 171082 856
rect 171250 800 171542 856
rect 171710 800 172002 856
rect 172170 800 172462 856
rect 172630 800 172830 856
rect 172998 800 173290 856
rect 173458 800 173750 856
rect 173918 800 174210 856
rect 174378 800 174670 856
rect 174838 800 175130 856
rect 175298 800 175498 856
rect 175666 800 175958 856
rect 176126 800 176418 856
rect 176586 800 176878 856
rect 177046 800 177338 856
rect 177506 800 177798 856
rect 177966 800 178258 856
rect 178426 800 178626 856
rect 178794 800 179086 856
rect 179254 800 179546 856
rect 179714 800 180006 856
rect 180174 800 180466 856
rect 180634 800 180926 856
rect 181094 800 181294 856
rect 181462 800 181754 856
rect 181922 800 182214 856
rect 182382 800 182674 856
rect 182842 800 183134 856
rect 183302 800 183594 856
rect 183762 800 183962 856
rect 184130 800 184422 856
rect 184590 800 184882 856
rect 185050 800 185342 856
rect 185510 800 185802 856
rect 185970 800 186262 856
rect 186430 800 186630 856
rect 186798 800 187090 856
rect 187258 800 187550 856
rect 187718 800 188010 856
rect 188178 800 188470 856
rect 188638 800 188930 856
rect 189098 800 189390 856
rect 189558 800 189758 856
rect 189926 800 190218 856
rect 190386 800 190678 856
rect 190846 800 191138 856
rect 191306 800 191598 856
rect 191766 800 192058 856
rect 192226 800 192426 856
rect 192594 800 192886 856
rect 193054 800 193346 856
rect 193514 800 193806 856
rect 193974 800 194266 856
rect 194434 800 194726 856
rect 194894 800 195094 856
rect 195262 800 195554 856
rect 195722 800 196014 856
rect 196182 800 196474 856
rect 196642 800 196934 856
rect 197102 800 197394 856
rect 197562 800 197762 856
rect 197930 800 198222 856
rect 198390 800 198682 856
rect 198850 800 199142 856
rect 199310 800 199602 856
rect 199770 800 200062 856
rect 200230 800 200522 856
rect 200690 800 200890 856
rect 201058 800 201350 856
rect 201518 800 201810 856
rect 201978 800 202270 856
rect 202438 800 202730 856
rect 202898 800 203190 856
rect 203358 800 203558 856
rect 203726 800 204018 856
rect 204186 800 204478 856
rect 204646 800 204938 856
rect 205106 800 205398 856
rect 205566 800 205858 856
rect 206026 800 206226 856
rect 206394 800 206686 856
rect 206854 800 207146 856
rect 207314 800 207606 856
rect 207774 800 208066 856
rect 208234 800 208526 856
rect 208694 800 208894 856
rect 209062 800 209354 856
rect 209522 800 209814 856
rect 209982 800 210274 856
rect 210442 800 210734 856
rect 210902 800 211194 856
rect 211362 800 211654 856
rect 211822 800 212022 856
rect 212190 800 212482 856
rect 212650 800 212942 856
rect 213110 800 213402 856
rect 213570 800 213862 856
rect 214030 800 214322 856
rect 214490 800 214690 856
rect 214858 800 215150 856
rect 215318 800 215610 856
rect 215778 800 216070 856
rect 216238 800 216530 856
rect 216698 800 216990 856
rect 217158 800 217358 856
rect 217526 800 217818 856
rect 217986 800 218278 856
rect 218446 800 218738 856
rect 218906 800 219198 856
rect 219366 800 219658 856
<< metal3 >>
rect 0 138456 800 138576
rect 219200 138456 220000 138576
rect 0 135872 800 135992
rect 219200 135872 220000 135992
rect 0 133288 800 133408
rect 219200 133152 220000 133272
rect 0 130704 800 130824
rect 219200 130568 220000 130688
rect 0 128120 800 128240
rect 219200 127848 220000 127968
rect 0 125536 800 125656
rect 219200 125264 220000 125384
rect 0 122952 800 123072
rect 219200 122680 220000 122800
rect 0 120368 800 120488
rect 219200 119960 220000 120080
rect 0 117784 800 117904
rect 219200 117376 220000 117496
rect 0 115200 800 115320
rect 219200 114656 220000 114776
rect 0 112616 800 112736
rect 219200 112072 220000 112192
rect 0 110032 800 110152
rect 219200 109488 220000 109608
rect 0 107448 800 107568
rect 219200 106768 220000 106888
rect 0 104864 800 104984
rect 219200 104184 220000 104304
rect 0 102280 800 102400
rect 219200 101464 220000 101584
rect 0 99696 800 99816
rect 219200 98880 220000 99000
rect 0 97112 800 97232
rect 219200 96160 220000 96280
rect 0 94528 800 94648
rect 219200 93576 220000 93696
rect 0 91808 800 91928
rect 219200 90992 220000 91112
rect 0 89224 800 89344
rect 219200 88272 220000 88392
rect 0 86640 800 86760
rect 219200 85688 220000 85808
rect 0 84056 800 84176
rect 219200 82968 220000 83088
rect 0 81472 800 81592
rect 219200 80384 220000 80504
rect 0 78888 800 79008
rect 219200 77800 220000 77920
rect 0 76304 800 76424
rect 219200 75080 220000 75200
rect 0 73720 800 73840
rect 219200 72496 220000 72616
rect 0 71136 800 71256
rect 219200 69776 220000 69896
rect 0 68552 800 68672
rect 219200 67192 220000 67312
rect 0 65968 800 66088
rect 219200 64472 220000 64592
rect 0 63384 800 63504
rect 219200 61888 220000 62008
rect 0 60800 800 60920
rect 219200 59304 220000 59424
rect 0 58216 800 58336
rect 219200 56584 220000 56704
rect 0 55632 800 55752
rect 219200 54000 220000 54120
rect 0 53048 800 53168
rect 219200 51280 220000 51400
rect 0 50464 800 50584
rect 219200 48696 220000 48816
rect 0 47880 800 48000
rect 219200 46112 220000 46232
rect 0 45160 800 45280
rect 219200 43392 220000 43512
rect 0 42576 800 42696
rect 219200 40808 220000 40928
rect 0 39992 800 40112
rect 219200 38088 220000 38208
rect 0 37408 800 37528
rect 219200 35504 220000 35624
rect 0 34824 800 34944
rect 219200 32784 220000 32904
rect 0 32240 800 32360
rect 219200 30200 220000 30320
rect 0 29656 800 29776
rect 219200 27616 220000 27736
rect 0 27072 800 27192
rect 219200 24896 220000 25016
rect 0 24488 800 24608
rect 219200 22312 220000 22432
rect 0 21904 800 22024
rect 219200 19592 220000 19712
rect 0 19320 800 19440
rect 219200 17008 220000 17128
rect 0 16736 800 16856
rect 219200 14424 220000 14544
rect 0 14152 800 14272
rect 0 11568 800 11688
rect 219200 11704 220000 11824
rect 0 8984 800 9104
rect 219200 9120 220000 9240
rect 0 6400 800 6520
rect 219200 6400 220000 6520
rect 0 3816 800 3936
rect 219200 3816 220000 3936
rect 0 1232 800 1352
rect 219200 1232 220000 1352
<< obsm3 >>
rect 880 138376 219120 138549
rect 800 136072 219200 138376
rect 880 135792 219120 136072
rect 800 133488 219200 135792
rect 880 133352 219200 133488
rect 880 133208 219120 133352
rect 800 133072 219120 133208
rect 800 130904 219200 133072
rect 880 130768 219200 130904
rect 880 130624 219120 130768
rect 800 130488 219120 130624
rect 800 128320 219200 130488
rect 880 128048 219200 128320
rect 880 128040 219120 128048
rect 800 127768 219120 128040
rect 800 125736 219200 127768
rect 880 125464 219200 125736
rect 880 125456 219120 125464
rect 800 125184 219120 125456
rect 800 123152 219200 125184
rect 880 122880 219200 123152
rect 880 122872 219120 122880
rect 800 122600 219120 122872
rect 800 120568 219200 122600
rect 880 120288 219200 120568
rect 800 120160 219200 120288
rect 800 119880 219120 120160
rect 800 117984 219200 119880
rect 880 117704 219200 117984
rect 800 117576 219200 117704
rect 800 117296 219120 117576
rect 800 115400 219200 117296
rect 880 115120 219200 115400
rect 800 114856 219200 115120
rect 800 114576 219120 114856
rect 800 112816 219200 114576
rect 880 112536 219200 112816
rect 800 112272 219200 112536
rect 800 111992 219120 112272
rect 800 110232 219200 111992
rect 880 109952 219200 110232
rect 800 109688 219200 109952
rect 800 109408 219120 109688
rect 800 107648 219200 109408
rect 880 107368 219200 107648
rect 800 106968 219200 107368
rect 800 106688 219120 106968
rect 800 105064 219200 106688
rect 880 104784 219200 105064
rect 800 104384 219200 104784
rect 800 104104 219120 104384
rect 800 102480 219200 104104
rect 880 102200 219200 102480
rect 800 101664 219200 102200
rect 800 101384 219120 101664
rect 800 99896 219200 101384
rect 880 99616 219200 99896
rect 800 99080 219200 99616
rect 800 98800 219120 99080
rect 800 97312 219200 98800
rect 880 97032 219200 97312
rect 800 96360 219200 97032
rect 800 96080 219120 96360
rect 800 94728 219200 96080
rect 880 94448 219200 94728
rect 800 93776 219200 94448
rect 800 93496 219120 93776
rect 800 92008 219200 93496
rect 880 91728 219200 92008
rect 800 91192 219200 91728
rect 800 90912 219120 91192
rect 800 89424 219200 90912
rect 880 89144 219200 89424
rect 800 88472 219200 89144
rect 800 88192 219120 88472
rect 800 86840 219200 88192
rect 880 86560 219200 86840
rect 800 85888 219200 86560
rect 800 85608 219120 85888
rect 800 84256 219200 85608
rect 880 83976 219200 84256
rect 800 83168 219200 83976
rect 800 82888 219120 83168
rect 800 81672 219200 82888
rect 880 81392 219200 81672
rect 800 80584 219200 81392
rect 800 80304 219120 80584
rect 800 79088 219200 80304
rect 880 78808 219200 79088
rect 800 78000 219200 78808
rect 800 77720 219120 78000
rect 800 76504 219200 77720
rect 880 76224 219200 76504
rect 800 75280 219200 76224
rect 800 75000 219120 75280
rect 800 73920 219200 75000
rect 880 73640 219200 73920
rect 800 72696 219200 73640
rect 800 72416 219120 72696
rect 800 71336 219200 72416
rect 880 71056 219200 71336
rect 800 69976 219200 71056
rect 800 69696 219120 69976
rect 800 68752 219200 69696
rect 880 68472 219200 68752
rect 800 67392 219200 68472
rect 800 67112 219120 67392
rect 800 66168 219200 67112
rect 880 65888 219200 66168
rect 800 64672 219200 65888
rect 800 64392 219120 64672
rect 800 63584 219200 64392
rect 880 63304 219200 63584
rect 800 62088 219200 63304
rect 800 61808 219120 62088
rect 800 61000 219200 61808
rect 880 60720 219200 61000
rect 800 59504 219200 60720
rect 800 59224 219120 59504
rect 800 58416 219200 59224
rect 880 58136 219200 58416
rect 800 56784 219200 58136
rect 800 56504 219120 56784
rect 800 55832 219200 56504
rect 880 55552 219200 55832
rect 800 54200 219200 55552
rect 800 53920 219120 54200
rect 800 53248 219200 53920
rect 880 52968 219200 53248
rect 800 51480 219200 52968
rect 800 51200 219120 51480
rect 800 50664 219200 51200
rect 880 50384 219200 50664
rect 800 48896 219200 50384
rect 800 48616 219120 48896
rect 800 48080 219200 48616
rect 880 47800 219200 48080
rect 800 46312 219200 47800
rect 800 46032 219120 46312
rect 800 45360 219200 46032
rect 880 45080 219200 45360
rect 800 43592 219200 45080
rect 800 43312 219120 43592
rect 800 42776 219200 43312
rect 880 42496 219200 42776
rect 800 41008 219200 42496
rect 800 40728 219120 41008
rect 800 40192 219200 40728
rect 880 39912 219200 40192
rect 800 38288 219200 39912
rect 800 38008 219120 38288
rect 800 37608 219200 38008
rect 880 37328 219200 37608
rect 800 35704 219200 37328
rect 800 35424 219120 35704
rect 800 35024 219200 35424
rect 880 34744 219200 35024
rect 800 32984 219200 34744
rect 800 32704 219120 32984
rect 800 32440 219200 32704
rect 880 32160 219200 32440
rect 800 30400 219200 32160
rect 800 30120 219120 30400
rect 800 29856 219200 30120
rect 880 29576 219200 29856
rect 800 27816 219200 29576
rect 800 27536 219120 27816
rect 800 27272 219200 27536
rect 880 26992 219200 27272
rect 800 25096 219200 26992
rect 800 24816 219120 25096
rect 800 24688 219200 24816
rect 880 24408 219200 24688
rect 800 22512 219200 24408
rect 800 22232 219120 22512
rect 800 22104 219200 22232
rect 880 21824 219200 22104
rect 800 19792 219200 21824
rect 800 19520 219120 19792
rect 880 19512 219120 19520
rect 880 19240 219200 19512
rect 800 17208 219200 19240
rect 800 16936 219120 17208
rect 880 16928 219120 16936
rect 880 16656 219200 16928
rect 800 14624 219200 16656
rect 800 14352 219120 14624
rect 880 14344 219120 14352
rect 880 14072 219200 14344
rect 800 11904 219200 14072
rect 800 11768 219120 11904
rect 880 11624 219120 11768
rect 880 11488 219200 11624
rect 800 9320 219200 11488
rect 800 9184 219120 9320
rect 880 9040 219120 9184
rect 880 8904 219200 9040
rect 800 6600 219200 8904
rect 880 6320 219120 6600
rect 800 4016 219200 6320
rect 880 3736 219120 4016
rect 800 1432 219200 3736
rect 880 1259 219120 1432
<< metal4 >>
rect 4018 156 4718 139652
rect 5058 -1164 5758 140972
rect 8518 156 9218 139652
rect 9558 -1164 10258 140972
rect 13018 156 13718 139652
rect 14058 -1164 14758 140972
rect 17518 156 18218 139652
rect 18558 16744 19258 140972
rect 22018 16696 22718 139652
rect 23058 16744 23758 140972
rect 26518 16696 27218 139652
rect 27558 16744 28258 140972
rect 31018 16696 31718 139652
rect 32058 16744 32758 140972
rect 35518 16696 36218 139652
rect 36558 16744 37258 140972
rect 18558 -1164 19258 1000
rect 22018 156 22718 1048
rect 23058 -1164 23758 1000
rect 26518 156 27218 1048
rect 27558 -1164 28258 1000
rect 31018 156 31718 1048
rect 32058 -1164 32758 1000
rect 35518 156 36218 1048
rect 36558 -1164 37258 1000
rect 40018 156 40718 139652
rect 41058 -1164 41758 140972
rect 44518 156 45218 139652
rect 45558 -1164 46258 140972
rect 49018 156 49718 139652
rect 50058 -1164 50758 140972
rect 53518 156 54218 139652
rect 54558 -1164 55258 140972
rect 58018 156 58718 139652
rect 59058 -1164 59758 140972
rect 62518 156 63218 139652
rect 63558 -1164 64258 140972
rect 67018 156 67718 139652
rect 68058 -1164 68758 140972
rect 71518 156 72218 139652
rect 72558 -1164 73258 140972
rect 76018 156 76718 139652
rect 77058 -1164 77758 140972
rect 80518 156 81218 139652
rect 81558 -1164 82258 140972
rect 85018 156 85718 139652
rect 86058 -1164 86758 140972
rect 89518 156 90218 139652
rect 90558 -1164 91258 140972
rect 94018 156 94718 139652
rect 95058 -1164 95758 140972
rect 98518 91064 99218 139652
rect 99558 91112 100258 140972
rect 103018 91064 103718 139652
rect 104058 91112 104758 140972
rect 107518 91064 108218 139652
rect 108558 91112 109258 140972
rect 112018 91064 112718 139652
rect 113058 91112 113758 140972
rect 116518 91064 117218 139652
rect 117558 91112 118258 140972
rect 121018 91064 121718 139652
rect 122058 91112 122758 140972
rect 125518 91064 126218 139652
rect 126558 91112 127258 140972
rect 130018 91064 130718 139652
rect 131058 91112 131758 140972
rect 134518 91064 135218 139652
rect 135558 91112 136258 140972
rect 139018 91064 139718 139652
rect 140058 91112 140758 140972
rect 143518 91064 144218 139652
rect 144558 91112 145258 140972
rect 148018 91064 148718 139652
rect 149058 91112 149758 140972
rect 152518 91064 153218 139652
rect 153558 91112 154258 140972
rect 157018 91064 157718 139652
rect 158058 91112 158758 140972
rect 161518 91064 162218 139652
rect 162558 91112 163258 140972
rect 166018 91064 166718 139652
rect 167058 91112 167758 140972
rect 170518 91064 171218 139652
rect 171558 91112 172258 140972
rect 175018 91064 175718 139652
rect 176058 91112 176758 140972
rect 179518 91064 180218 139652
rect 180558 91112 181258 140972
rect 184018 91064 184718 139652
rect 185058 91112 185758 140972
rect 188518 91064 189218 139652
rect 189558 91112 190258 140972
rect 193018 91064 193718 139652
rect 194058 91112 194758 140972
rect 197518 91064 198218 139652
rect 198558 91112 199258 140972
rect 202018 91064 202718 139652
rect 98518 156 99218 21048
rect 99558 -1164 100258 21000
rect 103018 156 103718 21048
rect 104058 -1164 104758 21000
rect 107518 156 108218 21048
rect 108558 -1164 109258 21000
rect 112018 156 112718 21048
rect 113058 -1164 113758 21000
rect 116518 156 117218 21048
rect 117558 -1164 118258 21000
rect 121018 156 121718 21048
rect 122058 -1164 122758 21000
rect 125518 156 126218 21048
rect 126558 -1164 127258 21000
rect 130018 156 130718 21048
rect 131058 -1164 131758 21000
rect 134518 156 135218 21048
rect 135558 -1164 136258 21000
rect 139018 156 139718 21048
rect 140058 -1164 140758 21000
rect 143518 156 144218 21048
rect 144558 -1164 145258 21000
rect 148018 156 148718 21048
rect 149058 -1164 149758 21000
rect 152518 156 153218 21048
rect 153558 -1164 154258 21000
rect 157018 156 157718 21048
rect 158058 -1164 158758 21000
rect 161518 156 162218 21048
rect 162558 -1164 163258 21000
rect 166018 156 166718 21048
rect 167058 -1164 167758 21000
rect 170518 156 171218 21048
rect 171558 -1164 172258 21000
rect 175018 156 175718 21048
rect 176058 -1164 176758 21000
rect 179518 156 180218 21048
rect 180558 -1164 181258 21000
rect 184018 156 184718 21048
rect 185058 -1164 185758 21000
rect 188518 156 189218 21048
rect 189558 -1164 190258 21000
rect 193018 156 193718 21048
rect 194058 -1164 194758 21000
rect 197518 156 198218 21048
rect 198558 -1164 199258 21000
rect 202018 156 202718 21048
rect 203058 -1164 203758 140972
rect 206518 156 207218 139652
rect 207558 -1164 208258 140972
rect 211018 156 211718 139652
rect 212058 -1164 212758 140972
rect 215518 156 216218 139652
rect 216558 -1164 217258 140972
<< obsm4 >>
rect 22798 16664 22978 79014
rect 23838 16664 26438 79014
rect 22798 16616 26438 16664
rect 27298 16664 27478 79014
rect 28338 16664 30938 79014
rect 27298 16616 30938 16664
rect 31798 16664 31978 79014
rect 32838 16664 35438 79014
rect 31798 16616 35438 16664
rect 36298 16664 36478 79014
rect 37338 16664 39938 79014
rect 36298 16616 39938 16664
rect 22000 4000 39938 16616
rect 40798 4000 40978 79014
rect 41838 4000 44438 79014
rect 45298 4000 45478 79014
rect 46338 4000 48938 79014
rect 49798 4000 49978 79014
rect 50838 4000 53438 79014
rect 54298 4000 54478 79014
rect 55338 4000 57938 79014
rect 58798 4000 58978 79014
rect 59838 4000 62438 79014
rect 63298 4000 63478 79014
rect 64338 4000 66938 79014
rect 67798 4000 67978 79014
rect 68838 4000 71438 79014
rect 72298 4000 72478 79014
rect 73338 4000 75938 79014
rect 76798 4000 76978 79014
rect 77838 4000 80438 79014
rect 81298 4000 81478 79014
rect 82338 4000 84938 79014
rect 85798 4000 85978 79014
rect 86838 4000 89438 79014
rect 90298 4000 90478 79014
rect 91338 4000 93938 79014
rect 94798 4000 94978 79014
rect 95838 21128 197798 79014
rect 95838 4000 98438 21128
rect 99298 21080 102938 21128
rect 99298 4000 99478 21080
rect 100338 4000 102938 21080
rect 103798 21080 107438 21128
rect 103798 4000 103978 21080
rect 104838 4000 107438 21080
rect 108298 21080 111938 21128
rect 108298 4000 108478 21080
rect 109338 4000 111938 21080
rect 112798 21080 116438 21128
rect 112798 4000 112978 21080
rect 113838 4000 116438 21080
rect 117298 21080 120938 21128
rect 117298 4000 117478 21080
rect 118338 4000 120938 21080
rect 121798 21080 125438 21128
rect 121798 4000 121978 21080
rect 122838 4000 125438 21080
rect 126298 21080 129938 21128
rect 126298 4000 126478 21080
rect 127338 4000 129938 21080
rect 130798 21080 134438 21128
rect 130798 4000 130978 21080
rect 131838 4000 134438 21080
rect 135298 21080 138938 21128
rect 135298 4000 135478 21080
rect 136338 4000 138938 21080
rect 139798 21080 143438 21128
rect 139798 4000 139978 21080
rect 140838 4000 143438 21080
rect 144298 21080 147938 21128
rect 144298 4000 144478 21080
rect 145338 4000 147938 21080
rect 148798 21080 152438 21128
rect 148798 4000 148978 21080
rect 149838 4000 152438 21080
rect 153298 21080 156938 21128
rect 153298 4000 153478 21080
rect 154338 4000 156938 21080
rect 157798 21080 161438 21128
rect 157798 4000 157978 21080
rect 158838 4000 161438 21080
rect 162298 21080 165938 21128
rect 162298 4000 162478 21080
rect 163338 4000 165938 21080
rect 166798 21080 170438 21128
rect 166798 4000 166978 21080
rect 167838 4000 170438 21080
rect 171298 21080 174938 21128
rect 171298 4000 171478 21080
rect 172338 4000 174938 21080
rect 175798 21080 179438 21128
rect 175798 4000 175978 21080
rect 176838 4000 179438 21080
rect 180298 21080 183938 21128
rect 180298 4000 180478 21080
rect 181338 4000 183938 21080
rect 184798 21080 188438 21128
rect 184798 4000 184978 21080
rect 185838 4000 188438 21080
rect 189298 21080 192938 21128
rect 189298 4000 189478 21080
rect 190338 4000 192938 21080
rect 193798 21080 197438 21128
rect 193798 4000 193978 21080
rect 194838 4000 197438 21080
<< metal5 >>
rect 1104 135608 218868 136308
rect 1104 132196 218868 132896
rect 1104 131108 218868 131808
rect 1104 127696 218868 128396
rect 1104 126608 218868 127308
rect 1104 123196 218868 123896
rect 1104 122108 218868 122808
rect 1104 118696 218868 119396
rect 1104 117608 218868 118308
rect 1104 114196 218868 114896
rect 1104 113108 218868 113808
rect 1104 109696 218868 110396
rect 1104 108608 218868 109308
rect 1104 105196 218868 105896
rect 1104 104108 218868 104808
rect 1104 100696 218868 101396
rect 1104 99608 218868 100308
rect 1104 96196 218868 96896
rect 1104 95108 218868 95808
rect 1104 91696 218868 92396
rect 1104 90608 218868 91308
rect 1104 87196 218868 87896
rect 1104 86108 218868 86808
rect 1104 82696 218868 83396
rect 1104 81608 218868 82308
rect 1104 78196 218868 78896
rect 1104 77108 218868 77808
rect 1104 73696 218868 74396
rect 1104 72608 218868 73308
rect 1104 69196 218868 69896
rect 1104 68108 218868 68808
rect 1104 64696 218868 65396
rect 1104 63608 218868 64308
rect 1104 60196 218868 60896
rect 1104 59108 218868 59808
rect 1104 55696 218868 56396
rect 1104 54608 218868 55308
rect 1104 51196 218868 51896
rect 1104 50108 218868 50808
rect 1104 46696 218868 47396
rect 1104 45608 218868 46308
rect 1104 42196 218868 42896
rect 1104 41108 218868 41808
rect 1104 37696 218868 38396
rect 1104 36608 218868 37308
rect 1104 33196 218868 33896
rect 1104 32108 218868 32808
rect 1104 28696 218868 29396
rect 1104 27608 218868 28308
rect 1104 24196 218868 24896
rect 1104 23108 218868 23808
rect 1104 19696 218868 20396
rect 1104 18608 218868 19308
rect 1104 15196 218868 15896
rect 1104 14108 218868 14808
rect 1104 10696 218868 11396
rect 1104 9608 218868 10308
rect 1104 6196 218868 6896
rect 1104 5108 218868 5808
<< labels >>
rlabel metal3 s 219200 56584 220000 56704 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 168010 139200 168066 140000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 143538 139200 143594 140000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 119066 139200 119122 140000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 94686 139200 94742 140000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 70214 139200 70270 140000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 45742 139200 45798 140000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 21362 139200 21418 140000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 138456 800 138576 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 128120 800 128240 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 117784 800 117904 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 219200 67192 220000 67312 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 107448 800 107568 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 97112 800 97232 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 86640 800 86760 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 76304 800 76424 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 65968 800 66088 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 55632 800 55752 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 45160 800 45280 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 34824 800 34944 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 24488 800 24608 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 219200 77800 220000 77920 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 219200 88272 220000 88392 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 219200 98880 220000 99000 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 219200 109488 220000 109608 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 219200 119960 220000 120080 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 219200 130568 220000 130688 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 216862 139200 216918 140000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 192390 139200 192446 140000 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 219200 1232 220000 1352 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 219200 90992 220000 91112 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 219200 101464 220000 101584 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 219200 112072 220000 112192 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 219200 122680 220000 122800 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 219200 133152 220000 133272 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 210790 139200 210846 140000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 186318 139200 186374 140000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 161846 139200 161902 140000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 137466 139200 137522 140000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 112994 139200 113050 140000 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 219200 9120 220000 9240 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 88522 139200 88578 140000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 64142 139200 64198 140000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 39670 139200 39726 140000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 15198 139200 15254 140000 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 135872 800 135992 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 115200 800 115320 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 219200 17008 220000 17128 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 219200 24896 220000 25016 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 219200 32784 220000 32904 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 219200 40808 220000 40928 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 219200 48696 220000 48816 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 219200 59304 220000 59424 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 219200 69776 220000 69896 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 219200 80384 220000 80504 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 219200 6400 220000 6520 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 219200 96160 220000 96280 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 219200 106768 220000 106888 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 219200 117376 220000 117496 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 219200 127848 220000 127968 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 219200 138456 220000 138576 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 198554 139200 198610 140000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 174082 139200 174138 140000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 149702 139200 149758 140000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 125230 139200 125286 140000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 100758 139200 100814 140000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 219200 14424 220000 14544 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 76378 139200 76434 140000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 51906 139200 51962 140000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 27434 139200 27490 140000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 3054 139200 3110 140000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 130704 800 130824 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 99696 800 99816 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 219200 22312 220000 22432 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 219200 30200 220000 30320 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 219200 38088 220000 38208 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 219200 46112 220000 46232 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 219200 54000 220000 54120 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 219200 64472 220000 64592 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 219200 75080 220000 75200 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 219200 85688 220000 85808 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 219200 3816 220000 3936 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 219200 93576 220000 93696 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 219200 104184 220000 104304 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 219200 114656 220000 114776 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 219200 125264 220000 125384 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 219200 135872 220000 135992 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 204626 139200 204682 140000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 180246 139200 180302 140000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 155774 139200 155830 140000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 131302 139200 131358 140000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 106922 139200 106978 140000 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 219200 11704 220000 11824 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 82450 139200 82506 140000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 57978 139200 58034 140000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 33598 139200 33654 140000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 9126 139200 9182 140000 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 219200 19592 220000 19712 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 71136 800 71256 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 60800 800 60920 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 219200 27616 220000 27736 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 219200 35504 220000 35624 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 219200 43392 220000 43512 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 219200 51280 220000 51400 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 219200 61888 220000 62008 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 219200 72496 220000 72616 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 219200 82968 220000 83088 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 183650 0 183706 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 196990 0 197046 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 202326 0 202382 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 181350 0 181406 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 184018 0 184074 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 190734 0 190790 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 192114 0 192170 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 193402 0 193458 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 194782 0 194838 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 196070 0 196126 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 198738 0 198794 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 200118 0 200174 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 201406 0 201462 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 202786 0 202842 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 208122 0 208178 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 210790 0 210846 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 212078 0 212134 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 213458 0 213514 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 214746 0 214802 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 216126 0 216182 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 217414 0 217470 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 63866 0 63922 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 127990 0 128046 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 141330 0 141386 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 153290 0 153346 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 164054 0 164110 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 165342 0 165398 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 173346 0 173402 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 176014 0 176070 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 180062 0 180118 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 216586 0 216642 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 120354 0 120410 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 169850 0 169906 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 179142 0 179198 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 219714 0 219770 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 532 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 211018 156 211718 139652 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 202018 91064 202718 139652 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 193018 91064 193718 139652 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 184018 91064 184718 139652 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 175018 91064 175718 139652 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 166018 91064 166718 139652 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 157018 91064 157718 139652 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 148018 91064 148718 139652 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 139018 91064 139718 139652 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 130018 91064 130718 139652 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 121018 91064 121718 139652 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 112018 91064 112718 139652 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 103018 91064 103718 139652 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 94018 156 94718 139652 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 85018 156 85718 139652 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 76018 156 76718 139652 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 67018 156 67718 139652 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 58018 156 58718 139652 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 49018 156 49718 139652 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 40018 156 40718 139652 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 31018 16696 31718 139652 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 22018 16696 22718 139652 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 13018 156 13718 139652 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 4018 156 4718 139652 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 202018 156 202718 21048 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 193018 156 193718 21048 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 184018 156 184718 21048 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 175018 156 175718 21048 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 166018 156 166718 21048 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 157018 156 157718 21048 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 148018 156 148718 21048 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 139018 156 139718 21048 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 130018 156 130718 21048 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 121018 156 121718 21048 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 112018 156 112718 21048 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 103018 156 103718 21048 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 31018 156 31718 1048 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s 22018 156 22718 1048 6 vccd1
port 675 nsew power bidirectional
rlabel metal5 s 1104 131108 218868 131808 6 vccd1
port 676 nsew power bidirectional
rlabel metal5 s 1104 122108 218868 122808 6 vccd1
port 677 nsew power bidirectional
rlabel metal5 s 1104 113108 218868 113808 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s 1104 104108 218868 104808 6 vccd1
port 679 nsew power bidirectional
rlabel metal5 s 1104 95108 218868 95808 6 vccd1
port 680 nsew power bidirectional
rlabel metal5 s 1104 86108 218868 86808 6 vccd1
port 681 nsew power bidirectional
rlabel metal5 s 1104 77108 218868 77808 6 vccd1
port 682 nsew power bidirectional
rlabel metal5 s 1104 68108 218868 68808 6 vccd1
port 683 nsew power bidirectional
rlabel metal5 s 1104 59108 218868 59808 6 vccd1
port 684 nsew power bidirectional
rlabel metal5 s 1104 50108 218868 50808 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s 1104 41108 218868 41808 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s 1104 32108 218868 32808 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s 1104 23108 218868 23808 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s 1104 14108 218868 14808 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s 1104 5108 218868 5808 6 vccd1
port 690 nsew power bidirectional
rlabel metal4 s 215518 156 216218 139652 6 vssd1
port 691 nsew ground bidirectional
rlabel metal4 s 206518 156 207218 139652 6 vssd1
port 692 nsew ground bidirectional
rlabel metal4 s 197518 91064 198218 139652 6 vssd1
port 693 nsew ground bidirectional
rlabel metal4 s 188518 91064 189218 139652 6 vssd1
port 694 nsew ground bidirectional
rlabel metal4 s 179518 91064 180218 139652 6 vssd1
port 695 nsew ground bidirectional
rlabel metal4 s 170518 91064 171218 139652 6 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s 161518 91064 162218 139652 6 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 152518 91064 153218 139652 6 vssd1
port 698 nsew ground bidirectional
rlabel metal4 s 143518 91064 144218 139652 6 vssd1
port 699 nsew ground bidirectional
rlabel metal4 s 134518 91064 135218 139652 6 vssd1
port 700 nsew ground bidirectional
rlabel metal4 s 125518 91064 126218 139652 6 vssd1
port 701 nsew ground bidirectional
rlabel metal4 s 116518 91064 117218 139652 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 107518 91064 108218 139652 6 vssd1
port 703 nsew ground bidirectional
rlabel metal4 s 98518 91064 99218 139652 6 vssd1
port 704 nsew ground bidirectional
rlabel metal4 s 89518 156 90218 139652 6 vssd1
port 705 nsew ground bidirectional
rlabel metal4 s 80518 156 81218 139652 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 71518 156 72218 139652 6 vssd1
port 707 nsew ground bidirectional
rlabel metal4 s 62518 156 63218 139652 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s 53518 156 54218 139652 6 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s 44518 156 45218 139652 6 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 35518 16696 36218 139652 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 26518 16696 27218 139652 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 17518 156 18218 139652 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 8518 156 9218 139652 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 197518 156 198218 21048 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 188518 156 189218 21048 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 179518 156 180218 21048 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 170518 156 171218 21048 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 161518 156 162218 21048 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 152518 156 153218 21048 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 143518 156 144218 21048 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 134518 156 135218 21048 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 125518 156 126218 21048 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 116518 156 117218 21048 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s 107518 156 108218 21048 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 98518 156 99218 21048 6 vssd1
port 726 nsew ground bidirectional
rlabel metal4 s 35518 156 36218 1048 6 vssd1
port 727 nsew ground bidirectional
rlabel metal4 s 26518 156 27218 1048 6 vssd1
port 728 nsew ground bidirectional
rlabel metal5 s 1104 135608 218868 136308 6 vssd1
port 729 nsew ground bidirectional
rlabel metal5 s 1104 126608 218868 127308 6 vssd1
port 730 nsew ground bidirectional
rlabel metal5 s 1104 117608 218868 118308 6 vssd1
port 731 nsew ground bidirectional
rlabel metal5 s 1104 108608 218868 109308 6 vssd1
port 732 nsew ground bidirectional
rlabel metal5 s 1104 99608 218868 100308 6 vssd1
port 733 nsew ground bidirectional
rlabel metal5 s 1104 90608 218868 91308 6 vssd1
port 734 nsew ground bidirectional
rlabel metal5 s 1104 81608 218868 82308 6 vssd1
port 735 nsew ground bidirectional
rlabel metal5 s 1104 72608 218868 73308 6 vssd1
port 736 nsew ground bidirectional
rlabel metal5 s 1104 63608 218868 64308 6 vssd1
port 737 nsew ground bidirectional
rlabel metal5 s 1104 54608 218868 55308 6 vssd1
port 738 nsew ground bidirectional
rlabel metal5 s 1104 45608 218868 46308 6 vssd1
port 739 nsew ground bidirectional
rlabel metal5 s 1104 36608 218868 37308 6 vssd1
port 740 nsew ground bidirectional
rlabel metal5 s 1104 27608 218868 28308 6 vssd1
port 741 nsew ground bidirectional
rlabel metal5 s 1104 18608 218868 19308 6 vssd1
port 742 nsew ground bidirectional
rlabel metal5 s 1104 9608 218868 10308 6 vssd1
port 743 nsew ground bidirectional
rlabel metal4 s 212058 -1164 212758 140972 6 vccd2
port 744 nsew power bidirectional
rlabel metal4 s 203058 -1164 203758 140972 6 vccd2
port 745 nsew power bidirectional
rlabel metal4 s 194058 91112 194758 140972 6 vccd2
port 746 nsew power bidirectional
rlabel metal4 s 185058 91112 185758 140972 6 vccd2
port 747 nsew power bidirectional
rlabel metal4 s 176058 91112 176758 140972 6 vccd2
port 748 nsew power bidirectional
rlabel metal4 s 167058 91112 167758 140972 6 vccd2
port 749 nsew power bidirectional
rlabel metal4 s 158058 91112 158758 140972 6 vccd2
port 750 nsew power bidirectional
rlabel metal4 s 149058 91112 149758 140972 6 vccd2
port 751 nsew power bidirectional
rlabel metal4 s 140058 91112 140758 140972 6 vccd2
port 752 nsew power bidirectional
rlabel metal4 s 131058 91112 131758 140972 6 vccd2
port 753 nsew power bidirectional
rlabel metal4 s 122058 91112 122758 140972 6 vccd2
port 754 nsew power bidirectional
rlabel metal4 s 113058 91112 113758 140972 6 vccd2
port 755 nsew power bidirectional
rlabel metal4 s 104058 91112 104758 140972 6 vccd2
port 756 nsew power bidirectional
rlabel metal4 s 95058 -1164 95758 140972 6 vccd2
port 757 nsew power bidirectional
rlabel metal4 s 86058 -1164 86758 140972 6 vccd2
port 758 nsew power bidirectional
rlabel metal4 s 77058 -1164 77758 140972 6 vccd2
port 759 nsew power bidirectional
rlabel metal4 s 68058 -1164 68758 140972 6 vccd2
port 760 nsew power bidirectional
rlabel metal4 s 59058 -1164 59758 140972 6 vccd2
port 761 nsew power bidirectional
rlabel metal4 s 50058 -1164 50758 140972 6 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 41058 -1164 41758 140972 6 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 32058 16744 32758 140972 6 vccd2
port 764 nsew power bidirectional
rlabel metal4 s 23058 16744 23758 140972 6 vccd2
port 765 nsew power bidirectional
rlabel metal4 s 14058 -1164 14758 140972 6 vccd2
port 766 nsew power bidirectional
rlabel metal4 s 5058 -1164 5758 140972 6 vccd2
port 767 nsew power bidirectional
rlabel metal4 s 194058 -1164 194758 21000 6 vccd2
port 768 nsew power bidirectional
rlabel metal4 s 185058 -1164 185758 21000 6 vccd2
port 769 nsew power bidirectional
rlabel metal4 s 176058 -1164 176758 21000 6 vccd2
port 770 nsew power bidirectional
rlabel metal4 s 167058 -1164 167758 21000 6 vccd2
port 771 nsew power bidirectional
rlabel metal4 s 158058 -1164 158758 21000 6 vccd2
port 772 nsew power bidirectional
rlabel metal4 s 149058 -1164 149758 21000 6 vccd2
port 773 nsew power bidirectional
rlabel metal4 s 140058 -1164 140758 21000 6 vccd2
port 774 nsew power bidirectional
rlabel metal4 s 131058 -1164 131758 21000 6 vccd2
port 775 nsew power bidirectional
rlabel metal4 s 122058 -1164 122758 21000 6 vccd2
port 776 nsew power bidirectional
rlabel metal4 s 113058 -1164 113758 21000 6 vccd2
port 777 nsew power bidirectional
rlabel metal4 s 104058 -1164 104758 21000 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 32058 -1164 32758 1000 8 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 23058 -1164 23758 1000 8 vccd2
port 780 nsew power bidirectional
rlabel metal5 s 1104 132196 218868 132896 6 vccd2
port 781 nsew power bidirectional
rlabel metal5 s 1104 123196 218868 123896 6 vccd2
port 782 nsew power bidirectional
rlabel metal5 s 1104 114196 218868 114896 6 vccd2
port 783 nsew power bidirectional
rlabel metal5 s 1104 105196 218868 105896 6 vccd2
port 784 nsew power bidirectional
rlabel metal5 s 1104 96196 218868 96896 6 vccd2
port 785 nsew power bidirectional
rlabel metal5 s 1104 87196 218868 87896 6 vccd2
port 786 nsew power bidirectional
rlabel metal5 s 1104 78196 218868 78896 6 vccd2
port 787 nsew power bidirectional
rlabel metal5 s 1104 69196 218868 69896 6 vccd2
port 788 nsew power bidirectional
rlabel metal5 s 1104 60196 218868 60896 6 vccd2
port 789 nsew power bidirectional
rlabel metal5 s 1104 51196 218868 51896 6 vccd2
port 790 nsew power bidirectional
rlabel metal5 s 1104 42196 218868 42896 6 vccd2
port 791 nsew power bidirectional
rlabel metal5 s 1104 33196 218868 33896 6 vccd2
port 792 nsew power bidirectional
rlabel metal5 s 1104 24196 218868 24896 6 vccd2
port 793 nsew power bidirectional
rlabel metal5 s 1104 15196 218868 15896 6 vccd2
port 794 nsew power bidirectional
rlabel metal5 s 1104 6196 218868 6896 6 vccd2
port 795 nsew power bidirectional
rlabel metal4 s 216558 -1164 217258 140972 6 vssd2
port 796 nsew ground bidirectional
rlabel metal4 s 207558 -1164 208258 140972 6 vssd2
port 797 nsew ground bidirectional
rlabel metal4 s 198558 91112 199258 140972 6 vssd2
port 798 nsew ground bidirectional
rlabel metal4 s 189558 91112 190258 140972 6 vssd2
port 799 nsew ground bidirectional
rlabel metal4 s 180558 91112 181258 140972 6 vssd2
port 800 nsew ground bidirectional
rlabel metal4 s 171558 91112 172258 140972 6 vssd2
port 801 nsew ground bidirectional
rlabel metal4 s 162558 91112 163258 140972 6 vssd2
port 802 nsew ground bidirectional
rlabel metal4 s 153558 91112 154258 140972 6 vssd2
port 803 nsew ground bidirectional
rlabel metal4 s 144558 91112 145258 140972 6 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 135558 91112 136258 140972 6 vssd2
port 805 nsew ground bidirectional
rlabel metal4 s 126558 91112 127258 140972 6 vssd2
port 806 nsew ground bidirectional
rlabel metal4 s 117558 91112 118258 140972 6 vssd2
port 807 nsew ground bidirectional
rlabel metal4 s 108558 91112 109258 140972 6 vssd2
port 808 nsew ground bidirectional
rlabel metal4 s 99558 91112 100258 140972 6 vssd2
port 809 nsew ground bidirectional
rlabel metal4 s 90558 -1164 91258 140972 6 vssd2
port 810 nsew ground bidirectional
rlabel metal4 s 81558 -1164 82258 140972 6 vssd2
port 811 nsew ground bidirectional
rlabel metal4 s 72558 -1164 73258 140972 6 vssd2
port 812 nsew ground bidirectional
rlabel metal4 s 63558 -1164 64258 140972 6 vssd2
port 813 nsew ground bidirectional
rlabel metal4 s 54558 -1164 55258 140972 6 vssd2
port 814 nsew ground bidirectional
rlabel metal4 s 45558 -1164 46258 140972 6 vssd2
port 815 nsew ground bidirectional
rlabel metal4 s 36558 16744 37258 140972 6 vssd2
port 816 nsew ground bidirectional
rlabel metal4 s 27558 16744 28258 140972 6 vssd2
port 817 nsew ground bidirectional
rlabel metal4 s 18558 16744 19258 140972 6 vssd2
port 818 nsew ground bidirectional
rlabel metal4 s 9558 -1164 10258 140972 6 vssd2
port 819 nsew ground bidirectional
rlabel metal4 s 198558 -1164 199258 21000 6 vssd2
port 820 nsew ground bidirectional
rlabel metal4 s 189558 -1164 190258 21000 6 vssd2
port 821 nsew ground bidirectional
rlabel metal4 s 180558 -1164 181258 21000 6 vssd2
port 822 nsew ground bidirectional
rlabel metal4 s 171558 -1164 172258 21000 6 vssd2
port 823 nsew ground bidirectional
rlabel metal4 s 162558 -1164 163258 21000 6 vssd2
port 824 nsew ground bidirectional
rlabel metal4 s 153558 -1164 154258 21000 6 vssd2
port 825 nsew ground bidirectional
rlabel metal4 s 144558 -1164 145258 21000 6 vssd2
port 826 nsew ground bidirectional
rlabel metal4 s 135558 -1164 136258 21000 6 vssd2
port 827 nsew ground bidirectional
rlabel metal4 s 126558 -1164 127258 21000 6 vssd2
port 828 nsew ground bidirectional
rlabel metal4 s 117558 -1164 118258 21000 6 vssd2
port 829 nsew ground bidirectional
rlabel metal4 s 108558 -1164 109258 21000 6 vssd2
port 830 nsew ground bidirectional
rlabel metal4 s 99558 -1164 100258 21000 6 vssd2
port 831 nsew ground bidirectional
rlabel metal4 s 36558 -1164 37258 1000 8 vssd2
port 832 nsew ground bidirectional
rlabel metal4 s 27558 -1164 28258 1000 8 vssd2
port 833 nsew ground bidirectional
rlabel metal4 s 18558 -1164 19258 1000 8 vssd2
port 834 nsew ground bidirectional
rlabel metal5 s 1104 127696 218868 128396 6 vssd2
port 835 nsew ground bidirectional
rlabel metal5 s 1104 118696 218868 119396 6 vssd2
port 836 nsew ground bidirectional
rlabel metal5 s 1104 109696 218868 110396 6 vssd2
port 837 nsew ground bidirectional
rlabel metal5 s 1104 100696 218868 101396 6 vssd2
port 838 nsew ground bidirectional
rlabel metal5 s 1104 91696 218868 92396 6 vssd2
port 839 nsew ground bidirectional
rlabel metal5 s 1104 82696 218868 83396 6 vssd2
port 840 nsew ground bidirectional
rlabel metal5 s 1104 73696 218868 74396 6 vssd2
port 841 nsew ground bidirectional
rlabel metal5 s 1104 64696 218868 65396 6 vssd2
port 842 nsew ground bidirectional
rlabel metal5 s 1104 55696 218868 56396 6 vssd2
port 843 nsew ground bidirectional
rlabel metal5 s 1104 46696 218868 47396 6 vssd2
port 844 nsew ground bidirectional
rlabel metal5 s 1104 37696 218868 38396 6 vssd2
port 845 nsew ground bidirectional
rlabel metal5 s 1104 28696 218868 29396 6 vssd2
port 846 nsew ground bidirectional
rlabel metal5 s 1104 19696 218868 20396 6 vssd2
port 847 nsew ground bidirectional
rlabel metal5 s 1104 10696 218868 11396 6 vssd2
port 848 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 140000
string LEFview TRUE
string GDS_FILE /project/openlane/adc_wrapper/runs/adc_wrapper/results/magic/adc_wrapper.gds
string GDS_END 13482398
string GDS_START 520188
<< end >>

