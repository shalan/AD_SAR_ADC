VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ACMP
  CLASS BLOCK ;
  FOREIGN ACMP ;
  ORIGIN 0.000 0.000 ;
  SIZE 62.820 BY 72.380 ;
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.630 35.380 53.130 36.500 ;
    END
  END INN
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.630 15.600 53.130 16.720 ;
    END
  END INP
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.630 55.160 53.130 56.280 ;
    END
  END Q
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.130 55.160 15.630 56.280 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.130 35.380 15.630 36.500 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.130 15.600 15.630 16.720 ;
    END
  END clk
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 40.235 0.000 42.335 72.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 30.580 0.000 32.680 72.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 20.925 0.000 23.025 72.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 56.520 4.000 58.820 68.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 4.000 4.000 6.300 68.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 4.000 66.080 58.820 68.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.875 62.820 49.675 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.130 62.820 36.930 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.385 62.820 24.185 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 4.000 4.000 58.820 6.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 60.520 0.000 62.820 72.380 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 35.405 0.000 37.505 72.380 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 25.755 0.000 27.855 72.380 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.000 2.300 72.380 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 62.820 72.380 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.505 62.820 43.305 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.755 62.820 30.555 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 62.820 2.300 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 17.150 17.065 45.670 55.315 ;
      LAYER met1 ;
        RECT 16.760 16.910 46.980 55.470 ;
      LAYER met2 ;
        RECT 15.630 56.560 20.645 72.380 ;
        RECT 15.910 54.880 20.645 56.560 ;
        RECT 15.630 36.780 20.645 54.880 ;
        RECT 15.910 35.100 20.645 36.780 ;
        RECT 15.630 17.000 20.645 35.100 ;
        RECT 15.910 15.320 20.645 17.000 ;
        RECT 15.630 0.000 20.645 15.320 ;
        RECT 23.305 0.000 25.475 72.380 ;
        RECT 28.135 0.000 30.300 72.380 ;
        RECT 32.960 0.000 35.125 72.380 ;
        RECT 37.785 0.000 39.955 72.380 ;
        RECT 42.615 56.560 47.630 72.380 ;
        RECT 42.615 54.880 47.350 56.560 ;
        RECT 42.615 36.780 47.630 54.880 ;
        RECT 42.615 35.100 47.350 36.780 ;
        RECT 42.615 17.000 47.630 35.100 ;
        RECT 42.615 15.320 47.350 17.000 ;
        RECT 42.615 0.000 47.630 15.320 ;
      LAYER met3 ;
        RECT 0.000 41.500 62.820 41.505 ;
        RECT 0.000 37.330 62.820 41.105 ;
        RECT 0.000 30.955 62.820 34.730 ;
        RECT 0.000 24.585 62.820 28.355 ;
        RECT 0.000 22.380 62.820 22.385 ;
  END
END ACMP
END LIBRARY

