magic
tech sky130A
magscale 1 2
timestamp 1626198473
<< checkpaint >>
rect -1260 -6322 101104 56510
<< locali >>
rect 45770 51554 90780 51562
rect 95360 51554 96184 51558
rect 45770 51520 96184 51554
rect 45770 51370 45824 51520
rect 95364 51516 96184 51520
rect 45770 51336 45777 51370
rect 45811 51336 45824 51370
rect 45770 51326 45824 51336
rect 96148 51466 96184 51516
rect 21190 51278 21746 51280
rect 21190 51274 37460 51278
rect 20370 51272 37460 51274
rect 20370 51255 48154 51272
rect 20370 51230 20399 51255
rect 20372 51221 20399 51230
rect 20433 51234 48154 51255
rect 20433 51230 21390 51234
rect 20433 51221 20452 51230
rect 20372 51210 20452 51221
rect 45768 51190 45818 51196
rect 45768 51156 45777 51190
rect 45811 51156 45818 51190
rect 796 50625 854 50672
rect 796 50591 811 50625
rect 845 50591 854 50625
rect 796 50586 854 50591
rect 808 50451 844 50452
rect 808 50417 809 50451
rect 843 50417 844 50451
rect 808 50416 844 50417
rect 20382 50411 20456 50432
rect 20382 50377 20399 50411
rect 20433 50377 20456 50411
rect 20382 49560 20456 50377
rect 45768 49816 45818 51156
rect 48098 50662 48154 51234
rect 48092 50643 48158 50662
rect 48092 50609 48111 50643
rect 48145 50609 48158 50643
rect 48092 50594 48158 50609
rect 48098 50590 48154 50594
rect 48114 50441 48158 50446
rect 48114 50407 48119 50441
rect 48153 50407 48158 50441
rect 48114 50402 48158 50407
rect 20380 26192 20460 49560
rect 45768 27474 45816 49816
rect 96148 49202 96190 51466
rect 96146 27622 96190 49202
rect 96146 27580 96196 27622
rect 43122 26731 43162 27404
rect 43122 26697 43124 26731
rect 43158 26697 43162 26731
rect 43122 26682 43162 26697
rect 90376 26755 90468 27392
rect 90376 26721 90401 26755
rect 90435 26721 90468 26755
rect 90376 26658 90468 26721
rect 43110 26517 43164 26526
rect 43110 26483 43120 26517
rect 43154 26483 43164 26517
rect 43110 26472 43164 26483
rect 20380 26162 20466 26192
rect 20386 2810 20466 26162
rect 43116 25406 43164 26472
rect 43110 24386 43164 25406
rect 43102 23928 43164 24386
rect 90376 26401 90434 26460
rect 90376 26367 90389 26401
rect 90423 26367 90434 26401
rect 20386 2312 20472 2810
rect 20382 2288 20472 2312
rect 20382 1880 20468 2288
rect 20600 2184 20702 2358
rect 20776 1880 20878 1974
rect 20382 1790 20884 1880
rect 20386 1788 20884 1790
rect 21292 -1170 21352 48
rect 24370 -1026 24430 192
rect 27710 -818 27770 440
rect 31104 -636 31164 734
rect 34346 -442 34406 1020
rect 37808 -300 37868 1456
rect 43102 1292 43154 23928
rect 67809 2339 68298 2354
rect 67809 2246 67830 2339
rect 68285 2280 68298 2339
rect 68286 2246 68298 2280
rect 67809 2221 68298 2246
rect 43092 -108 43158 1292
rect 48502 39 48572 54
rect 78542 50 78638 662
rect 81690 52 81788 1002
rect 85120 432 85182 1398
rect 85120 98 85190 432
rect 85120 72 85202 98
rect 85126 70 85202 72
rect 48502 5 48523 39
rect 48557 5 48572 39
rect 48502 -10 48572 5
rect 78540 23 78640 50
rect 78540 -11 78570 23
rect 78604 -11 78640 23
rect 81688 16 81790 52
rect 81688 8 81722 16
rect 78540 -38 78640 -11
rect 81690 -18 81722 8
rect 81756 8 81790 16
rect 85126 36 85142 70
rect 85176 36 85202 70
rect 85126 8 85202 36
rect 81756 -18 81788 8
rect 85126 -4 85190 8
rect 78542 -44 78638 -38
rect 81690 -48 81788 -18
rect 88292 -102 89642 -98
rect 90376 -102 90434 26367
rect 93032 26096 93112 27534
rect 96150 27322 96196 27580
rect 96320 27036 96520 27052
rect 96320 27002 96331 27036
rect 96365 27002 96520 27036
rect 96320 26988 96520 27002
rect 93930 26894 93980 26922
rect 93930 26860 93967 26894
rect 93930 26830 93980 26860
rect 96172 26364 96214 26570
rect 96172 26120 96218 26364
rect 96172 26100 96212 26120
rect 93540 26096 96212 26100
rect 93032 26030 96212 26096
rect 93032 26026 93562 26030
rect 88292 -108 90434 -102
rect 43090 -120 90434 -108
rect 43090 -154 44167 -120
rect 44201 -154 44219 -120
rect 44253 -154 44269 -120
rect 44303 -154 44321 -120
rect 44355 -154 90434 -120
rect 43090 -168 90434 -154
rect 43090 -172 85110 -168
rect 85226 -172 90434 -168
rect 43090 -186 43236 -172
rect 88292 -184 90434 -172
rect 85120 -264 85182 -238
rect 85120 -298 85134 -264
rect 85168 -272 85182 -264
rect 85168 -298 85194 -272
rect 37800 -304 63320 -300
rect 85120 -304 85194 -298
rect 37800 -316 85194 -304
rect 37800 -350 38678 -316
rect 38712 -350 38730 -316
rect 38764 -350 38780 -316
rect 38814 -350 38832 -316
rect 38866 -350 85194 -316
rect 37800 -362 85194 -350
rect 37800 -366 85178 -362
rect 37800 -372 63320 -366
rect 37808 -380 37868 -372
rect 34350 -468 34406 -442
rect 81688 -460 81790 -420
rect 44280 -462 81790 -460
rect 44280 -464 81724 -462
rect 39300 -468 81724 -464
rect 34350 -481 81724 -468
rect 34350 -515 35133 -481
rect 35167 -515 35185 -481
rect 35219 -515 35235 -481
rect 35269 -515 35287 -481
rect 35321 -496 81724 -481
rect 81758 -464 81790 -462
rect 81758 -496 81788 -464
rect 35321 -515 81788 -496
rect 34350 -520 81788 -515
rect 34350 -524 81758 -520
rect 34350 -528 70790 -524
rect 34350 -532 44304 -528
rect 34350 -534 39342 -532
rect 34448 -536 39342 -534
rect 31098 -644 36684 -636
rect 42164 -644 57422 -640
rect 31098 -648 65052 -644
rect 31098 -649 72694 -648
rect 31098 -683 31517 -649
rect 31551 -683 31569 -649
rect 31603 -683 31619 -649
rect 31653 -683 31671 -649
rect 31705 -660 72694 -649
rect 78542 -660 78638 -652
rect 31705 -675 78638 -660
rect 31705 -683 78574 -675
rect 31098 -696 78574 -683
rect 31104 -704 31164 -696
rect 36646 -704 78574 -696
rect 42164 -709 78574 -704
rect 78608 -709 78638 -675
rect 42164 -712 78638 -709
rect 57366 -716 78638 -712
rect 65008 -720 78638 -716
rect 78534 -730 78638 -720
rect 27698 -822 33728 -818
rect 27698 -829 75364 -822
rect 27698 -863 27851 -829
rect 27885 -863 27903 -829
rect 27937 -863 27953 -829
rect 27987 -863 28005 -829
rect 28039 -835 75364 -829
rect 28039 -863 75311 -835
rect 27698 -869 75311 -863
rect 75345 -866 75364 -835
rect 75345 -869 75362 -866
rect 27698 -876 75362 -869
rect 27710 -886 27770 -876
rect 75290 -884 75362 -876
rect 71794 -1026 71862 -1022
rect 24370 -1028 71862 -1026
rect 24370 -1030 71812 -1028
rect 24370 -1064 24779 -1030
rect 24813 -1064 24831 -1030
rect 24865 -1064 24881 -1030
rect 24915 -1064 24933 -1030
rect 24967 -1062 71812 -1030
rect 71846 -1062 71862 -1028
rect 24967 -1064 58626 -1062
rect 24370 -1068 58626 -1064
rect 24370 -1070 39590 -1068
rect 71794 -1072 71862 -1062
rect 46996 -1170 48574 -1160
rect 21286 -1172 27752 -1170
rect 40626 -1172 48574 -1170
rect 21286 -1177 48574 -1172
rect 21286 -1182 48521 -1177
rect 21286 -1216 21306 -1182
rect 21340 -1216 21358 -1182
rect 21392 -1216 21408 -1182
rect 21442 -1216 21460 -1182
rect 21494 -1211 48521 -1182
rect 48555 -1211 48574 -1177
rect 21494 -1216 48574 -1211
rect 21286 -1224 48574 -1216
rect 21286 -1230 47092 -1224
rect 21424 -1232 26450 -1230
rect 27734 -1232 40650 -1230
<< viali >>
rect 45777 51336 45811 51370
rect 20399 51221 20433 51255
rect 45777 51156 45811 51190
rect 811 50591 845 50625
rect 809 50417 843 50451
rect 20399 50377 20433 50411
rect 48111 50609 48145 50643
rect 48119 50407 48153 50441
rect 43124 26697 43158 26731
rect 90401 26721 90435 26755
rect 43120 26483 43154 26517
rect 90389 26367 90423 26401
rect 67830 2280 68285 2339
rect 67830 2246 68286 2280
rect 48523 5 48557 39
rect 78570 -11 78604 23
rect 81722 -18 81756 16
rect 85142 36 85176 70
rect 96331 27002 96365 27036
rect 93967 26860 94001 26894
rect 44167 -154 44201 -120
rect 44219 -154 44253 -120
rect 44269 -154 44303 -120
rect 44321 -154 44355 -120
rect 85134 -298 85168 -264
rect 38678 -350 38712 -316
rect 38730 -350 38764 -316
rect 38780 -350 38814 -316
rect 38832 -350 38866 -316
rect 35133 -515 35167 -481
rect 35185 -515 35219 -481
rect 35235 -515 35269 -481
rect 35287 -515 35321 -481
rect 81724 -496 81758 -462
rect 31517 -683 31551 -649
rect 31569 -683 31603 -649
rect 31619 -683 31653 -649
rect 31671 -683 31705 -649
rect 78574 -709 78608 -675
rect 27851 -863 27885 -829
rect 27903 -863 27937 -829
rect 27953 -863 27987 -829
rect 28005 -863 28039 -829
rect 75311 -869 75345 -835
rect 24779 -1064 24813 -1030
rect 24831 -1064 24865 -1030
rect 24881 -1064 24915 -1030
rect 24933 -1064 24967 -1030
rect 71812 -1062 71846 -1028
rect 21306 -1216 21340 -1182
rect 21358 -1216 21392 -1182
rect 21408 -1216 21442 -1182
rect 21460 -1216 21494 -1182
rect 48521 -1211 48555 -1177
<< metal1 >>
rect 45766 51372 45824 51384
rect 45764 51370 45824 51372
rect 45764 51336 45777 51370
rect 45811 51336 45824 51370
rect 45764 51326 45824 51336
rect 20376 51255 20450 51276
rect 20376 51221 20399 51255
rect 20433 51221 20450 51255
rect 625 50959 1053 50980
rect 625 50792 634 50959
rect 803 50958 1053 50959
rect 625 50791 806 50792
rect 1031 50791 1053 50958
rect 625 50785 1053 50791
rect 796 50625 854 50785
rect 796 50591 811 50625
rect 845 50591 854 50625
rect 796 50451 854 50591
rect 796 50417 809 50451
rect 843 50417 854 50451
rect 796 50404 854 50417
rect 20376 50411 20450 51221
rect 45768 51192 45822 51326
rect 45766 51190 45822 51192
rect 45766 51156 45777 51190
rect 45811 51156 45822 51190
rect 45766 51140 45822 51156
rect 48092 50658 48158 50662
rect 48092 50643 48168 50658
rect 48092 50609 48111 50643
rect 48145 50609 48168 50643
rect 48092 50594 48168 50609
rect 48100 50456 48168 50594
rect 20376 50377 20399 50411
rect 20433 50377 20450 50411
rect 48098 50441 48168 50456
rect 48098 50407 48119 50441
rect 48153 50412 48168 50441
rect 48153 50407 48164 50412
rect 48098 50388 48164 50407
rect 20376 50358 20450 50377
rect 94792 27354 94880 27366
rect 94792 27302 94825 27354
rect 94877 27302 94880 27354
rect 94792 27290 94880 27302
rect 96320 27047 96658 27053
rect 96320 27036 96390 27047
rect 96320 27002 96331 27036
rect 96365 27002 96390 27036
rect 96320 26995 96390 27002
rect 96572 26995 96573 27047
rect 96625 26995 96658 27047
rect 96320 26987 96658 26995
rect 96320 26986 96386 26987
rect 93703 26902 94020 26922
rect 93703 26850 93710 26902
rect 93813 26894 94020 26902
rect 93813 26860 93967 26894
rect 94001 26860 94020 26894
rect 93813 26850 94020 26860
rect 93703 26827 94020 26850
rect 43116 26742 43162 26758
rect 90362 26755 90468 26792
rect 43116 26731 43164 26742
rect 43116 26697 43124 26731
rect 43158 26697 43164 26731
rect 43116 26686 43164 26697
rect 90362 26721 90401 26755
rect 90435 26721 90468 26755
rect 43116 26526 43162 26686
rect 43110 26517 43162 26526
rect 43110 26483 43120 26517
rect 43154 26483 43162 26517
rect 43110 26472 43162 26483
rect 43116 26470 43162 26472
rect 90362 26401 90468 26721
rect 94048 26578 94160 26630
rect 94048 26526 94073 26578
rect 94125 26526 94160 26578
rect 94048 26492 94160 26526
rect 90362 26367 90389 26401
rect 90423 26367 90468 26401
rect 90362 26340 90468 26367
rect 67808 2339 68300 2411
rect 67808 2246 67830 2339
rect 68285 2280 68300 2339
rect 68286 2246 68300 2280
rect 48502 46 48572 54
rect 48502 39 48574 46
rect 48502 5 48523 39
rect 48557 5 48574 39
rect 48502 -10 48574 5
rect 44152 -120 44376 -99
rect 44152 -154 44167 -120
rect 44201 -154 44219 -120
rect 44253 -154 44269 -120
rect 44303 -154 44321 -120
rect 44355 -154 44376 -120
rect 38663 -316 38887 -300
rect 38663 -350 38678 -316
rect 38712 -350 38730 -316
rect 38764 -350 38780 -316
rect 38814 -350 38832 -316
rect 38866 -350 38887 -316
rect 35118 -481 35342 -468
rect 35118 -515 35133 -481
rect 35167 -515 35185 -481
rect 35219 -515 35235 -481
rect 35269 -515 35287 -481
rect 35321 -515 35342 -481
rect 31501 -649 31725 -636
rect 31501 -683 31517 -649
rect 31551 -683 31569 -649
rect 31603 -683 31619 -649
rect 31653 -683 31671 -649
rect 31705 -683 31725 -649
rect 27829 -829 28053 -818
rect 27829 -863 27851 -829
rect 27885 -863 27903 -829
rect 27937 -863 27953 -829
rect 27987 -863 28005 -829
rect 28039 -863 28053 -829
rect 24766 -1030 24990 -1020
rect 24766 -1064 24779 -1030
rect 24813 -1064 24831 -1030
rect 24865 -1064 24881 -1030
rect 24915 -1064 24933 -1030
rect 24967 -1064 24990 -1030
rect 21287 -1182 21511 -1170
rect 21287 -1216 21306 -1182
rect 21340 -1216 21358 -1182
rect 21392 -1216 21408 -1182
rect 21442 -1216 21460 -1182
rect 21494 -1216 21511 -1182
rect 21287 -2825 21511 -1216
rect 21287 -2992 21314 -2825
rect 21483 -2992 21511 -2825
rect 21287 -3006 21511 -2992
rect 24766 -2825 24990 -1064
rect 24766 -2992 24793 -2825
rect 24962 -2992 24990 -2825
rect 24766 -3006 24990 -2992
rect 27829 -2826 28053 -863
rect 27829 -2993 27856 -2826
rect 28025 -2993 28053 -2826
rect 27829 -3007 28053 -2993
rect 31501 -2826 31725 -683
rect 31501 -2993 31528 -2826
rect 31697 -2993 31725 -2826
rect 31501 -3007 31725 -2993
rect 35118 -2827 35342 -515
rect 35118 -2994 35145 -2827
rect 35314 -2994 35342 -2827
rect 35118 -3008 35342 -2994
rect 38663 -2827 38887 -350
rect 38663 -2994 38690 -2827
rect 38859 -2994 38887 -2827
rect 38663 -3008 38887 -2994
rect 44152 -2826 44376 -154
rect 48512 -1162 48574 -10
rect 48506 -1177 48574 -1162
rect 48506 -1211 48521 -1177
rect 48555 -1211 48574 -1177
rect 48506 -1224 48574 -1211
rect 44152 -2993 44179 -2826
rect 44348 -2993 44376 -2826
rect 44152 -3007 44376 -2993
rect 67808 -2848 68300 2246
rect 71798 -1022 71858 172
rect 75288 -780 75364 436
rect 85122 98 85186 126
rect 85122 70 85202 98
rect 78540 23 78640 50
rect 78540 -11 78570 23
rect 78604 -11 78640 23
rect 81688 42 81790 52
rect 81688 16 81792 42
rect 81688 8 81722 16
rect 78540 -38 78640 -11
rect 81694 -18 81722 8
rect 81756 -18 81792 16
rect 78542 -675 78638 -38
rect 81694 -462 81792 -18
rect 85122 36 85142 70
rect 85176 36 85202 70
rect 85122 8 85202 36
rect 85122 -206 85186 8
rect 85114 -264 85186 -206
rect 85114 -298 85134 -264
rect 85168 -272 85186 -264
rect 85168 -298 85194 -272
rect 85114 -362 85194 -298
rect 85114 -378 85178 -362
rect 81694 -496 81724 -462
rect 81758 -496 81792 -462
rect 81694 -534 81792 -496
rect 78542 -692 78574 -675
rect 78540 -709 78574 -692
rect 78608 -709 78638 -675
rect 78540 -730 78638 -709
rect 75288 -822 75360 -780
rect 75288 -835 75364 -822
rect 75288 -869 75311 -835
rect 75345 -866 75364 -835
rect 75345 -869 75362 -866
rect 75288 -872 75362 -869
rect 75290 -884 75362 -872
rect 71794 -1028 71862 -1022
rect 71794 -1062 71812 -1028
rect 71846 -1062 71862 -1028
rect 71794 -1072 71862 -1062
rect 67808 -3006 67823 -2848
rect 67875 -2849 68300 -2848
rect 67932 -2850 68053 -2849
rect 68105 -2850 68300 -2849
rect 67808 -3007 67880 -3006
rect 68039 -3007 68053 -2850
rect 68269 -3007 68300 -2850
rect 67808 -3009 68300 -3007
<< via1 >>
rect 634 50958 803 50959
rect 634 50792 1031 50958
rect 806 50791 1031 50792
rect 94825 27302 94877 27354
rect 96390 26995 96572 27047
rect 96573 26995 96625 27047
rect 93710 26850 93813 26902
rect 94073 26526 94125 26578
rect 21314 -2992 21483 -2825
rect 24793 -2992 24962 -2825
rect 27856 -2993 28025 -2826
rect 31528 -2993 31697 -2826
rect 35145 -2994 35314 -2827
rect 38690 -2994 38859 -2827
rect 44179 -2993 44348 -2826
rect 67823 -2849 67875 -2848
rect 67823 -2850 67932 -2849
rect 68053 -2850 68105 -2849
rect 67823 -3006 68039 -2850
rect 67880 -3007 68039 -3006
rect 68053 -3007 68269 -2850
<< metal2 >>
rect 759 54471 937 55250
rect 625 50959 1053 54471
rect 625 50792 634 50959
rect 803 50958 1053 50959
rect 625 50791 806 50792
rect 1031 50791 1053 50958
rect 24290 50910 25152 50920
rect 24290 50906 58282 50910
rect 24290 50854 58400 50906
rect 24290 50850 58282 50854
rect 25120 50848 58282 50850
rect 625 50785 1053 50791
rect 94810 27436 94880 27446
rect 94810 27380 94816 27436
rect 94872 27380 94880 27436
rect 94810 27354 94880 27380
rect 94810 27302 94825 27354
rect 94877 27302 94880 27354
rect 94810 27292 94880 27302
rect 96320 27048 97000 27053
rect 96320 27047 96619 27048
rect 96675 27047 97000 27048
rect 96320 26995 96390 27047
rect 96572 26995 96573 27047
rect 96320 26992 96619 26995
rect 96675 26992 96682 27047
rect 96320 26991 96682 26992
rect 96738 26991 96741 27047
rect 96852 26991 96854 27047
rect 96966 26991 97000 27047
rect 96320 26987 97000 26991
rect 93584 26903 93820 26922
rect 93584 26902 93658 26903
rect 93714 26902 93719 26903
rect 93775 26902 93820 26903
rect 93584 26846 93594 26902
rect 93650 26847 93658 26902
rect 93813 26850 93820 26902
rect 93714 26847 93719 26850
rect 93775 26847 93820 26850
rect 93650 26846 93820 26847
rect 93584 26827 93820 26846
rect 93934 26586 94146 26592
rect 93914 26578 94146 26586
rect 93914 26526 94073 26578
rect 94125 26526 94146 26578
rect 93914 26500 94146 26526
rect 93914 26240 93954 26500
rect 91012 26238 93958 26240
rect 90500 26202 93958 26238
rect 90500 26200 92030 26202
rect 90500 26198 91014 26200
rect 21288 -2825 21509 -2797
rect 21288 -2992 21314 -2825
rect 21483 -2992 21509 -2825
rect 21288 -3893 21509 -2992
rect 24767 -2825 24988 -2797
rect 24767 -2992 24793 -2825
rect 24962 -2992 24988 -2825
rect 24767 -3893 24988 -2992
rect 27830 -2826 28051 -2798
rect 27830 -2993 27856 -2826
rect 28025 -2993 28051 -2826
rect 27830 -3893 28051 -2993
rect 31502 -2826 31723 -2798
rect 31502 -2993 31528 -2826
rect 31697 -2993 31723 -2826
rect 31502 -3893 31723 -2993
rect 35119 -2827 35340 -2799
rect 35119 -2994 35145 -2827
rect 35314 -2994 35340 -2827
rect 35119 -3893 35340 -2994
rect 38664 -2827 38885 -2799
rect 38664 -2994 38690 -2827
rect 38859 -2994 38885 -2827
rect 38664 -3893 38885 -2994
rect 44153 -2826 44374 -2798
rect 44153 -2993 44179 -2826
rect 44348 -2993 44374 -2826
rect 44153 -3893 44374 -2993
rect 67808 -2848 68300 -2844
rect 67808 -3006 67823 -2848
rect 67875 -2849 68300 -2848
rect 67932 -2850 68053 -2849
rect 68105 -2850 68300 -2849
rect 67808 -3007 67880 -3006
rect 68039 -3007 68053 -2850
rect 68269 -3007 68300 -2850
rect 67808 -3890 68300 -3007
rect 21343 -4262 21458 -3893
rect 24820 -4262 24935 -3893
rect 21342 -5062 21458 -4262
rect 24819 -5062 24935 -4262
rect 27876 -5062 27992 -3893
rect 31555 -5062 31671 -3893
rect 35169 -5062 35285 -3893
rect 38704 -5062 38820 -3893
rect 44192 -5062 44308 -3893
rect 67957 -5062 68073 -3890
<< via2 >>
rect 11050 50850 11106 50906
rect 11112 50850 11168 50906
rect 11172 50850 11228 50906
rect 11234 50850 11290 50906
rect 11299 50850 11355 50906
rect 11361 50850 11417 50906
rect 11421 50850 11477 50906
rect 11483 50850 11539 50906
rect 11552 50850 11608 50906
rect 11614 50850 11670 50906
rect 11674 50850 11730 50906
rect 11736 50850 11792 50906
rect 11801 50850 11857 50906
rect 11863 50850 11919 50906
rect 11923 50850 11979 50906
rect 11985 50850 12041 50906
rect 94816 27380 94872 27436
rect 96619 27047 96675 27048
rect 96619 26995 96625 27047
rect 96625 26995 96675 27047
rect 96619 26992 96675 26995
rect 96682 26991 96738 27047
rect 96741 26991 96852 27047
rect 96854 26991 96966 27047
rect 93658 26902 93714 26903
rect 93719 26902 93775 26903
rect 93594 26846 93650 26902
rect 93658 26850 93710 26902
rect 93710 26850 93714 26902
rect 93719 26850 93775 26902
rect 93658 26847 93714 26850
rect 93719 26847 93775 26850
<< metal3 >>
rect 11020 51384 12070 51401
rect 11020 51383 11883 51384
rect 11020 51382 11818 51383
rect 11020 51381 11740 51382
rect 11020 51380 11609 51381
rect 11020 51379 11473 51380
rect 11020 51378 11408 51379
rect 11020 51377 11330 51378
rect 11020 51376 11194 51377
rect 11020 51307 11050 51376
rect 12018 51320 12070 51384
rect 11020 51240 11049 51307
rect 12017 51251 12070 51320
rect 11020 51176 11048 51240
rect 12016 51184 12070 51251
rect 11880 51183 12070 51184
rect 11802 51182 12070 51183
rect 11737 51181 12070 51182
rect 11606 51180 12070 51181
rect 11470 51179 12070 51180
rect 11392 51178 12070 51179
rect 11327 51177 12070 51178
rect 11191 51176 12070 51177
rect 11020 50906 12070 51176
rect 11020 50850 11050 50906
rect 11106 50850 11112 50906
rect 11168 50850 11172 50906
rect 11228 50850 11234 50906
rect 11290 50850 11299 50906
rect 11355 50850 11361 50906
rect 11417 50850 11421 50906
rect 11477 50850 11483 50906
rect 11539 50850 11552 50906
rect 11608 50850 11614 50906
rect 11670 50850 11674 50906
rect 11730 50850 11736 50906
rect 11792 50850 11801 50906
rect 11857 50850 11863 50906
rect 11919 50850 11923 50906
rect 11979 50850 11985 50906
rect 12041 50850 12070 50906
rect 11020 50840 12070 50850
rect 94810 27530 94890 27538
rect 94810 27466 94820 27530
rect 94884 27466 94890 27530
rect 94810 27456 94890 27466
rect 94810 27436 94880 27456
rect 94810 27380 94816 27436
rect 94872 27380 94880 27436
rect 94810 27372 94880 27380
rect 96515 27119 99401 28249
rect 96515 27048 99844 27119
rect 96515 26992 96619 27048
rect 96675 27047 99844 27048
rect 96675 26992 96682 27047
rect 96515 26991 96682 26992
rect 96738 26991 96741 27047
rect 96852 26991 96854 27047
rect 96966 26991 99844 27047
rect 96515 26959 99844 26991
rect 93584 26903 93817 26922
rect 93584 26902 93658 26903
rect 93584 26846 93594 26902
rect 93650 26847 93658 26902
rect 93714 26847 93719 26903
rect 93775 26847 93817 26903
rect 93650 26846 93817 26847
rect 93584 25195 93817 26846
rect 96515 25989 99401 26959
rect 93584 24952 99416 25195
rect 93584 24792 99844 24952
rect 93584 24621 99416 24792
rect 93584 24620 93817 24621
<< via3 >>
rect 11883 51383 12018 51384
rect 11818 51382 12018 51383
rect 11740 51381 12018 51382
rect 11609 51380 12018 51381
rect 11473 51379 12018 51380
rect 11408 51378 12018 51379
rect 11330 51377 12018 51378
rect 11194 51376 12018 51377
rect 11050 51320 12018 51376
rect 11050 51307 12017 51320
rect 11049 51251 12017 51307
rect 11049 51240 12016 51251
rect 11048 51184 12016 51240
rect 11048 51183 11880 51184
rect 11048 51182 11802 51183
rect 11048 51181 11737 51182
rect 11048 51180 11606 51181
rect 11048 51179 11470 51180
rect 11048 51178 11392 51179
rect 11048 51177 11327 51178
rect 11048 51176 11191 51177
rect 94820 27466 94884 27530
<< metal4 >>
rect 2836 50319 3900 55249
rect 11006 51384 12070 55250
rect 23762 51496 49764 51500
rect 22752 51434 49764 51496
rect 22752 51432 23808 51434
rect 11006 51383 11883 51384
rect 11006 51382 11818 51383
rect 11006 51381 11740 51382
rect 11006 51380 11609 51381
rect 11006 51379 11473 51380
rect 11006 51378 11408 51379
rect 11006 51377 11330 51378
rect 11006 51376 11194 51377
rect 11006 51307 11050 51376
rect 12018 51320 12070 51384
rect 11006 51240 11049 51307
rect 12017 51251 12070 51320
rect 11006 51176 11048 51240
rect 12016 51184 12070 51251
rect 11880 51183 12070 51184
rect 11802 51182 12070 51183
rect 11737 51181 12070 51182
rect 11606 51180 12070 51181
rect 11470 51179 12070 51180
rect 11392 51178 12070 51179
rect 11327 51177 12070 51178
rect 11191 51176 12070 51177
rect 11006 51139 12070 51176
rect 22764 50622 22848 51432
rect 49692 50314 49762 51434
rect 91334 28070 94890 28140
rect 94816 27590 94890 28070
rect 94810 27584 94890 27590
rect 94810 27530 94888 27584
rect 94810 27466 94820 27530
rect 94884 27466 94888 27530
rect 94810 27460 94888 27466
use res250_layout  res250_layout_0
timestamp 1626198473
transform 1 0 20392 0 1 2302
box 202 -342 510 -90
use 7bitdac_layout  7bitdac_layout_1
timestamp 1626198473
transform 1 0 252 0 1 2456
box -252 -2456 45562 48686
use 7bitdac_layout  7bitdac_layout_0
timestamp 1626198473
transform 1 0 47558 0 1 2444
box -252 -2456 45562 48686
use switch_layout  switch_layout_0
timestamp 1626198473
transform 1 0 93914 0 1 26310
box 40 154 2460 1180
<< labels >>
rlabel locali s 20652 2264 20652 2264 4 x1_vref5
port 1 nsew
rlabel locali s 20812 1868 20812 1868 4 x2_vref1
port 2 nsew
rlabel locali s 804 50664 804 50664 4 inp1
port 3 nsew
rlabel locali s 67994 2294 67994 2294 4 inp2
port 4 nsew
rlabel locali s 93952 26862 93952 26862 4 d7
port 5 nsew
rlabel locali s 96452 27014 96452 27014 4 out_v
port 6 nsew
rlabel locali s 96176 27544 96176 27544 4 x1_out_v
port 7 nsew
rlabel locali s 96200 26388 96200 26388 4 x2_out_v
port 8 nsew
rlabel locali s 43126 44 43126 44 4 d6
port 9 nsew
rlabel locali s 37842 -218 37842 -218 4 d5
port 10 nsew
rlabel locali s 34364 612 34364 612 4 d4
port 11 nsew
rlabel locali s 31132 486 31132 486 4 d3
port 12 nsew
rlabel locali s 27736 152 27736 152 4 d2
port 13 nsew
rlabel locali s 24396 40 24396 40 4 d1
port 14 nsew
rlabel locali s 21316 -64 21316 -64 4 d0
port 15 nsew
rlabel metal4 s 2836 50319 3900 55249 4 vdd
port 16 nsew
rlabel metal4 s 11006 51139 12070 55250 4 gnd
port 17 nsew
rlabel metal4 s 94864 27554 94864 27554 4 vdd!
port 18 nsew
rlabel metal2 s 44192 -5062 44308 -4262 4 d6
port 9 nsew
rlabel metal2 s 759 54450 937 55250 4 inp1
port 3 nsew
rlabel metal2 s 67957 -5062 68073 -4262 4 inp2
port 4 nsew
rlabel metal2 s 21342 -5062 21458 -4262 4 d0
port 15 nsew
rlabel metal2 s 24819 -5062 24935 -4262 4 d1
port 14 nsew
rlabel metal2 s 27876 -5062 27992 -4262 4 d2
port 13 nsew
rlabel metal2 s 31555 -5062 31671 -4262 4 d3
port 12 nsew
rlabel metal2 s 35169 -5062 35285 -4262 4 d4
port 11 nsew
rlabel metal2 s 38704 -5062 38820 -4262 4 d5
port 10 nsew
rlabel metal2 s 93978 26540 93978 26540 4 gnd!
port 19 nsew
rlabel metal3 s 99044 26959 99844 27119 4 out
port 20 nsew
rlabel metal3 s 99044 24792 99844 24952 4 d7
port 5 nsew
<< properties >>
string FIXED_BBOX -5878 -5062 99844 55250
string GDS_FILE 8bitdac_layout.gds
string GDS_START 76282
string GDS_END 111544
<< end >>
