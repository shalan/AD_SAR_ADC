magic
tech sky130A
magscale 1 2
timestamp 1626710249
<< checkpaint >>
rect -9836 -8766 593760 712702
<< locali >>
rect 389925 346307 389959 347225
rect 335185 336685 335277 336719
rect 335185 336583 335219 336685
rect 335277 336447 335311 336549
rect 335461 336311 335495 336685
rect 343557 336311 343591 336481
rect 343649 336039 343683 336277
rect 212733 323595 212767 326485
rect 223773 321963 223807 326485
rect 171793 3451 171827 4165
rect 182097 3723 182131 3825
rect 233893 3723 233927 3893
rect 182005 3451 182039 3689
rect 233985 3383 234019 3689
rect 92489 3179 92523 3281
rect 239321 3179 239355 3485
rect 239413 2975 239447 3621
rect 250361 3451 250395 4097
rect 250453 3995 250487 4097
rect 340797 3995 340831 4233
rect 250545 3859 250579 3961
rect 342269 3995 342303 4233
rect 248429 3281 248521 3315
rect 248429 3043 248463 3281
rect 285689 3179 285723 3485
rect 334081 3315 334115 3961
rect 357357 3927 357391 4233
rect 358829 3927 358863 4233
rect 125793 2839 125827 2873
rect 130485 2839 130519 2873
rect 132417 2839 132451 2873
rect 248521 2839 248555 3009
rect 125793 2805 125885 2839
rect 130485 2805 130703 2839
rect 132359 2805 132451 2839
rect 248463 2805 248555 2839
rect 390569 2839 390603 3485
rect 392041 2839 392075 3553
rect 390569 2805 390753 2839
rect 130669 2771 130703 2805
<< viali >>
rect 389925 347225 389959 347259
rect 389925 346273 389959 346307
rect 335277 336685 335311 336719
rect 335461 336685 335495 336719
rect 335185 336549 335219 336583
rect 335277 336549 335311 336583
rect 335277 336413 335311 336447
rect 335461 336277 335495 336311
rect 343557 336481 343591 336515
rect 343557 336277 343591 336311
rect 343649 336277 343683 336311
rect 343649 336005 343683 336039
rect 212733 326485 212767 326519
rect 212733 323561 212767 323595
rect 223773 326485 223807 326519
rect 223773 321929 223807 321963
rect 340797 4233 340831 4267
rect 171793 4165 171827 4199
rect 250361 4097 250395 4131
rect 233893 3893 233927 3927
rect 182097 3825 182131 3859
rect 171793 3417 171827 3451
rect 182005 3689 182039 3723
rect 182097 3689 182131 3723
rect 233893 3689 233927 3723
rect 233985 3689 234019 3723
rect 182005 3417 182039 3451
rect 239413 3621 239447 3655
rect 233985 3349 234019 3383
rect 239321 3485 239355 3519
rect 92489 3281 92523 3315
rect 92489 3145 92523 3179
rect 239321 3145 239355 3179
rect 250453 4097 250487 4131
rect 250453 3961 250487 3995
rect 250545 3961 250579 3995
rect 250545 3825 250579 3859
rect 334081 3961 334115 3995
rect 340797 3961 340831 3995
rect 342269 4233 342303 4267
rect 342269 3961 342303 3995
rect 357357 4233 357391 4267
rect 250361 3417 250395 3451
rect 285689 3485 285723 3519
rect 248521 3281 248555 3315
rect 357357 3893 357391 3927
rect 358829 4233 358863 4267
rect 358829 3893 358863 3927
rect 392041 3553 392075 3587
rect 334081 3281 334115 3315
rect 390569 3485 390603 3519
rect 285689 3145 285723 3179
rect 248429 3009 248463 3043
rect 248521 3009 248555 3043
rect 239413 2941 239447 2975
rect 125793 2873 125827 2907
rect 130485 2873 130519 2907
rect 132417 2873 132451 2907
rect 125885 2805 125919 2839
rect 132325 2805 132359 2839
rect 248429 2805 248463 2839
rect 390753 2805 390787 2839
rect 392041 2805 392075 2839
rect 130669 2737 130703 2771
<< metal1 >>
rect 324222 700952 324228 701004
rect 324280 700992 324286 701004
rect 413646 700992 413652 701004
rect 324280 700964 413652 700992
rect 324280 700952 324286 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 331122 700884 331128 700936
rect 331180 700924 331186 700936
rect 429838 700924 429844 700936
rect 331180 700896 429844 700924
rect 331180 700884 331186 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 336642 700816 336648 700868
rect 336700 700856 336706 700868
rect 446122 700856 446128 700868
rect 336700 700828 446128 700856
rect 336700 700816 336706 700828
rect 446122 700816 446128 700828
rect 446180 700816 446186 700868
rect 342162 700748 342168 700800
rect 342220 700788 342226 700800
rect 462314 700788 462320 700800
rect 342220 700760 462320 700788
rect 342220 700748 342226 700760
rect 462314 700748 462320 700760
rect 462372 700748 462378 700800
rect 349062 700680 349068 700732
rect 349120 700720 349126 700732
rect 478506 700720 478512 700732
rect 349120 700692 478512 700720
rect 349120 700680 349126 700692
rect 478506 700680 478512 700692
rect 478564 700680 478570 700732
rect 354582 700612 354588 700664
rect 354640 700652 354646 700664
rect 494790 700652 494796 700664
rect 354640 700624 494796 700652
rect 354640 700612 354646 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 288342 700544 288348 700596
rect 288400 700584 288406 700596
rect 316310 700584 316316 700596
rect 288400 700556 316316 700584
rect 288400 700544 288406 700556
rect 316310 700544 316316 700556
rect 316368 700544 316374 700596
rect 361482 700544 361488 700596
rect 361540 700584 361546 700596
rect 510982 700584 510988 700596
rect 361540 700556 510988 700584
rect 361540 700544 361546 700556
rect 510982 700544 510988 700556
rect 511040 700544 511046 700596
rect 293862 700476 293868 700528
rect 293920 700516 293926 700528
rect 332502 700516 332508 700528
rect 293920 700488 332508 700516
rect 293920 700476 293926 700488
rect 332502 700476 332508 700488
rect 332560 700476 332566 700528
rect 367002 700476 367008 700528
rect 367060 700516 367066 700528
rect 527174 700516 527180 700528
rect 367060 700488 527180 700516
rect 367060 700476 367066 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 299382 700408 299388 700460
rect 299440 700448 299446 700460
rect 348786 700448 348792 700460
rect 299440 700420 348792 700448
rect 299440 700408 299446 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 373902 700408 373908 700460
rect 373960 700448 373966 700460
rect 543458 700448 543464 700460
rect 373960 700420 543464 700448
rect 373960 700408 373966 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 106182 700380 106188 700392
rect 105504 700352 106188 700380
rect 105504 700340 105510 700352
rect 106182 700340 106188 700352
rect 106240 700340 106246 700392
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 235902 700380 235908 700392
rect 235224 700352 235908 700380
rect 235224 700340 235230 700352
rect 235902 700340 235908 700352
rect 235960 700340 235966 700392
rect 276658 700340 276664 700392
rect 276716 700380 276722 700392
rect 283834 700380 283840 700392
rect 276716 700352 283840 700380
rect 276716 700340 276722 700352
rect 283834 700340 283840 700352
rect 283892 700340 283898 700392
rect 306282 700340 306288 700392
rect 306340 700380 306346 700392
rect 364978 700380 364984 700392
rect 306340 700352 364984 700380
rect 306340 700340 306346 700352
rect 364978 700340 364984 700352
rect 365036 700340 365042 700392
rect 379422 700340 379428 700392
rect 379480 700380 379486 700392
rect 559650 700380 559656 700392
rect 379480 700352 559656 700380
rect 379480 700340 379486 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 281442 700272 281448 700324
rect 281500 700312 281506 700324
rect 300118 700312 300124 700324
rect 281500 700284 300124 700312
rect 281500 700272 281506 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 311802 700272 311808 700324
rect 311860 700312 311866 700324
rect 381170 700312 381176 700324
rect 311860 700284 381176 700312
rect 311860 700272 311866 700284
rect 381170 700272 381176 700284
rect 381228 700272 381234 700324
rect 384942 700272 384948 700324
rect 385000 700312 385006 700324
rect 575842 700312 575848 700324
rect 385000 700284 575848 700312
rect 385000 700272 385006 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 171042 700244 171048 700256
rect 170364 700216 171048 700244
rect 170364 700204 170370 700216
rect 171042 700204 171048 700216
rect 171100 700204 171106 700256
rect 318702 700204 318708 700256
rect 318760 700244 318766 700256
rect 397454 700244 397460 700256
rect 318760 700216 397460 700244
rect 318760 700204 318766 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 56778 700136 56784 700188
rect 56836 700176 56842 700188
rect 57882 700176 57888 700188
rect 56836 700148 57888 700176
rect 56836 700136 56842 700148
rect 57882 700136 57888 700148
rect 57940 700136 57946 700188
rect 186498 700136 186504 700188
rect 186556 700176 186562 700188
rect 187602 700176 187608 700188
rect 186556 700148 187608 700176
rect 186556 700136 186562 700148
rect 187602 700136 187608 700148
rect 187660 700136 187666 700188
rect 251450 700068 251456 700120
rect 251508 700108 251514 700120
rect 252462 700108 252468 700120
rect 251508 700080 252468 700108
rect 251508 700068 251514 700080
rect 252462 700068 252468 700080
rect 252520 700068 252526 700120
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 122742 699700 122748 699712
rect 121696 699672 122748 699700
rect 121696 699660 121702 699672
rect 122742 699660 122748 699672
rect 122800 699660 122806 699712
rect 3418 696940 3424 696992
rect 3476 696980 3482 696992
rect 86218 696980 86224 696992
rect 3476 696952 86224 696980
rect 3476 696940 3482 696952
rect 86218 696940 86224 696952
rect 86276 696940 86282 696992
rect 389818 696940 389824 696992
rect 389876 696980 389882 696992
rect 580166 696980 580172 696992
rect 389876 696952 580172 696980
rect 389876 696940 389882 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 389910 683136 389916 683188
rect 389968 683176 389974 683188
rect 580166 683176 580172 683188
rect 389968 683148 580172 683176
rect 389968 683136 389974 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 390002 670692 390008 670744
rect 390060 670732 390066 670744
rect 580166 670732 580172 670744
rect 390060 670704 580172 670732
rect 390060 670692 390066 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 2774 645056 2780 645108
rect 2832 645096 2838 645108
rect 4798 645096 4804 645108
rect 2832 645068 4804 645096
rect 2832 645056 2838 645068
rect 4798 645056 4804 645068
rect 4856 645056 4862 645108
rect 390094 643084 390100 643136
rect 390152 643124 390158 643136
rect 580166 643124 580172 643136
rect 390152 643096 580172 643124
rect 390152 643084 390158 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 390186 630640 390192 630692
rect 390244 630680 390250 630692
rect 579982 630680 579988 630692
rect 390244 630652 579988 630680
rect 390244 630640 390250 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 390278 616836 390284 616888
rect 390336 616876 390342 616888
rect 580166 616876 580172 616888
rect 390336 616848 580172 616876
rect 390336 616836 390342 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 390370 590656 390376 590708
rect 390428 590696 390434 590708
rect 579614 590696 579620 590708
rect 390428 590668 579620 590696
rect 390428 590656 390434 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 390462 576852 390468 576904
rect 390520 576892 390526 576904
rect 579614 576892 579620 576904
rect 390520 576864 579620 576892
rect 390520 576852 390526 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 389726 536800 389732 536852
rect 389784 536840 389790 536852
rect 579614 536840 579620 536852
rect 389784 536812 579620 536840
rect 389784 536800 389790 536812
rect 579614 536800 579620 536812
rect 579672 536800 579678 536852
rect 389634 524424 389640 524476
rect 389692 524464 389698 524476
rect 580166 524464 580172 524476
rect 389692 524436 580172 524464
rect 389692 524424 389698 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 389542 484372 389548 484424
rect 389600 484412 389606 484424
rect 580166 484412 580172 484424
rect 389600 484384 580172 484412
rect 389600 484372 389606 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 274910 481584 274916 481636
rect 274968 481624 274974 481636
rect 276658 481624 276664 481636
rect 274968 481596 276664 481624
rect 274968 481584 274974 481596
rect 276658 481584 276664 481596
rect 276716 481584 276722 481636
rect 305454 481584 305460 481636
rect 305512 481624 305518 481636
rect 306282 481624 306288 481636
rect 305512 481596 306288 481624
rect 305512 481584 305518 481596
rect 306282 481584 306288 481596
rect 306340 481584 306346 481636
rect 329834 481584 329840 481636
rect 329892 481624 329898 481636
rect 331122 481624 331128 481636
rect 329892 481596 331128 481624
rect 329892 481584 329898 481596
rect 331122 481584 331128 481596
rect 331180 481584 331186 481636
rect 154482 481516 154488 481568
rect 154540 481556 154546 481568
rect 225966 481556 225972 481568
rect 154540 481528 225972 481556
rect 154540 481516 154546 481528
rect 225966 481516 225972 481528
rect 226024 481516 226030 481568
rect 137922 481448 137928 481500
rect 137980 481488 137986 481500
rect 219894 481488 219900 481500
rect 137980 481460 219900 481488
rect 137980 481448 137986 481460
rect 219894 481448 219900 481460
rect 219952 481448 219958 481500
rect 122742 481380 122748 481432
rect 122800 481420 122806 481432
rect 213730 481420 213736 481432
rect 122800 481392 213736 481420
rect 122800 481380 122806 481392
rect 213730 481380 213736 481392
rect 213788 481380 213794 481432
rect 106182 481312 106188 481364
rect 106240 481352 106246 481364
rect 207658 481352 207664 481364
rect 106240 481324 207664 481352
rect 106240 481312 106246 481324
rect 207658 481312 207664 481324
rect 207716 481312 207722 481364
rect 287054 481312 287060 481364
rect 287112 481352 287118 481364
rect 288342 481352 288348 481364
rect 287112 481324 288348 481352
rect 287112 481312 287118 481324
rect 288342 481312 288348 481324
rect 288400 481312 288406 481364
rect 89622 481244 89628 481296
rect 89680 481284 89686 481296
rect 201586 481284 201592 481296
rect 89680 481256 201592 481284
rect 89680 481244 89686 481256
rect 201586 481244 201592 481256
rect 201644 481244 201650 481296
rect 73062 481176 73068 481228
rect 73120 481216 73126 481228
rect 195422 481216 195428 481228
rect 73120 481188 195428 481216
rect 73120 481176 73126 481188
rect 195422 481176 195428 481188
rect 195480 481176 195486 481228
rect 317690 481176 317696 481228
rect 317748 481216 317754 481228
rect 318702 481216 318708 481228
rect 317748 481188 318708 481216
rect 317748 481176 317754 481188
rect 318702 481176 318708 481188
rect 318760 481176 318766 481228
rect 57882 481108 57888 481160
rect 57940 481148 57946 481160
rect 189350 481148 189356 481160
rect 57940 481120 189356 481148
rect 57940 481108 57946 481120
rect 189350 481108 189356 481120
rect 189408 481108 189414 481160
rect 219342 481108 219348 481160
rect 219400 481148 219406 481160
rect 250438 481148 250444 481160
rect 219400 481120 250444 481148
rect 219400 481108 219406 481120
rect 250438 481108 250444 481120
rect 250496 481108 250502 481160
rect 360378 481108 360384 481160
rect 360436 481148 360442 481160
rect 361482 481148 361488 481160
rect 360436 481120 361488 481148
rect 360436 481108 360442 481120
rect 361482 481108 361488 481120
rect 361540 481108 361546 481160
rect 41322 481040 41328 481092
rect 41380 481080 41386 481092
rect 183186 481080 183192 481092
rect 41380 481052 183192 481080
rect 41380 481040 41386 481052
rect 183186 481040 183192 481052
rect 183244 481040 183250 481092
rect 202782 481040 202788 481092
rect 202840 481080 202846 481092
rect 244366 481080 244372 481092
rect 202840 481052 244372 481080
rect 202840 481040 202846 481052
rect 244366 481040 244372 481052
rect 244424 481040 244430 481092
rect 348234 481040 348240 481092
rect 348292 481080 348298 481092
rect 349062 481080 349068 481092
rect 348292 481052 349068 481080
rect 348292 481040 348298 481052
rect 349062 481040 349068 481052
rect 349120 481040 349126 481092
rect 24762 480972 24768 481024
rect 24820 481012 24826 481024
rect 177114 481012 177120 481024
rect 24820 480984 177120 481012
rect 24820 480972 24826 480984
rect 177114 480972 177120 480984
rect 177172 480972 177178 481024
rect 187602 480972 187608 481024
rect 187660 481012 187666 481024
rect 238202 481012 238208 481024
rect 187660 480984 238208 481012
rect 187660 480972 187666 480984
rect 238202 480972 238208 480984
rect 238260 480972 238266 481024
rect 252462 480972 252468 481024
rect 252520 481012 252526 481024
rect 262674 481012 262680 481024
rect 252520 480984 262680 481012
rect 252520 480972 252526 480984
rect 262674 480972 262680 480984
rect 262732 480972 262738 481024
rect 8202 480904 8208 480956
rect 8260 480944 8266 480956
rect 171042 480944 171048 480956
rect 8260 480916 171048 480944
rect 8260 480904 8266 480916
rect 171042 480904 171048 480916
rect 171100 480904 171106 480956
rect 232130 480944 232136 480956
rect 180766 480916 232136 480944
rect 170950 480836 170956 480888
rect 171008 480876 171014 480888
rect 180766 480876 180794 480916
rect 232130 480904 232136 480916
rect 232188 480904 232194 480956
rect 235902 480904 235908 480956
rect 235960 480944 235966 480956
rect 256510 480944 256516 480956
rect 235960 480916 256516 480944
rect 235960 480904 235966 480916
rect 256510 480904 256516 480916
rect 256568 480904 256574 480956
rect 171008 480848 180794 480876
rect 171008 480836 171014 480848
rect 372614 480768 372620 480820
rect 372672 480808 372678 480820
rect 373902 480808 373908 480820
rect 372672 480780 373908 480808
rect 372672 480768 372678 480780
rect 373902 480768 373908 480780
rect 373960 480768 373966 480820
rect 267642 480224 267648 480276
rect 267700 480264 267706 480276
rect 268746 480264 268752 480276
rect 267700 480236 268752 480264
rect 267700 480224 267706 480236
rect 268746 480224 268752 480236
rect 268804 480224 268810 480276
rect 86218 477436 86224 477488
rect 86276 477476 86282 477488
rect 165614 477476 165620 477488
rect 86276 477448 165620 477476
rect 86276 477436 86282 477448
rect 165614 477436 165620 477448
rect 165672 477436 165678 477488
rect 3418 471928 3424 471980
rect 3476 471968 3482 471980
rect 165614 471968 165620 471980
rect 3476 471940 165620 471968
rect 3476 471928 3482 471940
rect 165614 471928 165620 471940
rect 165672 471928 165678 471980
rect 389818 470568 389824 470620
rect 389876 470608 389882 470620
rect 579982 470608 579988 470620
rect 389876 470580 579988 470608
rect 389876 470568 389882 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 469140 3516 469192
rect 3568 469180 3574 469192
rect 165614 469180 165620 469192
rect 3568 469152 165620 469180
rect 3568 469140 3574 469152
rect 165614 469140 165620 469152
rect 165672 469140 165678 469192
rect 390094 469140 390100 469192
rect 390152 469180 390158 469192
rect 580258 469180 580264 469192
rect 390152 469152 580264 469180
rect 390152 469140 390158 469152
rect 580258 469140 580264 469152
rect 580316 469140 580322 469192
rect 4798 466352 4804 466404
rect 4856 466392 4862 466404
rect 165614 466392 165620 466404
rect 4856 466364 165620 466392
rect 4856 466352 4862 466364
rect 165614 466352 165620 466364
rect 165672 466352 165678 466404
rect 3602 463632 3608 463684
rect 3660 463672 3666 463684
rect 165614 463672 165620 463684
rect 3660 463644 165620 463672
rect 3660 463632 3666 463644
rect 165614 463632 165620 463644
rect 165672 463632 165678 463684
rect 3694 462272 3700 462324
rect 3752 462312 3758 462324
rect 165614 462312 165620 462324
rect 3752 462284 165620 462312
rect 3752 462272 3758 462284
rect 165614 462272 165620 462284
rect 165672 462272 165678 462324
rect 3786 459484 3792 459536
rect 3844 459524 3850 459536
rect 165614 459524 165620 459536
rect 3844 459496 165620 459524
rect 3844 459484 3850 459496
rect 165614 459484 165620 459496
rect 165672 459484 165678 459536
rect 390186 458124 390192 458176
rect 390244 458164 390250 458176
rect 580350 458164 580356 458176
rect 390244 458136 580356 458164
rect 390244 458124 390250 458136
rect 580350 458124 580356 458136
rect 580408 458124 580414 458176
rect 389910 456764 389916 456816
rect 389968 456804 389974 456816
rect 579798 456804 579804 456816
rect 389968 456776 579804 456804
rect 389968 456764 389974 456776
rect 579798 456764 579804 456776
rect 579856 456764 579862 456816
rect 3878 456696 3884 456748
rect 3936 456736 3942 456748
rect 165614 456736 165620 456748
rect 3936 456708 165620 456736
rect 3936 456696 3942 456708
rect 165614 456696 165620 456708
rect 165672 456696 165678 456748
rect 3970 453976 3976 454028
rect 4028 454016 4034 454028
rect 165614 454016 165620 454028
rect 4028 453988 165620 454016
rect 4028 453976 4034 453988
rect 165614 453976 165620 453988
rect 165672 453976 165678 454028
rect 4062 451188 4068 451240
rect 4120 451228 4126 451240
rect 165614 451228 165620 451240
rect 4120 451200 165620 451228
rect 4120 451188 4126 451200
rect 165614 451188 165620 451200
rect 165672 451188 165678 451240
rect 390186 451188 390192 451240
rect 390244 451228 390250 451240
rect 580442 451228 580448 451240
rect 390244 451200 580448 451228
rect 390244 451188 390250 451200
rect 580442 451188 580448 451200
rect 580500 451188 580506 451240
rect 3326 448468 3332 448520
rect 3384 448508 3390 448520
rect 165614 448508 165620 448520
rect 3384 448480 165620 448508
rect 3384 448468 3390 448480
rect 165614 448468 165620 448480
rect 165672 448468 165678 448520
rect 390186 448468 390192 448520
rect 390244 448508 390250 448520
rect 580534 448508 580540 448520
rect 390244 448480 580540 448508
rect 390244 448468 390250 448480
rect 580534 448468 580540 448480
rect 580592 448468 580598 448520
rect 3234 445680 3240 445732
rect 3292 445720 3298 445732
rect 165614 445720 165620 445732
rect 3292 445692 165620 445720
rect 3292 445680 3298 445692
rect 165614 445680 165620 445692
rect 165672 445680 165678 445732
rect 390002 444388 390008 444440
rect 390060 444428 390066 444440
rect 580166 444428 580172 444440
rect 390060 444400 580172 444428
rect 390060 444388 390066 444400
rect 580166 444388 580172 444400
rect 580224 444388 580230 444440
rect 3142 442892 3148 442944
rect 3200 442932 3206 442944
rect 165614 442932 165620 442944
rect 3200 442904 165620 442932
rect 3200 442892 3206 442904
rect 165614 442892 165620 442904
rect 165672 442892 165678 442944
rect 3050 441532 3056 441584
rect 3108 441572 3114 441584
rect 165614 441572 165620 441584
rect 3108 441544 165620 441572
rect 3108 441532 3114 441544
rect 165614 441532 165620 441544
rect 165672 441532 165678 441584
rect 390186 440172 390192 440224
rect 390244 440212 390250 440224
rect 580626 440212 580632 440224
rect 390244 440184 580632 440212
rect 390244 440172 390250 440184
rect 580626 440172 580632 440184
rect 580684 440172 580690 440224
rect 2958 438812 2964 438864
rect 3016 438852 3022 438864
rect 165614 438852 165620 438864
rect 3016 438824 165620 438852
rect 3016 438812 3022 438824
rect 165614 438812 165620 438824
rect 165672 438812 165678 438864
rect 390278 437384 390284 437436
rect 390336 437424 390342 437436
rect 580718 437424 580724 437436
rect 390336 437396 580724 437424
rect 390336 437384 390342 437396
rect 580718 437384 580724 437396
rect 580776 437384 580782 437436
rect 2866 436024 2872 436076
rect 2924 436064 2930 436076
rect 165614 436064 165620 436076
rect 2924 436036 165620 436064
rect 2924 436024 2930 436036
rect 165614 436024 165620 436036
rect 165672 436024 165678 436076
rect 2774 433236 2780 433288
rect 2832 433276 2838 433288
rect 165614 433276 165620 433288
rect 2832 433248 165620 433276
rect 2832 433236 2838 433248
rect 165614 433236 165620 433248
rect 165672 433236 165678 433288
rect 389818 430584 389824 430636
rect 389876 430624 389882 430636
rect 580166 430624 580172 430636
rect 389876 430596 580172 430624
rect 389876 430584 389882 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 430516 3424 430568
rect 3476 430556 3482 430568
rect 165614 430556 165620 430568
rect 3476 430528 165620 430556
rect 3476 430516 3482 430528
rect 165614 430516 165620 430528
rect 165672 430516 165678 430568
rect 3510 427728 3516 427780
rect 3568 427768 3574 427780
rect 165614 427768 165620 427780
rect 3568 427740 165620 427768
rect 3568 427728 3574 427740
rect 165614 427728 165620 427740
rect 165672 427728 165678 427780
rect 3602 425008 3608 425060
rect 3660 425048 3666 425060
rect 165614 425048 165620 425060
rect 3660 425020 165620 425048
rect 3660 425008 3666 425020
rect 165614 425008 165620 425020
rect 165672 425008 165678 425060
rect 3786 422220 3792 422272
rect 3844 422260 3850 422272
rect 165614 422260 165620 422272
rect 3844 422232 165620 422260
rect 3844 422220 3850 422232
rect 165614 422220 165620 422232
rect 165672 422220 165678 422272
rect 390094 419432 390100 419484
rect 390152 419472 390158 419484
rect 580166 419472 580172 419484
rect 390152 419444 580172 419472
rect 390152 419432 390158 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 3418 418140 3424 418192
rect 3476 418180 3482 418192
rect 165614 418180 165620 418192
rect 3476 418152 165620 418180
rect 3476 418140 3482 418152
rect 165614 418140 165620 418152
rect 165672 418140 165678 418192
rect 3786 416780 3792 416832
rect 3844 416820 3850 416832
rect 165614 416820 165620 416832
rect 3844 416792 165620 416820
rect 3844 416780 3850 416792
rect 165614 416780 165620 416792
rect 165672 416780 165678 416832
rect 3694 413992 3700 414044
rect 3752 414032 3758 414044
rect 165614 414032 165620 414044
rect 3752 414004 165620 414032
rect 3752 413992 3758 414004
rect 165614 413992 165620 414004
rect 165672 413992 165678 414044
rect 3602 411272 3608 411324
rect 3660 411312 3666 411324
rect 165614 411312 165620 411324
rect 3660 411284 165620 411312
rect 3660 411272 3666 411284
rect 165614 411272 165620 411284
rect 165672 411272 165678 411324
rect 3510 408484 3516 408536
rect 3568 408524 3574 408536
rect 165614 408524 165620 408536
rect 3568 408496 165620 408524
rect 3568 408484 3574 408496
rect 165614 408484 165620 408496
rect 165672 408484 165678 408536
rect 3418 405696 3424 405748
rect 3476 405736 3482 405748
rect 165614 405736 165620 405748
rect 3476 405708 165620 405736
rect 3476 405696 3482 405708
rect 165614 405696 165620 405708
rect 165672 405696 165678 405748
rect 390186 405628 390192 405680
rect 390244 405668 390250 405680
rect 580166 405668 580172 405680
rect 390244 405640 580172 405668
rect 390244 405628 390250 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 389174 404472 389180 404524
rect 389232 404512 389238 404524
rect 391198 404512 391204 404524
rect 389232 404484 391204 404512
rect 389232 404472 389238 404484
rect 391198 404472 391204 404484
rect 391256 404472 391262 404524
rect 3142 398828 3148 398880
rect 3200 398868 3206 398880
rect 165614 398868 165620 398880
rect 3200 398840 165620 398868
rect 3200 398828 3206 398840
rect 165614 398828 165620 398840
rect 165672 398828 165678 398880
rect 4798 396040 4804 396092
rect 4856 396080 4862 396092
rect 165614 396080 165620 396092
rect 4856 396052 165620 396080
rect 4856 396040 4862 396052
rect 165614 396040 165620 396052
rect 165672 396040 165678 396092
rect 390186 393320 390192 393372
rect 390244 393360 390250 393372
rect 396810 393360 396816 393372
rect 390244 393332 396816 393360
rect 390244 393320 390250 393332
rect 396810 393320 396816 393332
rect 396868 393320 396874 393372
rect 390186 391960 390192 392012
rect 390244 392000 390250 392012
rect 393958 392000 393964 392012
rect 390244 391972 393964 392000
rect 390244 391960 390250 391972
rect 393958 391960 393964 391972
rect 394016 391960 394022 392012
rect 390094 391892 390100 391944
rect 390152 391932 390158 391944
rect 580166 391932 580172 391944
rect 390152 391904 580172 391932
rect 390152 391892 390158 391904
rect 580166 391892 580172 391904
rect 580224 391892 580230 391944
rect 390186 389172 390192 389224
rect 390244 389212 390250 389224
rect 406378 389212 406384 389224
rect 390244 389184 406384 389212
rect 390244 389172 390250 389184
rect 406378 389172 406384 389184
rect 406436 389172 406442 389224
rect 21450 387812 21456 387864
rect 21508 387852 21514 387864
rect 165614 387852 165620 387864
rect 21508 387824 165620 387852
rect 21508 387812 21514 387824
rect 165614 387812 165620 387824
rect 165672 387812 165678 387864
rect 3234 385024 3240 385076
rect 3292 385064 3298 385076
rect 165614 385064 165620 385076
rect 3292 385036 165620 385064
rect 3292 385024 3298 385036
rect 165614 385024 165620 385036
rect 165672 385024 165678 385076
rect 390002 379448 390008 379500
rect 390060 379488 390066 379500
rect 580166 379488 580172 379500
rect 390060 379460 580172 379488
rect 390060 379448 390066 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 376728 3332 376780
rect 3384 376768 3390 376780
rect 165614 376768 165620 376780
rect 3384 376740 165620 376768
rect 3384 376728 3390 376740
rect 165614 376728 165620 376740
rect 165672 376728 165678 376780
rect 10318 375368 10324 375420
rect 10376 375408 10382 375420
rect 165614 375408 165620 375420
rect 10376 375380 165620 375408
rect 10376 375368 10382 375380
rect 165614 375368 165620 375380
rect 165672 375368 165678 375420
rect 390094 372580 390100 372632
rect 390152 372620 390158 372632
rect 403618 372620 403624 372632
rect 390152 372592 403624 372620
rect 390152 372580 390158 372592
rect 403618 372580 403624 372592
rect 403676 372580 403682 372632
rect 4062 369860 4068 369912
rect 4120 369900 4126 369912
rect 165614 369900 165620 369912
rect 4120 369872 165620 369900
rect 4120 369860 4126 369872
rect 165614 369860 165620 369872
rect 165672 369860 165678 369912
rect 28258 367072 28264 367124
rect 28316 367112 28322 367124
rect 165614 367112 165620 367124
rect 28316 367084 165620 367112
rect 28316 367072 28322 367084
rect 165614 367072 165620 367084
rect 165672 367072 165678 367124
rect 389910 365644 389916 365696
rect 389968 365684 389974 365696
rect 580166 365684 580172 365696
rect 389968 365656 580172 365684
rect 389968 365644 389974 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3970 364352 3976 364404
rect 4028 364392 4034 364404
rect 165614 364392 165620 364404
rect 4028 364364 165620 364392
rect 4028 364352 4034 364364
rect 165614 364352 165620 364364
rect 165672 364352 165678 364404
rect 3878 358776 3884 358828
rect 3936 358816 3942 358828
rect 165614 358816 165620 358828
rect 3936 358788 165620 358816
rect 3936 358776 3942 358788
rect 165614 358776 165620 358788
rect 165672 358776 165678 358828
rect 390094 357416 390100 357468
rect 390152 357456 390158 357468
rect 400858 357456 400864 357468
rect 390152 357428 400864 357456
rect 390152 357416 390158 357428
rect 400858 357416 400864 357428
rect 400916 357416 400922 357468
rect 389910 357280 389916 357332
rect 389968 357320 389974 357332
rect 390094 357320 390100 357332
rect 389968 357292 390100 357320
rect 389968 357280 389974 357292
rect 390094 357280 390100 357292
rect 390152 357280 390158 357332
rect 3786 356056 3792 356108
rect 3844 356096 3850 356108
rect 165614 356096 165620 356108
rect 3844 356068 165620 356096
rect 3844 356056 3850 356068
rect 165614 356056 165620 356068
rect 165672 356056 165678 356108
rect 11698 354696 11704 354748
rect 11756 354736 11762 354748
rect 165614 354736 165620 354748
rect 11756 354708 165620 354736
rect 11756 354696 11762 354708
rect 165614 354696 165620 354708
rect 165672 354696 165678 354748
rect 389910 354696 389916 354748
rect 389968 354736 389974 354748
rect 547138 354736 547144 354748
rect 389968 354708 547144 354736
rect 389968 354696 389974 354708
rect 547138 354696 547144 354708
rect 547196 354696 547202 354748
rect 389818 353200 389824 353252
rect 389876 353240 389882 353252
rect 580166 353240 580172 353252
rect 389876 353212 580172 353240
rect 389876 353200 389882 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3694 351908 3700 351960
rect 3752 351948 3758 351960
rect 165614 351948 165620 351960
rect 3752 351920 165620 351948
rect 3752 351908 3758 351920
rect 165614 351908 165620 351920
rect 165672 351908 165678 351960
rect 29638 349120 29644 349172
rect 29696 349160 29702 349172
rect 165614 349160 165620 349172
rect 29696 349132 165620 349160
rect 29696 349120 29702 349132
rect 165614 349120 165620 349132
rect 165672 349120 165678 349172
rect 389910 347256 389916 347268
rect 389871 347228 389916 347256
rect 389910 347216 389916 347228
rect 389968 347216 389974 347268
rect 3602 346400 3608 346452
rect 3660 346440 3666 346452
rect 165614 346440 165620 346452
rect 3660 346412 165620 346440
rect 3660 346400 3666 346412
rect 165614 346400 165620 346412
rect 165672 346400 165678 346452
rect 389910 346400 389916 346452
rect 389968 346440 389974 346452
rect 542998 346440 543004 346452
rect 389968 346412 543004 346440
rect 389968 346400 389974 346412
rect 542998 346400 543004 346412
rect 543056 346400 543062 346452
rect 389910 346304 389916 346316
rect 389871 346276 389916 346304
rect 389910 346264 389916 346276
rect 389968 346264 389974 346316
rect 3510 343612 3516 343664
rect 3568 343652 3574 343664
rect 165614 343652 165620 343664
rect 3568 343624 165620 343652
rect 3568 343612 3574 343624
rect 165614 343612 165620 343624
rect 165672 343612 165678 343664
rect 396810 341504 396816 341556
rect 396868 341544 396874 341556
rect 580258 341544 580264 341556
rect 396868 341516 580264 341544
rect 396868 341504 396874 341516
rect 580258 341504 580264 341516
rect 580316 341504 580322 341556
rect 3418 340892 3424 340944
rect 3476 340932 3482 340944
rect 165614 340932 165620 340944
rect 3476 340904 165620 340932
rect 3476 340892 3482 340904
rect 165614 340892 165620 340904
rect 165672 340892 165678 340944
rect 389082 340892 389088 340944
rect 389140 340932 389146 340944
rect 396718 340932 396724 340944
rect 389140 340904 396724 340932
rect 389140 340892 389146 340904
rect 396718 340892 396724 340904
rect 396776 340892 396782 340944
rect 391198 340144 391204 340196
rect 391256 340184 391262 340196
rect 580166 340184 580172 340196
rect 391256 340156 580172 340184
rect 391256 340144 391262 340156
rect 580166 340144 580172 340156
rect 580224 340144 580230 340196
rect 18598 338104 18604 338156
rect 18656 338144 18662 338156
rect 165614 338144 165620 338156
rect 18656 338116 165620 338144
rect 18656 338104 18662 338116
rect 165614 338104 165620 338116
rect 165672 338104 165678 338156
rect 389082 338104 389088 338156
rect 389140 338144 389146 338156
rect 519538 338144 519544 338156
rect 389140 338116 519544 338144
rect 389140 338104 389146 338116
rect 519538 338104 519544 338116
rect 519596 338104 519602 338156
rect 168374 336744 168380 336796
rect 168432 336784 168438 336796
rect 168742 336784 168748 336796
rect 168432 336756 168748 336784
rect 168432 336744 168438 336756
rect 168742 336744 168748 336756
rect 168800 336744 168806 336796
rect 189074 336744 189080 336796
rect 189132 336784 189138 336796
rect 189350 336784 189356 336796
rect 189132 336756 189356 336784
rect 189132 336744 189138 336756
rect 189350 336744 189356 336756
rect 189408 336744 189414 336796
rect 240134 336744 240140 336796
rect 240192 336784 240198 336796
rect 240410 336784 240416 336796
rect 240192 336756 240416 336784
rect 240192 336744 240198 336756
rect 240410 336744 240416 336756
rect 240468 336744 240474 336796
rect 118602 336676 118608 336728
rect 118660 336716 118666 336728
rect 212258 336716 212264 336728
rect 118660 336688 212264 336716
rect 118660 336676 118666 336688
rect 212258 336676 212264 336688
rect 212316 336676 212322 336728
rect 220814 336676 220820 336728
rect 220872 336716 220878 336728
rect 221182 336716 221188 336728
rect 220872 336688 221188 336716
rect 220872 336676 220878 336688
rect 221182 336676 221188 336688
rect 221240 336676 221246 336728
rect 233878 336676 233884 336728
rect 233936 336716 233942 336728
rect 237190 336716 237196 336728
rect 233936 336688 237196 336716
rect 233936 336676 233942 336688
rect 237190 336676 237196 336688
rect 237248 336676 237254 336728
rect 239398 336676 239404 336728
rect 239456 336716 239462 336728
rect 241606 336716 241612 336728
rect 239456 336688 241612 336716
rect 239456 336676 239462 336688
rect 241606 336676 241612 336688
rect 241664 336676 241670 336728
rect 242066 336676 242072 336728
rect 242124 336716 242130 336728
rect 255406 336716 255412 336728
rect 242124 336688 255412 336716
rect 242124 336676 242130 336688
rect 255406 336676 255412 336688
rect 255464 336676 255470 336728
rect 260650 336676 260656 336728
rect 260708 336716 260714 336728
rect 265618 336716 265624 336728
rect 260708 336688 265624 336716
rect 260708 336676 260714 336688
rect 265618 336676 265624 336688
rect 265676 336676 265682 336728
rect 271046 336676 271052 336728
rect 271104 336716 271110 336728
rect 271782 336716 271788 336728
rect 271104 336688 271788 336716
rect 271104 336676 271110 336688
rect 271782 336676 271788 336688
rect 271840 336676 271846 336728
rect 272242 336676 272248 336728
rect 272300 336716 272306 336728
rect 276198 336716 276204 336728
rect 272300 336688 276204 336716
rect 272300 336676 272306 336688
rect 276198 336676 276204 336688
rect 276256 336676 276262 336728
rect 276382 336676 276388 336728
rect 276440 336716 276446 336728
rect 277210 336716 277216 336728
rect 276440 336688 277216 336716
rect 276440 336676 276446 336688
rect 277210 336676 277216 336688
rect 277268 336676 277274 336728
rect 279050 336676 279056 336728
rect 279108 336716 279114 336728
rect 280062 336716 280068 336728
rect 279108 336688 280068 336716
rect 279108 336676 279114 336688
rect 280062 336676 280068 336688
rect 280120 336676 280126 336728
rect 280338 336676 280344 336728
rect 280396 336716 280402 336728
rect 281350 336716 281356 336728
rect 280396 336688 281356 336716
rect 280396 336676 280402 336688
rect 281350 336676 281356 336688
rect 281408 336676 281414 336728
rect 281718 336676 281724 336728
rect 281776 336716 281782 336728
rect 282822 336716 282828 336728
rect 281776 336688 282828 336716
rect 281776 336676 281782 336688
rect 282822 336676 282828 336688
rect 282880 336676 282886 336728
rect 286134 336676 286140 336728
rect 286192 336716 286198 336728
rect 286870 336716 286876 336728
rect 286192 336688 286876 336716
rect 286192 336676 286198 336688
rect 286870 336676 286876 336688
rect 286928 336676 286934 336728
rect 289722 336676 289728 336728
rect 289780 336716 289786 336728
rect 290458 336716 290464 336728
rect 289780 336688 290464 336716
rect 289780 336676 289786 336688
rect 290458 336676 290464 336688
rect 290516 336676 290522 336728
rect 291470 336676 291476 336728
rect 291528 336716 291534 336728
rect 292482 336716 292488 336728
rect 291528 336688 292488 336716
rect 291528 336676 291534 336688
rect 292482 336676 292488 336688
rect 292540 336676 292546 336728
rect 292850 336676 292856 336728
rect 292908 336716 292914 336728
rect 293770 336716 293776 336728
rect 292908 336688 293776 336716
rect 292908 336676 292914 336688
rect 293770 336676 293776 336688
rect 293828 336676 293834 336728
rect 294598 336676 294604 336728
rect 294656 336716 294662 336728
rect 295242 336716 295248 336728
rect 294656 336688 295248 336716
rect 294656 336676 294662 336688
rect 295242 336676 295248 336688
rect 295300 336676 295306 336728
rect 295978 336676 295984 336728
rect 296036 336716 296042 336728
rect 296622 336716 296628 336728
rect 296036 336688 296628 336716
rect 296036 336676 296042 336688
rect 296622 336676 296628 336688
rect 296680 336676 296686 336728
rect 298646 336676 298652 336728
rect 298704 336716 298710 336728
rect 299382 336716 299388 336728
rect 298704 336688 299388 336716
rect 298704 336676 298710 336688
rect 299382 336676 299388 336688
rect 299440 336676 299446 336728
rect 299934 336676 299940 336728
rect 299992 336716 299998 336728
rect 300762 336716 300768 336728
rect 299992 336688 300768 336716
rect 299992 336676 299998 336688
rect 300762 336676 300768 336688
rect 300820 336676 300826 336728
rect 300854 336676 300860 336728
rect 300912 336716 300918 336728
rect 301958 336716 301964 336728
rect 300912 336688 301964 336716
rect 300912 336676 300918 336688
rect 301958 336676 301964 336688
rect 302016 336676 302022 336728
rect 303982 336676 303988 336728
rect 304040 336716 304046 336728
rect 304718 336716 304724 336728
rect 304040 336688 304724 336716
rect 304040 336676 304046 336688
rect 304718 336676 304724 336688
rect 304776 336676 304782 336728
rect 305270 336676 305276 336728
rect 305328 336716 305334 336728
rect 306098 336716 306104 336728
rect 305328 336688 306104 336716
rect 305328 336676 305334 336688
rect 306098 336676 306104 336688
rect 306156 336676 306162 336728
rect 306650 336676 306656 336728
rect 306708 336716 306714 336728
rect 307478 336716 307484 336728
rect 306708 336688 307484 336716
rect 306708 336676 306714 336688
rect 307478 336676 307484 336688
rect 307536 336676 307542 336728
rect 307938 336676 307944 336728
rect 307996 336716 308002 336728
rect 308858 336716 308864 336728
rect 307996 336688 308864 336716
rect 307996 336676 308002 336688
rect 308858 336676 308864 336688
rect 308916 336676 308922 336728
rect 309318 336676 309324 336728
rect 309376 336716 309382 336728
rect 310238 336716 310244 336728
rect 309376 336688 310244 336716
rect 309376 336676 309382 336688
rect 310238 336676 310244 336688
rect 310296 336676 310302 336728
rect 310606 336676 310612 336728
rect 310664 336716 310670 336728
rect 311618 336716 311624 336728
rect 310664 336688 311624 336716
rect 310664 336676 310670 336688
rect 311618 336676 311624 336688
rect 311676 336676 311682 336728
rect 312446 336676 312452 336728
rect 312504 336716 312510 336728
rect 313182 336716 313188 336728
rect 312504 336688 313188 336716
rect 312504 336676 312510 336688
rect 313182 336676 313188 336688
rect 313240 336676 313246 336728
rect 313274 336676 313280 336728
rect 313332 336716 313338 336728
rect 314470 336716 314476 336728
rect 313332 336688 314476 336716
rect 313332 336676 313338 336688
rect 314470 336676 314476 336688
rect 314528 336676 314534 336728
rect 314654 336676 314660 336728
rect 314712 336716 314718 336728
rect 315850 336716 315856 336728
rect 314712 336688 315856 336716
rect 314712 336676 314718 336688
rect 315850 336676 315856 336688
rect 315908 336676 315914 336728
rect 316402 336676 316408 336728
rect 316460 336716 316466 336728
rect 317322 336716 317328 336728
rect 316460 336688 317328 336716
rect 316460 336676 316466 336688
rect 317322 336676 317328 336688
rect 317380 336676 317386 336728
rect 319070 336676 319076 336728
rect 319128 336716 319134 336728
rect 320082 336716 320088 336728
rect 319128 336688 320088 336716
rect 319128 336676 319134 336688
rect 320082 336676 320088 336688
rect 320140 336676 320146 336728
rect 320450 336676 320456 336728
rect 320508 336716 320514 336728
rect 321462 336716 321468 336728
rect 320508 336688 321468 336716
rect 320508 336676 320514 336688
rect 321462 336676 321468 336688
rect 321520 336676 321526 336728
rect 324406 336676 324412 336728
rect 324464 336716 324470 336728
rect 325602 336716 325608 336728
rect 324464 336688 325608 336716
rect 324464 336676 324470 336688
rect 325602 336676 325608 336688
rect 325660 336676 325666 336728
rect 327534 336676 327540 336728
rect 327592 336716 327598 336728
rect 328270 336716 328276 336728
rect 327592 336688 328276 336716
rect 327592 336676 327598 336688
rect 328270 336676 328276 336688
rect 328328 336676 328334 336728
rect 328914 336676 328920 336728
rect 328972 336716 328978 336728
rect 329650 336716 329656 336728
rect 328972 336688 329656 336716
rect 328972 336676 328978 336688
rect 329650 336676 329656 336688
rect 329708 336676 329714 336728
rect 330202 336676 330208 336728
rect 330260 336716 330266 336728
rect 331122 336716 331128 336728
rect 330260 336688 331128 336716
rect 330260 336676 330266 336688
rect 331122 336676 331128 336688
rect 331180 336676 331186 336728
rect 331582 336676 331588 336728
rect 331640 336716 331646 336728
rect 332410 336716 332416 336728
rect 331640 336688 332416 336716
rect 331640 336676 331646 336688
rect 332410 336676 332416 336688
rect 332468 336676 332474 336728
rect 332870 336676 332876 336728
rect 332928 336716 332934 336728
rect 333882 336716 333888 336728
rect 332928 336688 333888 336716
rect 332928 336676 332934 336688
rect 333882 336676 333888 336688
rect 333940 336676 333946 336728
rect 334250 336676 334256 336728
rect 334308 336716 334314 336728
rect 335170 336716 335176 336728
rect 334308 336688 335176 336716
rect 334308 336676 334314 336688
rect 335170 336676 335176 336688
rect 335228 336676 335234 336728
rect 335265 336719 335323 336725
rect 335265 336685 335277 336719
rect 335311 336716 335323 336719
rect 335449 336719 335507 336725
rect 335449 336716 335461 336719
rect 335311 336688 335461 336716
rect 335311 336685 335323 336688
rect 335265 336679 335323 336685
rect 335449 336685 335461 336688
rect 335495 336685 335507 336719
rect 335449 336679 335507 336685
rect 335538 336676 335544 336728
rect 335596 336716 335602 336728
rect 336642 336716 336648 336728
rect 335596 336688 336648 336716
rect 335596 336676 335602 336688
rect 336642 336676 336648 336688
rect 336700 336676 336706 336728
rect 336918 336676 336924 336728
rect 336976 336716 336982 336728
rect 337930 336716 337936 336728
rect 336976 336688 337936 336716
rect 336976 336676 336982 336688
rect 337930 336676 337936 336688
rect 337988 336676 337994 336728
rect 338206 336676 338212 336728
rect 338264 336716 338270 336728
rect 339402 336716 339408 336728
rect 338264 336688 339408 336716
rect 338264 336676 338270 336688
rect 339402 336676 339408 336688
rect 339460 336676 339466 336728
rect 339586 336676 339592 336728
rect 339644 336716 339650 336728
rect 340690 336716 340696 336728
rect 339644 336688 340696 336716
rect 339644 336676 339650 336688
rect 340690 336676 340696 336688
rect 340748 336676 340754 336728
rect 340874 336676 340880 336728
rect 340932 336716 340938 336728
rect 342162 336716 342168 336728
rect 340932 336688 342168 336716
rect 340932 336676 340938 336688
rect 342162 336676 342168 336688
rect 342220 336676 342226 336728
rect 343174 336676 343180 336728
rect 343232 336716 343238 336728
rect 343542 336716 343548 336728
rect 343232 336688 343548 336716
rect 343232 336676 343238 336688
rect 343542 336676 343548 336688
rect 343600 336676 343606 336728
rect 345382 336676 345388 336728
rect 345440 336716 345446 336728
rect 346118 336716 346124 336728
rect 345440 336688 346124 336716
rect 345440 336676 345446 336688
rect 346118 336676 346124 336688
rect 346176 336676 346182 336728
rect 348050 336676 348056 336728
rect 348108 336716 348114 336728
rect 348878 336716 348884 336728
rect 348108 336688 348884 336716
rect 348108 336676 348114 336688
rect 348878 336676 348884 336688
rect 348936 336676 348942 336728
rect 350718 336676 350724 336728
rect 350776 336716 350782 336728
rect 351822 336716 351828 336728
rect 350776 336688 351828 336716
rect 350776 336676 350782 336688
rect 351822 336676 351828 336688
rect 351880 336676 351886 336728
rect 352006 336676 352012 336728
rect 352064 336716 352070 336728
rect 353110 336716 353116 336728
rect 352064 336688 353116 336716
rect 352064 336676 352070 336688
rect 353110 336676 353116 336688
rect 353168 336676 353174 336728
rect 355134 336676 355140 336728
rect 355192 336716 355198 336728
rect 355870 336716 355876 336728
rect 355192 336688 355876 336716
rect 355192 336676 355198 336688
rect 355870 336676 355876 336688
rect 355928 336676 355934 336728
rect 356054 336676 356060 336728
rect 356112 336716 356118 336728
rect 357342 336716 357348 336728
rect 356112 336688 357348 336716
rect 356112 336676 356118 336688
rect 357342 336676 357348 336688
rect 357400 336676 357406 336728
rect 357802 336676 357808 336728
rect 357860 336716 357866 336728
rect 358630 336716 358636 336728
rect 357860 336688 358636 336716
rect 357860 336676 357866 336688
rect 358630 336676 358636 336688
rect 358688 336676 358694 336728
rect 359182 336676 359188 336728
rect 359240 336716 359246 336728
rect 360010 336716 360016 336728
rect 359240 336688 360016 336716
rect 359240 336676 359246 336688
rect 360010 336676 360016 336688
rect 360068 336676 360074 336728
rect 360470 336676 360476 336728
rect 360528 336716 360534 336728
rect 361390 336716 361396 336728
rect 360528 336688 361396 336716
rect 360528 336676 360534 336688
rect 361390 336676 361396 336688
rect 361448 336676 361454 336728
rect 361850 336676 361856 336728
rect 361908 336716 361914 336728
rect 362678 336716 362684 336728
rect 361908 336688 362684 336716
rect 361908 336676 361914 336688
rect 362678 336676 362684 336688
rect 362736 336676 362742 336728
rect 363138 336676 363144 336728
rect 363196 336716 363202 336728
rect 364058 336716 364064 336728
rect 363196 336688 364064 336716
rect 363196 336676 363202 336688
rect 364058 336676 364064 336688
rect 364116 336676 364122 336728
rect 364518 336676 364524 336728
rect 364576 336716 364582 336728
rect 365438 336716 365444 336728
rect 364576 336688 365444 336716
rect 364576 336676 364582 336688
rect 365438 336676 365444 336688
rect 365496 336676 365502 336728
rect 365806 336676 365812 336728
rect 365864 336716 365870 336728
rect 366818 336716 366824 336728
rect 365864 336688 366824 336716
rect 365864 336676 365870 336688
rect 366818 336676 366824 336688
rect 366876 336676 366882 336728
rect 367186 336676 367192 336728
rect 367244 336716 367250 336728
rect 368198 336716 368204 336728
rect 367244 336688 368204 336716
rect 367244 336676 367250 336688
rect 368198 336676 368204 336688
rect 368256 336676 368262 336728
rect 368934 336676 368940 336728
rect 368992 336716 368998 336728
rect 369762 336716 369768 336728
rect 368992 336688 369768 336716
rect 368992 336676 368998 336688
rect 369762 336676 369768 336688
rect 369820 336676 369826 336728
rect 369854 336676 369860 336728
rect 369912 336716 369918 336728
rect 370958 336716 370964 336728
rect 369912 336688 370964 336716
rect 369912 336676 369918 336688
rect 370958 336676 370964 336688
rect 371016 336676 371022 336728
rect 372062 336676 372068 336728
rect 372120 336716 372126 336728
rect 372430 336716 372436 336728
rect 372120 336688 372436 336716
rect 372120 336676 372126 336688
rect 372430 336676 372436 336688
rect 372488 336676 372494 336728
rect 373442 336676 373448 336728
rect 373500 336716 373506 336728
rect 373810 336716 373816 336728
rect 373500 336688 373816 336716
rect 373500 336676 373506 336688
rect 373810 336676 373816 336688
rect 373868 336676 373874 336728
rect 374730 336676 374736 336728
rect 374788 336716 374794 336728
rect 375190 336716 375196 336728
rect 374788 336688 375196 336716
rect 374788 336676 374794 336688
rect 375190 336676 375196 336688
rect 375248 336676 375254 336728
rect 375650 336676 375656 336728
rect 375708 336716 375714 336728
rect 376662 336716 376668 336728
rect 375708 336688 376668 336716
rect 375708 336676 375714 336688
rect 376662 336676 376668 336688
rect 376720 336676 376726 336728
rect 376938 336676 376944 336728
rect 376996 336716 377002 336728
rect 378042 336716 378048 336728
rect 376996 336688 378048 336716
rect 376996 336676 377002 336688
rect 378042 336676 378048 336688
rect 378100 336676 378106 336728
rect 378778 336676 378784 336728
rect 378836 336716 378842 336728
rect 379330 336716 379336 336728
rect 378836 336688 379336 336716
rect 378836 336676 378842 336688
rect 379330 336676 379336 336688
rect 379388 336676 379394 336728
rect 380066 336676 380072 336728
rect 380124 336716 380130 336728
rect 380710 336716 380716 336728
rect 380124 336688 380716 336716
rect 380124 336676 380130 336688
rect 380710 336676 380716 336688
rect 380768 336676 380774 336728
rect 380986 336676 380992 336728
rect 381044 336716 381050 336728
rect 382090 336716 382096 336728
rect 381044 336688 382096 336716
rect 381044 336676 381050 336688
rect 382090 336676 382096 336688
rect 382148 336676 382154 336728
rect 383654 336676 383660 336728
rect 383712 336716 383718 336728
rect 384850 336716 384856 336728
rect 383712 336688 384856 336716
rect 383712 336676 383718 336688
rect 384850 336676 384856 336688
rect 384908 336676 384914 336728
rect 385862 336676 385868 336728
rect 385920 336716 385926 336728
rect 386322 336716 386328 336728
rect 385920 336688 386328 336716
rect 385920 336676 385926 336688
rect 386322 336676 386328 336688
rect 386380 336676 386386 336728
rect 386782 336676 386788 336728
rect 386840 336716 386846 336728
rect 387518 336716 387524 336728
rect 386840 336688 387524 336716
rect 386840 336676 386846 336688
rect 387518 336676 387524 336688
rect 387576 336676 387582 336728
rect 111702 336608 111708 336660
rect 111760 336648 111766 336660
rect 209590 336648 209596 336660
rect 111760 336620 209596 336648
rect 111760 336608 111766 336620
rect 209590 336608 209596 336620
rect 209648 336608 209654 336660
rect 231854 336648 231860 336660
rect 222856 336620 231860 336648
rect 222856 336592 222884 336620
rect 231854 336608 231860 336620
rect 231912 336608 231918 336660
rect 235902 336608 235908 336660
rect 235960 336648 235966 336660
rect 256786 336648 256792 336660
rect 235960 336620 256792 336648
rect 235960 336608 235966 336620
rect 256786 336608 256792 336620
rect 256844 336608 256850 336660
rect 258718 336608 258724 336660
rect 258776 336648 258782 336660
rect 264790 336648 264796 336660
rect 258776 336620 264796 336648
rect 258776 336608 258782 336620
rect 264790 336608 264796 336620
rect 264848 336608 264854 336660
rect 270586 336608 270592 336660
rect 270644 336648 270650 336660
rect 271874 336648 271880 336660
rect 270644 336620 271880 336648
rect 270644 336608 270650 336620
rect 271874 336608 271880 336620
rect 271932 336608 271938 336660
rect 277670 336608 277676 336660
rect 277728 336648 277734 336660
rect 278590 336648 278596 336660
rect 277728 336620 278596 336648
rect 277728 336608 277734 336620
rect 278590 336608 278596 336620
rect 278648 336608 278654 336660
rect 299474 336608 299480 336660
rect 299532 336648 299538 336660
rect 300670 336648 300676 336660
rect 299532 336620 300676 336648
rect 299532 336608 299538 336620
rect 300670 336608 300676 336620
rect 300728 336608 300734 336660
rect 301314 336608 301320 336660
rect 301372 336648 301378 336660
rect 302142 336648 302148 336660
rect 301372 336620 302148 336648
rect 301372 336608 301378 336620
rect 302142 336608 302148 336620
rect 302200 336608 302206 336660
rect 304442 336608 304448 336660
rect 304500 336648 304506 336660
rect 304902 336648 304908 336660
rect 304500 336620 304908 336648
rect 304500 336608 304506 336620
rect 304902 336608 304908 336620
rect 304960 336608 304966 336660
rect 305730 336608 305736 336660
rect 305788 336648 305794 336660
rect 306282 336648 306288 336660
rect 305788 336620 306288 336648
rect 305788 336608 305794 336620
rect 306282 336608 306288 336620
rect 306340 336608 306346 336660
rect 307110 336608 307116 336660
rect 307168 336648 307174 336660
rect 307662 336648 307668 336660
rect 307168 336620 307668 336648
rect 307168 336608 307174 336620
rect 307662 336608 307668 336620
rect 307720 336608 307726 336660
rect 308398 336608 308404 336660
rect 308456 336648 308462 336660
rect 309042 336648 309048 336660
rect 308456 336620 309048 336648
rect 308456 336608 308462 336620
rect 309042 336608 309048 336620
rect 309100 336608 309106 336660
rect 309778 336608 309784 336660
rect 309836 336648 309842 336660
rect 310422 336648 310428 336660
rect 309836 336620 310428 336648
rect 309836 336608 309842 336620
rect 310422 336608 310428 336620
rect 310480 336608 310486 336660
rect 311066 336608 311072 336660
rect 311124 336648 311130 336660
rect 311802 336648 311808 336660
rect 311124 336620 311808 336648
rect 311124 336608 311130 336620
rect 311802 336608 311808 336620
rect 311860 336608 311866 336660
rect 315114 336608 315120 336660
rect 315172 336648 315178 336660
rect 315942 336648 315948 336660
rect 315172 336620 315948 336648
rect 315172 336608 315178 336620
rect 315942 336608 315948 336620
rect 316000 336608 316006 336660
rect 323118 336608 323124 336660
rect 323176 336648 323182 336660
rect 411254 336648 411260 336660
rect 323176 336620 411260 336648
rect 323176 336608 323182 336620
rect 411254 336608 411260 336620
rect 411312 336608 411318 336660
rect 103422 336540 103428 336592
rect 103480 336580 103486 336592
rect 103480 336552 202092 336580
rect 103480 336540 103486 336552
rect 50338 336472 50344 336524
rect 50396 336512 50402 336524
rect 185486 336512 185492 336524
rect 50396 336484 185492 336512
rect 50396 336472 50402 336484
rect 185486 336472 185492 336484
rect 185544 336472 185550 336524
rect 202064 336512 202092 336552
rect 202138 336540 202144 336592
rect 202196 336580 202202 336592
rect 205082 336580 205088 336592
rect 202196 336552 205088 336580
rect 202196 336540 202202 336552
rect 205082 336540 205088 336552
rect 205140 336540 205146 336592
rect 222838 336540 222844 336592
rect 222896 336540 222902 336592
rect 231118 336540 231124 336592
rect 231176 336580 231182 336592
rect 254118 336580 254124 336592
rect 231176 336552 254124 336580
rect 231176 336540 231182 336552
rect 254118 336540 254124 336552
rect 254176 336540 254182 336592
rect 296806 336540 296812 336592
rect 296864 336580 296870 336592
rect 297910 336580 297916 336592
rect 296864 336552 297916 336580
rect 296864 336540 296870 336552
rect 297910 336540 297916 336552
rect 297968 336540 297974 336592
rect 313734 336540 313740 336592
rect 313792 336580 313798 336592
rect 314562 336580 314568 336592
rect 313792 336552 314568 336580
rect 313792 336540 313798 336552
rect 314562 336540 314568 336552
rect 314620 336540 314626 336592
rect 328454 336540 328460 336592
rect 328512 336580 328518 336592
rect 335173 336583 335231 336589
rect 335173 336580 335185 336583
rect 328512 336552 335185 336580
rect 328512 336540 328518 336552
rect 335173 336549 335185 336552
rect 335219 336549 335231 336583
rect 335173 336543 335231 336549
rect 335265 336583 335323 336589
rect 335265 336549 335277 336583
rect 335311 336580 335323 336583
rect 418154 336580 418160 336592
rect 335311 336552 418160 336580
rect 335311 336549 335323 336552
rect 335265 336543 335323 336549
rect 418154 336540 418160 336552
rect 418212 336540 418218 336592
rect 206922 336512 206928 336524
rect 202064 336484 206928 336512
rect 206922 336472 206928 336484
rect 206980 336472 206986 336524
rect 226978 336472 226984 336524
rect 227036 336512 227042 336524
rect 252738 336512 252744 336524
rect 227036 336484 252744 336512
rect 227036 336472 227042 336484
rect 252738 336472 252744 336484
rect 252796 336472 252802 336524
rect 331214 336472 331220 336524
rect 331272 336512 331278 336524
rect 331272 336484 340184 336512
rect 331272 336472 331278 336484
rect 43438 336404 43444 336456
rect 43496 336444 43502 336456
rect 182818 336444 182824 336456
rect 43496 336416 182824 336444
rect 43496 336404 43502 336416
rect 182818 336404 182824 336416
rect 182876 336404 182882 336456
rect 220722 336404 220728 336456
rect 220780 336444 220786 336456
rect 250990 336444 250996 336456
rect 220780 336416 250996 336444
rect 220780 336404 220786 336416
rect 250990 336404 250996 336416
rect 251048 336404 251054 336456
rect 298094 336404 298100 336456
rect 298152 336444 298158 336456
rect 318058 336444 318064 336456
rect 298152 336416 318064 336444
rect 298152 336404 298158 336416
rect 318058 336404 318064 336416
rect 318116 336404 318122 336456
rect 325786 336404 325792 336456
rect 325844 336444 325850 336456
rect 335265 336447 335323 336453
rect 335265 336444 335277 336447
rect 325844 336416 335277 336444
rect 325844 336404 325850 336416
rect 335265 336413 335277 336416
rect 335311 336413 335323 336447
rect 340156 336444 340184 336484
rect 342254 336472 342260 336524
rect 342312 336512 342318 336524
rect 343450 336512 343456 336524
rect 342312 336484 343456 336512
rect 342312 336472 342318 336484
rect 343450 336472 343456 336484
rect 343508 336472 343514 336524
rect 343545 336515 343603 336521
rect 343545 336481 343557 336515
rect 343591 336512 343603 336515
rect 425054 336512 425060 336524
rect 343591 336484 425060 336512
rect 343591 336481 343603 336484
rect 343545 336475 343603 336481
rect 425054 336472 425060 336484
rect 425112 336472 425118 336524
rect 431954 336444 431960 336456
rect 340156 336416 431960 336444
rect 335265 336407 335323 336413
rect 431954 336404 431960 336416
rect 432012 336404 432018 336456
rect 35158 336336 35164 336388
rect 35216 336376 35222 336388
rect 177022 336376 177028 336388
rect 35216 336348 177028 336376
rect 35216 336336 35222 336348
rect 177022 336336 177028 336348
rect 177080 336336 177086 336388
rect 213822 336336 213828 336388
rect 213880 336376 213886 336388
rect 248322 336376 248328 336388
rect 213880 336348 248328 336376
rect 213880 336336 213886 336348
rect 248322 336336 248328 336348
rect 248380 336336 248386 336388
rect 253290 336336 253296 336388
rect 253348 336376 253354 336388
rect 262122 336376 262128 336388
rect 253348 336348 262128 336376
rect 253348 336336 253354 336348
rect 262122 336336 262128 336348
rect 262180 336336 262186 336388
rect 287054 336336 287060 336388
rect 287112 336376 287118 336388
rect 288250 336376 288256 336388
rect 287112 336348 288256 336376
rect 287112 336336 287118 336348
rect 288250 336336 288256 336348
rect 288308 336336 288314 336388
rect 290642 336336 290648 336388
rect 290700 336376 290706 336388
rect 316678 336376 316684 336388
rect 290700 336348 316684 336376
rect 290700 336336 290706 336348
rect 316678 336336 316684 336348
rect 316736 336336 316742 336388
rect 333790 336336 333796 336388
rect 333848 336376 333854 336388
rect 440234 336376 440240 336388
rect 333848 336348 440240 336376
rect 333848 336336 333854 336348
rect 440234 336336 440240 336348
rect 440292 336336 440298 336388
rect 36538 336268 36544 336320
rect 36596 336308 36602 336320
rect 180150 336308 180156 336320
rect 36596 336280 180156 336308
rect 36596 336268 36602 336280
rect 180150 336268 180156 336280
rect 180208 336268 180214 336320
rect 219342 336268 219348 336320
rect 219400 336308 219406 336320
rect 250070 336308 250076 336320
rect 219400 336280 250076 336308
rect 219400 336268 219406 336280
rect 250070 336268 250076 336280
rect 250128 336268 250134 336320
rect 251818 336268 251824 336320
rect 251876 336308 251882 336320
rect 260742 336308 260748 336320
rect 251876 336280 260748 336308
rect 251876 336268 251882 336280
rect 260742 336268 260748 336280
rect 260800 336268 260806 336320
rect 278130 336268 278136 336320
rect 278188 336308 278194 336320
rect 291838 336308 291844 336320
rect 278188 336280 291844 336308
rect 278188 336268 278194 336280
rect 291838 336268 291844 336280
rect 291896 336268 291902 336320
rect 293310 336268 293316 336320
rect 293368 336308 293374 336320
rect 320818 336308 320824 336320
rect 293368 336280 320824 336308
rect 293368 336268 293374 336280
rect 320818 336268 320824 336280
rect 320876 336268 320882 336320
rect 335449 336311 335507 336317
rect 335449 336277 335461 336311
rect 335495 336308 335507 336311
rect 343545 336311 343603 336317
rect 343545 336308 343557 336311
rect 335495 336280 343557 336308
rect 335495 336277 335507 336280
rect 335449 336271 335507 336277
rect 343545 336277 343557 336280
rect 343591 336277 343603 336311
rect 343545 336271 343603 336277
rect 343637 336311 343695 336317
rect 343637 336277 343649 336311
rect 343683 336308 343695 336311
rect 447134 336308 447140 336320
rect 343683 336280 447140 336308
rect 343683 336277 343695 336280
rect 343637 336271 343695 336277
rect 447134 336268 447140 336280
rect 447192 336268 447198 336320
rect 32398 336200 32404 336252
rect 32456 336240 32462 336252
rect 177114 336240 177120 336252
rect 32456 336212 177120 336240
rect 32456 336200 32462 336212
rect 177114 336200 177120 336212
rect 177172 336200 177178 336252
rect 183554 336200 183560 336252
rect 183612 336240 183618 336252
rect 183830 336240 183836 336252
rect 183612 336212 183836 336240
rect 183612 336200 183618 336212
rect 183830 336200 183836 336212
rect 183888 336200 183894 336252
rect 212442 336200 212448 336252
rect 212500 336240 212506 336252
rect 247494 336240 247500 336252
rect 212500 336212 247500 336240
rect 212500 336200 212506 336212
rect 247494 336200 247500 336212
rect 247552 336200 247558 336252
rect 247678 336200 247684 336252
rect 247736 336240 247742 336252
rect 251450 336240 251456 336252
rect 247736 336212 251456 336240
rect 247736 336200 247742 336212
rect 251450 336200 251456 336212
rect 251508 336200 251514 336252
rect 253842 336200 253848 336252
rect 253900 336240 253906 336252
rect 263410 336240 263416 336252
rect 253900 336212 263416 336240
rect 253900 336200 253906 336212
rect 263410 336200 263416 336212
rect 263468 336200 263474 336252
rect 275462 336200 275468 336252
rect 275520 336240 275526 336252
rect 282178 336240 282184 336252
rect 275520 336212 282184 336240
rect 275520 336200 275526 336212
rect 282178 336200 282184 336212
rect 282236 336200 282242 336252
rect 286594 336200 286600 336252
rect 286652 336240 286658 336252
rect 313918 336240 313924 336252
rect 286652 336212 313924 336240
rect 286652 336200 286658 336212
rect 313918 336200 313924 336212
rect 313976 336200 313982 336252
rect 315574 336200 315580 336252
rect 315632 336240 315638 336252
rect 335998 336240 336004 336252
rect 315632 336212 336004 336240
rect 315632 336200 315638 336212
rect 335998 336200 336004 336212
rect 336056 336200 336062 336252
rect 341334 336200 341340 336252
rect 341392 336240 341398 336252
rect 342070 336240 342076 336252
rect 341392 336212 342076 336240
rect 341392 336200 341398 336212
rect 342070 336200 342076 336212
rect 342128 336200 342134 336252
rect 454034 336240 454040 336252
rect 342180 336212 454040 336240
rect 22738 336132 22744 336184
rect 22796 336172 22802 336184
rect 173894 336172 173900 336184
rect 22796 336144 173900 336172
rect 22796 336132 22802 336144
rect 173894 336132 173900 336144
rect 173952 336132 173958 336184
rect 210970 336132 210976 336184
rect 211028 336172 211034 336184
rect 246942 336172 246948 336184
rect 211028 336144 246948 336172
rect 211028 336132 211034 336144
rect 246942 336132 246948 336144
rect 247000 336132 247006 336184
rect 250530 336132 250536 336184
rect 250588 336172 250594 336184
rect 259454 336172 259460 336184
rect 250588 336144 259460 336172
rect 250588 336132 250594 336144
rect 259454 336132 259460 336144
rect 259512 336132 259518 336184
rect 260742 336132 260748 336184
rect 260800 336172 260806 336184
rect 266078 336172 266084 336184
rect 260800 336144 266084 336172
rect 260800 336132 260806 336144
rect 266078 336132 266084 336144
rect 266136 336132 266142 336184
rect 274542 336132 274548 336184
rect 274600 336172 274606 336184
rect 283190 336172 283196 336184
rect 274600 336144 283196 336172
rect 274600 336132 274606 336144
rect 283190 336132 283196 336144
rect 283248 336132 283254 336184
rect 287882 336132 287888 336184
rect 287940 336172 287946 336184
rect 317690 336172 317696 336184
rect 287940 336144 317696 336172
rect 287940 336132 287946 336144
rect 317690 336132 317696 336144
rect 317748 336132 317754 336184
rect 323578 336172 323584 336184
rect 319824 336144 323584 336172
rect 17218 336064 17224 336116
rect 17276 336104 17282 336116
rect 173526 336104 173532 336116
rect 17276 336076 173532 336104
rect 17276 336064 17282 336076
rect 173526 336064 173532 336076
rect 173584 336064 173590 336116
rect 177298 336064 177304 336116
rect 177356 336104 177362 336116
rect 202414 336104 202420 336116
rect 177356 336076 202420 336104
rect 177356 336064 177362 336076
rect 202414 336064 202420 336076
rect 202472 336064 202478 336116
rect 209682 336064 209688 336116
rect 209740 336104 209746 336116
rect 246482 336104 246488 336116
rect 209740 336076 246488 336104
rect 209740 336064 209746 336076
rect 246482 336064 246488 336076
rect 246540 336064 246546 336116
rect 249058 336064 249064 336116
rect 249116 336104 249122 336116
rect 258074 336104 258080 336116
rect 249116 336076 258080 336104
rect 249116 336064 249122 336076
rect 258074 336064 258080 336076
rect 258132 336064 258138 336116
rect 275002 336064 275008 336116
rect 275060 336104 275066 336116
rect 284478 336104 284484 336116
rect 275060 336076 284484 336104
rect 275060 336064 275066 336076
rect 284478 336064 284484 336076
rect 284536 336064 284542 336116
rect 290182 336064 290188 336116
rect 290240 336104 290246 336116
rect 319824 336104 319852 336144
rect 323578 336132 323584 336144
rect 323636 336132 323642 336184
rect 290240 336076 319852 336104
rect 290240 336064 290246 336076
rect 321738 336064 321744 336116
rect 321796 336104 321802 336116
rect 322842 336104 322848 336116
rect 321796 336076 322848 336104
rect 321796 336064 321802 336076
rect 322842 336064 322848 336076
rect 322900 336064 322906 336116
rect 339126 336064 339132 336116
rect 339184 336104 339190 336116
rect 342180 336104 342208 336212
rect 454034 336200 454040 336212
rect 454092 336200 454098 336252
rect 460934 336172 460940 336184
rect 339184 336076 342208 336104
rect 343744 336144 460940 336172
rect 339184 336064 339190 336076
rect 7558 335996 7564 336048
rect 7616 336036 7622 336048
rect 170398 336036 170404 336048
rect 7616 336008 170404 336036
rect 7616 335996 7622 336008
rect 170398 335996 170404 336008
rect 170456 335996 170462 336048
rect 173158 335996 173164 336048
rect 173216 336036 173222 336048
rect 199746 336036 199752 336048
rect 173216 336008 199752 336036
rect 173216 335996 173222 336008
rect 199746 335996 199752 336008
rect 199804 335996 199810 336048
rect 206922 335996 206928 336048
rect 206980 336036 206986 336048
rect 245654 336036 245660 336048
rect 206980 336008 245660 336036
rect 206980 335996 206986 336008
rect 245654 335996 245660 336008
rect 245712 335996 245718 336048
rect 248322 335996 248328 336048
rect 248380 336036 248386 336048
rect 261202 336036 261208 336048
rect 248380 336008 261208 336036
rect 248380 335996 248386 336008
rect 261202 335996 261208 336008
rect 261260 335996 261266 336048
rect 275922 335996 275928 336048
rect 275980 336036 275986 336048
rect 275980 336008 277394 336036
rect 275980 335996 275986 336008
rect 121362 335928 121368 335980
rect 121420 335968 121426 335980
rect 213546 335968 213552 335980
rect 121420 335940 213552 335968
rect 121420 335928 121426 335940
rect 213546 335928 213552 335940
rect 213604 335928 213610 335980
rect 229738 335928 229744 335980
rect 229796 335968 229802 335980
rect 231394 335968 231400 335980
rect 229796 335940 231400 335968
rect 229796 335928 229802 335940
rect 231394 335928 231400 335940
rect 231452 335928 231458 335980
rect 250438 335928 250444 335980
rect 250496 335968 250502 335980
rect 257246 335968 257252 335980
rect 250496 335940 257252 335968
rect 250496 335928 250502 335940
rect 257246 335928 257252 335940
rect 257304 335928 257310 335980
rect 265710 335928 265716 335980
rect 265768 335968 265774 335980
rect 266630 335968 266636 335980
rect 265768 335940 266636 335968
rect 265768 335928 265774 335940
rect 266630 335928 266636 335940
rect 266688 335928 266694 335980
rect 277366 335968 277394 336008
rect 285674 335996 285680 336048
rect 285732 336036 285738 336048
rect 286962 336036 286968 336048
rect 285732 336008 286968 336036
rect 285732 335996 285738 336008
rect 286962 335996 286968 336008
rect 287020 335996 287026 336048
rect 291930 335996 291936 336048
rect 291988 336036 291994 336048
rect 328546 336036 328552 336048
rect 291988 336008 328552 336036
rect 291988 335996 291994 336008
rect 328546 335996 328552 336008
rect 328604 335996 328610 336048
rect 336458 335996 336464 336048
rect 336516 336036 336522 336048
rect 343637 336039 343695 336045
rect 343637 336036 343649 336039
rect 336516 336008 343649 336036
rect 336516 335996 336522 336008
rect 343637 336005 343649 336008
rect 343683 336005 343695 336039
rect 343637 335999 343695 336005
rect 285766 335968 285772 335980
rect 277366 335940 285772 335968
rect 285766 335928 285772 335940
rect 285824 335928 285830 335980
rect 294138 335928 294144 335980
rect 294196 335968 294202 335980
rect 295058 335968 295064 335980
rect 294196 335940 295064 335968
rect 294196 335928 294202 335940
rect 295058 335928 295064 335940
rect 295116 335928 295122 335980
rect 341794 335928 341800 335980
rect 341852 335968 341858 335980
rect 343744 335968 343772 336144
rect 460934 336132 460940 336144
rect 460992 336132 460998 336184
rect 344462 336064 344468 336116
rect 344520 336104 344526 336116
rect 467834 336104 467840 336116
rect 344520 336076 467840 336104
rect 344520 336064 344526 336076
rect 467834 336064 467840 336076
rect 467892 336064 467898 336116
rect 345842 335996 345848 336048
rect 345900 336036 345906 336048
rect 346302 336036 346308 336048
rect 345900 336008 346308 336036
rect 345900 335996 345906 336008
rect 346302 335996 346308 336008
rect 346360 335996 346366 336048
rect 348510 335996 348516 336048
rect 348568 336036 348574 336048
rect 349062 336036 349068 336048
rect 348568 336008 349068 336036
rect 348568 335996 348574 336008
rect 349062 335996 349068 336008
rect 349120 335996 349126 336048
rect 353386 335996 353392 336048
rect 353444 336036 353450 336048
rect 354490 336036 354496 336048
rect 353444 336008 354496 336036
rect 353444 335996 353450 336008
rect 354490 335996 354496 336008
rect 354548 335996 354554 336048
rect 474734 336036 474740 336048
rect 354646 336008 474740 336036
rect 341852 335940 343772 335968
rect 341852 335928 341858 335940
rect 347130 335928 347136 335980
rect 347188 335968 347194 335980
rect 354646 335968 354674 336008
rect 474734 335996 474740 336008
rect 474792 335996 474798 336048
rect 347188 335940 354674 335968
rect 347188 335928 347194 335940
rect 360930 335928 360936 335980
rect 360988 335968 360994 335980
rect 361482 335968 361488 335980
rect 360988 335940 361488 335968
rect 360988 335928 360994 335940
rect 361482 335928 361488 335940
rect 361540 335928 361546 335980
rect 363598 335928 363604 335980
rect 363656 335968 363662 335980
rect 364242 335968 364248 335980
rect 363656 335940 364248 335968
rect 363656 335928 363662 335940
rect 364242 335928 364248 335940
rect 364300 335928 364306 335980
rect 364978 335928 364984 335980
rect 365036 335968 365042 335980
rect 365622 335968 365628 335980
rect 365036 335940 365628 335968
rect 365036 335928 365042 335940
rect 365622 335928 365628 335940
rect 365680 335928 365686 335980
rect 366266 335928 366272 335980
rect 366324 335968 366330 335980
rect 367002 335968 367008 335980
rect 366324 335940 367008 335968
rect 366324 335928 366330 335940
rect 367002 335928 367008 335940
rect 367060 335928 367066 335980
rect 367646 335928 367652 335980
rect 367704 335968 367710 335980
rect 368382 335968 368388 335980
rect 367704 335940 368388 335968
rect 367704 335928 367710 335940
rect 368382 335928 368388 335940
rect 368440 335928 368446 335980
rect 368566 335928 368572 335980
rect 368624 335968 368630 335980
rect 369578 335968 369584 335980
rect 368624 335940 369584 335968
rect 368624 335928 368630 335940
rect 369578 335928 369584 335940
rect 369636 335928 369642 335980
rect 370314 335928 370320 335980
rect 370372 335968 370378 335980
rect 371142 335968 371148 335980
rect 370372 335940 371148 335968
rect 370372 335928 370378 335940
rect 371142 335928 371148 335940
rect 371200 335928 371206 335980
rect 378318 335928 378324 335980
rect 378376 335968 378382 335980
rect 379422 335968 379428 335980
rect 378376 335940 379428 335968
rect 378376 335928 378382 335940
rect 379422 335928 379428 335940
rect 379480 335928 379486 335980
rect 379698 335928 379704 335980
rect 379756 335968 379762 335980
rect 380802 335968 380808 335980
rect 379756 335940 380808 335968
rect 379756 335928 379762 335940
rect 380802 335928 380808 335940
rect 380860 335928 380866 335980
rect 385034 335928 385040 335980
rect 385092 335968 385098 335980
rect 386138 335968 386144 335980
rect 385092 335940 386144 335968
rect 385092 335928 385098 335940
rect 386138 335928 386144 335940
rect 386196 335928 386202 335980
rect 288802 335860 288808 335912
rect 288860 335900 288866 335912
rect 289722 335900 289728 335912
rect 288860 335872 289728 335900
rect 288860 335860 288866 335872
rect 289722 335860 289728 335872
rect 289780 335860 289786 335912
rect 311986 335860 311992 335912
rect 312044 335900 312050 335912
rect 312998 335900 313004 335912
rect 312044 335872 313004 335900
rect 312044 335860 312050 335872
rect 312998 335860 313004 335872
rect 313056 335860 313062 335912
rect 344002 335860 344008 335912
rect 344060 335900 344066 335912
rect 344830 335900 344836 335912
rect 344060 335872 344836 335900
rect 344060 335860 344066 335872
rect 344830 335860 344836 335872
rect 344888 335860 344894 335912
rect 354674 335860 354680 335912
rect 354732 335900 354738 335912
rect 355778 335900 355784 335912
rect 354732 335872 355784 335900
rect 354732 335860 354738 335872
rect 355778 335860 355784 335872
rect 355836 335860 355842 335912
rect 358262 335860 358268 335912
rect 358320 335900 358326 335912
rect 358722 335900 358728 335912
rect 358320 335872 358728 335900
rect 358320 335860 358326 335872
rect 358722 335860 358728 335872
rect 358780 335860 358786 335912
rect 382366 335860 382372 335912
rect 382424 335900 382430 335912
rect 383470 335900 383476 335912
rect 382424 335872 383476 335900
rect 382424 335860 382430 335872
rect 383470 335860 383476 335872
rect 383528 335860 383534 335912
rect 265618 335792 265624 335844
rect 265676 335832 265682 335844
rect 266538 335832 266544 335844
rect 265676 335804 266544 335832
rect 265676 335792 265682 335804
rect 266538 335792 266544 335804
rect 266596 335792 266602 335844
rect 327074 335792 327080 335844
rect 327132 335832 327138 335844
rect 328362 335832 328368 335844
rect 327132 335804 328368 335832
rect 327132 335792 327138 335804
rect 328362 335792 328368 335804
rect 328420 335792 328426 335844
rect 266998 335724 267004 335776
rect 267056 335764 267062 335776
rect 267918 335764 267924 335776
rect 267056 335736 267924 335764
rect 267056 335724 267062 335736
rect 267918 335724 267924 335736
rect 267976 335724 267982 335776
rect 272334 335656 272340 335708
rect 272392 335696 272398 335708
rect 275278 335696 275284 335708
rect 272392 335668 275284 335696
rect 272392 335656 272398 335668
rect 275278 335656 275284 335668
rect 275336 335656 275342 335708
rect 302602 335656 302608 335708
rect 302660 335696 302666 335708
rect 303522 335696 303528 335708
rect 302660 335668 303528 335696
rect 302660 335656 302666 335668
rect 303522 335656 303528 335668
rect 303580 335656 303586 335708
rect 242250 335588 242256 335640
rect 242308 335628 242314 335640
rect 242986 335628 242992 335640
rect 242308 335600 242992 335628
rect 242308 335588 242314 335600
rect 242986 335588 242992 335600
rect 243044 335588 243050 335640
rect 252002 335588 252008 335640
rect 252060 335628 252066 335640
rect 258534 335628 258540 335640
rect 252060 335600 258540 335628
rect 252060 335588 252066 335600
rect 258534 335588 258540 335600
rect 258592 335588 258598 335640
rect 259362 335588 259368 335640
rect 259420 335628 259426 335640
rect 265250 335628 265256 335640
rect 259420 335600 265256 335628
rect 259420 335588 259426 335600
rect 265250 335588 265256 335600
rect 265308 335588 265314 335640
rect 362310 335588 362316 335640
rect 362368 335628 362374 335640
rect 362862 335628 362868 335640
rect 362368 335600 362868 335628
rect 362368 335588 362374 335600
rect 362862 335588 362868 335600
rect 362920 335588 362926 335640
rect 376110 335588 376116 335640
rect 376168 335628 376174 335640
rect 376570 335628 376576 335640
rect 376168 335600 376576 335628
rect 376168 335588 376174 335600
rect 376570 335588 376576 335600
rect 376628 335588 376634 335640
rect 272794 335520 272800 335572
rect 272852 335560 272858 335572
rect 277578 335560 277584 335572
rect 272852 335532 277584 335560
rect 272852 335520 272858 335532
rect 277578 335520 277584 335532
rect 277636 335520 277642 335572
rect 284386 335520 284392 335572
rect 284444 335560 284450 335572
rect 285582 335560 285588 335572
rect 284444 335532 285588 335560
rect 284444 335520 284450 335532
rect 285582 335520 285588 335532
rect 285640 335520 285646 335572
rect 295518 335520 295524 335572
rect 295576 335560 295582 335572
rect 296438 335560 296444 335572
rect 295576 335532 296444 335560
rect 295576 335520 295582 335532
rect 296438 335520 296444 335532
rect 296496 335520 296502 335572
rect 298186 335520 298192 335572
rect 298244 335560 298250 335572
rect 299290 335560 299296 335572
rect 298244 335532 299296 335560
rect 298244 335520 298250 335532
rect 299290 335520 299296 335532
rect 299348 335520 299354 335572
rect 374270 335520 374276 335572
rect 374328 335560 374334 335572
rect 375282 335560 375288 335572
rect 374328 335532 375288 335560
rect 374328 335520 374334 335532
rect 375282 335520 375288 335532
rect 375340 335520 375346 335572
rect 273254 335452 273260 335504
rect 273312 335492 273318 335504
rect 274542 335492 274548 335504
rect 273312 335464 274548 335492
rect 273312 335452 273318 335464
rect 274542 335452 274548 335464
rect 274600 335452 274606 335504
rect 236638 335384 236644 335436
rect 236696 335424 236702 335436
rect 239858 335424 239864 335436
rect 236696 335396 239864 335424
rect 236696 335384 236702 335396
rect 239858 335384 239864 335396
rect 239916 335384 239922 335436
rect 283006 335384 283012 335436
rect 283064 335424 283070 335436
rect 284202 335424 284208 335436
rect 283064 335396 284208 335424
rect 283064 335384 283070 335396
rect 284202 335384 284208 335396
rect 284260 335384 284266 335436
rect 346670 335384 346676 335436
rect 346728 335424 346734 335436
rect 347590 335424 347596 335436
rect 346728 335396 347596 335424
rect 346728 335384 346734 335396
rect 347590 335384 347596 335396
rect 347648 335384 347654 335436
rect 349338 335384 349344 335436
rect 349396 335424 349402 335436
rect 350258 335424 350264 335436
rect 349396 335396 350264 335424
rect 349396 335384 349402 335396
rect 350258 335384 350264 335396
rect 350316 335384 350322 335436
rect 246298 335316 246304 335368
rect 246356 335356 246362 335368
rect 248782 335356 248788 335368
rect 246356 335328 248788 335356
rect 246356 335316 246362 335328
rect 248782 335316 248788 335328
rect 248840 335316 248846 335368
rect 253198 335316 253204 335368
rect 253256 335356 253262 335368
rect 259914 335356 259920 335368
rect 253256 335328 259920 335356
rect 253256 335316 253262 335328
rect 259914 335316 259920 335328
rect 259972 335316 259978 335368
rect 126882 334636 126888 334688
rect 126940 334676 126946 334688
rect 215386 334676 215392 334688
rect 126940 334648 215392 334676
rect 126940 334636 126946 334648
rect 215386 334636 215392 334648
rect 215444 334636 215450 334688
rect 318610 334636 318616 334688
rect 318668 334676 318674 334688
rect 398834 334676 398840 334688
rect 318668 334648 398840 334676
rect 318668 334636 318674 334648
rect 398834 334636 398840 334648
rect 398892 334636 398898 334688
rect 25498 334568 25504 334620
rect 25556 334608 25562 334620
rect 176562 334608 176568 334620
rect 25556 334580 176568 334608
rect 25556 334568 25562 334580
rect 176562 334568 176568 334580
rect 176620 334568 176626 334620
rect 180702 334568 180708 334620
rect 180760 334608 180766 334620
rect 235810 334608 235816 334620
rect 180760 334580 235816 334608
rect 180760 334568 180766 334580
rect 235810 334568 235816 334580
rect 235868 334568 235874 334620
rect 350442 334568 350448 334620
rect 350500 334608 350506 334620
rect 483014 334608 483020 334620
rect 350500 334580 483020 334608
rect 350500 334568 350506 334580
rect 483014 334568 483020 334580
rect 483072 334568 483078 334620
rect 161382 333276 161388 333328
rect 161440 333316 161446 333328
rect 228726 333316 228732 333328
rect 161440 333288 228732 333316
rect 161440 333276 161446 333288
rect 228726 333276 228732 333288
rect 228784 333276 228790 333328
rect 352926 333276 352932 333328
rect 352984 333316 352990 333328
rect 489914 333316 489920 333328
rect 352984 333288 489920 333316
rect 352984 333276 352990 333288
rect 489914 333276 489920 333288
rect 489972 333276 489978 333328
rect 135162 333208 135168 333260
rect 135220 333248 135226 333260
rect 218422 333248 218428 333260
rect 135220 333220 218428 333248
rect 135220 333208 135226 333220
rect 218422 333208 218428 333220
rect 218480 333208 218486 333260
rect 539594 333248 539600 333260
rect 373966 333220 539600 333248
rect 371234 333140 371240 333192
rect 371292 333180 371298 333192
rect 373966 333180 373994 333220
rect 539594 333208 539600 333220
rect 539652 333208 539658 333260
rect 371292 333152 373994 333180
rect 371292 333140 371298 333152
rect 3050 332528 3056 332580
rect 3108 332568 3114 332580
rect 166902 332568 166908 332580
rect 3108 332540 166908 332568
rect 3108 332528 3114 332540
rect 166902 332528 166908 332540
rect 166960 332528 166966 332580
rect 356974 331916 356980 331968
rect 357032 331956 357038 331968
rect 500954 331956 500960 331968
rect 357032 331928 500960 331956
rect 357032 331916 357038 331928
rect 500954 331916 500960 331928
rect 501012 331916 501018 331968
rect 136542 331848 136548 331900
rect 136600 331888 136606 331900
rect 218974 331888 218980 331900
rect 136600 331860 218980 331888
rect 136600 331848 136606 331860
rect 218974 331848 218980 331860
rect 219032 331848 219038 331900
rect 377858 331848 377864 331900
rect 377916 331888 377922 331900
rect 556154 331888 556160 331900
rect 377916 331860 556160 331888
rect 377916 331848 377922 331860
rect 556154 331848 556160 331860
rect 556212 331848 556218 331900
rect 187878 331168 187884 331220
rect 187936 331208 187942 331220
rect 188062 331208 188068 331220
rect 187936 331180 188068 331208
rect 187936 331168 187942 331180
rect 188062 331168 188068 331180
rect 188120 331168 188126 331220
rect 200390 331168 200396 331220
rect 200448 331208 200454 331220
rect 200574 331208 200580 331220
rect 200448 331180 200580 331208
rect 200448 331168 200454 331180
rect 200574 331168 200580 331180
rect 200632 331168 200638 331220
rect 203150 331168 203156 331220
rect 203208 331208 203214 331220
rect 203334 331208 203340 331220
rect 203208 331180 203340 331208
rect 203208 331168 203214 331180
rect 203334 331168 203340 331180
rect 203392 331168 203398 331220
rect 373258 330692 373264 330744
rect 373316 330732 373322 330744
rect 373902 330732 373908 330744
rect 373316 330704 373908 330732
rect 373316 330692 373322 330704
rect 373902 330692 373908 330704
rect 373960 330692 373966 330744
rect 165522 330624 165528 330676
rect 165580 330664 165586 330676
rect 230014 330664 230020 330676
rect 165580 330636 230020 330664
rect 165580 330624 165586 330636
rect 230014 330624 230020 330636
rect 230072 330624 230078 330676
rect 155862 330556 155868 330608
rect 155920 330596 155926 330608
rect 226334 330596 226340 330608
rect 155920 330568 226340 330596
rect 155920 330556 155926 330568
rect 226334 330556 226340 330568
rect 226392 330556 226398 330608
rect 15838 330488 15844 330540
rect 15896 330528 15902 330540
rect 171686 330528 171692 330540
rect 15896 330500 171692 330528
rect 15896 330488 15902 330500
rect 171686 330488 171692 330500
rect 171744 330488 171750 330540
rect 172606 330488 172612 330540
rect 172664 330528 172670 330540
rect 172790 330528 172796 330540
rect 172664 330500 172796 330528
rect 172664 330488 172670 330500
rect 172790 330488 172796 330500
rect 172848 330488 172854 330540
rect 173986 330488 173992 330540
rect 174044 330528 174050 330540
rect 174446 330528 174452 330540
rect 174044 330500 174452 330528
rect 174044 330488 174050 330500
rect 174446 330488 174452 330500
rect 174504 330488 174510 330540
rect 175458 330488 175464 330540
rect 175516 330528 175522 330540
rect 175918 330528 175924 330540
rect 175516 330500 175924 330528
rect 175516 330488 175522 330500
rect 175918 330488 175924 330500
rect 175976 330488 175982 330540
rect 178126 330488 178132 330540
rect 178184 330528 178190 330540
rect 179046 330528 179052 330540
rect 178184 330500 179052 330528
rect 178184 330488 178190 330500
rect 179046 330488 179052 330500
rect 179104 330488 179110 330540
rect 248506 330488 248512 330540
rect 248564 330528 248570 330540
rect 249334 330528 249340 330540
rect 248564 330500 249340 330528
rect 248564 330488 248570 330500
rect 249334 330488 249340 330500
rect 249392 330488 249398 330540
rect 251266 330488 251272 330540
rect 251324 330528 251330 330540
rect 251910 330528 251916 330540
rect 251324 330500 251916 330528
rect 251324 330488 251330 330500
rect 251910 330488 251916 330500
rect 251968 330488 251974 330540
rect 252646 330488 252652 330540
rect 252704 330528 252710 330540
rect 253382 330528 253388 330540
rect 252704 330500 253388 330528
rect 252704 330488 252710 330500
rect 253382 330488 253388 330500
rect 253440 330488 253446 330540
rect 301774 330488 301780 330540
rect 301832 330528 301838 330540
rect 354674 330528 354680 330540
rect 301832 330500 354680 330528
rect 301832 330488 301838 330500
rect 354674 330488 354680 330500
rect 354732 330488 354738 330540
rect 359642 330488 359648 330540
rect 359700 330528 359706 330540
rect 507854 330528 507860 330540
rect 359700 330500 507860 330528
rect 359700 330488 359706 330500
rect 507854 330488 507860 330500
rect 507912 330488 507918 330540
rect 169846 330420 169852 330472
rect 169904 330460 169910 330472
rect 170582 330460 170588 330472
rect 169904 330432 170588 330460
rect 169904 330420 169910 330432
rect 170582 330420 170588 330432
rect 170640 330420 170646 330472
rect 133782 329128 133788 329180
rect 133840 329168 133846 329180
rect 218054 329168 218060 329180
rect 133840 329140 218060 329168
rect 133840 329128 133846 329140
rect 218054 329128 218060 329140
rect 218112 329128 218118 329180
rect 314194 329128 314200 329180
rect 314252 329168 314258 329180
rect 387794 329168 387800 329180
rect 314252 329140 387800 329168
rect 314252 329128 314258 329140
rect 387794 329128 387800 329140
rect 387852 329128 387858 329180
rect 113082 329060 113088 329112
rect 113140 329100 113146 329112
rect 210418 329100 210424 329112
rect 113140 329072 210424 329100
rect 113140 329060 113146 329072
rect 210418 329060 210424 329072
rect 210476 329060 210482 329112
rect 357434 329060 357440 329112
rect 357492 329100 357498 329112
rect 502334 329100 502340 329112
rect 357492 329072 502340 329100
rect 357492 329060 357498 329072
rect 502334 329060 502340 329072
rect 502392 329060 502398 329112
rect 180886 328924 180892 328976
rect 180944 328964 180950 328976
rect 181622 328964 181628 328976
rect 180944 328936 181628 328964
rect 180944 328924 180950 328936
rect 181622 328924 181628 328936
rect 181680 328924 181686 328976
rect 129642 327768 129648 327820
rect 129700 327808 129706 327820
rect 216674 327808 216680 327820
rect 129700 327780 216680 327808
rect 129700 327768 129706 327780
rect 216674 327768 216680 327780
rect 216732 327768 216738 327820
rect 317138 327768 317144 327820
rect 317196 327808 317202 327820
rect 394694 327808 394700 327820
rect 317196 327780 394700 327808
rect 317196 327768 317202 327780
rect 394694 327768 394700 327780
rect 394752 327768 394758 327820
rect 46198 327700 46204 327752
rect 46256 327740 46262 327752
rect 183738 327740 183744 327752
rect 46256 327712 183744 327740
rect 46256 327700 46262 327712
rect 183738 327700 183744 327712
rect 183796 327700 183802 327752
rect 351546 327700 351552 327752
rect 351604 327740 351610 327752
rect 485774 327740 485780 327752
rect 351604 327712 485780 327740
rect 351604 327700 351610 327712
rect 485774 327700 485780 327712
rect 485832 327700 485838 327752
rect 212718 326516 212724 326528
rect 212679 326488 212724 326516
rect 212718 326476 212724 326488
rect 212776 326476 212782 326528
rect 223758 326516 223764 326528
rect 223719 326488 223764 326516
rect 223758 326476 223764 326488
rect 223816 326476 223822 326528
rect 140682 326408 140688 326460
rect 140740 326448 140746 326460
rect 220354 326448 220360 326460
rect 140740 326420 220360 326448
rect 140740 326408 140746 326420
rect 220354 326408 220360 326420
rect 220412 326408 220418 326460
rect 224954 326408 224960 326460
rect 225012 326448 225018 326460
rect 225782 326448 225788 326460
rect 225012 326420 225788 326448
rect 225012 326408 225018 326420
rect 225782 326408 225788 326420
rect 225840 326408 225846 326460
rect 229278 326408 229284 326460
rect 229336 326408 229342 326460
rect 262398 326408 262404 326460
rect 262456 326408 262462 326460
rect 269206 326408 269212 326460
rect 269264 326408 269270 326460
rect 318518 326408 318524 326460
rect 318576 326448 318582 326460
rect 398926 326448 398932 326460
rect 318576 326420 398932 326448
rect 318576 326408 318582 326420
rect 398926 326408 398932 326420
rect 398984 326408 398990 326460
rect 39298 326340 39304 326392
rect 39356 326380 39362 326392
rect 180978 326380 180984 326392
rect 39356 326352 180984 326380
rect 39356 326340 39362 326352
rect 180978 326340 180984 326352
rect 181036 326340 181042 326392
rect 186314 326340 186320 326392
rect 186372 326380 186378 326392
rect 186958 326380 186964 326392
rect 186372 326352 186964 326380
rect 186372 326340 186378 326352
rect 186958 326340 186964 326352
rect 187016 326340 187022 326392
rect 187786 326340 187792 326392
rect 187844 326380 187850 326392
rect 188246 326380 188252 326392
rect 187844 326352 188252 326380
rect 187844 326340 187850 326352
rect 188246 326340 188252 326352
rect 188304 326340 188310 326392
rect 189166 326340 189172 326392
rect 189224 326380 189230 326392
rect 189718 326380 189724 326392
rect 189224 326352 189724 326380
rect 189224 326340 189230 326352
rect 189718 326340 189724 326352
rect 189776 326340 189782 326392
rect 190454 326340 190460 326392
rect 190512 326380 190518 326392
rect 190730 326380 190736 326392
rect 190512 326352 190736 326380
rect 190512 326340 190518 326352
rect 190730 326340 190736 326352
rect 190788 326340 190794 326392
rect 200298 326340 200304 326392
rect 200356 326380 200362 326392
rect 200758 326380 200764 326392
rect 200356 326352 200764 326380
rect 200356 326340 200362 326352
rect 200758 326340 200764 326352
rect 200816 326340 200822 326392
rect 203058 326340 203064 326392
rect 203116 326380 203122 326392
rect 203518 326380 203524 326392
rect 203116 326352 203524 326380
rect 203116 326340 203122 326352
rect 203518 326340 203524 326352
rect 203576 326340 203582 326392
rect 204346 326340 204352 326392
rect 204404 326380 204410 326392
rect 205174 326380 205180 326392
rect 204404 326352 205180 326380
rect 204404 326340 204410 326352
rect 205174 326340 205180 326352
rect 205232 326340 205238 326392
rect 205726 326340 205732 326392
rect 205784 326380 205790 326392
rect 206094 326380 206100 326392
rect 205784 326352 206100 326380
rect 205784 326340 205790 326352
rect 206094 326340 206100 326352
rect 206152 326340 206158 326392
rect 211246 326340 211252 326392
rect 211304 326380 211310 326392
rect 211430 326380 211436 326392
rect 211304 326352 211436 326380
rect 211304 326340 211310 326352
rect 211430 326340 211436 326352
rect 211488 326340 211494 326392
rect 215386 326340 215392 326392
rect 215444 326380 215450 326392
rect 215846 326380 215852 326392
rect 215444 326352 215852 326380
rect 215444 326340 215450 326352
rect 215846 326340 215852 326352
rect 215904 326340 215910 326392
rect 219434 326340 219440 326392
rect 219492 326380 219498 326392
rect 219894 326380 219900 326392
rect 219492 326352 219900 326380
rect 219492 326340 219498 326352
rect 219894 326340 219900 326352
rect 219952 326340 219958 326392
rect 223574 326340 223580 326392
rect 223632 326380 223638 326392
rect 224310 326380 224316 326392
rect 223632 326352 224316 326380
rect 223632 326340 223638 326352
rect 224310 326340 224316 326352
rect 224368 326340 224374 326392
rect 225046 326340 225052 326392
rect 225104 326380 225110 326392
rect 225230 326380 225236 326392
rect 225104 326352 225236 326380
rect 225104 326340 225110 326352
rect 225230 326340 225236 326352
rect 225288 326340 225294 326392
rect 227806 326340 227812 326392
rect 227864 326380 227870 326392
rect 227990 326380 227996 326392
rect 227864 326352 227996 326380
rect 227864 326340 227870 326352
rect 227990 326340 227996 326352
rect 228048 326340 228054 326392
rect 204438 326272 204444 326324
rect 204496 326312 204502 326324
rect 204622 326312 204628 326324
rect 204496 326284 204628 326312
rect 204496 326272 204502 326284
rect 204622 326272 204628 326284
rect 204680 326272 204686 326324
rect 229296 326256 229324 326408
rect 230566 326340 230572 326392
rect 230624 326380 230630 326392
rect 230750 326380 230756 326392
rect 230624 326352 230756 326380
rect 230624 326340 230630 326352
rect 230750 326340 230756 326352
rect 230808 326340 230814 326392
rect 231946 326340 231952 326392
rect 232004 326380 232010 326392
rect 232406 326380 232412 326392
rect 232004 326352 232412 326380
rect 232004 326340 232010 326352
rect 232406 326340 232412 326352
rect 232464 326340 232470 326392
rect 233418 326340 233424 326392
rect 233476 326380 233482 326392
rect 234246 326380 234252 326392
rect 233476 326352 234252 326380
rect 233476 326340 233482 326352
rect 234246 326340 234252 326352
rect 234304 326340 234310 326392
rect 241606 326340 241612 326392
rect 241664 326380 241670 326392
rect 242158 326380 242164 326392
rect 241664 326352 242164 326380
rect 241664 326340 241670 326352
rect 242158 326340 242164 326352
rect 242216 326340 242222 326392
rect 242986 326340 242992 326392
rect 243044 326380 243050 326392
rect 243446 326380 243452 326392
rect 243044 326352 243452 326380
rect 243044 326340 243050 326352
rect 243446 326340 243452 326352
rect 243504 326340 243510 326392
rect 255406 326340 255412 326392
rect 255464 326380 255470 326392
rect 255958 326380 255964 326392
rect 255464 326352 255964 326380
rect 255464 326340 255470 326352
rect 255958 326340 255964 326352
rect 256016 326340 256022 326392
rect 262416 326256 262444 326408
rect 267826 326340 267832 326392
rect 267884 326380 267890 326392
rect 268470 326380 268476 326392
rect 267884 326352 268476 326380
rect 267884 326340 267890 326352
rect 268470 326340 268476 326352
rect 268528 326340 268534 326392
rect 269224 326256 269252 326408
rect 354214 326340 354220 326392
rect 354272 326380 354278 326392
rect 492674 326380 492680 326392
rect 354272 326352 492680 326380
rect 354272 326340 354278 326352
rect 492674 326340 492680 326352
rect 492732 326340 492738 326392
rect 190546 326204 190552 326256
rect 190604 326244 190610 326256
rect 191006 326244 191012 326256
rect 190604 326216 191012 326244
rect 190604 326204 190610 326216
rect 191006 326204 191012 326216
rect 191064 326204 191070 326256
rect 229278 326204 229284 326256
rect 229336 326204 229342 326256
rect 262398 326204 262404 326256
rect 262456 326204 262462 326256
rect 269206 326204 269212 326256
rect 269264 326204 269270 326256
rect 232038 325864 232044 325916
rect 232096 325904 232102 325916
rect 232774 325904 232780 325916
rect 232096 325876 232780 325904
rect 232096 325864 232102 325876
rect 232774 325864 232780 325876
rect 232832 325864 232838 325916
rect 389174 325592 389180 325644
rect 389232 325632 389238 325644
rect 579890 325632 579896 325644
rect 389232 325604 579896 325632
rect 389232 325592 389238 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 144822 324980 144828 325032
rect 144880 325020 144886 325032
rect 221642 325020 221648 325032
rect 144880 324992 221648 325020
rect 144880 324980 144886 324992
rect 221642 324980 221648 324992
rect 221700 324980 221706 325032
rect 33778 324912 33784 324964
rect 33836 324952 33842 324964
rect 179506 324952 179512 324964
rect 33836 324924 179512 324952
rect 33836 324912 33842 324924
rect 179506 324912 179512 324924
rect 179564 324912 179570 324964
rect 317230 324912 317236 324964
rect 317288 324952 317294 324964
rect 396074 324952 396080 324964
rect 317288 324924 396080 324952
rect 317288 324912 317294 324924
rect 396074 324912 396080 324924
rect 396132 324912 396138 324964
rect 208486 324368 208492 324420
rect 208544 324408 208550 324420
rect 208762 324408 208768 324420
rect 208544 324380 208768 324408
rect 208544 324368 208550 324380
rect 208762 324368 208768 324380
rect 208820 324368 208826 324420
rect 222194 324232 222200 324284
rect 222252 324272 222258 324284
rect 222654 324272 222660 324284
rect 222252 324244 222660 324272
rect 222252 324232 222258 324244
rect 222654 324232 222660 324244
rect 222712 324232 222718 324284
rect 236086 323688 236092 323740
rect 236144 323728 236150 323740
rect 236362 323728 236368 323740
rect 236144 323700 236368 323728
rect 236144 323688 236150 323700
rect 236362 323688 236368 323700
rect 236420 323688 236426 323740
rect 147582 323620 147588 323672
rect 147640 323660 147646 323672
rect 222746 323660 222752 323672
rect 147640 323632 222752 323660
rect 147640 323620 147646 323632
rect 222746 323620 222752 323632
rect 222804 323620 222810 323672
rect 324130 323620 324136 323672
rect 324188 323660 324194 323672
rect 412634 323660 412640 323672
rect 324188 323632 412640 323660
rect 324188 323620 324194 323632
rect 412634 323620 412640 323632
rect 412692 323620 412698 323672
rect 28902 323552 28908 323604
rect 28960 323592 28966 323604
rect 178218 323592 178224 323604
rect 28960 323564 178224 323592
rect 28960 323552 28966 323564
rect 178218 323552 178224 323564
rect 178276 323552 178282 323604
rect 212718 323592 212724 323604
rect 212679 323564 212724 323592
rect 212718 323552 212724 323564
rect 212776 323552 212782 323604
rect 229186 323552 229192 323604
rect 229244 323592 229250 323604
rect 229370 323592 229376 323604
rect 229244 323564 229376 323592
rect 229244 323552 229250 323564
rect 229370 323552 229376 323564
rect 229428 323552 229434 323604
rect 234706 323552 234712 323604
rect 234764 323592 234770 323604
rect 234890 323592 234896 323604
rect 234764 323564 234896 323592
rect 234764 323552 234770 323564
rect 234890 323552 234896 323564
rect 234948 323552 234954 323604
rect 365438 323552 365444 323604
rect 365496 323592 365502 323604
rect 521654 323592 521660 323604
rect 365496 323564 521660 323592
rect 365496 323552 365502 323564
rect 521654 323552 521660 323564
rect 521712 323552 521718 323604
rect 131022 322260 131028 322312
rect 131080 322300 131086 322312
rect 216766 322300 216772 322312
rect 131080 322272 216772 322300
rect 131080 322260 131086 322272
rect 216766 322260 216772 322272
rect 216824 322260 216830 322312
rect 319898 322260 319904 322312
rect 319956 322300 319962 322312
rect 401594 322300 401600 322312
rect 319956 322272 401600 322300
rect 319956 322260 319962 322272
rect 401594 322260 401600 322272
rect 401652 322260 401658 322312
rect 51718 322192 51724 322244
rect 51776 322232 51782 322244
rect 186498 322232 186504 322244
rect 51776 322204 186504 322232
rect 51776 322192 51782 322204
rect 186498 322192 186504 322204
rect 186556 322192 186562 322244
rect 362678 322192 362684 322244
rect 362736 322232 362742 322244
rect 514754 322232 514760 322244
rect 362736 322204 514760 322232
rect 362736 322192 362742 322204
rect 514754 322192 514760 322204
rect 514812 322192 514818 322244
rect 223758 321960 223764 321972
rect 223719 321932 223764 321960
rect 223758 321920 223764 321932
rect 223816 321920 223822 321972
rect 321278 320900 321284 320952
rect 321336 320940 321342 320952
rect 405734 320940 405740 320952
rect 321336 320912 405740 320940
rect 321336 320900 321342 320912
rect 405734 320900 405740 320912
rect 405792 320900 405798 320952
rect 14458 320832 14464 320884
rect 14516 320872 14522 320884
rect 172606 320872 172612 320884
rect 14516 320844 172612 320872
rect 14516 320832 14522 320844
rect 172606 320832 172612 320844
rect 172664 320832 172670 320884
rect 177942 320832 177948 320884
rect 178000 320872 178006 320884
rect 233418 320872 233424 320884
rect 178000 320844 233424 320872
rect 178000 320832 178006 320844
rect 233418 320832 233424 320844
rect 233476 320832 233482 320884
rect 364058 320832 364064 320884
rect 364116 320872 364122 320884
rect 517514 320872 517520 320884
rect 364116 320844 517520 320872
rect 364116 320832 364122 320844
rect 517514 320832 517520 320844
rect 517572 320832 517578 320884
rect 3050 320084 3056 320136
rect 3108 320124 3114 320136
rect 166810 320124 166816 320136
rect 3108 320096 166816 320124
rect 3108 320084 3114 320096
rect 166810 320084 166816 320096
rect 166868 320084 166874 320136
rect 326890 319472 326896 319524
rect 326948 319512 326954 319524
rect 419534 319512 419540 319524
rect 326948 319484 419540 319512
rect 326948 319472 326954 319484
rect 419534 319472 419540 319484
rect 419592 319472 419598 319524
rect 153102 319404 153108 319456
rect 153160 319444 153166 319456
rect 225138 319444 225144 319456
rect 153160 319416 225144 319444
rect 153160 319404 153166 319416
rect 225138 319404 225144 319416
rect 225196 319404 225202 319456
rect 370958 319404 370964 319456
rect 371016 319444 371022 319456
rect 535454 319444 535460 319456
rect 371016 319416 535460 319444
rect 371016 319404 371022 319416
rect 535454 319404 535460 319416
rect 535512 319404 535518 319456
rect 262306 319336 262312 319388
rect 262364 319376 262370 319388
rect 262490 319376 262496 319388
rect 262364 319348 262496 319376
rect 262364 319336 262370 319348
rect 262490 319336 262496 319348
rect 262548 319336 262554 319388
rect 269114 319336 269120 319388
rect 269172 319376 269178 319388
rect 269298 319376 269304 319388
rect 269172 319348 269304 319376
rect 269172 319336 269178 319348
rect 269298 319336 269304 319348
rect 269356 319336 269362 319388
rect 142062 318044 142068 318096
rect 142120 318084 142126 318096
rect 220906 318084 220912 318096
rect 142120 318056 220912 318084
rect 142120 318044 142126 318056
rect 220906 318044 220912 318056
rect 220964 318044 220970 318096
rect 353110 318044 353116 318096
rect 353168 318084 353174 318096
rect 488534 318084 488540 318096
rect 353168 318056 488540 318084
rect 353168 318044 353174 318056
rect 488534 318044 488540 318056
rect 488592 318044 488598 318096
rect 137922 316684 137928 316736
rect 137980 316724 137986 316736
rect 219526 316724 219532 316736
rect 137980 316696 219532 316724
rect 137980 316684 137986 316696
rect 219526 316684 219532 316696
rect 219584 316684 219590 316736
rect 355778 316684 355784 316736
rect 355836 316724 355842 316736
rect 495434 316724 495440 316736
rect 355836 316696 495440 316724
rect 355836 316684 355842 316696
rect 495434 316684 495440 316696
rect 495492 316684 495498 316736
rect 144730 315256 144736 315308
rect 144788 315296 144794 315308
rect 222286 315296 222292 315308
rect 144788 315268 222292 315296
rect 144788 315256 144794 315268
rect 222286 315256 222292 315268
rect 222344 315256 222350 315308
rect 358538 315256 358544 315308
rect 358596 315296 358602 315308
rect 506474 315296 506480 315308
rect 358596 315268 506480 315296
rect 358596 315256 358602 315268
rect 506474 315256 506480 315268
rect 506532 315256 506538 315308
rect 198826 313964 198832 314016
rect 198884 314004 198890 314016
rect 199010 314004 199016 314016
rect 198884 313976 199016 314004
rect 198884 313964 198890 313976
rect 199010 313964 199016 313976
rect 199068 313964 199074 314016
rect 148962 313896 148968 313948
rect 149020 313936 149026 313948
rect 223758 313936 223764 313948
rect 149020 313908 223764 313936
rect 149020 313896 149026 313908
rect 223758 313896 223764 313908
rect 223816 313896 223822 313948
rect 361298 313896 361304 313948
rect 361356 313936 361362 313948
rect 513374 313936 513380 313948
rect 361356 313908 513380 313936
rect 361356 313896 361362 313908
rect 513374 313896 513380 313908
rect 513432 313896 513438 313948
rect 201586 313828 201592 313880
rect 201644 313868 201650 313880
rect 201770 313868 201776 313880
rect 201644 313840 201776 313868
rect 201644 313828 201650 313840
rect 201770 313828 201776 313840
rect 201828 313828 201834 313880
rect 389266 313216 389272 313268
rect 389324 313256 389330 313268
rect 580166 313256 580172 313268
rect 389324 313228 580172 313256
rect 389324 313216 389330 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 88242 312536 88248 312588
rect 88300 312576 88306 312588
rect 200298 312576 200304 312588
rect 88300 312548 200304 312576
rect 88300 312536 88306 312548
rect 200298 312536 200304 312548
rect 200356 312536 200362 312588
rect 95142 311108 95148 311160
rect 95200 311148 95206 311160
rect 203058 311148 203064 311160
rect 95200 311120 203064 311148
rect 95200 311108 95206 311120
rect 203058 311108 203064 311120
rect 203116 311108 203122 311160
rect 348878 311108 348884 311160
rect 348936 311148 348942 311160
rect 477494 311148 477500 311160
rect 348936 311120 477500 311148
rect 348936 311108 348942 311120
rect 477494 311108 477500 311120
rect 477552 311108 477558 311160
rect 106182 309748 106188 309800
rect 106240 309788 106246 309800
rect 207198 309788 207204 309800
rect 106240 309760 207204 309788
rect 106240 309748 106246 309760
rect 207198 309748 207204 309760
rect 207256 309748 207262 309800
rect 355870 309748 355876 309800
rect 355928 309788 355934 309800
rect 496814 309788 496820 309800
rect 355928 309760 496820 309788
rect 355928 309748 355934 309760
rect 496814 309748 496820 309760
rect 496872 309748 496878 309800
rect 117222 308388 117228 308440
rect 117280 308428 117286 308440
rect 211246 308428 211252 308440
rect 117280 308400 211252 308428
rect 117280 308388 117286 308400
rect 211246 308388 211252 308400
rect 211304 308388 211310 308440
rect 350350 308388 350356 308440
rect 350408 308428 350414 308440
rect 481634 308428 481640 308440
rect 350408 308400 481640 308428
rect 350408 308388 350414 308400
rect 481634 308388 481640 308400
rect 481692 308388 481698 308440
rect 99282 307028 99288 307080
rect 99340 307068 99346 307080
rect 202138 307068 202144 307080
rect 99340 307040 202144 307068
rect 99340 307028 99346 307040
rect 202138 307028 202144 307040
rect 202196 307028 202202 307080
rect 357250 307028 357256 307080
rect 357308 307068 357314 307080
rect 499574 307068 499580 307080
rect 357308 307040 499580 307068
rect 357308 307028 357314 307040
rect 499574 307028 499580 307040
rect 499632 307028 499638 307080
rect 119982 305600 119988 305652
rect 120040 305640 120046 305652
rect 212626 305640 212632 305652
rect 120040 305612 212632 305640
rect 120040 305600 120046 305612
rect 212626 305600 212632 305612
rect 212684 305600 212690 305652
rect 303338 305600 303344 305652
rect 303396 305640 303402 305652
rect 357434 305640 357440 305652
rect 303396 305612 357440 305640
rect 303396 305600 303402 305612
rect 357434 305600 357440 305612
rect 357492 305600 357498 305652
rect 358630 305600 358636 305652
rect 358688 305640 358694 305652
rect 503714 305640 503720 305652
rect 358688 305612 503720 305640
rect 358688 305600 358694 305612
rect 503714 305600 503720 305612
rect 503772 305600 503778 305652
rect 124122 304240 124128 304292
rect 124180 304280 124186 304292
rect 214098 304280 214104 304292
rect 124180 304252 214104 304280
rect 124180 304240 124186 304252
rect 214098 304240 214104 304252
rect 214156 304240 214162 304292
rect 366818 304240 366824 304292
rect 366876 304280 366882 304292
rect 524414 304280 524420 304292
rect 366876 304252 524420 304280
rect 366876 304240 366882 304252
rect 524414 304240 524420 304252
rect 524472 304240 524478 304292
rect 47578 302880 47584 302932
rect 47636 302920 47642 302932
rect 185026 302920 185032 302932
rect 47636 302892 185032 302920
rect 47636 302880 47642 302892
rect 185026 302880 185032 302892
rect 185084 302880 185090 302932
rect 361390 302880 361396 302932
rect 361448 302920 361454 302932
rect 510614 302920 510620 302932
rect 361448 302892 510620 302920
rect 361448 302880 361454 302892
rect 510614 302880 510620 302892
rect 510672 302880 510678 302932
rect 40678 301452 40684 301504
rect 40736 301492 40742 301504
rect 182266 301492 182272 301504
rect 40736 301464 182272 301492
rect 40736 301452 40742 301464
rect 182266 301452 182272 301464
rect 182324 301452 182330 301504
rect 368198 301452 368204 301504
rect 368256 301492 368262 301504
rect 528554 301492 528560 301504
rect 368256 301464 528560 301492
rect 368256 301452 368262 301464
rect 528554 301452 528560 301464
rect 528612 301452 528618 301504
rect 372338 300092 372344 300144
rect 372396 300132 372402 300144
rect 542354 300132 542360 300144
rect 372396 300104 542360 300132
rect 372396 300092 372402 300104
rect 542354 300092 542360 300104
rect 542412 300092 542418 300144
rect 389358 299412 389364 299464
rect 389416 299452 389422 299464
rect 579614 299452 579620 299464
rect 389416 299424 579620 299452
rect 389416 299412 389422 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 369578 297372 369584 297424
rect 369636 297412 369642 297424
rect 531314 297412 531320 297424
rect 369636 297384 531320 297412
rect 369636 297372 369642 297384
rect 531314 297372 531320 297384
rect 531372 297372 531378 297424
rect 373718 295944 373724 295996
rect 373776 295984 373782 295996
rect 546494 295984 546500 295996
rect 373776 295956 546500 295984
rect 373776 295944 373782 295956
rect 546494 295944 546500 295956
rect 546552 295944 546558 295996
rect 376478 294584 376484 294636
rect 376536 294624 376542 294636
rect 553394 294624 553400 294636
rect 376536 294596 553400 294624
rect 376536 294584 376542 294596
rect 553394 294584 553400 294596
rect 553452 294584 553458 294636
rect 2774 293564 2780 293616
rect 2832 293604 2838 293616
rect 4798 293604 4804 293616
rect 2832 293576 4804 293604
rect 2832 293564 2838 293576
rect 4798 293564 4804 293576
rect 4856 293564 4862 293616
rect 375098 293224 375104 293276
rect 375156 293264 375162 293276
rect 549254 293264 549260 293276
rect 375156 293236 549260 293264
rect 375156 293224 375162 293236
rect 549254 293224 549260 293236
rect 549312 293224 549318 293276
rect 379238 291796 379244 291848
rect 379296 291836 379302 291848
rect 560294 291836 560300 291848
rect 379296 291808 560300 291836
rect 379296 291796 379302 291808
rect 560294 291796 560300 291808
rect 560352 291796 560358 291848
rect 380618 290436 380624 290488
rect 380676 290476 380682 290488
rect 564434 290476 564440 290488
rect 380676 290448 564440 290476
rect 380676 290436 380682 290448
rect 564434 290436 564440 290448
rect 564492 290436 564498 290488
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 166718 280140 166724 280152
rect 3200 280112 166724 280140
rect 3200 280100 3206 280112
rect 166718 280100 166724 280112
rect 166776 280100 166782 280152
rect 393958 273164 393964 273216
rect 394016 273204 394022 273216
rect 580166 273204 580172 273216
rect 394016 273176 580172 273204
rect 394016 273164 394022 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 166626 267696 166632 267708
rect 3016 267668 166632 267696
rect 3016 267656 3022 267668
rect 166626 267656 166632 267668
rect 166684 267656 166690 267708
rect 406378 259360 406384 259412
rect 406436 259400 406442 259412
rect 580166 259400 580172 259412
rect 406436 259372 580172 259400
rect 406436 259360 406442 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 21450 255252 21456 255264
rect 3200 255224 21456 255252
rect 3200 255212 3206 255224
rect 21450 255212 21456 255224
rect 21508 255212 21514 255264
rect 21358 254532 21364 254584
rect 21416 254572 21422 254584
rect 173986 254572 173992 254584
rect 21416 254544 173992 254572
rect 21416 254532 21422 254544
rect 173986 254532 173992 254544
rect 174044 254532 174050 254584
rect 389450 245556 389456 245608
rect 389508 245596 389514 245608
rect 580166 245596 580172 245608
rect 389508 245568 580172 245596
rect 389508 245556 389514 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 389542 233180 389548 233232
rect 389600 233220 389606 233232
rect 579982 233220 579988 233232
rect 389600 233192 579988 233220
rect 389600 233180 389606 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3234 229032 3240 229084
rect 3292 229072 3298 229084
rect 166534 229072 166540 229084
rect 3292 229044 166540 229072
rect 3292 229032 3298 229044
rect 166534 229032 166540 229044
rect 166592 229032 166598 229084
rect 290458 224204 290464 224256
rect 290516 224244 290522 224256
rect 322934 224244 322940 224256
rect 290516 224216 322940 224244
rect 290516 224204 290522 224216
rect 322934 224204 322940 224216
rect 322992 224204 322998 224256
rect 319990 222844 319996 222896
rect 320048 222884 320054 222896
rect 402974 222884 402980 222896
rect 320048 222856 402980 222884
rect 320048 222844 320054 222856
rect 402974 222844 402980 222856
rect 403032 222844 403038 222896
rect 153010 221416 153016 221468
rect 153068 221456 153074 221468
rect 225046 221456 225052 221468
rect 153068 221428 225052 221456
rect 153068 221416 153074 221428
rect 225046 221416 225052 221428
rect 225104 221416 225110 221468
rect 297910 221416 297916 221468
rect 297968 221456 297974 221468
rect 340874 221456 340880 221468
rect 297968 221428 340880 221456
rect 297968 221416 297974 221428
rect 340874 221416 340880 221428
rect 340932 221416 340938 221468
rect 143442 220056 143448 220108
rect 143500 220096 143506 220108
rect 220814 220096 220820 220108
rect 143500 220068 220820 220096
rect 143500 220056 143506 220068
rect 220814 220056 220820 220068
rect 220872 220056 220878 220108
rect 296438 220056 296444 220108
rect 296496 220096 296502 220108
rect 338114 220096 338120 220108
rect 296496 220068 338120 220096
rect 296496 220056 296502 220068
rect 338114 220056 338120 220068
rect 338172 220056 338178 220108
rect 362770 220056 362776 220108
rect 362828 220096 362834 220108
rect 516134 220096 516140 220108
rect 362828 220068 516140 220096
rect 362828 220056 362834 220068
rect 516134 220056 516140 220068
rect 516192 220056 516198 220108
rect 389634 219376 389640 219428
rect 389692 219416 389698 219428
rect 580166 219416 580172 219428
rect 389692 219388 580172 219416
rect 389692 219376 389698 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 202782 218696 202788 218748
rect 202840 218736 202846 218748
rect 242986 218736 242992 218748
rect 202840 218708 242992 218736
rect 202840 218696 202846 218708
rect 242986 218696 242992 218708
rect 243044 218696 243050 218748
rect 284018 218696 284024 218748
rect 284076 218736 284082 218748
rect 306374 218736 306380 218748
rect 284076 218708 306380 218736
rect 284076 218696 284082 218708
rect 306374 218696 306380 218708
rect 306432 218696 306438 218748
rect 279878 217336 279884 217388
rect 279936 217376 279942 217388
rect 295334 217376 295340 217388
rect 279936 217348 295340 217376
rect 279936 217336 279942 217348
rect 295334 217336 295340 217348
rect 295392 217336 295398 217388
rect 183462 217268 183468 217320
rect 183520 217308 183526 217320
rect 236086 217308 236092 217320
rect 183520 217280 236092 217308
rect 183520 217268 183526 217280
rect 236086 217268 236092 217280
rect 236144 217268 236150 217320
rect 293770 217268 293776 217320
rect 293828 217308 293834 217320
rect 331214 217308 331220 217320
rect 293828 217280 331220 217308
rect 293828 217268 293834 217280
rect 331214 217268 331220 217280
rect 331272 217268 331278 217320
rect 351730 217268 351736 217320
rect 351788 217308 351794 217320
rect 487154 217308 487160 217320
rect 351788 217280 487160 217308
rect 351788 217268 351794 217280
rect 487154 217268 487160 217280
rect 487212 217268 487218 217320
rect 195882 215908 195888 215960
rect 195940 215948 195946 215960
rect 239398 215948 239404 215960
rect 195940 215920 239404 215948
rect 195940 215908 195946 215920
rect 239398 215908 239404 215920
rect 239456 215908 239462 215960
rect 282638 215908 282644 215960
rect 282696 215948 282702 215960
rect 302234 215948 302240 215960
rect 282696 215920 302240 215948
rect 282696 215908 282702 215920
rect 302234 215908 302240 215920
rect 302292 215908 302298 215960
rect 355962 215908 355968 215960
rect 356020 215948 356026 215960
rect 498194 215948 498200 215960
rect 356020 215920 498200 215948
rect 356020 215908 356026 215920
rect 498194 215908 498200 215920
rect 498252 215908 498258 215960
rect 3234 215228 3240 215280
rect 3292 215268 3298 215280
rect 166442 215268 166448 215280
rect 3292 215240 166448 215268
rect 3292 215228 3298 215240
rect 166442 215228 166448 215240
rect 166500 215228 166506 215280
rect 389726 206932 389732 206984
rect 389784 206972 389790 206984
rect 579798 206972 579804 206984
rect 389784 206944 579804 206972
rect 389784 206932 389790 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 390462 193128 390468 193180
rect 390520 193168 390526 193180
rect 580166 193168 580172 193180
rect 390520 193140 580172 193168
rect 390520 193128 390526 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 10318 189020 10324 189032
rect 3384 188992 10324 189020
rect 3384 188980 3390 188992
rect 10318 188980 10324 188992
rect 10376 188980 10382 189032
rect 403618 179324 403624 179376
rect 403676 179364 403682 179376
rect 580166 179364 580172 179376
rect 403676 179336 580172 179364
rect 403676 179324 403682 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 3326 176604 3332 176656
rect 3384 176644 3390 176656
rect 166350 176644 166356 176656
rect 3384 176616 166356 176644
rect 3384 176604 3390 176616
rect 166350 176604 166356 176616
rect 166408 176604 166414 176656
rect 390370 166948 390376 167000
rect 390428 166988 390434 167000
rect 580166 166988 580172 167000
rect 390428 166960 580172 166988
rect 390428 166948 390434 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 390278 153144 390284 153196
rect 390336 153184 390342 153196
rect 580166 153184 580172 153196
rect 390336 153156 580172 153184
rect 390336 153144 390342 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 28258 150396 28264 150408
rect 3384 150368 28264 150396
rect 3384 150356 3390 150368
rect 28258 150356 28264 150368
rect 28316 150356 28322 150408
rect 390186 139340 390192 139392
rect 390244 139380 390250 139392
rect 580166 139380 580172 139392
rect 390244 139352 580172 139380
rect 390244 139340 390250 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 390094 126896 390100 126948
rect 390152 126936 390158 126948
rect 580166 126936 580172 126948
rect 390152 126908 580172 126936
rect 390152 126896 390158 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 3142 124108 3148 124160
rect 3200 124148 3206 124160
rect 166258 124148 166264 124160
rect 3200 124120 166264 124148
rect 3200 124108 3206 124120
rect 166258 124108 166264 124120
rect 166316 124108 166322 124160
rect 390002 113092 390008 113144
rect 390060 113132 390066 113144
rect 579798 113132 579804 113144
rect 390060 113104 579804 113132
rect 390060 113092 390066 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 400858 100648 400864 100700
rect 400916 100688 400922 100700
rect 580166 100688 580172 100700
rect 400916 100660 580172 100688
rect 400916 100648 400922 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 547138 86912 547144 86964
rect 547196 86952 547202 86964
rect 580166 86952 580172 86964
rect 547196 86924 580172 86952
rect 547196 86912 547202 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 11698 85524 11704 85536
rect 3200 85496 11704 85524
rect 3200 85484 3206 85496
rect 11698 85484 11704 85496
rect 11756 85484 11762 85536
rect 389910 73108 389916 73160
rect 389968 73148 389974 73160
rect 580166 73148 580172 73160
rect 389968 73120 580172 73148
rect 389968 73108 389974 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 389818 60664 389824 60716
rect 389876 60704 389882 60716
rect 580166 60704 580172 60716
rect 389876 60676 580172 60704
rect 389876 60664 389882 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 2866 59304 2872 59356
rect 2924 59344 2930 59356
rect 29638 59344 29644 59356
rect 2924 59316 29644 59344
rect 2924 59304 2930 59316
rect 29638 59304 29644 59316
rect 29696 59304 29702 59356
rect 542998 46860 543004 46912
rect 543056 46900 543062 46912
rect 580166 46900 580172 46912
rect 543056 46872 580172 46900
rect 543056 46860 543062 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 358722 42032 358728 42084
rect 358780 42072 358786 42084
rect 505094 42072 505100 42084
rect 358780 42044 505100 42072
rect 358780 42032 358786 42044
rect 505094 42032 505100 42044
rect 505152 42032 505158 42084
rect 81342 28228 81348 28280
rect 81400 28268 81406 28280
rect 197538 28268 197544 28280
rect 81400 28240 197544 28268
rect 81400 28228 81406 28240
rect 197538 28228 197544 28240
rect 197596 28228 197602 28280
rect 157242 26868 157248 26920
rect 157300 26908 157306 26920
rect 226426 26908 226432 26920
rect 157300 26880 226432 26908
rect 157300 26868 157306 26880
rect 226426 26868 226432 26880
rect 226484 26868 226490 26920
rect 150342 25508 150348 25560
rect 150400 25548 150406 25560
rect 223666 25548 223672 25560
rect 150400 25520 223672 25548
rect 150400 25508 150406 25520
rect 223666 25508 223672 25520
rect 223724 25508 223730 25560
rect 146202 24080 146208 24132
rect 146260 24120 146266 24132
rect 222194 24120 222200 24132
rect 146260 24092 222200 24120
rect 146260 24080 146266 24092
rect 222194 24080 222200 24092
rect 222252 24080 222258 24132
rect 360010 24080 360016 24132
rect 360068 24120 360074 24132
rect 506566 24120 506572 24132
rect 360068 24092 506572 24120
rect 360068 24080 360074 24092
rect 506566 24080 506572 24092
rect 506624 24080 506630 24132
rect 136450 22720 136456 22772
rect 136508 22760 136514 22772
rect 218330 22760 218336 22772
rect 136508 22732 218336 22760
rect 136508 22720 136514 22732
rect 218330 22720 218336 22732
rect 218388 22720 218394 22772
rect 299198 22720 299204 22772
rect 299256 22760 299262 22772
rect 347774 22760 347780 22772
rect 299256 22732 347780 22760
rect 299256 22720 299262 22732
rect 347774 22720 347780 22732
rect 347832 22720 347838 22772
rect 353018 22720 353024 22772
rect 353076 22760 353082 22772
rect 490006 22760 490012 22772
rect 353076 22732 490012 22760
rect 353076 22720 353082 22732
rect 490006 22720 490012 22732
rect 490064 22720 490070 22772
rect 194410 21428 194416 21480
rect 194468 21468 194474 21480
rect 240318 21468 240324 21480
rect 194468 21440 240324 21468
rect 194468 21428 194474 21440
rect 240318 21428 240324 21440
rect 240376 21428 240382 21480
rect 110322 21360 110328 21412
rect 110380 21400 110386 21412
rect 208486 21400 208492 21412
rect 110380 21372 208492 21400
rect 110380 21360 110386 21372
rect 208486 21360 208492 21372
rect 208544 21360 208550 21412
rect 296530 21360 296536 21412
rect 296588 21400 296594 21412
rect 340966 21400 340972 21412
rect 296588 21372 340972 21400
rect 296588 21360 296594 21372
rect 340966 21360 340972 21372
rect 341024 21360 341030 21412
rect 347590 21360 347596 21412
rect 347648 21400 347654 21412
rect 473354 21400 473360 21412
rect 347648 21372 473360 21400
rect 347648 21360 347654 21372
rect 473354 21360 473360 21372
rect 473412 21360 473418 21412
rect 396718 20612 396724 20664
rect 396776 20652 396782 20664
rect 579982 20652 579988 20664
rect 396776 20624 579988 20652
rect 396776 20612 396782 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 187602 19932 187608 19984
rect 187660 19972 187666 19984
rect 237558 19972 237564 19984
rect 187660 19944 237564 19972
rect 187660 19932 187666 19944
rect 237558 19932 237564 19944
rect 237616 19932 237622 19984
rect 292390 19932 292396 19984
rect 292448 19972 292454 19984
rect 329834 19972 329840 19984
rect 292448 19944 329840 19972
rect 292448 19932 292454 19944
rect 329834 19932 329840 19944
rect 329892 19932 329898 19984
rect 286870 18640 286876 18692
rect 286928 18680 286934 18692
rect 313274 18680 313280 18692
rect 286928 18652 313280 18680
rect 286928 18640 286934 18652
rect 313274 18640 313280 18652
rect 313332 18640 313338 18692
rect 184842 18572 184848 18624
rect 184900 18612 184906 18624
rect 233878 18612 233884 18624
rect 184900 18584 233884 18612
rect 184900 18572 184906 18584
rect 233878 18572 233884 18584
rect 233936 18572 233942 18624
rect 300578 18572 300584 18624
rect 300636 18612 300642 18624
rect 350534 18612 350540 18624
rect 300636 18584 350540 18612
rect 300636 18572 300642 18584
rect 350534 18572 350540 18584
rect 350592 18572 350598 18624
rect 360102 18572 360108 18624
rect 360160 18612 360166 18624
rect 509234 18612 509240 18624
rect 360160 18584 509240 18612
rect 360160 18572 360166 18584
rect 509234 18572 509240 18584
rect 509292 18572 509298 18624
rect 316678 17892 316684 17944
rect 316736 17932 316742 17944
rect 324314 17932 324320 17944
rect 316736 17904 324320 17932
rect 316736 17892 316742 17904
rect 324314 17892 324320 17904
rect 324372 17892 324378 17944
rect 173802 17212 173808 17264
rect 173860 17252 173866 17264
rect 232038 17252 232044 17264
rect 173860 17224 232044 17252
rect 173860 17212 173866 17224
rect 232038 17212 232044 17224
rect 232096 17212 232102 17264
rect 325418 17212 325424 17264
rect 325476 17252 325482 17264
rect 415486 17252 415492 17264
rect 325476 17224 415492 17252
rect 325476 17212 325482 17224
rect 415486 17212 415492 17224
rect 415544 17212 415550 17264
rect 169570 15852 169576 15904
rect 169628 15892 169634 15904
rect 222838 15892 222844 15904
rect 169628 15864 222844 15892
rect 169628 15852 169634 15864
rect 222838 15852 222844 15864
rect 222896 15852 222902 15904
rect 289630 15852 289636 15904
rect 289688 15892 289694 15904
rect 322106 15892 322112 15904
rect 289688 15864 322112 15892
rect 289688 15852 289694 15864
rect 322106 15852 322112 15864
rect 322164 15852 322170 15904
rect 322658 15852 322664 15904
rect 322716 15892 322722 15904
rect 409598 15892 409604 15904
rect 322716 15864 409604 15892
rect 322716 15852 322722 15864
rect 409598 15852 409604 15864
rect 409656 15852 409662 15904
rect 215202 14560 215208 14612
rect 215260 14600 215266 14612
rect 246298 14600 246304 14612
rect 215260 14572 246304 14600
rect 215260 14560 215266 14572
rect 246298 14560 246304 14572
rect 246356 14560 246362 14612
rect 191742 14492 191748 14544
rect 191800 14532 191806 14544
rect 236638 14532 236644 14544
rect 191800 14504 236644 14532
rect 191800 14492 191806 14504
rect 236638 14492 236644 14504
rect 236696 14492 236702 14544
rect 132218 14424 132224 14476
rect 132276 14464 132282 14476
rect 216674 14464 216680 14476
rect 132276 14436 216680 14464
rect 132276 14424 132282 14436
rect 216674 14424 216680 14436
rect 216732 14424 216738 14476
rect 299290 14424 299296 14476
rect 299348 14464 299354 14476
rect 345750 14464 345756 14476
rect 299348 14436 345756 14464
rect 299348 14424 299354 14436
rect 345750 14424 345756 14436
rect 345808 14424 345814 14476
rect 354490 14424 354496 14476
rect 354548 14464 354554 14476
rect 492306 14464 492312 14476
rect 354548 14436 492312 14464
rect 354548 14424 354554 14436
rect 492306 14424 492312 14436
rect 492364 14424 492370 14476
rect 179046 13132 179052 13184
rect 179104 13172 179110 13184
rect 234706 13172 234712 13184
rect 179104 13144 234712 13172
rect 179104 13132 179110 13144
rect 234706 13132 234712 13144
rect 234764 13132 234770 13184
rect 335998 13132 336004 13184
rect 336056 13172 336062 13184
rect 390646 13172 390652 13184
rect 336056 13144 390652 13172
rect 336056 13132 336062 13144
rect 390646 13132 390652 13144
rect 390704 13132 390710 13184
rect 138842 13064 138848 13116
rect 138900 13104 138906 13116
rect 219434 13104 219440 13116
rect 138900 13076 219440 13104
rect 138900 13064 138906 13076
rect 219434 13064 219440 13076
rect 219492 13064 219498 13116
rect 295058 13064 295064 13116
rect 295116 13104 295122 13116
rect 334986 13104 334992 13116
rect 295116 13076 334992 13104
rect 295116 13064 295122 13076
rect 334986 13064 334992 13076
rect 335044 13064 335050 13116
rect 357342 13064 357348 13116
rect 357400 13104 357406 13116
rect 499390 13104 499396 13116
rect 357400 13076 499396 13104
rect 357400 13064 357406 13076
rect 499390 13064 499396 13076
rect 499448 13064 499454 13116
rect 200022 11840 200028 11892
rect 200080 11880 200086 11892
rect 242250 11880 242256 11892
rect 200080 11852 242256 11880
rect 200080 11840 200086 11852
rect 242250 11840 242256 11852
rect 242308 11840 242314 11892
rect 176562 11772 176568 11824
rect 176620 11812 176626 11824
rect 233326 11812 233332 11824
rect 176620 11784 233332 11812
rect 176620 11772 176626 11784
rect 233326 11772 233332 11784
rect 233384 11772 233390 11824
rect 292482 11772 292488 11824
rect 292540 11812 292546 11824
rect 327994 11812 328000 11824
rect 292540 11784 328000 11812
rect 292540 11772 292546 11784
rect 327994 11772 328000 11784
rect 328052 11772 328058 11824
rect 103238 11704 103244 11756
rect 103296 11744 103302 11756
rect 205726 11744 205732 11756
rect 103296 11716 205732 11744
rect 103296 11704 103302 11716
rect 205726 11704 205732 11716
rect 205784 11704 205790 11756
rect 293862 11704 293868 11756
rect 293920 11744 293926 11756
rect 332594 11744 332600 11756
rect 293920 11716 332600 11744
rect 293920 11704 293926 11716
rect 332594 11704 332600 11716
rect 332652 11704 332658 11756
rect 348970 11704 348976 11756
rect 349028 11744 349034 11756
rect 480530 11744 480536 11756
rect 349028 11716 480536 11744
rect 349028 11704 349034 11716
rect 480530 11704 480536 11716
rect 480588 11704 480594 11756
rect 318058 10480 318064 10532
rect 318116 10520 318122 10532
rect 344554 10520 344560 10532
rect 318116 10492 344560 10520
rect 318116 10480 318122 10492
rect 344554 10480 344560 10492
rect 344612 10480 344618 10532
rect 289722 10412 289728 10464
rect 289780 10452 289786 10464
rect 320726 10452 320732 10464
rect 289780 10424 320732 10452
rect 289780 10412 289786 10424
rect 320726 10412 320732 10424
rect 320784 10412 320790 10464
rect 172422 10344 172428 10396
rect 172480 10384 172486 10396
rect 231946 10384 231952 10396
rect 172480 10356 231952 10384
rect 172480 10344 172486 10356
rect 231946 10344 231952 10356
rect 232004 10344 232010 10396
rect 291102 10344 291108 10396
rect 291160 10384 291166 10396
rect 326798 10384 326804 10396
rect 291160 10356 326804 10384
rect 291160 10344 291166 10356
rect 326798 10344 326804 10356
rect 326856 10344 326862 10396
rect 92382 10276 92388 10328
rect 92440 10316 92446 10328
rect 177298 10316 177304 10328
rect 92440 10288 177304 10316
rect 92440 10276 92446 10288
rect 177298 10276 177304 10288
rect 177356 10276 177362 10328
rect 205542 10276 205548 10328
rect 205600 10316 205606 10328
rect 244458 10316 244464 10328
rect 205600 10288 244464 10316
rect 205600 10276 205606 10288
rect 244458 10276 244464 10288
rect 244516 10276 244522 10328
rect 295150 10276 295156 10328
rect 295208 10316 295214 10328
rect 337470 10316 337476 10328
rect 295208 10288 337476 10316
rect 295208 10276 295214 10288
rect 337470 10276 337476 10288
rect 337528 10276 337534 10328
rect 354582 10276 354588 10328
rect 354640 10316 354646 10328
rect 494698 10316 494704 10328
rect 354640 10288 494704 10316
rect 354640 10276 354646 10288
rect 494698 10276 494704 10288
rect 494756 10276 494762 10328
rect 332318 9596 332324 9648
rect 332376 9636 332382 9648
rect 435542 9636 435548 9648
rect 332376 9608 435548 9636
rect 332376 9596 332382 9608
rect 435542 9596 435548 9608
rect 435600 9596 435606 9648
rect 333790 9528 333796 9580
rect 333848 9568 333854 9580
rect 439130 9568 439136 9580
rect 333848 9540 439136 9568
rect 333848 9528 333854 9540
rect 439130 9528 439136 9540
rect 439188 9528 439194 9580
rect 335078 9460 335084 9512
rect 335136 9500 335142 9512
rect 442626 9500 442632 9512
rect 335136 9472 442632 9500
rect 335136 9460 335142 9472
rect 442626 9460 442632 9472
rect 442684 9460 442690 9512
rect 336550 9392 336556 9444
rect 336608 9432 336614 9444
rect 446214 9432 446220 9444
rect 336608 9404 446220 9432
rect 336608 9392 336614 9404
rect 446214 9392 446220 9404
rect 446272 9392 446278 9444
rect 337838 9324 337844 9376
rect 337896 9364 337902 9376
rect 449802 9364 449808 9376
rect 337896 9336 449808 9364
rect 337896 9324 337902 9336
rect 449802 9324 449808 9336
rect 449860 9324 449866 9376
rect 339310 9256 339316 9308
rect 339368 9296 339374 9308
rect 453298 9296 453304 9308
rect 339368 9268 453304 9296
rect 339368 9256 339374 9268
rect 453298 9256 453304 9268
rect 453356 9256 453362 9308
rect 340598 9188 340604 9240
rect 340656 9228 340662 9240
rect 456886 9228 456892 9240
rect 340656 9200 456892 9228
rect 340656 9188 340662 9200
rect 456886 9188 456892 9200
rect 456944 9188 456950 9240
rect 342070 9120 342076 9172
rect 342128 9160 342134 9172
rect 460382 9160 460388 9172
rect 342128 9132 460388 9160
rect 342128 9120 342134 9132
rect 460382 9120 460388 9132
rect 460440 9120 460446 9172
rect 343266 9052 343272 9104
rect 343324 9092 343330 9104
rect 463970 9092 463976 9104
rect 343324 9064 463976 9092
rect 343324 9052 343330 9064
rect 463970 9052 463976 9064
rect 464028 9052 464034 9104
rect 168650 8984 168656 9036
rect 168708 9024 168714 9036
rect 229738 9024 229744 9036
rect 168708 8996 229744 9024
rect 168708 8984 168714 8996
rect 229738 8984 229744 8996
rect 229796 8984 229802 9036
rect 344830 8984 344836 9036
rect 344888 9024 344894 9036
rect 467466 9024 467472 9036
rect 344888 8996 467472 9024
rect 344888 8984 344894 8996
rect 467466 8984 467472 8996
rect 467524 8984 467530 9036
rect 84470 8916 84476 8968
rect 84528 8956 84534 8968
rect 173158 8956 173164 8968
rect 84528 8928 173164 8956
rect 84528 8916 84534 8928
rect 173158 8916 173164 8928
rect 173216 8916 173222 8968
rect 186130 8916 186136 8968
rect 186188 8956 186194 8968
rect 237466 8956 237472 8968
rect 186188 8928 237472 8956
rect 186188 8916 186194 8928
rect 237466 8916 237472 8928
rect 237524 8916 237530 8968
rect 285398 8916 285404 8968
rect 285456 8956 285462 8968
rect 310238 8956 310244 8968
rect 285456 8928 310244 8956
rect 285456 8916 285462 8928
rect 310238 8916 310244 8928
rect 310296 8916 310302 8968
rect 346118 8916 346124 8968
rect 346176 8956 346182 8968
rect 471054 8956 471060 8968
rect 346176 8928 471060 8956
rect 346176 8916 346182 8928
rect 471054 8916 471060 8928
rect 471112 8916 471118 8968
rect 331030 8848 331036 8900
rect 331088 8888 331094 8900
rect 432046 8888 432052 8900
rect 331088 8860 432052 8888
rect 331088 8848 331094 8860
rect 432046 8848 432052 8860
rect 432104 8848 432110 8900
rect 329558 8780 329564 8832
rect 329616 8820 329622 8832
rect 428458 8820 428464 8832
rect 329616 8792 428464 8820
rect 329616 8780 329622 8792
rect 428458 8780 428464 8792
rect 428516 8780 428522 8832
rect 328178 8712 328184 8764
rect 328236 8752 328242 8764
rect 424962 8752 424968 8764
rect 328236 8724 424968 8752
rect 328236 8712 328242 8724
rect 424962 8712 424968 8724
rect 425020 8712 425026 8764
rect 326982 8644 326988 8696
rect 327040 8684 327046 8696
rect 421374 8684 421380 8696
rect 327040 8656 421380 8684
rect 327040 8644 327046 8656
rect 421374 8644 421380 8656
rect 421432 8644 421438 8696
rect 325510 8576 325516 8628
rect 325568 8616 325574 8628
rect 417878 8616 417884 8628
rect 325568 8588 417884 8616
rect 325568 8576 325574 8588
rect 417878 8576 417884 8588
rect 417936 8576 417942 8628
rect 324222 8508 324228 8560
rect 324280 8548 324286 8560
rect 414290 8548 414296 8560
rect 324280 8520 414296 8548
rect 324280 8508 324286 8520
rect 414290 8508 414296 8520
rect 414348 8508 414354 8560
rect 322750 8440 322756 8492
rect 322808 8480 322814 8492
rect 410794 8480 410800 8492
rect 322808 8452 410800 8480
rect 322808 8440 322814 8452
rect 410794 8440 410800 8452
rect 410852 8440 410858 8492
rect 321370 8372 321376 8424
rect 321428 8412 321434 8424
rect 407206 8412 407212 8424
rect 321428 8384 407212 8412
rect 321428 8372 321434 8384
rect 407206 8372 407212 8384
rect 407264 8372 407270 8424
rect 97442 8236 97448 8288
rect 97500 8276 97506 8288
rect 204438 8276 204444 8288
rect 97500 8248 204444 8276
rect 97500 8236 97506 8248
rect 204438 8236 204444 8248
rect 204496 8236 204502 8288
rect 372430 8236 372436 8288
rect 372488 8276 372494 8288
rect 541986 8276 541992 8288
rect 372488 8248 541992 8276
rect 372488 8236 372494 8248
rect 541986 8236 541992 8248
rect 542044 8236 542050 8288
rect 93946 8168 93952 8220
rect 94004 8208 94010 8220
rect 202966 8208 202972 8220
rect 94004 8180 202972 8208
rect 94004 8168 94010 8180
rect 202966 8168 202972 8180
rect 203024 8168 203030 8220
rect 373810 8168 373816 8220
rect 373868 8208 373874 8220
rect 545482 8208 545488 8220
rect 373868 8180 545488 8208
rect 373868 8168 373874 8180
rect 545482 8168 545488 8180
rect 545540 8168 545546 8220
rect 90358 8100 90364 8152
rect 90416 8140 90422 8152
rect 201586 8140 201592 8152
rect 90416 8112 201592 8140
rect 90416 8100 90422 8112
rect 201586 8100 201592 8112
rect 201644 8100 201650 8152
rect 375190 8100 375196 8152
rect 375248 8140 375254 8152
rect 549070 8140 549076 8152
rect 375248 8112 549076 8140
rect 375248 8100 375254 8112
rect 549070 8100 549076 8112
rect 549128 8100 549134 8152
rect 86862 8032 86868 8084
rect 86920 8072 86926 8084
rect 200206 8072 200212 8084
rect 86920 8044 200212 8072
rect 86920 8032 86926 8044
rect 200206 8032 200212 8044
rect 200264 8032 200270 8084
rect 376570 8032 376576 8084
rect 376628 8072 376634 8084
rect 552658 8072 552664 8084
rect 376628 8044 552664 8072
rect 376628 8032 376634 8044
rect 552658 8032 552664 8044
rect 552716 8032 552722 8084
rect 83274 7964 83280 8016
rect 83332 8004 83338 8016
rect 198826 8004 198832 8016
rect 83332 7976 198832 8004
rect 83332 7964 83338 7976
rect 198826 7964 198832 7976
rect 198884 7964 198890 8016
rect 304718 7964 304724 8016
rect 304776 8004 304782 8016
rect 361114 8004 361120 8016
rect 304776 7976 361120 8004
rect 304776 7964 304782 7976
rect 361114 7964 361120 7976
rect 361172 7964 361178 8016
rect 377950 7964 377956 8016
rect 378008 8004 378014 8016
rect 556246 8004 556252 8016
rect 378008 7976 556252 8004
rect 378008 7964 378014 7976
rect 556246 7964 556252 7976
rect 556304 7964 556310 8016
rect 79686 7896 79692 7948
rect 79744 7936 79750 7948
rect 197446 7936 197452 7948
rect 79744 7908 197452 7936
rect 79744 7896 79750 7908
rect 197446 7896 197452 7908
rect 197504 7896 197510 7948
rect 306098 7896 306104 7948
rect 306156 7936 306162 7948
rect 364610 7936 364616 7948
rect 306156 7908 364616 7936
rect 306156 7896 306162 7908
rect 364610 7896 364616 7908
rect 364668 7896 364674 7948
rect 379330 7896 379336 7948
rect 379388 7936 379394 7948
rect 559742 7936 559748 7948
rect 379388 7908 559748 7936
rect 379388 7896 379394 7908
rect 559742 7896 559748 7908
rect 559800 7896 559806 7948
rect 77386 7828 77392 7880
rect 77444 7868 77450 7880
rect 196158 7868 196164 7880
rect 77444 7840 196164 7868
rect 77444 7828 77450 7840
rect 196158 7828 196164 7840
rect 196216 7828 196222 7880
rect 307478 7828 307484 7880
rect 307536 7868 307542 7880
rect 368198 7868 368204 7880
rect 307536 7840 368204 7868
rect 307536 7828 307542 7840
rect 368198 7828 368204 7840
rect 368256 7828 368262 7880
rect 380710 7828 380716 7880
rect 380768 7868 380774 7880
rect 563238 7868 563244 7880
rect 380768 7840 563244 7868
rect 380768 7828 380774 7840
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 73798 7760 73804 7812
rect 73856 7800 73862 7812
rect 194778 7800 194784 7812
rect 73856 7772 194784 7800
rect 73856 7760 73862 7772
rect 194778 7760 194784 7772
rect 194836 7760 194842 7812
rect 308858 7760 308864 7812
rect 308916 7800 308922 7812
rect 371694 7800 371700 7812
rect 308916 7772 371700 7800
rect 308916 7760 308922 7772
rect 371694 7760 371700 7772
rect 371752 7760 371758 7812
rect 381998 7760 382004 7812
rect 382056 7800 382062 7812
rect 566826 7800 566832 7812
rect 382056 7772 566832 7800
rect 382056 7760 382062 7772
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 70302 7692 70308 7744
rect 70360 7732 70366 7744
rect 193398 7732 193404 7744
rect 70360 7704 193404 7732
rect 70360 7692 70366 7704
rect 193398 7692 193404 7704
rect 193456 7692 193462 7744
rect 310146 7692 310152 7744
rect 310204 7732 310210 7744
rect 375190 7732 375196 7744
rect 310204 7704 375196 7732
rect 310204 7692 310210 7704
rect 375190 7692 375196 7704
rect 375248 7692 375254 7744
rect 383378 7692 383384 7744
rect 383436 7732 383442 7744
rect 570322 7732 570328 7744
rect 383436 7704 570328 7732
rect 383436 7692 383442 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 66714 7624 66720 7676
rect 66772 7664 66778 7676
rect 192018 7664 192024 7676
rect 66772 7636 192024 7664
rect 66772 7624 66778 7636
rect 192018 7624 192024 7636
rect 192076 7624 192082 7676
rect 311618 7624 311624 7676
rect 311676 7664 311682 7676
rect 378870 7664 378876 7676
rect 311676 7636 378876 7664
rect 311676 7624 311682 7636
rect 378870 7624 378876 7636
rect 378928 7624 378934 7676
rect 384758 7624 384764 7676
rect 384816 7664 384822 7676
rect 573910 7664 573916 7676
rect 384816 7636 573916 7664
rect 384816 7624 384822 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 63218 7556 63224 7608
rect 63276 7596 63282 7608
rect 190730 7596 190736 7608
rect 63276 7568 190736 7596
rect 63276 7556 63282 7568
rect 190730 7556 190736 7568
rect 190788 7556 190794 7608
rect 221550 7556 221556 7608
rect 221608 7596 221614 7608
rect 247678 7596 247684 7608
rect 221608 7568 247684 7596
rect 221608 7556 221614 7568
rect 247678 7556 247684 7568
rect 247736 7556 247742 7608
rect 312998 7556 313004 7608
rect 313056 7596 313062 7608
rect 382366 7596 382372 7608
rect 313056 7568 382372 7596
rect 313056 7556 313062 7568
rect 382366 7556 382372 7568
rect 382424 7556 382430 7608
rect 386046 7556 386052 7608
rect 386104 7596 386110 7608
rect 577406 7596 577412 7608
rect 386104 7568 577412 7596
rect 386104 7556 386110 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 101030 7488 101036 7540
rect 101088 7528 101094 7540
rect 205818 7528 205824 7540
rect 101088 7500 205824 7528
rect 101088 7488 101094 7500
rect 205818 7488 205824 7500
rect 205876 7488 205882 7540
rect 371050 7488 371056 7540
rect 371108 7528 371114 7540
rect 538398 7528 538404 7540
rect 371108 7500 538404 7528
rect 371108 7488 371114 7500
rect 538398 7488 538404 7500
rect 538456 7488 538462 7540
rect 104526 7420 104532 7472
rect 104584 7460 104590 7472
rect 207106 7460 207112 7472
rect 104584 7432 207112 7460
rect 104584 7420 104590 7432
rect 207106 7420 207112 7432
rect 207164 7420 207170 7472
rect 369670 7420 369676 7472
rect 369728 7460 369734 7472
rect 534902 7460 534908 7472
rect 369728 7432 534908 7460
rect 369728 7420 369734 7432
rect 534902 7420 534908 7432
rect 534960 7420 534966 7472
rect 108114 7352 108120 7404
rect 108172 7392 108178 7404
rect 208578 7392 208584 7404
rect 108172 7364 208584 7392
rect 108172 7352 108178 7364
rect 208578 7352 208584 7364
rect 208636 7352 208642 7404
rect 368290 7352 368296 7404
rect 368348 7392 368354 7404
rect 531406 7392 531412 7404
rect 368348 7364 531412 7392
rect 368348 7352 368354 7364
rect 531406 7352 531412 7364
rect 531464 7352 531470 7404
rect 111610 7284 111616 7336
rect 111668 7324 111674 7336
rect 209866 7324 209872 7336
rect 111668 7296 209872 7324
rect 111668 7284 111674 7296
rect 209866 7284 209872 7296
rect 209924 7284 209930 7336
rect 366910 7284 366916 7336
rect 366968 7324 366974 7336
rect 527818 7324 527824 7336
rect 366968 7296 527824 7324
rect 366968 7284 366974 7296
rect 527818 7284 527824 7296
rect 527876 7284 527882 7336
rect 115198 7216 115204 7268
rect 115256 7256 115262 7268
rect 211338 7256 211344 7268
rect 115256 7228 211344 7256
rect 115256 7216 115262 7228
rect 211338 7216 211344 7228
rect 211396 7216 211402 7268
rect 365530 7216 365536 7268
rect 365588 7256 365594 7268
rect 524230 7256 524236 7268
rect 365588 7228 524236 7256
rect 365588 7216 365594 7228
rect 524230 7216 524236 7228
rect 524288 7216 524294 7268
rect 118786 7148 118792 7200
rect 118844 7188 118850 7200
rect 212718 7188 212724 7200
rect 118844 7160 212724 7188
rect 118844 7148 118850 7160
rect 212718 7148 212724 7160
rect 212776 7148 212782 7200
rect 364150 7148 364156 7200
rect 364208 7188 364214 7200
rect 520734 7188 520740 7200
rect 364208 7160 520740 7188
rect 364208 7148 364214 7160
rect 520734 7148 520740 7160
rect 520792 7148 520798 7200
rect 122282 7080 122288 7132
rect 122340 7120 122346 7132
rect 214006 7120 214012 7132
rect 122340 7092 214012 7120
rect 122340 7080 122346 7092
rect 214006 7080 214012 7092
rect 214064 7080 214070 7132
rect 315758 7080 315764 7132
rect 315816 7120 315822 7132
rect 393038 7120 393044 7132
rect 315816 7092 393044 7120
rect 315816 7080 315822 7092
rect 393038 7080 393044 7092
rect 393096 7080 393102 7132
rect 160094 7012 160100 7064
rect 160152 7052 160158 7064
rect 227806 7052 227812 7064
rect 160152 7024 227812 7052
rect 160152 7012 160158 7024
rect 227806 7012 227812 7024
rect 227864 7012 227870 7064
rect 315850 7012 315856 7064
rect 315908 7052 315914 7064
rect 389450 7052 389456 7064
rect 315908 7024 389456 7052
rect 315908 7012 315914 7024
rect 389450 7012 389456 7024
rect 389508 7012 389514 7064
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 18598 6848 18604 6860
rect 3476 6820 18604 6848
rect 3476 6808 3482 6820
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 48958 6808 48964 6860
rect 49016 6848 49022 6860
rect 186406 6848 186412 6860
rect 49016 6820 186412 6848
rect 49016 6808 49022 6820
rect 186406 6808 186412 6820
rect 186464 6808 186470 6860
rect 337930 6808 337936 6860
rect 337988 6848 337994 6860
rect 448606 6848 448612 6860
rect 337988 6820 448612 6848
rect 337988 6808 337994 6820
rect 448606 6808 448612 6820
rect 448664 6808 448670 6860
rect 519538 6808 519544 6860
rect 519596 6848 519602 6860
rect 580166 6848 580172 6860
rect 519596 6820 580172 6848
rect 519596 6808 519602 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 44266 6740 44272 6792
rect 44324 6780 44330 6792
rect 183646 6780 183652 6792
rect 44324 6752 183652 6780
rect 44324 6740 44330 6752
rect 183646 6740 183652 6752
rect 183704 6740 183710 6792
rect 339402 6740 339408 6792
rect 339460 6780 339466 6792
rect 452102 6780 452108 6792
rect 339460 6752 452108 6780
rect 339460 6740 339466 6752
rect 452102 6740 452108 6752
rect 452160 6740 452166 6792
rect 40770 6672 40776 6724
rect 40828 6712 40834 6724
rect 182358 6712 182364 6724
rect 40828 6684 182364 6712
rect 40828 6672 40834 6684
rect 182358 6672 182364 6684
rect 182416 6672 182422 6724
rect 340690 6672 340696 6724
rect 340748 6712 340754 6724
rect 455690 6712 455696 6724
rect 340748 6684 455696 6712
rect 340748 6672 340754 6684
rect 455690 6672 455696 6684
rect 455748 6672 455754 6724
rect 37182 6604 37188 6656
rect 37240 6644 37246 6656
rect 180886 6644 180892 6656
rect 37240 6616 180892 6644
rect 37240 6604 37246 6616
rect 180886 6604 180892 6616
rect 180944 6604 180950 6656
rect 197906 6604 197912 6656
rect 197964 6644 197970 6656
rect 241606 6644 241612 6656
rect 197964 6616 241612 6644
rect 197964 6604 197970 6616
rect 241606 6604 241612 6616
rect 241664 6604 241670 6656
rect 342162 6604 342168 6656
rect 342220 6644 342226 6656
rect 459186 6644 459192 6656
rect 342220 6616 459192 6644
rect 342220 6604 342226 6616
rect 459186 6604 459192 6616
rect 459244 6604 459250 6656
rect 33594 6536 33600 6588
rect 33652 6576 33658 6588
rect 179598 6576 179604 6588
rect 33652 6548 179604 6576
rect 33652 6536 33658 6548
rect 179598 6536 179604 6548
rect 179656 6536 179662 6588
rect 192018 6536 192024 6588
rect 192076 6576 192082 6588
rect 240226 6576 240232 6588
rect 192076 6548 240232 6576
rect 192076 6536 192082 6548
rect 240226 6536 240232 6548
rect 240284 6536 240290 6588
rect 343450 6536 343456 6588
rect 343508 6576 343514 6588
rect 462774 6576 462780 6588
rect 343508 6548 462780 6576
rect 343508 6536 343514 6548
rect 462774 6536 462780 6548
rect 462832 6536 462838 6588
rect 30098 6468 30104 6520
rect 30156 6508 30162 6520
rect 178126 6508 178132 6520
rect 30156 6480 178132 6508
rect 30156 6468 30162 6480
rect 178126 6468 178132 6480
rect 178184 6468 178190 6520
rect 188522 6468 188528 6520
rect 188580 6508 188586 6520
rect 238846 6508 238852 6520
rect 188580 6480 238852 6508
rect 188580 6468 188586 6480
rect 238846 6468 238852 6480
rect 238904 6468 238910 6520
rect 343358 6468 343364 6520
rect 343416 6508 343422 6520
rect 466270 6508 466276 6520
rect 343416 6480 466276 6508
rect 343416 6468 343422 6480
rect 466270 6468 466276 6480
rect 466328 6468 466334 6520
rect 26510 6400 26516 6452
rect 26568 6440 26574 6452
rect 176746 6440 176752 6452
rect 26568 6412 176752 6440
rect 26568 6400 26574 6412
rect 176746 6400 176752 6412
rect 176804 6400 176810 6452
rect 184934 6400 184940 6452
rect 184992 6440 184998 6452
rect 237374 6440 237380 6452
rect 184992 6412 237380 6440
rect 184992 6400 184998 6412
rect 237374 6400 237380 6412
rect 237432 6400 237438 6452
rect 344922 6400 344928 6452
rect 344980 6440 344986 6452
rect 469858 6440 469864 6452
rect 344980 6412 469864 6440
rect 344980 6400 344986 6412
rect 469858 6400 469864 6412
rect 469916 6400 469922 6452
rect 21818 6332 21824 6384
rect 21876 6372 21882 6384
rect 175458 6372 175464 6384
rect 21876 6344 175464 6372
rect 21876 6332 21882 6344
rect 175458 6332 175464 6344
rect 175516 6332 175522 6384
rect 181438 6332 181444 6384
rect 181496 6372 181502 6384
rect 236178 6372 236184 6384
rect 181496 6344 236184 6372
rect 181496 6332 181502 6344
rect 236178 6332 236184 6344
rect 236236 6332 236242 6384
rect 346210 6332 346216 6384
rect 346268 6372 346274 6384
rect 473446 6372 473452 6384
rect 346268 6344 473452 6372
rect 346268 6332 346274 6344
rect 473446 6332 473452 6344
rect 473504 6332 473510 6384
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 174078 6304 174084 6316
rect 17092 6276 174084 6304
rect 17092 6264 17098 6276
rect 174078 6264 174084 6276
rect 174136 6264 174142 6316
rect 177850 6264 177856 6316
rect 177908 6304 177914 6316
rect 234798 6304 234804 6316
rect 177908 6276 234804 6304
rect 177908 6264 177914 6276
rect 234798 6264 234804 6276
rect 234856 6264 234862 6316
rect 347682 6264 347688 6316
rect 347740 6304 347746 6316
rect 476942 6304 476948 6316
rect 347740 6276 476948 6304
rect 347740 6264 347746 6276
rect 476942 6264 476948 6276
rect 477000 6264 477006 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 171226 6236 171232 6248
rect 8812 6208 171232 6236
rect 8812 6196 8818 6208
rect 171226 6196 171232 6208
rect 171284 6196 171290 6248
rect 174262 6196 174268 6248
rect 174320 6236 174326 6248
rect 233234 6236 233240 6248
rect 174320 6208 233240 6236
rect 174320 6196 174326 6208
rect 233234 6196 233240 6208
rect 233292 6196 233298 6248
rect 281258 6196 281264 6248
rect 281316 6236 281322 6248
rect 299658 6236 299664 6248
rect 281316 6208 299664 6236
rect 281316 6196 281322 6208
rect 299658 6196 299664 6208
rect 299716 6196 299722 6248
rect 350258 6196 350264 6248
rect 350316 6236 350322 6248
rect 481726 6236 481732 6248
rect 350316 6208 481732 6236
rect 350316 6196 350322 6208
rect 481726 6196 481732 6208
rect 481784 6196 481790 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 168558 6168 168564 6180
rect 4120 6140 168564 6168
rect 4120 6128 4126 6140
rect 168558 6128 168564 6140
rect 168616 6128 168622 6180
rect 170766 6128 170772 6180
rect 170824 6168 170830 6180
rect 232130 6168 232136 6180
rect 170824 6140 232136 6168
rect 170824 6128 170830 6140
rect 232130 6128 232136 6140
rect 232188 6128 232194 6180
rect 288158 6128 288164 6180
rect 288216 6168 288222 6180
rect 317322 6168 317328 6180
rect 288216 6140 317328 6168
rect 288216 6128 288222 6140
rect 317322 6128 317328 6140
rect 317380 6128 317386 6180
rect 320818 6128 320824 6180
rect 320876 6168 320882 6180
rect 332686 6168 332692 6180
rect 320876 6140 332692 6168
rect 320876 6128 320882 6140
rect 332686 6128 332692 6140
rect 332744 6128 332750 6180
rect 351822 6128 351828 6180
rect 351880 6168 351886 6180
rect 485222 6168 485228 6180
rect 351880 6140 485228 6168
rect 351880 6128 351886 6140
rect 485222 6128 485228 6140
rect 485280 6128 485286 6180
rect 52546 6060 52552 6112
rect 52604 6100 52610 6112
rect 187878 6100 187884 6112
rect 52604 6072 187884 6100
rect 52604 6060 52610 6072
rect 187878 6060 187884 6072
rect 187936 6060 187942 6112
rect 336642 6060 336648 6112
rect 336700 6100 336706 6112
rect 445018 6100 445024 6112
rect 336700 6072 445024 6100
rect 336700 6060 336706 6072
rect 445018 6060 445024 6072
rect 445076 6060 445082 6112
rect 56042 5992 56048 6044
rect 56100 6032 56106 6044
rect 189258 6032 189264 6044
rect 56100 6004 189264 6032
rect 56100 5992 56106 6004
rect 189258 5992 189264 6004
rect 189316 5992 189322 6044
rect 335170 5992 335176 6044
rect 335228 6032 335234 6044
rect 441522 6032 441528 6044
rect 335228 6004 441528 6032
rect 335228 5992 335234 6004
rect 441522 5992 441528 6004
rect 441580 5992 441586 6044
rect 59630 5924 59636 5976
rect 59688 5964 59694 5976
rect 190638 5964 190644 5976
rect 59688 5936 190644 5964
rect 59688 5924 59694 5936
rect 190638 5924 190644 5936
rect 190696 5924 190702 5976
rect 333882 5924 333888 5976
rect 333940 5964 333946 5976
rect 437934 5964 437940 5976
rect 333940 5936 437940 5964
rect 333940 5924 333946 5936
rect 437934 5924 437940 5936
rect 437992 5924 437998 5976
rect 76190 5856 76196 5908
rect 76248 5896 76254 5908
rect 196066 5896 196072 5908
rect 76248 5868 196072 5896
rect 76248 5856 76254 5868
rect 196066 5856 196072 5868
rect 196124 5856 196130 5908
rect 332410 5856 332416 5908
rect 332468 5896 332474 5908
rect 434438 5896 434444 5908
rect 332468 5868 434444 5896
rect 332468 5856 332474 5868
rect 434438 5856 434444 5868
rect 434496 5856 434502 5908
rect 128170 5788 128176 5840
rect 128228 5828 128234 5840
rect 215386 5828 215392 5840
rect 128228 5800 215392 5828
rect 128228 5788 128234 5800
rect 215386 5788 215392 5800
rect 215444 5788 215450 5840
rect 331122 5788 331128 5840
rect 331180 5828 331186 5840
rect 430850 5828 430856 5840
rect 331180 5800 430856 5828
rect 331180 5788 331186 5800
rect 430850 5788 430856 5800
rect 430908 5788 430914 5840
rect 158898 5720 158904 5772
rect 158956 5760 158962 5772
rect 227898 5760 227904 5772
rect 158956 5732 227904 5760
rect 158956 5720 158962 5732
rect 227898 5720 227904 5732
rect 227956 5720 227962 5772
rect 329650 5720 329656 5772
rect 329708 5760 329714 5772
rect 427262 5760 427268 5772
rect 329708 5732 427268 5760
rect 329708 5720 329714 5732
rect 427262 5720 427268 5732
rect 427320 5720 427326 5772
rect 163682 5652 163688 5704
rect 163740 5692 163746 5704
rect 229186 5692 229192 5704
rect 163740 5664 229192 5692
rect 163740 5652 163746 5664
rect 229186 5652 229192 5664
rect 229244 5652 229250 5704
rect 328270 5652 328276 5704
rect 328328 5692 328334 5704
rect 423766 5692 423772 5704
rect 328328 5664 423772 5692
rect 328328 5652 328334 5664
rect 423766 5652 423772 5664
rect 423824 5652 423830 5704
rect 167178 5584 167184 5636
rect 167236 5624 167242 5636
rect 230566 5624 230572 5636
rect 167236 5596 230572 5624
rect 167236 5584 167242 5596
rect 230566 5584 230572 5596
rect 230624 5584 230630 5636
rect 313918 5516 313924 5568
rect 313976 5556 313982 5568
rect 315022 5556 315028 5568
rect 313976 5528 315028 5556
rect 313976 5516 313982 5528
rect 315022 5516 315028 5528
rect 315080 5516 315086 5568
rect 323578 5516 323584 5568
rect 323636 5556 323642 5568
rect 324406 5556 324412 5568
rect 323636 5528 324412 5556
rect 323636 5516 323642 5528
rect 324406 5516 324412 5528
rect 324464 5516 324470 5568
rect 65518 5448 65524 5500
rect 65576 5488 65582 5500
rect 191926 5488 191932 5500
rect 65576 5460 191932 5488
rect 65576 5448 65582 5460
rect 191926 5448 191932 5460
rect 191984 5448 191990 5500
rect 302142 5448 302148 5500
rect 302200 5488 302206 5500
rect 354030 5488 354036 5500
rect 302200 5460 354036 5488
rect 302200 5448 302206 5460
rect 354030 5448 354036 5460
rect 354088 5448 354094 5500
rect 372246 5448 372252 5500
rect 372304 5488 372310 5500
rect 540790 5488 540796 5500
rect 372304 5460 540796 5488
rect 372304 5448 372310 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 62022 5380 62028 5432
rect 62080 5420 62086 5432
rect 190546 5420 190552 5432
rect 62080 5392 190552 5420
rect 62080 5380 62086 5392
rect 190546 5380 190552 5392
rect 190604 5380 190610 5432
rect 302050 5380 302056 5432
rect 302108 5420 302114 5432
rect 356330 5420 356336 5432
rect 302108 5392 356336 5420
rect 302108 5380 302114 5392
rect 356330 5380 356336 5392
rect 356388 5380 356394 5432
rect 373902 5380 373908 5432
rect 373960 5420 373966 5432
rect 544378 5420 544384 5432
rect 373960 5392 544384 5420
rect 373960 5380 373966 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 58434 5312 58440 5364
rect 58492 5352 58498 5364
rect 189166 5352 189172 5364
rect 58492 5324 189172 5352
rect 58492 5312 58498 5324
rect 189166 5312 189172 5324
rect 189224 5312 189230 5364
rect 303522 5312 303528 5364
rect 303580 5352 303586 5364
rect 357526 5352 357532 5364
rect 303580 5324 357532 5352
rect 303580 5312 303586 5324
rect 357526 5312 357532 5324
rect 357584 5312 357590 5364
rect 375282 5312 375288 5364
rect 375340 5352 375346 5364
rect 547874 5352 547880 5364
rect 375340 5324 547880 5352
rect 375340 5312 375346 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 54938 5244 54944 5296
rect 54996 5284 55002 5296
rect 187786 5284 187792 5296
rect 54996 5256 187792 5284
rect 54996 5244 55002 5256
rect 187786 5244 187792 5256
rect 187844 5244 187850 5296
rect 303430 5244 303436 5296
rect 303488 5284 303494 5296
rect 359918 5284 359924 5296
rect 303488 5256 359924 5284
rect 303488 5244 303494 5256
rect 359918 5244 359924 5256
rect 359976 5244 359982 5296
rect 376662 5244 376668 5296
rect 376720 5284 376726 5296
rect 551462 5284 551468 5296
rect 376720 5256 551468 5284
rect 376720 5244 376726 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 51350 5176 51356 5228
rect 51408 5216 51414 5228
rect 186314 5216 186320 5228
rect 51408 5188 186320 5216
rect 51408 5176 51414 5188
rect 186314 5176 186320 5188
rect 186372 5176 186378 5228
rect 211062 5176 211068 5228
rect 211120 5216 211126 5228
rect 247126 5216 247132 5228
rect 211120 5188 247132 5216
rect 211120 5176 211126 5188
rect 247126 5176 247132 5188
rect 247184 5176 247190 5228
rect 304810 5176 304816 5228
rect 304868 5216 304874 5228
rect 363506 5216 363512 5228
rect 304868 5188 363512 5216
rect 304868 5176 304874 5188
rect 363506 5176 363512 5188
rect 363564 5176 363570 5228
rect 378042 5176 378048 5228
rect 378100 5216 378106 5228
rect 554958 5216 554964 5228
rect 378100 5188 554964 5216
rect 378100 5176 378106 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 47854 5108 47860 5160
rect 47912 5148 47918 5160
rect 185118 5148 185124 5160
rect 47912 5120 185124 5148
rect 47912 5108 47918 5120
rect 185118 5108 185124 5120
rect 185176 5108 185182 5160
rect 207382 5108 207388 5160
rect 207440 5148 207446 5160
rect 245838 5148 245844 5160
rect 207440 5120 245844 5148
rect 207440 5108 207446 5120
rect 245838 5108 245844 5120
rect 245896 5108 245902 5160
rect 306190 5108 306196 5160
rect 306248 5148 306254 5160
rect 367002 5148 367008 5160
rect 306248 5120 367008 5148
rect 306248 5108 306254 5120
rect 367002 5108 367008 5120
rect 367060 5108 367066 5160
rect 379422 5108 379428 5160
rect 379480 5148 379486 5160
rect 558546 5148 558552 5160
rect 379480 5120 558552 5148
rect 379480 5108 379486 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 172698 5080 172704 5092
rect 12400 5052 172704 5080
rect 12400 5040 12406 5052
rect 172698 5040 172704 5052
rect 172756 5040 172762 5092
rect 203886 5040 203892 5092
rect 203944 5080 203950 5092
rect 244366 5080 244372 5092
rect 203944 5052 244372 5080
rect 203944 5040 203950 5052
rect 244366 5040 244372 5052
rect 244424 5040 244430 5092
rect 307570 5040 307576 5092
rect 307628 5080 307634 5092
rect 370590 5080 370596 5092
rect 307628 5052 370596 5080
rect 307628 5040 307634 5052
rect 370590 5040 370596 5052
rect 370648 5040 370654 5092
rect 380802 5040 380808 5092
rect 380860 5080 380866 5092
rect 562042 5080 562048 5092
rect 380860 5052 562048 5080
rect 380860 5040 380866 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 169846 5012 169852 5024
rect 7708 4984 169852 5012
rect 7708 4972 7714 4984
rect 169846 4972 169852 4984
rect 169904 4972 169910 5024
rect 200298 4972 200304 5024
rect 200356 5012 200362 5024
rect 243078 5012 243084 5024
rect 200356 4984 243084 5012
rect 200356 4972 200362 4984
rect 243078 4972 243084 4984
rect 243136 4972 243142 5024
rect 308950 4972 308956 5024
rect 309008 5012 309014 5024
rect 374086 5012 374092 5024
rect 309008 4984 374092 5012
rect 309008 4972 309014 4984
rect 374086 4972 374092 4984
rect 374144 4972 374150 5024
rect 382090 4972 382096 5024
rect 382148 5012 382154 5024
rect 565630 5012 565636 5024
rect 382148 4984 565636 5012
rect 382148 4972 382154 4984
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 168374 4944 168380 4956
rect 2924 4916 168380 4944
rect 2924 4904 2930 4916
rect 168374 4904 168380 4916
rect 168432 4904 168438 4956
rect 196802 4904 196808 4956
rect 196860 4944 196866 4956
rect 241698 4944 241704 4956
rect 196860 4916 241704 4944
rect 196860 4904 196866 4916
rect 241698 4904 241704 4916
rect 241756 4904 241762 4956
rect 310330 4904 310336 4956
rect 310388 4944 310394 4956
rect 377674 4944 377680 4956
rect 310388 4916 377680 4944
rect 310388 4904 310394 4916
rect 377674 4904 377680 4916
rect 377732 4904 377738 4956
rect 383470 4904 383476 4956
rect 383528 4944 383534 4956
rect 569126 4944 569132 4956
rect 383528 4916 569132 4944
rect 383528 4904 383534 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 166994 4876 167000 4888
rect 624 4848 167000 4876
rect 624 4836 630 4848
rect 166994 4836 167000 4848
rect 167052 4836 167058 4888
rect 193214 4836 193220 4888
rect 193272 4876 193278 4888
rect 240134 4876 240140 4888
rect 193272 4848 240140 4876
rect 193272 4836 193278 4848
rect 240134 4836 240140 4848
rect 240192 4836 240198 4888
rect 311710 4836 311716 4888
rect 311768 4876 311774 4888
rect 381170 4876 381176 4888
rect 311768 4848 381176 4876
rect 311768 4836 311774 4848
rect 381170 4836 381176 4848
rect 381228 4836 381234 4888
rect 384850 4836 384856 4888
rect 384908 4876 384914 4888
rect 572714 4876 572720 4888
rect 384908 4848 572720 4876
rect 384908 4836 384914 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 168466 4808 168472 4820
rect 1728 4780 168472 4808
rect 1728 4768 1734 4780
rect 168466 4768 168472 4780
rect 168524 4768 168530 4820
rect 189718 4768 189724 4820
rect 189776 4808 189782 4820
rect 238938 4808 238944 4820
rect 189776 4780 238944 4808
rect 189776 4768 189782 4780
rect 238938 4768 238944 4780
rect 238996 4768 239002 4820
rect 277118 4768 277124 4820
rect 277176 4808 277182 4820
rect 288986 4808 288992 4820
rect 277176 4780 288992 4808
rect 277176 4768 277182 4780
rect 288986 4768 288992 4780
rect 289044 4768 289050 4820
rect 313090 4768 313096 4820
rect 313148 4808 313154 4820
rect 384758 4808 384764 4820
rect 313148 4780 384764 4808
rect 313148 4768 313154 4780
rect 384758 4768 384764 4780
rect 384816 4768 384822 4820
rect 386138 4768 386144 4820
rect 386196 4808 386202 4820
rect 576302 4808 576308 4820
rect 386196 4780 576308 4808
rect 386196 4768 386202 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 69106 4700 69112 4752
rect 69164 4740 69170 4752
rect 193306 4740 193312 4752
rect 69164 4712 193312 4740
rect 69164 4700 69170 4712
rect 193306 4700 193312 4712
rect 193364 4700 193370 4752
rect 301958 4700 301964 4752
rect 302016 4740 302022 4752
rect 352834 4740 352840 4752
rect 302016 4712 352840 4740
rect 302016 4700 302022 4712
rect 352834 4700 352840 4712
rect 352892 4700 352898 4752
rect 371142 4700 371148 4752
rect 371200 4740 371206 4752
rect 537202 4740 537208 4752
rect 371200 4712 537208 4740
rect 371200 4700 371206 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 72602 4632 72608 4684
rect 72660 4672 72666 4684
rect 194686 4672 194692 4684
rect 72660 4644 194692 4672
rect 72660 4632 72666 4644
rect 194686 4632 194692 4644
rect 194744 4632 194750 4684
rect 300670 4632 300676 4684
rect 300728 4672 300734 4684
rect 349246 4672 349252 4684
rect 300728 4644 349252 4672
rect 300728 4632 300734 4644
rect 349246 4632 349252 4644
rect 349304 4632 349310 4684
rect 369762 4632 369768 4684
rect 369820 4672 369826 4684
rect 533706 4672 533712 4684
rect 369820 4644 533712 4672
rect 369820 4632 369826 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 126974 4564 126980 4616
rect 127032 4604 127038 4616
rect 215478 4604 215484 4616
rect 127032 4576 215484 4604
rect 127032 4564 127038 4576
rect 215478 4564 215484 4576
rect 215536 4564 215542 4616
rect 300762 4564 300768 4616
rect 300820 4604 300826 4616
rect 350442 4604 350448 4616
rect 300820 4576 350448 4604
rect 300820 4564 300826 4576
rect 350442 4564 350448 4576
rect 350500 4564 350506 4616
rect 368382 4564 368388 4616
rect 368440 4604 368446 4616
rect 530118 4604 530124 4616
rect 368440 4576 530124 4604
rect 368440 4564 368446 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 150618 4496 150624 4548
rect 150676 4536 150682 4548
rect 223574 4536 223580 4548
rect 150676 4508 223580 4536
rect 150676 4496 150682 4508
rect 223574 4496 223580 4508
rect 223632 4496 223638 4548
rect 299382 4496 299388 4548
rect 299440 4536 299446 4548
rect 299440 4508 345014 4536
rect 299440 4496 299446 4508
rect 154206 4428 154212 4480
rect 154264 4468 154270 4480
rect 224954 4468 224960 4480
rect 154264 4440 224960 4468
rect 154264 4428 154270 4440
rect 224954 4428 224960 4440
rect 225012 4428 225018 4480
rect 298002 4428 298008 4480
rect 298060 4468 298066 4480
rect 343358 4468 343364 4480
rect 298060 4440 343364 4468
rect 298060 4428 298066 4440
rect 343358 4428 343364 4440
rect 343416 4428 343422 4480
rect 157794 4360 157800 4412
rect 157852 4400 157858 4412
rect 226518 4400 226524 4412
rect 157852 4372 226524 4400
rect 157852 4360 157858 4372
rect 226518 4360 226524 4372
rect 226576 4360 226582 4412
rect 296622 4360 296628 4412
rect 296680 4400 296686 4412
rect 339862 4400 339868 4412
rect 296680 4372 339868 4400
rect 296680 4360 296686 4372
rect 339862 4360 339868 4372
rect 339920 4360 339926 4412
rect 344986 4400 345014 4508
rect 366910 4496 366916 4548
rect 366968 4536 366974 4548
rect 526622 4536 526628 4548
rect 366968 4508 526628 4536
rect 366968 4496 366974 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 365622 4428 365628 4480
rect 365680 4468 365686 4480
rect 523034 4468 523040 4480
rect 365680 4440 523040 4468
rect 365680 4428 365686 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 346946 4400 346952 4412
rect 344986 4372 346952 4400
rect 346946 4360 346952 4372
rect 347004 4360 347010 4412
rect 364242 4360 364248 4412
rect 364300 4400 364306 4412
rect 519538 4400 519544 4412
rect 364300 4372 519544 4400
rect 364300 4360 364306 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 162486 4292 162492 4344
rect 162544 4332 162550 4344
rect 229278 4332 229284 4344
rect 162544 4304 229284 4332
rect 162544 4292 162550 4304
rect 229278 4292 229284 4304
rect 229336 4292 229342 4344
rect 295242 4292 295248 4344
rect 295300 4332 295306 4344
rect 336274 4332 336280 4344
rect 295300 4304 336280 4332
rect 295300 4292 295306 4304
rect 336274 4292 336280 4304
rect 336332 4292 336338 4344
rect 362862 4292 362868 4344
rect 362920 4332 362926 4344
rect 515950 4332 515956 4344
rect 362920 4304 515956 4332
rect 362920 4292 362926 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 166074 4224 166080 4276
rect 166132 4264 166138 4276
rect 230658 4264 230664 4276
rect 166132 4236 230664 4264
rect 166132 4224 166138 4236
rect 230658 4224 230664 4236
rect 230716 4224 230722 4276
rect 340785 4267 340843 4273
rect 340785 4233 340797 4267
rect 340831 4264 340843 4267
rect 342257 4267 342315 4273
rect 342257 4264 342269 4267
rect 340831 4236 342269 4264
rect 340831 4233 340843 4236
rect 340785 4227 340843 4233
rect 342257 4233 342269 4236
rect 342303 4233 342315 4267
rect 342257 4227 342315 4233
rect 357345 4267 357403 4273
rect 357345 4233 357357 4267
rect 357391 4264 357403 4267
rect 358817 4267 358875 4273
rect 358817 4264 358829 4267
rect 357391 4236 358829 4264
rect 357391 4233 357403 4236
rect 357345 4227 357403 4233
rect 358817 4233 358829 4236
rect 358863 4233 358875 4267
rect 358817 4227 358875 4233
rect 361482 4224 361488 4276
rect 361540 4264 361546 4276
rect 512454 4264 512460 4276
rect 361540 4236 512460 4264
rect 361540 4224 361546 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 135254 4156 135260 4208
rect 135312 4196 135318 4208
rect 136450 4196 136456 4208
rect 135312 4168 136456 4196
rect 135312 4156 135318 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 144822 4196 144828 4208
rect 143592 4168 144828 4196
rect 143592 4156 143598 4168
rect 144822 4156 144828 4168
rect 144880 4156 144886 4208
rect 151814 4156 151820 4208
rect 151872 4196 151878 4208
rect 153102 4196 153108 4208
rect 151872 4168 153108 4196
rect 151872 4156 151878 4168
rect 153102 4156 153108 4168
rect 153160 4156 153166 4208
rect 171781 4199 171839 4205
rect 171781 4165 171793 4199
rect 171827 4196 171839 4199
rect 178310 4196 178316 4208
rect 171827 4168 178316 4196
rect 171827 4165 171839 4168
rect 171781 4159 171839 4165
rect 178310 4156 178316 4168
rect 178368 4156 178374 4208
rect 291838 4156 291844 4208
rect 291896 4196 291902 4208
rect 292574 4196 292580 4208
rect 291896 4168 292580 4196
rect 291896 4156 291902 4168
rect 292574 4156 292580 4168
rect 292632 4156 292638 4208
rect 314470 4156 314476 4208
rect 314528 4196 314534 4208
rect 385954 4196 385960 4208
rect 314528 4168 385960 4196
rect 314528 4156 314534 4168
rect 385954 4156 385960 4168
rect 386012 4156 386018 4208
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 7558 4128 7564 4140
rect 6512 4100 7564 4128
rect 6512 4088 6518 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 78582 4088 78588 4140
rect 78640 4128 78646 4140
rect 197354 4128 197360 4140
rect 78640 4100 197360 4128
rect 78640 4088 78646 4100
rect 197354 4088 197360 4100
rect 197412 4088 197418 4140
rect 233418 4088 233424 4140
rect 233476 4128 233482 4140
rect 250349 4131 250407 4137
rect 250349 4128 250361 4131
rect 233476 4100 250361 4128
rect 233476 4088 233482 4100
rect 250349 4097 250361 4100
rect 250395 4097 250407 4131
rect 250349 4091 250407 4097
rect 250441 4131 250499 4137
rect 250441 4097 250453 4131
rect 250487 4128 250499 4131
rect 254026 4128 254032 4140
rect 250487 4100 254032 4128
rect 250487 4097 250499 4100
rect 250441 4091 250499 4097
rect 254026 4088 254032 4100
rect 254084 4088 254090 4140
rect 279970 4088 279976 4140
rect 280028 4128 280034 4140
rect 297266 4128 297272 4140
rect 280028 4100 297272 4128
rect 280028 4088 280034 4100
rect 297266 4088 297272 4100
rect 297324 4088 297330 4140
rect 332502 4088 332508 4140
rect 332560 4128 332566 4140
rect 436738 4128 436744 4140
rect 332560 4100 436744 4128
rect 332560 4088 332566 4100
rect 436738 4088 436744 4100
rect 436796 4088 436802 4140
rect 74994 4020 75000 4072
rect 75052 4060 75058 4072
rect 195974 4060 195980 4072
rect 75052 4032 195980 4060
rect 75052 4020 75058 4032
rect 195974 4020 195980 4032
rect 196032 4020 196038 4072
rect 231026 4020 231032 4072
rect 231084 4060 231090 4072
rect 254118 4060 254124 4072
rect 231084 4032 254124 4060
rect 231084 4020 231090 4032
rect 254118 4020 254124 4032
rect 254176 4020 254182 4072
rect 288250 4020 288256 4072
rect 288308 4060 288314 4072
rect 316218 4060 316224 4072
rect 288308 4032 316224 4060
rect 288308 4020 288314 4032
rect 316218 4020 316224 4032
rect 316276 4020 316282 4072
rect 335262 4020 335268 4072
rect 335320 4060 335326 4072
rect 443822 4060 443828 4072
rect 335320 4032 443828 4060
rect 335320 4020 335326 4032
rect 443822 4020 443828 4032
rect 443880 4020 443886 4072
rect 71498 3952 71504 4004
rect 71556 3992 71562 4004
rect 194594 3992 194600 4004
rect 71556 3964 194600 3992
rect 71556 3952 71562 3964
rect 194594 3952 194600 3964
rect 194652 3952 194658 4004
rect 229830 3952 229836 4004
rect 229888 3992 229894 4004
rect 250441 3995 250499 4001
rect 250441 3992 250453 3995
rect 229888 3964 250453 3992
rect 229888 3952 229894 3964
rect 250441 3961 250453 3964
rect 250487 3961 250499 3995
rect 250441 3955 250499 3961
rect 250533 3995 250591 4001
rect 250533 3961 250545 3995
rect 250579 3992 250591 3995
rect 252646 3992 252652 4004
rect 250579 3964 252652 3992
rect 250579 3961 250591 3964
rect 250533 3955 250591 3961
rect 252646 3952 252652 3964
rect 252704 3952 252710 4004
rect 277210 3952 277216 4004
rect 277268 3992 277274 4004
rect 287790 3992 287796 4004
rect 277268 3964 287796 3992
rect 277268 3952 277274 3964
rect 287790 3952 287796 3964
rect 287848 3952 287854 4004
rect 288342 3952 288348 4004
rect 288400 3992 288406 4004
rect 319714 3992 319720 4004
rect 288400 3964 319720 3992
rect 288400 3952 288406 3964
rect 319714 3952 319720 3964
rect 319772 3952 319778 4004
rect 328362 3952 328368 4004
rect 328420 3992 328426 4004
rect 334069 3995 334127 4001
rect 334069 3992 334081 3995
rect 328420 3964 334081 3992
rect 328420 3952 328426 3964
rect 334069 3961 334081 3964
rect 334115 3961 334127 3995
rect 334069 3955 334127 3961
rect 338022 3952 338028 4004
rect 338080 3992 338086 4004
rect 340785 3995 340843 4001
rect 340785 3992 340797 3995
rect 338080 3964 340797 3992
rect 338080 3952 338086 3964
rect 340785 3961 340797 3964
rect 340831 3961 340843 3995
rect 340785 3955 340843 3961
rect 340874 3952 340880 4004
rect 340932 3992 340938 4004
rect 342162 3992 342168 4004
rect 340932 3964 342168 3992
rect 340932 3952 340938 3964
rect 342162 3952 342168 3964
rect 342220 3952 342226 4004
rect 342257 3995 342315 4001
rect 342257 3961 342269 3995
rect 342303 3992 342315 3995
rect 450906 3992 450912 4004
rect 342303 3964 450912 3992
rect 342303 3961 342315 3964
rect 342257 3955 342315 3961
rect 450906 3952 450912 3964
rect 450964 3952 450970 4004
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 17218 3924 17224 3936
rect 14792 3896 17224 3924
rect 14792 3884 14798 3896
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 67910 3884 67916 3936
rect 67968 3924 67974 3936
rect 193122 3924 193128 3936
rect 67968 3896 193128 3924
rect 67968 3884 67974 3896
rect 193122 3884 193128 3896
rect 193180 3884 193186 3936
rect 228726 3884 228732 3936
rect 228784 3924 228790 3936
rect 231118 3924 231124 3936
rect 228784 3896 231124 3924
rect 228784 3884 228790 3896
rect 231118 3884 231124 3896
rect 231176 3884 231182 3936
rect 233881 3927 233939 3933
rect 233881 3893 233893 3927
rect 233927 3924 233939 3927
rect 252738 3924 252744 3936
rect 233927 3896 252744 3924
rect 233927 3893 233939 3896
rect 233881 3887 233939 3893
rect 252738 3884 252744 3896
rect 252796 3884 252802 3936
rect 281442 3884 281448 3936
rect 281500 3924 281506 3936
rect 300762 3924 300768 3936
rect 281500 3896 300768 3924
rect 281500 3884 281506 3896
rect 300762 3884 300768 3896
rect 300820 3884 300826 3936
rect 304902 3884 304908 3936
rect 304960 3924 304966 3936
rect 357345 3927 357403 3933
rect 357345 3924 357357 3927
rect 304960 3896 357357 3924
rect 304960 3884 304966 3896
rect 357345 3893 357357 3896
rect 357391 3893 357403 3927
rect 357345 3887 357403 3893
rect 357434 3884 357440 3936
rect 357492 3924 357498 3936
rect 358722 3924 358728 3936
rect 357492 3896 358728 3924
rect 357492 3884 357498 3896
rect 358722 3884 358728 3896
rect 358780 3884 358786 3936
rect 358817 3927 358875 3933
rect 358817 3893 358829 3927
rect 358863 3924 358875 3927
rect 362310 3924 362316 3936
rect 358863 3896 362316 3924
rect 358863 3893 358875 3896
rect 358817 3887 358875 3893
rect 362310 3884 362316 3896
rect 362368 3884 362374 3936
rect 382182 3884 382188 3936
rect 382240 3924 382246 3936
rect 568022 3924 568028 3936
rect 382240 3896 568028 3924
rect 382240 3884 382246 3896
rect 568022 3884 568028 3896
rect 568080 3884 568086 3936
rect 45462 3816 45468 3868
rect 45520 3856 45526 3868
rect 47578 3856 47584 3868
rect 45520 3828 47584 3856
rect 45520 3816 45526 3828
rect 47578 3816 47584 3828
rect 47636 3816 47642 3868
rect 64322 3816 64328 3868
rect 64380 3856 64386 3868
rect 182085 3859 182143 3865
rect 182085 3856 182097 3859
rect 64380 3828 182097 3856
rect 64380 3816 64386 3828
rect 182085 3825 182097 3828
rect 182131 3825 182143 3859
rect 190454 3856 190460 3868
rect 182085 3819 182143 3825
rect 182192 3828 190460 3856
rect 60826 3748 60832 3800
rect 60884 3788 60890 3800
rect 182192 3788 182220 3828
rect 190454 3816 190460 3828
rect 190512 3816 190518 3868
rect 227530 3816 227536 3868
rect 227588 3856 227594 3868
rect 250533 3859 250591 3865
rect 250533 3856 250545 3859
rect 227588 3828 250545 3856
rect 227588 3816 227594 3828
rect 250533 3825 250545 3828
rect 250579 3825 250591 3859
rect 259638 3856 259644 3868
rect 250533 3819 250591 3825
rect 252204 3828 259644 3856
rect 191834 3788 191840 3800
rect 60884 3760 182220 3788
rect 190426 3760 191840 3788
rect 60884 3748 60890 3760
rect 57238 3680 57244 3732
rect 57296 3720 57302 3732
rect 181993 3723 182051 3729
rect 181993 3720 182005 3723
rect 57296 3692 182005 3720
rect 57296 3680 57302 3692
rect 181993 3689 182005 3692
rect 182039 3689 182051 3723
rect 181993 3683 182051 3689
rect 182085 3723 182143 3729
rect 182085 3689 182097 3723
rect 182131 3720 182143 3723
rect 190426 3720 190454 3760
rect 191834 3748 191840 3760
rect 191892 3748 191898 3800
rect 223942 3748 223948 3800
rect 224000 3788 224006 3800
rect 251266 3788 251272 3800
rect 224000 3760 251272 3788
rect 224000 3748 224006 3760
rect 251266 3748 251272 3760
rect 251324 3748 251330 3800
rect 182131 3692 190454 3720
rect 182131 3689 182143 3692
rect 182085 3683 182143 3689
rect 226334 3680 226340 3732
rect 226392 3720 226398 3732
rect 233881 3723 233939 3729
rect 233881 3720 233893 3723
rect 226392 3692 233893 3720
rect 226392 3680 226398 3692
rect 233881 3689 233893 3692
rect 233927 3689 233939 3723
rect 233881 3683 233939 3689
rect 233973 3723 234031 3729
rect 233973 3689 233985 3723
rect 234019 3720 234031 3723
rect 251358 3720 251364 3732
rect 234019 3692 251364 3720
rect 234019 3689 234031 3692
rect 233973 3683 234031 3689
rect 251358 3680 251364 3692
rect 251416 3680 251422 3732
rect 53742 3612 53748 3664
rect 53800 3652 53806 3664
rect 187694 3652 187700 3664
rect 53800 3624 187700 3652
rect 53800 3612 53806 3624
rect 187694 3612 187700 3624
rect 187752 3612 187758 3664
rect 219250 3612 219256 3664
rect 219308 3652 219314 3664
rect 239401 3655 239459 3661
rect 239401 3652 239413 3655
rect 219308 3624 239413 3652
rect 219308 3612 219314 3624
rect 239401 3621 239413 3624
rect 239447 3621 239459 3655
rect 239401 3615 239459 3621
rect 247586 3612 247592 3664
rect 247644 3652 247650 3664
rect 248322 3652 248328 3664
rect 247644 3624 248328 3652
rect 247644 3612 247650 3624
rect 248322 3612 248328 3624
rect 248380 3612 248386 3664
rect 250530 3652 250536 3664
rect 248616 3624 250536 3652
rect 25314 3544 25320 3596
rect 25372 3584 25378 3596
rect 32398 3584 32404 3596
rect 25372 3556 32404 3584
rect 25372 3544 25378 3556
rect 32398 3544 32404 3556
rect 32456 3544 32462 3596
rect 34790 3544 34796 3596
rect 34848 3584 34854 3596
rect 39298 3584 39304 3596
rect 34848 3556 39304 3584
rect 34848 3544 34854 3556
rect 39298 3544 39304 3556
rect 39356 3544 39362 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 183554 3584 183560 3596
rect 43128 3556 183560 3584
rect 43128 3544 43134 3556
rect 183554 3544 183560 3556
rect 183612 3544 183618 3596
rect 216858 3544 216864 3596
rect 216916 3584 216922 3596
rect 216916 3556 239444 3584
rect 216916 3544 216922 3556
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14458 3516 14464 3528
rect 13596 3488 14464 3516
rect 13596 3476 13602 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 21358 3516 21364 3528
rect 18288 3488 21364 3516
rect 18288 3476 18294 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24268 3488 26234 3516
rect 24268 3476 24274 3488
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 22738 3448 22744 3460
rect 15988 3420 22744 3448
rect 15988 3408 15994 3420
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 26206 3448 26234 3488
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28902 3516 28908 3528
rect 27764 3488 28908 3516
rect 27764 3476 27770 3488
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 39574 3476 39580 3528
rect 39632 3516 39638 3528
rect 43438 3516 43444 3528
rect 39632 3488 43444 3516
rect 39632 3476 39638 3488
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 43640 3488 171916 3516
rect 35158 3448 35164 3460
rect 26206 3420 35164 3448
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 35986 3340 35992 3392
rect 36044 3380 36050 3392
rect 43640 3380 43668 3488
rect 171781 3451 171839 3457
rect 171781 3448 171793 3451
rect 36044 3352 43668 3380
rect 45526 3420 171793 3448
rect 36044 3340 36050 3352
rect 9950 3272 9956 3324
rect 10008 3312 10014 3324
rect 15838 3312 15844 3324
rect 10008 3284 15844 3312
rect 10008 3272 10014 3284
rect 15838 3272 15844 3284
rect 15896 3272 15902 3324
rect 28902 3272 28908 3324
rect 28960 3312 28966 3324
rect 45526 3312 45554 3420
rect 171781 3417 171793 3420
rect 171827 3417 171839 3451
rect 171888 3448 171916 3488
rect 171962 3476 171968 3528
rect 172020 3516 172026 3528
rect 172422 3516 172428 3528
rect 172020 3488 172428 3516
rect 172020 3476 172026 3488
rect 172422 3476 172428 3488
rect 172480 3476 172486 3528
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 173802 3516 173808 3528
rect 173216 3488 173808 3516
rect 173216 3476 173222 3488
rect 173802 3476 173808 3488
rect 173860 3476 173866 3528
rect 175458 3476 175464 3528
rect 175516 3516 175522 3528
rect 176562 3516 176568 3528
rect 175516 3488 176568 3516
rect 175516 3476 175522 3488
rect 176562 3476 176568 3488
rect 176620 3476 176626 3528
rect 176654 3476 176660 3528
rect 176712 3516 176718 3528
rect 177942 3516 177948 3528
rect 176712 3488 177948 3516
rect 176712 3476 176718 3488
rect 177942 3476 177948 3488
rect 178000 3476 178006 3528
rect 180242 3476 180248 3528
rect 180300 3516 180306 3528
rect 180702 3516 180708 3528
rect 180300 3488 180708 3516
rect 180300 3476 180306 3488
rect 180702 3476 180708 3488
rect 180760 3476 180766 3528
rect 182542 3476 182548 3528
rect 182600 3516 182606 3528
rect 183462 3516 183468 3528
rect 182600 3488 183468 3516
rect 182600 3476 182606 3488
rect 183462 3476 183468 3488
rect 183520 3476 183526 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191742 3516 191748 3528
rect 190880 3488 191748 3516
rect 190880 3476 190886 3488
rect 191742 3476 191748 3488
rect 191800 3476 191806 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 200022 3516 200028 3528
rect 199160 3488 200028 3516
rect 199160 3476 199166 3488
rect 200022 3476 200028 3488
rect 200080 3476 200086 3528
rect 201494 3476 201500 3528
rect 201552 3516 201558 3528
rect 202782 3516 202788 3528
rect 201552 3488 202788 3516
rect 201552 3476 201558 3488
rect 202782 3476 202788 3488
rect 202840 3476 202846 3528
rect 205082 3476 205088 3528
rect 205140 3516 205146 3528
rect 205542 3516 205548 3528
rect 205140 3488 205548 3516
rect 205140 3476 205146 3488
rect 205542 3476 205548 3488
rect 205600 3476 205606 3528
rect 206186 3476 206192 3528
rect 206244 3516 206250 3528
rect 206922 3516 206928 3528
rect 206244 3488 206928 3516
rect 206244 3476 206250 3488
rect 206922 3476 206928 3488
rect 206980 3476 206986 3528
rect 208578 3476 208584 3528
rect 208636 3516 208642 3528
rect 209682 3516 209688 3528
rect 208636 3488 209688 3516
rect 208636 3476 208642 3488
rect 209682 3476 209688 3488
rect 209740 3476 209746 3528
rect 209774 3476 209780 3528
rect 209832 3516 209838 3528
rect 210970 3516 210976 3528
rect 209832 3488 210976 3516
rect 209832 3476 209838 3488
rect 210970 3476 210976 3488
rect 211028 3476 211034 3528
rect 213362 3476 213368 3528
rect 213420 3516 213426 3528
rect 213822 3516 213828 3528
rect 213420 3488 213828 3516
rect 213420 3476 213426 3488
rect 213822 3476 213828 3488
rect 213880 3476 213886 3528
rect 214466 3476 214472 3528
rect 214524 3516 214530 3528
rect 215202 3516 215208 3528
rect 214524 3488 215208 3516
rect 214524 3476 214530 3488
rect 215202 3476 215208 3488
rect 215260 3476 215266 3528
rect 215662 3476 215668 3528
rect 215720 3516 215726 3528
rect 239309 3519 239367 3525
rect 239309 3516 239321 3519
rect 215720 3488 239321 3516
rect 215720 3476 215726 3488
rect 239309 3485 239321 3488
rect 239355 3485 239367 3519
rect 239416 3516 239444 3556
rect 242894 3544 242900 3596
rect 242952 3584 242958 3596
rect 248616 3584 248644 3624
rect 250530 3612 250536 3624
rect 250588 3612 250594 3664
rect 252204 3584 252232 3828
rect 259638 3816 259644 3828
rect 259696 3816 259702 3868
rect 282822 3816 282828 3868
rect 282880 3856 282886 3868
rect 301958 3856 301964 3868
rect 282880 3828 301964 3856
rect 282880 3816 282886 3828
rect 301958 3816 301964 3828
rect 302016 3816 302022 3868
rect 306282 3816 306288 3868
rect 306340 3856 306346 3868
rect 365806 3856 365812 3868
rect 306340 3828 365812 3856
rect 306340 3816 306346 3828
rect 365806 3816 365812 3828
rect 365864 3816 365870 3868
rect 383562 3816 383568 3868
rect 383620 3856 383626 3868
rect 571518 3856 571524 3868
rect 383620 3828 571524 3856
rect 383620 3816 383626 3828
rect 571518 3816 571524 3828
rect 571576 3816 571582 3868
rect 255866 3748 255872 3800
rect 255924 3788 255930 3800
rect 263778 3788 263784 3800
rect 255924 3760 263784 3788
rect 255924 3748 255930 3760
rect 263778 3748 263784 3760
rect 263836 3748 263842 3800
rect 284202 3748 284208 3800
rect 284260 3788 284266 3800
rect 305546 3788 305552 3800
rect 284260 3760 305552 3788
rect 284260 3748 284266 3760
rect 305546 3748 305552 3760
rect 305604 3748 305610 3800
rect 369394 3788 369400 3800
rect 309244 3760 369400 3788
rect 257062 3680 257068 3732
rect 257120 3720 257126 3732
rect 258718 3720 258724 3732
rect 257120 3692 258724 3720
rect 257120 3680 257126 3692
rect 258718 3680 258724 3692
rect 258776 3680 258782 3732
rect 263686 3720 263692 3732
rect 259288 3692 263692 3720
rect 254670 3612 254676 3664
rect 254728 3652 254734 3664
rect 259288 3652 259316 3692
rect 263686 3680 263692 3692
rect 263744 3680 263750 3732
rect 285582 3680 285588 3732
rect 285640 3720 285646 3732
rect 309042 3720 309048 3732
rect 285640 3692 309048 3720
rect 285640 3680 285646 3692
rect 309042 3680 309048 3692
rect 309100 3680 309106 3732
rect 262306 3652 262312 3664
rect 254728 3624 259316 3652
rect 259380 3624 262312 3652
rect 254728 3612 254734 3624
rect 242952 3556 248644 3584
rect 248708 3556 252232 3584
rect 242952 3544 242958 3556
rect 248506 3516 248512 3528
rect 239416 3488 248512 3516
rect 239309 3479 239367 3485
rect 248506 3476 248512 3488
rect 248564 3476 248570 3528
rect 181070 3448 181076 3460
rect 171888 3420 181076 3448
rect 171781 3411 171839 3417
rect 181070 3408 181076 3420
rect 181128 3408 181134 3460
rect 181993 3451 182051 3457
rect 181993 3417 182005 3451
rect 182039 3448 182051 3451
rect 189074 3448 189080 3460
rect 182039 3420 189080 3448
rect 182039 3417 182051 3420
rect 181993 3411 182051 3417
rect 189074 3408 189080 3420
rect 189132 3408 189138 3460
rect 202690 3408 202696 3460
rect 202748 3448 202754 3460
rect 244182 3448 244188 3460
rect 202748 3420 244188 3448
rect 202748 3408 202754 3420
rect 244182 3408 244188 3420
rect 244240 3408 244246 3460
rect 245194 3408 245200 3460
rect 245252 3448 245258 3460
rect 248708 3448 248736 3556
rect 252370 3544 252376 3596
rect 252428 3584 252434 3596
rect 259380 3584 259408 3624
rect 262306 3612 262312 3624
rect 262364 3612 262370 3664
rect 282730 3612 282736 3664
rect 282788 3652 282794 3664
rect 304350 3652 304356 3664
rect 282788 3624 304356 3652
rect 282788 3612 282794 3624
rect 304350 3612 304356 3624
rect 304408 3612 304414 3664
rect 307662 3612 307668 3664
rect 307720 3652 307726 3664
rect 309244 3652 309272 3760
rect 369394 3748 369400 3760
rect 369452 3748 369458 3800
rect 384942 3748 384948 3800
rect 385000 3788 385006 3800
rect 575106 3788 575112 3800
rect 385000 3760 575112 3788
rect 385000 3748 385006 3760
rect 575106 3748 575112 3760
rect 575164 3748 575170 3800
rect 372890 3720 372896 3732
rect 307720 3624 309272 3652
rect 309336 3692 372896 3720
rect 307720 3612 307726 3624
rect 252428 3556 259408 3584
rect 252428 3544 252434 3556
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 260650 3584 260656 3596
rect 259512 3556 260656 3584
rect 259512 3544 259518 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 261754 3544 261760 3596
rect 261812 3584 261818 3596
rect 265618 3584 265624 3596
rect 261812 3556 265624 3584
rect 261812 3544 261818 3556
rect 265618 3544 265624 3556
rect 265676 3544 265682 3596
rect 269114 3544 269120 3596
rect 269172 3584 269178 3596
rect 270034 3584 270040 3596
rect 269172 3556 270040 3584
rect 269172 3544 269178 3556
rect 270034 3544 270040 3556
rect 270092 3544 270098 3596
rect 274358 3544 274364 3596
rect 274416 3584 274422 3596
rect 280706 3584 280712 3596
rect 274416 3556 280712 3584
rect 274416 3544 274422 3556
rect 280706 3544 280712 3556
rect 280764 3544 280770 3596
rect 284110 3544 284116 3596
rect 284168 3584 284174 3596
rect 307938 3584 307944 3596
rect 284168 3556 307944 3584
rect 284168 3544 284174 3556
rect 307938 3544 307944 3556
rect 307996 3544 308002 3596
rect 308950 3544 308956 3596
rect 309008 3584 309014 3596
rect 309336 3584 309364 3692
rect 372890 3680 372896 3692
rect 372948 3680 372954 3732
rect 386322 3680 386328 3732
rect 386380 3720 386386 3732
rect 578602 3720 578608 3732
rect 386380 3692 578608 3720
rect 386380 3680 386386 3692
rect 578602 3680 578608 3692
rect 578660 3680 578666 3732
rect 310422 3612 310428 3664
rect 310480 3652 310486 3664
rect 376478 3652 376484 3664
rect 310480 3624 376484 3652
rect 310480 3612 310486 3624
rect 376478 3612 376484 3624
rect 376536 3612 376542 3664
rect 387610 3612 387616 3664
rect 387668 3652 387674 3664
rect 582190 3652 582196 3664
rect 387668 3624 582196 3652
rect 387668 3612 387674 3624
rect 582190 3612 582196 3624
rect 582248 3612 582254 3664
rect 309008 3556 309364 3584
rect 309008 3544 309014 3556
rect 311802 3544 311808 3596
rect 311860 3584 311866 3596
rect 379974 3584 379980 3596
rect 311860 3556 379980 3584
rect 311860 3544 311866 3556
rect 379974 3544 379980 3556
rect 380032 3544 380038 3596
rect 387518 3544 387524 3596
rect 387576 3584 387582 3596
rect 392029 3587 392087 3593
rect 387576 3556 391980 3584
rect 387576 3544 387582 3556
rect 248782 3476 248788 3528
rect 248840 3516 248846 3528
rect 248840 3488 258074 3516
rect 248840 3476 248846 3488
rect 245252 3420 248736 3448
rect 250349 3451 250407 3457
rect 245252 3408 245258 3420
rect 250349 3417 250361 3451
rect 250395 3448 250407 3451
rect 255498 3448 255504 3460
rect 250395 3420 255504 3448
rect 250395 3417 250407 3420
rect 250349 3411 250407 3417
rect 255498 3408 255504 3420
rect 255556 3408 255562 3460
rect 258046 3448 258074 3488
rect 258258 3476 258264 3528
rect 258316 3516 258322 3528
rect 259362 3516 259368 3528
rect 258316 3488 259368 3516
rect 258316 3476 258322 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 265342 3476 265348 3528
rect 265400 3516 265406 3528
rect 266998 3516 267004 3528
rect 265400 3488 267004 3516
rect 265400 3476 265406 3488
rect 266998 3476 267004 3488
rect 267056 3476 267062 3528
rect 271690 3476 271696 3528
rect 271748 3516 271754 3528
rect 274818 3516 274824 3528
rect 271748 3488 274824 3516
rect 271748 3476 271754 3488
rect 274818 3476 274824 3488
rect 274876 3476 274882 3528
rect 278590 3476 278596 3528
rect 278648 3516 278654 3528
rect 285677 3519 285735 3525
rect 285677 3516 285689 3519
rect 278648 3488 285689 3516
rect 278648 3476 278654 3488
rect 285677 3485 285689 3488
rect 285723 3485 285735 3519
rect 285677 3479 285735 3485
rect 286962 3476 286968 3528
rect 287020 3516 287026 3528
rect 312630 3516 312636 3528
rect 287020 3488 312636 3516
rect 287020 3476 287026 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 313182 3476 313188 3528
rect 313240 3516 313246 3528
rect 383562 3516 383568 3528
rect 313240 3488 383568 3516
rect 313240 3476 313246 3488
rect 383562 3476 383568 3488
rect 383620 3476 383626 3528
rect 386230 3476 386236 3528
rect 386288 3516 386294 3528
rect 390557 3519 390615 3525
rect 390557 3516 390569 3519
rect 386288 3488 390569 3516
rect 386288 3476 386294 3488
rect 390557 3485 390569 3488
rect 390603 3485 390615 3519
rect 390557 3479 390615 3485
rect 390646 3476 390652 3528
rect 390704 3516 390710 3528
rect 391842 3516 391848 3528
rect 390704 3488 391848 3516
rect 390704 3476 390710 3488
rect 391842 3476 391848 3488
rect 391900 3476 391906 3528
rect 391952 3516 391980 3556
rect 392029 3553 392041 3587
rect 392075 3584 392087 3587
rect 579798 3584 579804 3596
rect 392075 3556 579804 3584
rect 392075 3553 392087 3556
rect 392029 3547 392087 3553
rect 579798 3544 579804 3556
rect 579856 3544 579862 3596
rect 580994 3516 581000 3528
rect 391952 3488 581000 3516
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 261018 3448 261024 3460
rect 258046 3420 261024 3448
rect 261018 3408 261024 3420
rect 261076 3408 261082 3460
rect 262950 3408 262956 3460
rect 263008 3448 263014 3460
rect 265710 3448 265716 3460
rect 263008 3420 265716 3448
rect 263008 3408 263014 3420
rect 265710 3408 265716 3420
rect 265768 3408 265774 3460
rect 274450 3408 274456 3460
rect 274508 3448 274514 3460
rect 281902 3448 281908 3460
rect 274508 3420 281908 3448
rect 274508 3408 274514 3420
rect 281902 3408 281908 3420
rect 281960 3408 281966 3460
rect 285490 3408 285496 3460
rect 285548 3448 285554 3460
rect 311434 3448 311440 3460
rect 285548 3420 311440 3448
rect 285548 3408 285554 3420
rect 311434 3408 311440 3420
rect 311492 3408 311498 3460
rect 314562 3408 314568 3460
rect 314620 3448 314626 3460
rect 387150 3448 387156 3460
rect 314620 3420 387156 3448
rect 314620 3408 314626 3420
rect 387150 3408 387156 3420
rect 387208 3408 387214 3460
rect 387702 3408 387708 3460
rect 387760 3448 387766 3460
rect 583386 3448 583392 3460
rect 387760 3420 583392 3448
rect 387760 3408 387766 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 50154 3340 50160 3392
rect 50212 3380 50218 3392
rect 51718 3380 51724 3392
rect 50212 3352 51724 3380
rect 50212 3340 50218 3352
rect 51718 3340 51724 3352
rect 51776 3340 51782 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 82078 3340 82084 3392
rect 82136 3380 82142 3392
rect 198918 3380 198924 3392
rect 82136 3352 198924 3380
rect 82136 3340 82142 3352
rect 198918 3340 198924 3352
rect 198976 3340 198982 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219342 3380 219348 3392
rect 218112 3352 219348 3380
rect 218112 3340 218118 3352
rect 219342 3340 219348 3352
rect 219400 3340 219406 3392
rect 225138 3340 225144 3392
rect 225196 3380 225202 3392
rect 226978 3380 226984 3392
rect 225196 3352 226984 3380
rect 225196 3340 225202 3352
rect 226978 3340 226984 3352
rect 227036 3340 227042 3392
rect 233973 3383 234031 3389
rect 233973 3380 233985 3383
rect 229066 3352 233985 3380
rect 28960 3284 45554 3312
rect 28960 3272 28966 3284
rect 91554 3272 91560 3324
rect 91612 3312 91618 3324
rect 92382 3312 92388 3324
rect 91612 3284 92388 3312
rect 91612 3272 91618 3284
rect 92382 3272 92388 3284
rect 92440 3272 92446 3324
rect 92477 3315 92535 3321
rect 92477 3281 92489 3315
rect 92523 3312 92535 3315
rect 200390 3312 200396 3324
rect 92523 3284 200396 3312
rect 92523 3281 92535 3284
rect 92477 3275 92535 3281
rect 200390 3272 200396 3284
rect 200448 3272 200454 3324
rect 222746 3272 222752 3324
rect 222804 3312 222810 3324
rect 229066 3312 229094 3352
rect 233973 3349 233985 3352
rect 234019 3349 234031 3383
rect 233973 3343 234031 3349
rect 234614 3340 234620 3392
rect 234672 3380 234678 3392
rect 255406 3380 255412 3392
rect 234672 3352 255412 3380
rect 234672 3340 234678 3352
rect 255406 3340 255412 3352
rect 255464 3340 255470 3392
rect 281350 3340 281356 3392
rect 281408 3380 281414 3392
rect 298462 3380 298468 3392
rect 281408 3352 298468 3380
rect 281408 3340 281414 3352
rect 298462 3340 298468 3352
rect 298520 3340 298526 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 429654 3380 429660 3392
rect 333992 3352 429660 3380
rect 222804 3284 229094 3312
rect 222804 3272 222810 3284
rect 238110 3272 238116 3324
rect 238168 3312 238174 3324
rect 248414 3312 248420 3324
rect 238168 3284 248420 3312
rect 238168 3272 238174 3284
rect 248414 3272 248420 3284
rect 248472 3272 248478 3324
rect 248509 3315 248567 3321
rect 248509 3281 248521 3315
rect 248555 3312 248567 3315
rect 253198 3312 253204 3324
rect 248555 3284 253204 3312
rect 248555 3281 248567 3284
rect 248509 3275 248567 3281
rect 253198 3272 253204 3284
rect 253256 3272 253262 3324
rect 282178 3272 282184 3324
rect 282236 3312 282242 3324
rect 285398 3312 285404 3324
rect 282236 3284 285404 3312
rect 282236 3272 282242 3284
rect 285398 3272 285404 3284
rect 285456 3272 285462 3324
rect 294874 3312 294880 3324
rect 285508 3284 294880 3312
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 201678 3244 201684 3256
rect 89220 3216 201684 3244
rect 89220 3204 89226 3216
rect 201678 3204 201684 3216
rect 201736 3204 201742 3256
rect 241698 3204 241704 3256
rect 241756 3244 241762 3256
rect 258166 3244 258172 3256
rect 241756 3216 258172 3244
rect 241756 3204 241762 3216
rect 258166 3204 258172 3216
rect 258224 3204 258230 3256
rect 280062 3204 280068 3256
rect 280120 3244 280126 3256
rect 285508 3244 285536 3284
rect 294874 3272 294880 3284
rect 294932 3272 294938 3324
rect 329742 3272 329748 3324
rect 329800 3312 329806 3324
rect 333992 3312 334020 3352
rect 429654 3340 429660 3352
rect 429712 3340 429718 3392
rect 431954 3340 431960 3392
rect 432012 3380 432018 3392
rect 433242 3380 433248 3392
rect 432012 3352 433248 3380
rect 432012 3340 432018 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474550 3380 474556 3392
rect 473412 3352 474556 3380
rect 473412 3340 473418 3352
rect 474550 3340 474556 3352
rect 474608 3340 474614 3392
rect 481634 3340 481640 3392
rect 481692 3380 481698 3392
rect 482830 3380 482836 3392
rect 481692 3352 482836 3380
rect 481692 3340 481698 3352
rect 482830 3340 482836 3352
rect 482888 3340 482894 3392
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 491110 3380 491116 3392
rect 489972 3352 491116 3380
rect 489972 3340 489978 3352
rect 491110 3340 491116 3352
rect 491168 3340 491174 3392
rect 531314 3340 531320 3392
rect 531372 3380 531378 3392
rect 532510 3380 532516 3392
rect 531372 3352 532516 3380
rect 531372 3340 531378 3352
rect 532510 3340 532516 3352
rect 532568 3340 532574 3392
rect 556154 3340 556160 3392
rect 556212 3380 556218 3392
rect 557350 3380 557356 3392
rect 556212 3352 557356 3380
rect 556212 3340 556218 3352
rect 557350 3340 557356 3352
rect 557408 3340 557414 3392
rect 329800 3284 334020 3312
rect 334069 3315 334127 3321
rect 329800 3272 329806 3284
rect 334069 3281 334081 3315
rect 334115 3312 334127 3315
rect 422570 3312 422576 3324
rect 334115 3284 422576 3312
rect 334115 3281 334127 3284
rect 334069 3275 334127 3281
rect 422570 3272 422576 3284
rect 422628 3272 422634 3324
rect 293678 3244 293684 3256
rect 280120 3216 285536 3244
rect 285600 3216 293684 3244
rect 280120 3204 280126 3216
rect 23014 3136 23020 3188
rect 23072 3176 23078 3188
rect 25498 3176 25504 3188
rect 23072 3148 25504 3176
rect 23072 3136 23078 3148
rect 25498 3136 25504 3148
rect 25556 3136 25562 3188
rect 31294 3136 31300 3188
rect 31352 3176 31358 3188
rect 33778 3176 33784 3188
rect 31352 3148 33784 3176
rect 31352 3136 31358 3148
rect 33778 3136 33784 3148
rect 33836 3136 33842 3188
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 40678 3176 40684 3188
rect 38436 3148 40684 3176
rect 38436 3136 38442 3148
rect 40678 3136 40684 3148
rect 40736 3136 40742 3188
rect 46658 3136 46664 3188
rect 46716 3176 46722 3188
rect 50338 3176 50344 3188
rect 46716 3148 50344 3176
rect 46716 3136 46722 3148
rect 50338 3136 50344 3148
rect 50396 3136 50402 3188
rect 85666 3136 85672 3188
rect 85724 3176 85730 3188
rect 92477 3179 92535 3185
rect 92477 3176 92489 3179
rect 85724 3148 92489 3176
rect 85724 3136 85730 3148
rect 92477 3145 92489 3148
rect 92523 3145 92535 3179
rect 92477 3139 92535 3145
rect 92750 3136 92756 3188
rect 92808 3176 92814 3188
rect 203150 3176 203156 3188
rect 92808 3148 203156 3176
rect 92808 3136 92814 3148
rect 203150 3136 203156 3148
rect 203208 3136 203214 3188
rect 239309 3179 239367 3185
rect 239309 3145 239321 3179
rect 239355 3176 239367 3179
rect 248690 3176 248696 3188
rect 239355 3148 248696 3176
rect 239355 3145 239367 3148
rect 239309 3139 239367 3145
rect 248690 3136 248696 3148
rect 248748 3136 248754 3188
rect 251174 3136 251180 3188
rect 251232 3176 251238 3188
rect 262398 3176 262404 3188
rect 251232 3148 262404 3176
rect 251232 3136 251238 3148
rect 262398 3136 262404 3148
rect 262456 3136 262462 3188
rect 264146 3136 264152 3188
rect 264204 3176 264210 3188
rect 266446 3176 266452 3188
rect 264204 3148 266452 3176
rect 264204 3136 264210 3148
rect 266446 3136 266452 3148
rect 266504 3136 266510 3188
rect 278682 3136 278688 3188
rect 278740 3176 278746 3188
rect 285600 3176 285628 3216
rect 293678 3204 293684 3216
rect 293736 3204 293742 3256
rect 325510 3204 325516 3256
rect 325568 3244 325574 3256
rect 415394 3244 415400 3256
rect 325568 3216 415400 3244
rect 325568 3204 325574 3216
rect 415394 3204 415400 3216
rect 415452 3204 415458 3256
rect 415486 3204 415492 3256
rect 415544 3244 415550 3256
rect 416682 3244 416688 3256
rect 415544 3216 416688 3244
rect 415544 3204 415550 3216
rect 416682 3204 416688 3216
rect 416740 3204 416746 3256
rect 278740 3148 285628 3176
rect 285677 3179 285735 3185
rect 278740 3136 278746 3148
rect 285677 3145 285689 3179
rect 285723 3176 285735 3179
rect 291378 3176 291384 3188
rect 285723 3148 291384 3176
rect 285723 3145 285735 3148
rect 285677 3139 285735 3145
rect 291378 3136 291384 3148
rect 291436 3136 291442 3188
rect 322842 3136 322848 3188
rect 322900 3176 322906 3188
rect 408402 3176 408408 3188
rect 322900 3148 408408 3176
rect 322900 3136 322906 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 98638 3068 98644 3120
rect 98696 3108 98702 3120
rect 99282 3108 99288 3120
rect 98696 3080 99288 3108
rect 98696 3068 98702 3080
rect 99282 3068 99288 3080
rect 99340 3068 99346 3120
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 103238 3108 103244 3120
rect 102284 3080 103244 3108
rect 102284 3068 102290 3080
rect 103238 3068 103244 3080
rect 103296 3068 103302 3120
rect 105722 3068 105728 3120
rect 105780 3108 105786 3120
rect 106182 3108 106188 3120
rect 105780 3080 106188 3108
rect 105780 3068 105786 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 109310 3068 109316 3120
rect 109368 3108 109374 3120
rect 110322 3108 110328 3120
rect 109368 3080 110328 3108
rect 109368 3068 109374 3080
rect 110322 3068 110328 3080
rect 110380 3068 110386 3120
rect 204530 3108 204536 3120
rect 110432 3080 204536 3108
rect 41874 3000 41880 3052
rect 41932 3040 41938 3052
rect 46198 3040 46204 3052
rect 41932 3012 46204 3040
rect 41932 3000 41938 3012
rect 46198 3000 46204 3012
rect 46256 3000 46262 3052
rect 96246 3000 96252 3052
rect 96304 3040 96310 3052
rect 110432 3040 110460 3080
rect 204530 3068 204536 3080
rect 204588 3068 204594 3120
rect 240502 3068 240508 3120
rect 240560 3108 240566 3120
rect 251910 3108 251916 3120
rect 240560 3080 251916 3108
rect 240560 3068 240566 3080
rect 251910 3068 251916 3080
rect 251968 3068 251974 3120
rect 266538 3068 266544 3120
rect 266596 3108 266602 3120
rect 268010 3108 268016 3120
rect 266596 3080 268016 3108
rect 266596 3068 266602 3080
rect 268010 3068 268016 3080
rect 268068 3068 268074 3120
rect 274542 3068 274548 3120
rect 274600 3108 274606 3120
rect 274600 3080 277256 3108
rect 274600 3068 274606 3080
rect 204346 3040 204352 3052
rect 96304 3012 110460 3040
rect 110524 3012 204352 3040
rect 96304 3000 96310 3012
rect 32398 2932 32404 2984
rect 32456 2972 32462 2984
rect 36538 2972 36544 2984
rect 32456 2944 36544 2972
rect 32456 2932 32462 2944
rect 36538 2932 36544 2944
rect 36596 2932 36602 2984
rect 99834 2932 99840 2984
rect 99892 2972 99898 2984
rect 110524 2972 110552 3012
rect 204346 3000 204352 3012
rect 204404 3000 204410 3052
rect 232222 3000 232228 3052
rect 232280 3040 232286 3052
rect 242158 3040 242164 3052
rect 232280 3012 242164 3040
rect 232280 3000 232286 3012
rect 242158 3000 242164 3012
rect 242216 3000 242222 3052
rect 244090 3000 244096 3052
rect 244148 3040 244154 3052
rect 248417 3043 248475 3049
rect 248417 3040 248429 3043
rect 244148 3012 248429 3040
rect 244148 3000 244154 3012
rect 248417 3009 248429 3012
rect 248463 3009 248475 3043
rect 248417 3003 248475 3009
rect 248509 3043 248567 3049
rect 248509 3009 248521 3043
rect 248555 3040 248567 3043
rect 251818 3040 251824 3052
rect 248555 3012 251824 3040
rect 248555 3009 248567 3012
rect 248509 3003 248567 3009
rect 251818 3000 251824 3012
rect 251876 3000 251882 3052
rect 275278 3000 275284 3052
rect 275336 3040 275342 3052
rect 277118 3040 277124 3052
rect 275336 3012 277124 3040
rect 275336 3000 275342 3012
rect 277118 3000 277124 3012
rect 277176 3000 277182 3052
rect 277228 3040 277256 3080
rect 277302 3068 277308 3120
rect 277360 3108 277366 3120
rect 290182 3108 290188 3120
rect 277360 3080 290188 3108
rect 277360 3068 277366 3080
rect 290182 3068 290188 3080
rect 290240 3068 290246 3120
rect 321462 3068 321468 3120
rect 321520 3108 321526 3120
rect 404814 3108 404820 3120
rect 321520 3080 404820 3108
rect 321520 3068 321526 3080
rect 404814 3068 404820 3080
rect 404872 3068 404878 3120
rect 279510 3040 279516 3052
rect 277228 3012 279516 3040
rect 279510 3000 279516 3012
rect 279568 3000 279574 3052
rect 320082 3000 320088 3052
rect 320140 3040 320146 3052
rect 320140 3012 398788 3040
rect 320140 3000 320146 3012
rect 207290 2972 207296 2984
rect 99892 2944 110552 2972
rect 113146 2944 207296 2972
rect 99892 2932 99898 2944
rect 110506 2864 110512 2916
rect 110564 2904 110570 2916
rect 111702 2904 111708 2916
rect 110564 2876 111708 2904
rect 110564 2864 110570 2876
rect 111702 2864 111708 2876
rect 111760 2864 111766 2916
rect 106918 2796 106924 2848
rect 106976 2836 106982 2848
rect 113146 2836 113174 2944
rect 207290 2932 207296 2944
rect 207348 2932 207354 2984
rect 239401 2975 239459 2981
rect 239401 2941 239413 2975
rect 239447 2972 239459 2975
rect 249886 2972 249892 2984
rect 239447 2944 249892 2972
rect 239447 2941 239459 2944
rect 239401 2935 239459 2941
rect 249886 2932 249892 2944
rect 249944 2932 249950 2984
rect 271782 2932 271788 2984
rect 271840 2972 271846 2984
rect 273622 2972 273628 2984
rect 271840 2944 273628 2972
rect 271840 2932 271846 2944
rect 273622 2932 273628 2944
rect 273680 2932 273686 2984
rect 318610 2932 318616 2984
rect 318668 2972 318674 2984
rect 397730 2972 397736 2984
rect 318668 2944 397736 2972
rect 318668 2932 318674 2944
rect 397730 2932 397736 2944
rect 397788 2932 397794 2984
rect 398760 2972 398788 3012
rect 398834 3000 398840 3052
rect 398892 3040 398898 3052
rect 400122 3040 400128 3052
rect 398892 3012 400128 3040
rect 398892 3000 398898 3012
rect 400122 3000 400128 3012
rect 400180 3000 400186 3052
rect 401318 2972 401324 2984
rect 398760 2944 401324 2972
rect 401318 2932 401324 2944
rect 401376 2932 401382 2984
rect 116394 2864 116400 2916
rect 116452 2904 116458 2916
rect 117222 2904 117228 2916
rect 116452 2876 117228 2904
rect 116452 2864 116458 2876
rect 117222 2864 117228 2876
rect 117280 2864 117286 2916
rect 117590 2864 117596 2916
rect 117648 2904 117654 2916
rect 118602 2904 118608 2916
rect 117648 2876 118608 2904
rect 117648 2864 117654 2876
rect 118602 2864 118608 2876
rect 118660 2864 118666 2916
rect 123478 2864 123484 2916
rect 123536 2904 123542 2916
rect 124122 2904 124128 2916
rect 123536 2876 124128 2904
rect 123536 2864 123542 2876
rect 124122 2864 124128 2876
rect 124180 2864 124186 2916
rect 124674 2864 124680 2916
rect 124732 2904 124738 2916
rect 125781 2907 125839 2913
rect 125781 2904 125793 2907
rect 124732 2876 125793 2904
rect 124732 2864 124738 2876
rect 125781 2873 125793 2876
rect 125827 2873 125839 2907
rect 125781 2867 125839 2873
rect 125962 2864 125968 2916
rect 126020 2904 126026 2916
rect 126882 2904 126888 2916
rect 126020 2876 126888 2904
rect 126020 2864 126026 2876
rect 126882 2864 126888 2876
rect 126940 2864 126946 2916
rect 130473 2907 130531 2913
rect 130473 2904 130485 2907
rect 126992 2876 130485 2904
rect 106976 2808 113174 2836
rect 106976 2796 106982 2808
rect 114002 2796 114008 2848
rect 114060 2836 114066 2848
rect 125873 2839 125931 2845
rect 114060 2808 125732 2836
rect 114060 2796 114066 2808
rect 125704 2768 125732 2808
rect 125873 2805 125885 2839
rect 125919 2836 125931 2839
rect 126992 2836 127020 2876
rect 130473 2873 130485 2876
rect 130519 2873 130531 2907
rect 130473 2867 130531 2873
rect 130562 2864 130568 2916
rect 130620 2904 130626 2916
rect 131022 2904 131028 2916
rect 130620 2876 131028 2904
rect 130620 2864 130626 2876
rect 131022 2864 131028 2876
rect 131080 2864 131086 2916
rect 131758 2864 131764 2916
rect 131816 2904 131822 2916
rect 132218 2904 132224 2916
rect 131816 2876 132224 2904
rect 131816 2864 131822 2876
rect 132218 2864 132224 2876
rect 132276 2864 132282 2916
rect 132405 2907 132463 2913
rect 132405 2873 132417 2907
rect 132451 2904 132463 2907
rect 210050 2904 210056 2916
rect 132451 2876 210056 2904
rect 132451 2873 132463 2876
rect 132405 2867 132463 2873
rect 210050 2864 210056 2876
rect 210108 2864 210114 2916
rect 237006 2864 237012 2916
rect 237064 2904 237070 2916
rect 237064 2876 249472 2904
rect 237064 2864 237070 2876
rect 132313 2839 132371 2845
rect 132313 2836 132325 2839
rect 125919 2808 127020 2836
rect 127084 2808 130332 2836
rect 125919 2805 125931 2808
rect 125873 2799 125931 2805
rect 127084 2768 127112 2808
rect 125704 2740 127112 2768
rect 130304 2700 130332 2808
rect 130580 2808 132325 2836
rect 130580 2700 130608 2808
rect 132313 2805 132325 2808
rect 132359 2805 132371 2839
rect 214190 2836 214196 2848
rect 132313 2799 132371 2805
rect 132466 2808 214196 2836
rect 130657 2771 130715 2777
rect 130657 2737 130669 2771
rect 130703 2768 130715 2771
rect 132466 2768 132494 2808
rect 214190 2796 214196 2808
rect 214248 2796 214254 2848
rect 239306 2796 239312 2848
rect 239364 2836 239370 2848
rect 239364 2808 246344 2836
rect 239364 2796 239370 2808
rect 130703 2740 132494 2768
rect 246316 2768 246344 2808
rect 246390 2796 246396 2848
rect 246448 2836 246454 2848
rect 248417 2839 248475 2845
rect 248417 2836 248429 2839
rect 246448 2808 248429 2836
rect 246448 2796 246454 2808
rect 248417 2805 248429 2808
rect 248463 2805 248475 2839
rect 249058 2836 249064 2848
rect 248417 2799 248475 2805
rect 248524 2808 249064 2836
rect 248524 2768 248552 2808
rect 249058 2796 249064 2808
rect 249116 2796 249122 2848
rect 249444 2836 249472 2876
rect 249978 2864 249984 2916
rect 250036 2904 250042 2916
rect 253290 2904 253296 2916
rect 250036 2876 253296 2904
rect 250036 2864 250042 2876
rect 253290 2864 253296 2876
rect 253348 2864 253354 2916
rect 317230 2864 317236 2916
rect 317288 2904 317294 2916
rect 394234 2904 394240 2916
rect 317288 2876 394240 2904
rect 317288 2864 317294 2876
rect 394234 2864 394240 2876
rect 394292 2864 394298 2916
rect 250438 2836 250444 2848
rect 249444 2808 250444 2836
rect 250438 2796 250444 2808
rect 250496 2796 250502 2848
rect 256878 2836 256884 2848
rect 250548 2808 256884 2836
rect 246316 2740 248552 2768
rect 130703 2737 130715 2740
rect 130657 2731 130715 2737
rect 248598 2728 248604 2780
rect 248656 2768 248662 2780
rect 250548 2768 250576 2808
rect 256878 2796 256884 2808
rect 256936 2796 256942 2848
rect 315942 2796 315948 2848
rect 316000 2836 316006 2848
rect 390646 2836 390652 2848
rect 316000 2808 390652 2836
rect 316000 2796 316006 2808
rect 390646 2796 390652 2808
rect 390704 2796 390710 2848
rect 390741 2839 390799 2845
rect 390741 2805 390753 2839
rect 390787 2836 390799 2839
rect 392029 2839 392087 2845
rect 392029 2836 392041 2839
rect 390787 2808 392041 2836
rect 390787 2805 390799 2808
rect 390741 2799 390799 2805
rect 392029 2805 392041 2808
rect 392075 2805 392087 2839
rect 392029 2799 392087 2805
rect 248656 2740 250576 2768
rect 248656 2728 248662 2740
rect 130304 2672 130608 2700
<< via1 >>
rect 324228 700952 324280 701004
rect 413652 700952 413704 701004
rect 331128 700884 331180 700936
rect 429844 700884 429896 700936
rect 336648 700816 336700 700868
rect 446128 700816 446180 700868
rect 342168 700748 342220 700800
rect 462320 700748 462372 700800
rect 349068 700680 349120 700732
rect 478512 700680 478564 700732
rect 354588 700612 354640 700664
rect 494796 700612 494848 700664
rect 288348 700544 288400 700596
rect 316316 700544 316368 700596
rect 361488 700544 361540 700596
rect 510988 700544 511040 700596
rect 293868 700476 293920 700528
rect 332508 700476 332560 700528
rect 367008 700476 367060 700528
rect 527180 700476 527232 700528
rect 299388 700408 299440 700460
rect 348792 700408 348844 700460
rect 373908 700408 373960 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 105452 700340 105504 700392
rect 106188 700340 106240 700392
rect 235172 700340 235224 700392
rect 235908 700340 235960 700392
rect 276664 700340 276716 700392
rect 283840 700340 283892 700392
rect 306288 700340 306340 700392
rect 364984 700340 365036 700392
rect 379428 700340 379480 700392
rect 559656 700340 559708 700392
rect 281448 700272 281500 700324
rect 300124 700272 300176 700324
rect 311808 700272 311860 700324
rect 381176 700272 381228 700324
rect 384948 700272 385000 700324
rect 575848 700272 575900 700324
rect 170312 700204 170364 700256
rect 171048 700204 171100 700256
rect 318708 700204 318760 700256
rect 397460 700204 397512 700256
rect 56784 700136 56836 700188
rect 57888 700136 57940 700188
rect 186504 700136 186556 700188
rect 187608 700136 187660 700188
rect 251456 700068 251508 700120
rect 252468 700068 252520 700120
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 121644 699660 121696 699712
rect 122748 699660 122800 699712
rect 3424 696940 3476 696992
rect 86224 696940 86276 696992
rect 389824 696940 389876 696992
rect 580172 696940 580224 696992
rect 389916 683136 389968 683188
rect 580172 683136 580224 683188
rect 390008 670692 390060 670744
rect 580172 670692 580224 670744
rect 2780 645056 2832 645108
rect 4804 645056 4856 645108
rect 390100 643084 390152 643136
rect 580172 643084 580224 643136
rect 390192 630640 390244 630692
rect 579988 630640 580040 630692
rect 390284 616836 390336 616888
rect 580172 616836 580224 616888
rect 390376 590656 390428 590708
rect 579620 590656 579672 590708
rect 390468 576852 390520 576904
rect 579620 576852 579672 576904
rect 389732 536800 389784 536852
rect 579620 536800 579672 536852
rect 389640 524424 389692 524476
rect 580172 524424 580224 524476
rect 389548 484372 389600 484424
rect 580172 484372 580224 484424
rect 274916 481584 274968 481636
rect 276664 481584 276716 481636
rect 305460 481584 305512 481636
rect 306288 481584 306340 481636
rect 329840 481584 329892 481636
rect 331128 481584 331180 481636
rect 154488 481516 154540 481568
rect 225972 481516 226024 481568
rect 137928 481448 137980 481500
rect 219900 481448 219952 481500
rect 122748 481380 122800 481432
rect 213736 481380 213788 481432
rect 106188 481312 106240 481364
rect 207664 481312 207716 481364
rect 287060 481312 287112 481364
rect 288348 481312 288400 481364
rect 89628 481244 89680 481296
rect 201592 481244 201644 481296
rect 73068 481176 73120 481228
rect 195428 481176 195480 481228
rect 317696 481176 317748 481228
rect 318708 481176 318760 481228
rect 57888 481108 57940 481160
rect 189356 481108 189408 481160
rect 219348 481108 219400 481160
rect 250444 481108 250496 481160
rect 360384 481108 360436 481160
rect 361488 481108 361540 481160
rect 41328 481040 41380 481092
rect 183192 481040 183244 481092
rect 202788 481040 202840 481092
rect 244372 481040 244424 481092
rect 348240 481040 348292 481092
rect 349068 481040 349120 481092
rect 24768 480972 24820 481024
rect 177120 480972 177172 481024
rect 187608 480972 187660 481024
rect 238208 480972 238260 481024
rect 252468 480972 252520 481024
rect 262680 480972 262732 481024
rect 8208 480904 8260 480956
rect 171048 480904 171100 480956
rect 170956 480836 171008 480888
rect 232136 480904 232188 480956
rect 235908 480904 235960 480956
rect 256516 480904 256568 480956
rect 372620 480768 372672 480820
rect 373908 480768 373960 480820
rect 267648 480224 267700 480276
rect 268752 480224 268804 480276
rect 86224 477436 86276 477488
rect 165620 477436 165672 477488
rect 3424 471928 3476 471980
rect 165620 471928 165672 471980
rect 389824 470568 389876 470620
rect 579988 470568 580040 470620
rect 3516 469140 3568 469192
rect 165620 469140 165672 469192
rect 390100 469140 390152 469192
rect 580264 469140 580316 469192
rect 4804 466352 4856 466404
rect 165620 466352 165672 466404
rect 3608 463632 3660 463684
rect 165620 463632 165672 463684
rect 3700 462272 3752 462324
rect 165620 462272 165672 462324
rect 3792 459484 3844 459536
rect 165620 459484 165672 459536
rect 390192 458124 390244 458176
rect 580356 458124 580408 458176
rect 389916 456764 389968 456816
rect 579804 456764 579856 456816
rect 3884 456696 3936 456748
rect 165620 456696 165672 456748
rect 3976 453976 4028 454028
rect 165620 453976 165672 454028
rect 4068 451188 4120 451240
rect 165620 451188 165672 451240
rect 390192 451188 390244 451240
rect 580448 451188 580500 451240
rect 3332 448468 3384 448520
rect 165620 448468 165672 448520
rect 390192 448468 390244 448520
rect 580540 448468 580592 448520
rect 3240 445680 3292 445732
rect 165620 445680 165672 445732
rect 390008 444388 390060 444440
rect 580172 444388 580224 444440
rect 3148 442892 3200 442944
rect 165620 442892 165672 442944
rect 3056 441532 3108 441584
rect 165620 441532 165672 441584
rect 390192 440172 390244 440224
rect 580632 440172 580684 440224
rect 2964 438812 3016 438864
rect 165620 438812 165672 438864
rect 390284 437384 390336 437436
rect 580724 437384 580776 437436
rect 2872 436024 2924 436076
rect 165620 436024 165672 436076
rect 2780 433236 2832 433288
rect 165620 433236 165672 433288
rect 389824 430584 389876 430636
rect 580172 430584 580224 430636
rect 3424 430516 3476 430568
rect 165620 430516 165672 430568
rect 3516 427728 3568 427780
rect 165620 427728 165672 427780
rect 3608 425008 3660 425060
rect 165620 425008 165672 425060
rect 3792 422220 3844 422272
rect 165620 422220 165672 422272
rect 390100 419432 390152 419484
rect 580172 419432 580224 419484
rect 3424 418140 3476 418192
rect 165620 418140 165672 418192
rect 3792 416780 3844 416832
rect 165620 416780 165672 416832
rect 3700 413992 3752 414044
rect 165620 413992 165672 414044
rect 3608 411272 3660 411324
rect 165620 411272 165672 411324
rect 3516 408484 3568 408536
rect 165620 408484 165672 408536
rect 3424 405696 3476 405748
rect 165620 405696 165672 405748
rect 390192 405628 390244 405680
rect 580172 405628 580224 405680
rect 389180 404472 389232 404524
rect 391204 404472 391256 404524
rect 3148 398828 3200 398880
rect 165620 398828 165672 398880
rect 4804 396040 4856 396092
rect 165620 396040 165672 396092
rect 390192 393320 390244 393372
rect 396816 393320 396868 393372
rect 390192 391960 390244 392012
rect 393964 391960 394016 392012
rect 390100 391892 390152 391944
rect 580172 391892 580224 391944
rect 390192 389172 390244 389224
rect 406384 389172 406436 389224
rect 21456 387812 21508 387864
rect 165620 387812 165672 387864
rect 3240 385024 3292 385076
rect 165620 385024 165672 385076
rect 390008 379448 390060 379500
rect 580172 379448 580224 379500
rect 3332 376728 3384 376780
rect 165620 376728 165672 376780
rect 10324 375368 10376 375420
rect 165620 375368 165672 375420
rect 390100 372580 390152 372632
rect 403624 372580 403676 372632
rect 4068 369860 4120 369912
rect 165620 369860 165672 369912
rect 28264 367072 28316 367124
rect 165620 367072 165672 367124
rect 389916 365644 389968 365696
rect 580172 365644 580224 365696
rect 3976 364352 4028 364404
rect 165620 364352 165672 364404
rect 3884 358776 3936 358828
rect 165620 358776 165672 358828
rect 390100 357416 390152 357468
rect 400864 357416 400916 357468
rect 389916 357280 389968 357332
rect 390100 357280 390152 357332
rect 3792 356056 3844 356108
rect 165620 356056 165672 356108
rect 11704 354696 11756 354748
rect 165620 354696 165672 354748
rect 389916 354696 389968 354748
rect 547144 354696 547196 354748
rect 389824 353200 389876 353252
rect 580172 353200 580224 353252
rect 3700 351908 3752 351960
rect 165620 351908 165672 351960
rect 29644 349120 29696 349172
rect 165620 349120 165672 349172
rect 389916 347259 389968 347268
rect 389916 347225 389925 347259
rect 389925 347225 389959 347259
rect 389959 347225 389968 347259
rect 389916 347216 389968 347225
rect 3608 346400 3660 346452
rect 165620 346400 165672 346452
rect 389916 346400 389968 346452
rect 543004 346400 543056 346452
rect 389916 346307 389968 346316
rect 389916 346273 389925 346307
rect 389925 346273 389959 346307
rect 389959 346273 389968 346307
rect 389916 346264 389968 346273
rect 3516 343612 3568 343664
rect 165620 343612 165672 343664
rect 396816 341504 396868 341556
rect 580264 341504 580316 341556
rect 3424 340892 3476 340944
rect 165620 340892 165672 340944
rect 389088 340892 389140 340944
rect 396724 340892 396776 340944
rect 391204 340144 391256 340196
rect 580172 340144 580224 340196
rect 18604 338104 18656 338156
rect 165620 338104 165672 338156
rect 389088 338104 389140 338156
rect 519544 338104 519596 338156
rect 168380 336744 168432 336796
rect 168748 336744 168800 336796
rect 189080 336744 189132 336796
rect 189356 336744 189408 336796
rect 240140 336744 240192 336796
rect 240416 336744 240468 336796
rect 118608 336676 118660 336728
rect 212264 336676 212316 336728
rect 220820 336676 220872 336728
rect 221188 336676 221240 336728
rect 233884 336676 233936 336728
rect 237196 336676 237248 336728
rect 239404 336676 239456 336728
rect 241612 336676 241664 336728
rect 242072 336676 242124 336728
rect 255412 336676 255464 336728
rect 260656 336676 260708 336728
rect 265624 336676 265676 336728
rect 271052 336676 271104 336728
rect 271788 336676 271840 336728
rect 272248 336676 272300 336728
rect 276204 336676 276256 336728
rect 276388 336676 276440 336728
rect 277216 336676 277268 336728
rect 279056 336676 279108 336728
rect 280068 336676 280120 336728
rect 280344 336676 280396 336728
rect 281356 336676 281408 336728
rect 281724 336676 281776 336728
rect 282828 336676 282880 336728
rect 286140 336676 286192 336728
rect 286876 336676 286928 336728
rect 289728 336676 289780 336728
rect 290464 336676 290516 336728
rect 291476 336676 291528 336728
rect 292488 336676 292540 336728
rect 292856 336676 292908 336728
rect 293776 336676 293828 336728
rect 294604 336676 294656 336728
rect 295248 336676 295300 336728
rect 295984 336676 296036 336728
rect 296628 336676 296680 336728
rect 298652 336676 298704 336728
rect 299388 336676 299440 336728
rect 299940 336676 299992 336728
rect 300768 336676 300820 336728
rect 300860 336676 300912 336728
rect 301964 336676 302016 336728
rect 303988 336676 304040 336728
rect 304724 336676 304776 336728
rect 305276 336676 305328 336728
rect 306104 336676 306156 336728
rect 306656 336676 306708 336728
rect 307484 336676 307536 336728
rect 307944 336676 307996 336728
rect 308864 336676 308916 336728
rect 309324 336676 309376 336728
rect 310244 336676 310296 336728
rect 310612 336676 310664 336728
rect 311624 336676 311676 336728
rect 312452 336676 312504 336728
rect 313188 336676 313240 336728
rect 313280 336676 313332 336728
rect 314476 336676 314528 336728
rect 314660 336676 314712 336728
rect 315856 336676 315908 336728
rect 316408 336676 316460 336728
rect 317328 336676 317380 336728
rect 319076 336676 319128 336728
rect 320088 336676 320140 336728
rect 320456 336676 320508 336728
rect 321468 336676 321520 336728
rect 324412 336676 324464 336728
rect 325608 336676 325660 336728
rect 327540 336676 327592 336728
rect 328276 336676 328328 336728
rect 328920 336676 328972 336728
rect 329656 336676 329708 336728
rect 330208 336676 330260 336728
rect 331128 336676 331180 336728
rect 331588 336676 331640 336728
rect 332416 336676 332468 336728
rect 332876 336676 332928 336728
rect 333888 336676 333940 336728
rect 334256 336676 334308 336728
rect 335176 336676 335228 336728
rect 335544 336676 335596 336728
rect 336648 336676 336700 336728
rect 336924 336676 336976 336728
rect 337936 336676 337988 336728
rect 338212 336676 338264 336728
rect 339408 336676 339460 336728
rect 339592 336676 339644 336728
rect 340696 336676 340748 336728
rect 340880 336676 340932 336728
rect 342168 336676 342220 336728
rect 343180 336676 343232 336728
rect 343548 336676 343600 336728
rect 345388 336676 345440 336728
rect 346124 336676 346176 336728
rect 348056 336676 348108 336728
rect 348884 336676 348936 336728
rect 350724 336676 350776 336728
rect 351828 336676 351880 336728
rect 352012 336676 352064 336728
rect 353116 336676 353168 336728
rect 355140 336676 355192 336728
rect 355876 336676 355928 336728
rect 356060 336676 356112 336728
rect 357348 336676 357400 336728
rect 357808 336676 357860 336728
rect 358636 336676 358688 336728
rect 359188 336676 359240 336728
rect 360016 336676 360068 336728
rect 360476 336676 360528 336728
rect 361396 336676 361448 336728
rect 361856 336676 361908 336728
rect 362684 336676 362736 336728
rect 363144 336676 363196 336728
rect 364064 336676 364116 336728
rect 364524 336676 364576 336728
rect 365444 336676 365496 336728
rect 365812 336676 365864 336728
rect 366824 336676 366876 336728
rect 367192 336676 367244 336728
rect 368204 336676 368256 336728
rect 368940 336676 368992 336728
rect 369768 336676 369820 336728
rect 369860 336676 369912 336728
rect 370964 336676 371016 336728
rect 372068 336676 372120 336728
rect 372436 336676 372488 336728
rect 373448 336676 373500 336728
rect 373816 336676 373868 336728
rect 374736 336676 374788 336728
rect 375196 336676 375248 336728
rect 375656 336676 375708 336728
rect 376668 336676 376720 336728
rect 376944 336676 376996 336728
rect 378048 336676 378100 336728
rect 378784 336676 378836 336728
rect 379336 336676 379388 336728
rect 380072 336676 380124 336728
rect 380716 336676 380768 336728
rect 380992 336676 381044 336728
rect 382096 336676 382148 336728
rect 383660 336676 383712 336728
rect 384856 336676 384908 336728
rect 385868 336676 385920 336728
rect 386328 336676 386380 336728
rect 386788 336676 386840 336728
rect 387524 336676 387576 336728
rect 111708 336608 111760 336660
rect 209596 336608 209648 336660
rect 231860 336608 231912 336660
rect 235908 336608 235960 336660
rect 256792 336608 256844 336660
rect 258724 336608 258776 336660
rect 264796 336608 264848 336660
rect 270592 336608 270644 336660
rect 271880 336608 271932 336660
rect 277676 336608 277728 336660
rect 278596 336608 278648 336660
rect 299480 336608 299532 336660
rect 300676 336608 300728 336660
rect 301320 336608 301372 336660
rect 302148 336608 302200 336660
rect 304448 336608 304500 336660
rect 304908 336608 304960 336660
rect 305736 336608 305788 336660
rect 306288 336608 306340 336660
rect 307116 336608 307168 336660
rect 307668 336608 307720 336660
rect 308404 336608 308456 336660
rect 309048 336608 309100 336660
rect 309784 336608 309836 336660
rect 310428 336608 310480 336660
rect 311072 336608 311124 336660
rect 311808 336608 311860 336660
rect 315120 336608 315172 336660
rect 315948 336608 316000 336660
rect 323124 336608 323176 336660
rect 411260 336608 411312 336660
rect 103428 336540 103480 336592
rect 50344 336472 50396 336524
rect 185492 336472 185544 336524
rect 202144 336540 202196 336592
rect 205088 336540 205140 336592
rect 222844 336540 222896 336592
rect 231124 336540 231176 336592
rect 254124 336540 254176 336592
rect 296812 336540 296864 336592
rect 297916 336540 297968 336592
rect 313740 336540 313792 336592
rect 314568 336540 314620 336592
rect 328460 336540 328512 336592
rect 418160 336540 418212 336592
rect 206928 336472 206980 336524
rect 226984 336472 227036 336524
rect 252744 336472 252796 336524
rect 331220 336472 331272 336524
rect 43444 336404 43496 336456
rect 182824 336404 182876 336456
rect 220728 336404 220780 336456
rect 250996 336404 251048 336456
rect 298100 336404 298152 336456
rect 318064 336404 318116 336456
rect 325792 336404 325844 336456
rect 342260 336472 342312 336524
rect 343456 336472 343508 336524
rect 425060 336472 425112 336524
rect 431960 336404 432012 336456
rect 35164 336336 35216 336388
rect 177028 336336 177080 336388
rect 213828 336336 213880 336388
rect 248328 336336 248380 336388
rect 253296 336336 253348 336388
rect 262128 336336 262180 336388
rect 287060 336336 287112 336388
rect 288256 336336 288308 336388
rect 290648 336336 290700 336388
rect 316684 336336 316736 336388
rect 333796 336336 333848 336388
rect 440240 336336 440292 336388
rect 36544 336268 36596 336320
rect 180156 336268 180208 336320
rect 219348 336268 219400 336320
rect 250076 336268 250128 336320
rect 251824 336268 251876 336320
rect 260748 336268 260800 336320
rect 278136 336268 278188 336320
rect 291844 336268 291896 336320
rect 293316 336268 293368 336320
rect 320824 336268 320876 336320
rect 447140 336268 447192 336320
rect 32404 336200 32456 336252
rect 177120 336200 177172 336252
rect 183560 336200 183612 336252
rect 183836 336200 183888 336252
rect 212448 336200 212500 336252
rect 247500 336200 247552 336252
rect 247684 336200 247736 336252
rect 251456 336200 251508 336252
rect 253848 336200 253900 336252
rect 263416 336200 263468 336252
rect 275468 336200 275520 336252
rect 282184 336200 282236 336252
rect 286600 336200 286652 336252
rect 313924 336200 313976 336252
rect 315580 336200 315632 336252
rect 336004 336200 336056 336252
rect 341340 336200 341392 336252
rect 342076 336200 342128 336252
rect 22744 336132 22796 336184
rect 173900 336132 173952 336184
rect 210976 336132 211028 336184
rect 246948 336132 247000 336184
rect 250536 336132 250588 336184
rect 259460 336132 259512 336184
rect 260748 336132 260800 336184
rect 266084 336132 266136 336184
rect 274548 336132 274600 336184
rect 283196 336132 283248 336184
rect 287888 336132 287940 336184
rect 317696 336132 317748 336184
rect 17224 336064 17276 336116
rect 173532 336064 173584 336116
rect 177304 336064 177356 336116
rect 202420 336064 202472 336116
rect 209688 336064 209740 336116
rect 246488 336064 246540 336116
rect 249064 336064 249116 336116
rect 258080 336064 258132 336116
rect 275008 336064 275060 336116
rect 284484 336064 284536 336116
rect 290188 336064 290240 336116
rect 323584 336132 323636 336184
rect 321744 336064 321796 336116
rect 322848 336064 322900 336116
rect 339132 336064 339184 336116
rect 454040 336200 454092 336252
rect 7564 335996 7616 336048
rect 170404 335996 170456 336048
rect 173164 335996 173216 336048
rect 199752 335996 199804 336048
rect 206928 335996 206980 336048
rect 245660 335996 245712 336048
rect 248328 335996 248380 336048
rect 261208 335996 261260 336048
rect 275928 335996 275980 336048
rect 121368 335928 121420 335980
rect 213552 335928 213604 335980
rect 229744 335928 229796 335980
rect 231400 335928 231452 335980
rect 250444 335928 250496 335980
rect 257252 335928 257304 335980
rect 265716 335928 265768 335980
rect 266636 335928 266688 335980
rect 285680 335996 285732 336048
rect 286968 335996 287020 336048
rect 291936 335996 291988 336048
rect 328552 335996 328604 336048
rect 336464 335996 336516 336048
rect 285772 335928 285824 335980
rect 294144 335928 294196 335980
rect 295064 335928 295116 335980
rect 341800 335928 341852 335980
rect 460940 336132 460992 336184
rect 344468 336064 344520 336116
rect 467840 336064 467892 336116
rect 345848 335996 345900 336048
rect 346308 335996 346360 336048
rect 348516 335996 348568 336048
rect 349068 335996 349120 336048
rect 353392 335996 353444 336048
rect 354496 335996 354548 336048
rect 347136 335928 347188 335980
rect 474740 335996 474792 336048
rect 360936 335928 360988 335980
rect 361488 335928 361540 335980
rect 363604 335928 363656 335980
rect 364248 335928 364300 335980
rect 364984 335928 365036 335980
rect 365628 335928 365680 335980
rect 366272 335928 366324 335980
rect 367008 335928 367060 335980
rect 367652 335928 367704 335980
rect 368388 335928 368440 335980
rect 368572 335928 368624 335980
rect 369584 335928 369636 335980
rect 370320 335928 370372 335980
rect 371148 335928 371200 335980
rect 378324 335928 378376 335980
rect 379428 335928 379480 335980
rect 379704 335928 379756 335980
rect 380808 335928 380860 335980
rect 385040 335928 385092 335980
rect 386144 335928 386196 335980
rect 288808 335860 288860 335912
rect 289728 335860 289780 335912
rect 311992 335860 312044 335912
rect 313004 335860 313056 335912
rect 344008 335860 344060 335912
rect 344836 335860 344888 335912
rect 354680 335860 354732 335912
rect 355784 335860 355836 335912
rect 358268 335860 358320 335912
rect 358728 335860 358780 335912
rect 382372 335860 382424 335912
rect 383476 335860 383528 335912
rect 265624 335792 265676 335844
rect 266544 335792 266596 335844
rect 327080 335792 327132 335844
rect 328368 335792 328420 335844
rect 267004 335724 267056 335776
rect 267924 335724 267976 335776
rect 272340 335656 272392 335708
rect 275284 335656 275336 335708
rect 302608 335656 302660 335708
rect 303528 335656 303580 335708
rect 242256 335588 242308 335640
rect 242992 335588 243044 335640
rect 252008 335588 252060 335640
rect 258540 335588 258592 335640
rect 259368 335588 259420 335640
rect 265256 335588 265308 335640
rect 362316 335588 362368 335640
rect 362868 335588 362920 335640
rect 376116 335588 376168 335640
rect 376576 335588 376628 335640
rect 272800 335520 272852 335572
rect 277584 335520 277636 335572
rect 284392 335520 284444 335572
rect 285588 335520 285640 335572
rect 295524 335520 295576 335572
rect 296444 335520 296496 335572
rect 298192 335520 298244 335572
rect 299296 335520 299348 335572
rect 374276 335520 374328 335572
rect 375288 335520 375340 335572
rect 273260 335452 273312 335504
rect 274548 335452 274600 335504
rect 236644 335384 236696 335436
rect 239864 335384 239916 335436
rect 283012 335384 283064 335436
rect 284208 335384 284260 335436
rect 346676 335384 346728 335436
rect 347596 335384 347648 335436
rect 349344 335384 349396 335436
rect 350264 335384 350316 335436
rect 246304 335316 246356 335368
rect 248788 335316 248840 335368
rect 253204 335316 253256 335368
rect 259920 335316 259972 335368
rect 126888 334636 126940 334688
rect 215392 334636 215444 334688
rect 318616 334636 318668 334688
rect 398840 334636 398892 334688
rect 25504 334568 25556 334620
rect 176568 334568 176620 334620
rect 180708 334568 180760 334620
rect 235816 334568 235868 334620
rect 350448 334568 350500 334620
rect 483020 334568 483072 334620
rect 161388 333276 161440 333328
rect 228732 333276 228784 333328
rect 352932 333276 352984 333328
rect 489920 333276 489972 333328
rect 135168 333208 135220 333260
rect 218428 333208 218480 333260
rect 371240 333140 371292 333192
rect 539600 333208 539652 333260
rect 3056 332528 3108 332580
rect 166908 332528 166960 332580
rect 356980 331916 357032 331968
rect 500960 331916 501012 331968
rect 136548 331848 136600 331900
rect 218980 331848 219032 331900
rect 377864 331848 377916 331900
rect 556160 331848 556212 331900
rect 187884 331168 187936 331220
rect 188068 331168 188120 331220
rect 200396 331168 200448 331220
rect 200580 331168 200632 331220
rect 203156 331168 203208 331220
rect 203340 331168 203392 331220
rect 373264 330692 373316 330744
rect 373908 330692 373960 330744
rect 165528 330624 165580 330676
rect 230020 330624 230072 330676
rect 155868 330556 155920 330608
rect 226340 330556 226392 330608
rect 15844 330488 15896 330540
rect 171692 330488 171744 330540
rect 172612 330488 172664 330540
rect 172796 330488 172848 330540
rect 173992 330488 174044 330540
rect 174452 330488 174504 330540
rect 175464 330488 175516 330540
rect 175924 330488 175976 330540
rect 178132 330488 178184 330540
rect 179052 330488 179104 330540
rect 248512 330488 248564 330540
rect 249340 330488 249392 330540
rect 251272 330488 251324 330540
rect 251916 330488 251968 330540
rect 252652 330488 252704 330540
rect 253388 330488 253440 330540
rect 301780 330488 301832 330540
rect 354680 330488 354732 330540
rect 359648 330488 359700 330540
rect 507860 330488 507912 330540
rect 169852 330420 169904 330472
rect 170588 330420 170640 330472
rect 133788 329128 133840 329180
rect 218060 329128 218112 329180
rect 314200 329128 314252 329180
rect 387800 329128 387852 329180
rect 113088 329060 113140 329112
rect 210424 329060 210476 329112
rect 357440 329060 357492 329112
rect 502340 329060 502392 329112
rect 180892 328924 180944 328976
rect 181628 328924 181680 328976
rect 129648 327768 129700 327820
rect 216680 327768 216732 327820
rect 317144 327768 317196 327820
rect 394700 327768 394752 327820
rect 46204 327700 46256 327752
rect 183744 327700 183796 327752
rect 351552 327700 351604 327752
rect 485780 327700 485832 327752
rect 212724 326519 212776 326528
rect 212724 326485 212733 326519
rect 212733 326485 212767 326519
rect 212767 326485 212776 326519
rect 212724 326476 212776 326485
rect 223764 326519 223816 326528
rect 223764 326485 223773 326519
rect 223773 326485 223807 326519
rect 223807 326485 223816 326519
rect 223764 326476 223816 326485
rect 140688 326408 140740 326460
rect 220360 326408 220412 326460
rect 224960 326408 225012 326460
rect 225788 326408 225840 326460
rect 229284 326408 229336 326460
rect 262404 326408 262456 326460
rect 269212 326408 269264 326460
rect 318524 326408 318576 326460
rect 398932 326408 398984 326460
rect 39304 326340 39356 326392
rect 180984 326340 181036 326392
rect 186320 326340 186372 326392
rect 186964 326340 187016 326392
rect 187792 326340 187844 326392
rect 188252 326340 188304 326392
rect 189172 326340 189224 326392
rect 189724 326340 189776 326392
rect 190460 326340 190512 326392
rect 190736 326340 190788 326392
rect 200304 326340 200356 326392
rect 200764 326340 200816 326392
rect 203064 326340 203116 326392
rect 203524 326340 203576 326392
rect 204352 326340 204404 326392
rect 205180 326340 205232 326392
rect 205732 326340 205784 326392
rect 206100 326340 206152 326392
rect 211252 326340 211304 326392
rect 211436 326340 211488 326392
rect 215392 326340 215444 326392
rect 215852 326340 215904 326392
rect 219440 326340 219492 326392
rect 219900 326340 219952 326392
rect 223580 326340 223632 326392
rect 224316 326340 224368 326392
rect 225052 326340 225104 326392
rect 225236 326340 225288 326392
rect 227812 326340 227864 326392
rect 227996 326340 228048 326392
rect 204444 326272 204496 326324
rect 204628 326272 204680 326324
rect 230572 326340 230624 326392
rect 230756 326340 230808 326392
rect 231952 326340 232004 326392
rect 232412 326340 232464 326392
rect 233424 326340 233476 326392
rect 234252 326340 234304 326392
rect 241612 326340 241664 326392
rect 242164 326340 242216 326392
rect 242992 326340 243044 326392
rect 243452 326340 243504 326392
rect 255412 326340 255464 326392
rect 255964 326340 256016 326392
rect 267832 326340 267884 326392
rect 268476 326340 268528 326392
rect 354220 326340 354272 326392
rect 492680 326340 492732 326392
rect 190552 326204 190604 326256
rect 191012 326204 191064 326256
rect 229284 326204 229336 326256
rect 262404 326204 262456 326256
rect 269212 326204 269264 326256
rect 232044 325864 232096 325916
rect 232780 325864 232832 325916
rect 389180 325592 389232 325644
rect 579896 325592 579948 325644
rect 144828 324980 144880 325032
rect 221648 324980 221700 325032
rect 33784 324912 33836 324964
rect 179512 324912 179564 324964
rect 317236 324912 317288 324964
rect 396080 324912 396132 324964
rect 208492 324368 208544 324420
rect 208768 324368 208820 324420
rect 222200 324232 222252 324284
rect 222660 324232 222712 324284
rect 236092 323688 236144 323740
rect 236368 323688 236420 323740
rect 147588 323620 147640 323672
rect 222752 323620 222804 323672
rect 324136 323620 324188 323672
rect 412640 323620 412692 323672
rect 28908 323552 28960 323604
rect 178224 323552 178276 323604
rect 212724 323595 212776 323604
rect 212724 323561 212733 323595
rect 212733 323561 212767 323595
rect 212767 323561 212776 323595
rect 212724 323552 212776 323561
rect 229192 323552 229244 323604
rect 229376 323552 229428 323604
rect 234712 323552 234764 323604
rect 234896 323552 234948 323604
rect 365444 323552 365496 323604
rect 521660 323552 521712 323604
rect 131028 322260 131080 322312
rect 216772 322260 216824 322312
rect 319904 322260 319956 322312
rect 401600 322260 401652 322312
rect 51724 322192 51776 322244
rect 186504 322192 186556 322244
rect 362684 322192 362736 322244
rect 514760 322192 514812 322244
rect 223764 321963 223816 321972
rect 223764 321929 223773 321963
rect 223773 321929 223807 321963
rect 223807 321929 223816 321963
rect 223764 321920 223816 321929
rect 321284 320900 321336 320952
rect 405740 320900 405792 320952
rect 14464 320832 14516 320884
rect 172612 320832 172664 320884
rect 177948 320832 178000 320884
rect 233424 320832 233476 320884
rect 364064 320832 364116 320884
rect 517520 320832 517572 320884
rect 3056 320084 3108 320136
rect 166816 320084 166868 320136
rect 326896 319472 326948 319524
rect 419540 319472 419592 319524
rect 153108 319404 153160 319456
rect 225144 319404 225196 319456
rect 370964 319404 371016 319456
rect 535460 319404 535512 319456
rect 262312 319336 262364 319388
rect 262496 319336 262548 319388
rect 269120 319336 269172 319388
rect 269304 319336 269356 319388
rect 142068 318044 142120 318096
rect 220912 318044 220964 318096
rect 353116 318044 353168 318096
rect 488540 318044 488592 318096
rect 137928 316684 137980 316736
rect 219532 316684 219584 316736
rect 355784 316684 355836 316736
rect 495440 316684 495492 316736
rect 144736 315256 144788 315308
rect 222292 315256 222344 315308
rect 358544 315256 358596 315308
rect 506480 315256 506532 315308
rect 198832 313964 198884 314016
rect 199016 313964 199068 314016
rect 148968 313896 149020 313948
rect 223764 313896 223816 313948
rect 361304 313896 361356 313948
rect 513380 313896 513432 313948
rect 201592 313828 201644 313880
rect 201776 313828 201828 313880
rect 389272 313216 389324 313268
rect 580172 313216 580224 313268
rect 88248 312536 88300 312588
rect 200304 312536 200356 312588
rect 95148 311108 95200 311160
rect 203064 311108 203116 311160
rect 348884 311108 348936 311160
rect 477500 311108 477552 311160
rect 106188 309748 106240 309800
rect 207204 309748 207256 309800
rect 355876 309748 355928 309800
rect 496820 309748 496872 309800
rect 117228 308388 117280 308440
rect 211252 308388 211304 308440
rect 350356 308388 350408 308440
rect 481640 308388 481692 308440
rect 99288 307028 99340 307080
rect 202144 307028 202196 307080
rect 357256 307028 357308 307080
rect 499580 307028 499632 307080
rect 119988 305600 120040 305652
rect 212632 305600 212684 305652
rect 303344 305600 303396 305652
rect 357440 305600 357492 305652
rect 358636 305600 358688 305652
rect 503720 305600 503772 305652
rect 124128 304240 124180 304292
rect 214104 304240 214156 304292
rect 366824 304240 366876 304292
rect 524420 304240 524472 304292
rect 47584 302880 47636 302932
rect 185032 302880 185084 302932
rect 361396 302880 361448 302932
rect 510620 302880 510672 302932
rect 40684 301452 40736 301504
rect 182272 301452 182324 301504
rect 368204 301452 368256 301504
rect 528560 301452 528612 301504
rect 372344 300092 372396 300144
rect 542360 300092 542412 300144
rect 389364 299412 389416 299464
rect 579620 299412 579672 299464
rect 369584 297372 369636 297424
rect 531320 297372 531372 297424
rect 373724 295944 373776 295996
rect 546500 295944 546552 295996
rect 376484 294584 376536 294636
rect 553400 294584 553452 294636
rect 2780 293564 2832 293616
rect 4804 293564 4856 293616
rect 375104 293224 375156 293276
rect 549260 293224 549312 293276
rect 379244 291796 379296 291848
rect 560300 291796 560352 291848
rect 380624 290436 380676 290488
rect 564440 290436 564492 290488
rect 3148 280100 3200 280152
rect 166724 280100 166776 280152
rect 393964 273164 394016 273216
rect 580172 273164 580224 273216
rect 2964 267656 3016 267708
rect 166632 267656 166684 267708
rect 406384 259360 406436 259412
rect 580172 259360 580224 259412
rect 3148 255212 3200 255264
rect 21456 255212 21508 255264
rect 21364 254532 21416 254584
rect 173992 254532 174044 254584
rect 389456 245556 389508 245608
rect 580172 245556 580224 245608
rect 389548 233180 389600 233232
rect 579988 233180 580040 233232
rect 3240 229032 3292 229084
rect 166540 229032 166592 229084
rect 290464 224204 290516 224256
rect 322940 224204 322992 224256
rect 319996 222844 320048 222896
rect 402980 222844 403032 222896
rect 153016 221416 153068 221468
rect 225052 221416 225104 221468
rect 297916 221416 297968 221468
rect 340880 221416 340932 221468
rect 143448 220056 143500 220108
rect 220820 220056 220872 220108
rect 296444 220056 296496 220108
rect 338120 220056 338172 220108
rect 362776 220056 362828 220108
rect 516140 220056 516192 220108
rect 389640 219376 389692 219428
rect 580172 219376 580224 219428
rect 202788 218696 202840 218748
rect 242992 218696 243044 218748
rect 284024 218696 284076 218748
rect 306380 218696 306432 218748
rect 279884 217336 279936 217388
rect 295340 217336 295392 217388
rect 183468 217268 183520 217320
rect 236092 217268 236144 217320
rect 293776 217268 293828 217320
rect 331220 217268 331272 217320
rect 351736 217268 351788 217320
rect 487160 217268 487212 217320
rect 195888 215908 195940 215960
rect 239404 215908 239456 215960
rect 282644 215908 282696 215960
rect 302240 215908 302292 215960
rect 355968 215908 356020 215960
rect 498200 215908 498252 215960
rect 3240 215228 3292 215280
rect 166448 215228 166500 215280
rect 389732 206932 389784 206984
rect 579804 206932 579856 206984
rect 390468 193128 390520 193180
rect 580172 193128 580224 193180
rect 3332 188980 3384 189032
rect 10324 188980 10376 189032
rect 403624 179324 403676 179376
rect 580172 179324 580224 179376
rect 3332 176604 3384 176656
rect 166356 176604 166408 176656
rect 390376 166948 390428 167000
rect 580172 166948 580224 167000
rect 390284 153144 390336 153196
rect 580172 153144 580224 153196
rect 3332 150356 3384 150408
rect 28264 150356 28316 150408
rect 390192 139340 390244 139392
rect 580172 139340 580224 139392
rect 390100 126896 390152 126948
rect 580172 126896 580224 126948
rect 3148 124108 3200 124160
rect 166264 124108 166316 124160
rect 390008 113092 390060 113144
rect 579804 113092 579856 113144
rect 400864 100648 400916 100700
rect 580172 100648 580224 100700
rect 547144 86912 547196 86964
rect 580172 86912 580224 86964
rect 3148 85484 3200 85536
rect 11704 85484 11756 85536
rect 389916 73108 389968 73160
rect 580172 73108 580224 73160
rect 389824 60664 389876 60716
rect 580172 60664 580224 60716
rect 2872 59304 2924 59356
rect 29644 59304 29696 59356
rect 543004 46860 543056 46912
rect 580172 46860 580224 46912
rect 358728 42032 358780 42084
rect 505100 42032 505152 42084
rect 81348 28228 81400 28280
rect 197544 28228 197596 28280
rect 157248 26868 157300 26920
rect 226432 26868 226484 26920
rect 150348 25508 150400 25560
rect 223672 25508 223724 25560
rect 146208 24080 146260 24132
rect 222200 24080 222252 24132
rect 360016 24080 360068 24132
rect 506572 24080 506624 24132
rect 136456 22720 136508 22772
rect 218336 22720 218388 22772
rect 299204 22720 299256 22772
rect 347780 22720 347832 22772
rect 353024 22720 353076 22772
rect 490012 22720 490064 22772
rect 194416 21428 194468 21480
rect 240324 21428 240376 21480
rect 110328 21360 110380 21412
rect 208492 21360 208544 21412
rect 296536 21360 296588 21412
rect 340972 21360 341024 21412
rect 347596 21360 347648 21412
rect 473360 21360 473412 21412
rect 396724 20612 396776 20664
rect 579988 20612 580040 20664
rect 187608 19932 187660 19984
rect 237564 19932 237616 19984
rect 292396 19932 292448 19984
rect 329840 19932 329892 19984
rect 286876 18640 286928 18692
rect 313280 18640 313332 18692
rect 184848 18572 184900 18624
rect 233884 18572 233936 18624
rect 300584 18572 300636 18624
rect 350540 18572 350592 18624
rect 360108 18572 360160 18624
rect 509240 18572 509292 18624
rect 316684 17892 316736 17944
rect 324320 17892 324372 17944
rect 173808 17212 173860 17264
rect 232044 17212 232096 17264
rect 325424 17212 325476 17264
rect 415492 17212 415544 17264
rect 169576 15852 169628 15904
rect 222844 15852 222896 15904
rect 289636 15852 289688 15904
rect 322112 15852 322164 15904
rect 322664 15852 322716 15904
rect 409604 15852 409656 15904
rect 215208 14560 215260 14612
rect 246304 14560 246356 14612
rect 191748 14492 191800 14544
rect 236644 14492 236696 14544
rect 132224 14424 132276 14476
rect 216680 14424 216732 14476
rect 299296 14424 299348 14476
rect 345756 14424 345808 14476
rect 354496 14424 354548 14476
rect 492312 14424 492364 14476
rect 179052 13132 179104 13184
rect 234712 13132 234764 13184
rect 336004 13132 336056 13184
rect 390652 13132 390704 13184
rect 138848 13064 138900 13116
rect 219440 13064 219492 13116
rect 295064 13064 295116 13116
rect 334992 13064 335044 13116
rect 357348 13064 357400 13116
rect 499396 13064 499448 13116
rect 200028 11840 200080 11892
rect 242256 11840 242308 11892
rect 176568 11772 176620 11824
rect 233332 11772 233384 11824
rect 292488 11772 292540 11824
rect 328000 11772 328052 11824
rect 103244 11704 103296 11756
rect 205732 11704 205784 11756
rect 293868 11704 293920 11756
rect 332600 11704 332652 11756
rect 348976 11704 349028 11756
rect 480536 11704 480588 11756
rect 318064 10480 318116 10532
rect 344560 10480 344612 10532
rect 289728 10412 289780 10464
rect 320732 10412 320784 10464
rect 172428 10344 172480 10396
rect 231952 10344 232004 10396
rect 291108 10344 291160 10396
rect 326804 10344 326856 10396
rect 92388 10276 92440 10328
rect 177304 10276 177356 10328
rect 205548 10276 205600 10328
rect 244464 10276 244516 10328
rect 295156 10276 295208 10328
rect 337476 10276 337528 10328
rect 354588 10276 354640 10328
rect 494704 10276 494756 10328
rect 332324 9596 332376 9648
rect 435548 9596 435600 9648
rect 333796 9528 333848 9580
rect 439136 9528 439188 9580
rect 335084 9460 335136 9512
rect 442632 9460 442684 9512
rect 336556 9392 336608 9444
rect 446220 9392 446272 9444
rect 337844 9324 337896 9376
rect 449808 9324 449860 9376
rect 339316 9256 339368 9308
rect 453304 9256 453356 9308
rect 340604 9188 340656 9240
rect 456892 9188 456944 9240
rect 342076 9120 342128 9172
rect 460388 9120 460440 9172
rect 343272 9052 343324 9104
rect 463976 9052 464028 9104
rect 168656 8984 168708 9036
rect 229744 8984 229796 9036
rect 344836 8984 344888 9036
rect 467472 8984 467524 9036
rect 84476 8916 84528 8968
rect 173164 8916 173216 8968
rect 186136 8916 186188 8968
rect 237472 8916 237524 8968
rect 285404 8916 285456 8968
rect 310244 8916 310296 8968
rect 346124 8916 346176 8968
rect 471060 8916 471112 8968
rect 331036 8848 331088 8900
rect 432052 8848 432104 8900
rect 329564 8780 329616 8832
rect 428464 8780 428516 8832
rect 328184 8712 328236 8764
rect 424968 8712 425020 8764
rect 326988 8644 327040 8696
rect 421380 8644 421432 8696
rect 325516 8576 325568 8628
rect 417884 8576 417936 8628
rect 324228 8508 324280 8560
rect 414296 8508 414348 8560
rect 322756 8440 322808 8492
rect 410800 8440 410852 8492
rect 321376 8372 321428 8424
rect 407212 8372 407264 8424
rect 97448 8236 97500 8288
rect 204444 8236 204496 8288
rect 372436 8236 372488 8288
rect 541992 8236 542044 8288
rect 93952 8168 94004 8220
rect 202972 8168 203024 8220
rect 373816 8168 373868 8220
rect 545488 8168 545540 8220
rect 90364 8100 90416 8152
rect 201592 8100 201644 8152
rect 375196 8100 375248 8152
rect 549076 8100 549128 8152
rect 86868 8032 86920 8084
rect 200212 8032 200264 8084
rect 376576 8032 376628 8084
rect 552664 8032 552716 8084
rect 83280 7964 83332 8016
rect 198832 7964 198884 8016
rect 304724 7964 304776 8016
rect 361120 7964 361172 8016
rect 377956 7964 378008 8016
rect 556252 7964 556304 8016
rect 79692 7896 79744 7948
rect 197452 7896 197504 7948
rect 306104 7896 306156 7948
rect 364616 7896 364668 7948
rect 379336 7896 379388 7948
rect 559748 7896 559800 7948
rect 77392 7828 77444 7880
rect 196164 7828 196216 7880
rect 307484 7828 307536 7880
rect 368204 7828 368256 7880
rect 380716 7828 380768 7880
rect 563244 7828 563296 7880
rect 73804 7760 73856 7812
rect 194784 7760 194836 7812
rect 308864 7760 308916 7812
rect 371700 7760 371752 7812
rect 382004 7760 382056 7812
rect 566832 7760 566884 7812
rect 70308 7692 70360 7744
rect 193404 7692 193456 7744
rect 310152 7692 310204 7744
rect 375196 7692 375248 7744
rect 383384 7692 383436 7744
rect 570328 7692 570380 7744
rect 66720 7624 66772 7676
rect 192024 7624 192076 7676
rect 311624 7624 311676 7676
rect 378876 7624 378928 7676
rect 384764 7624 384816 7676
rect 573916 7624 573968 7676
rect 63224 7556 63276 7608
rect 190736 7556 190788 7608
rect 221556 7556 221608 7608
rect 247684 7556 247736 7608
rect 313004 7556 313056 7608
rect 382372 7556 382424 7608
rect 386052 7556 386104 7608
rect 577412 7556 577464 7608
rect 101036 7488 101088 7540
rect 205824 7488 205876 7540
rect 371056 7488 371108 7540
rect 538404 7488 538456 7540
rect 104532 7420 104584 7472
rect 207112 7420 207164 7472
rect 369676 7420 369728 7472
rect 534908 7420 534960 7472
rect 108120 7352 108172 7404
rect 208584 7352 208636 7404
rect 368296 7352 368348 7404
rect 531412 7352 531464 7404
rect 111616 7284 111668 7336
rect 209872 7284 209924 7336
rect 366916 7284 366968 7336
rect 527824 7284 527876 7336
rect 115204 7216 115256 7268
rect 211344 7216 211396 7268
rect 365536 7216 365588 7268
rect 524236 7216 524288 7268
rect 118792 7148 118844 7200
rect 212724 7148 212776 7200
rect 364156 7148 364208 7200
rect 520740 7148 520792 7200
rect 122288 7080 122340 7132
rect 214012 7080 214064 7132
rect 315764 7080 315816 7132
rect 393044 7080 393096 7132
rect 160100 7012 160152 7064
rect 227812 7012 227864 7064
rect 315856 7012 315908 7064
rect 389456 7012 389508 7064
rect 3424 6808 3476 6860
rect 18604 6808 18656 6860
rect 48964 6808 49016 6860
rect 186412 6808 186464 6860
rect 337936 6808 337988 6860
rect 448612 6808 448664 6860
rect 519544 6808 519596 6860
rect 580172 6808 580224 6860
rect 44272 6740 44324 6792
rect 183652 6740 183704 6792
rect 339408 6740 339460 6792
rect 452108 6740 452160 6792
rect 40776 6672 40828 6724
rect 182364 6672 182416 6724
rect 340696 6672 340748 6724
rect 455696 6672 455748 6724
rect 37188 6604 37240 6656
rect 180892 6604 180944 6656
rect 197912 6604 197964 6656
rect 241612 6604 241664 6656
rect 342168 6604 342220 6656
rect 459192 6604 459244 6656
rect 33600 6536 33652 6588
rect 179604 6536 179656 6588
rect 192024 6536 192076 6588
rect 240232 6536 240284 6588
rect 343456 6536 343508 6588
rect 462780 6536 462832 6588
rect 30104 6468 30156 6520
rect 178132 6468 178184 6520
rect 188528 6468 188580 6520
rect 238852 6468 238904 6520
rect 343364 6468 343416 6520
rect 466276 6468 466328 6520
rect 26516 6400 26568 6452
rect 176752 6400 176804 6452
rect 184940 6400 184992 6452
rect 237380 6400 237432 6452
rect 344928 6400 344980 6452
rect 469864 6400 469916 6452
rect 21824 6332 21876 6384
rect 175464 6332 175516 6384
rect 181444 6332 181496 6384
rect 236184 6332 236236 6384
rect 346216 6332 346268 6384
rect 473452 6332 473504 6384
rect 17040 6264 17092 6316
rect 174084 6264 174136 6316
rect 177856 6264 177908 6316
rect 234804 6264 234856 6316
rect 347688 6264 347740 6316
rect 476948 6264 477000 6316
rect 8760 6196 8812 6248
rect 171232 6196 171284 6248
rect 174268 6196 174320 6248
rect 233240 6196 233292 6248
rect 281264 6196 281316 6248
rect 299664 6196 299716 6248
rect 350264 6196 350316 6248
rect 481732 6196 481784 6248
rect 4068 6128 4120 6180
rect 168564 6128 168616 6180
rect 170772 6128 170824 6180
rect 232136 6128 232188 6180
rect 288164 6128 288216 6180
rect 317328 6128 317380 6180
rect 320824 6128 320876 6180
rect 332692 6128 332744 6180
rect 351828 6128 351880 6180
rect 485228 6128 485280 6180
rect 52552 6060 52604 6112
rect 187884 6060 187936 6112
rect 336648 6060 336700 6112
rect 445024 6060 445076 6112
rect 56048 5992 56100 6044
rect 189264 5992 189316 6044
rect 335176 5992 335228 6044
rect 441528 5992 441580 6044
rect 59636 5924 59688 5976
rect 190644 5924 190696 5976
rect 333888 5924 333940 5976
rect 437940 5924 437992 5976
rect 76196 5856 76248 5908
rect 196072 5856 196124 5908
rect 332416 5856 332468 5908
rect 434444 5856 434496 5908
rect 128176 5788 128228 5840
rect 215392 5788 215444 5840
rect 331128 5788 331180 5840
rect 430856 5788 430908 5840
rect 158904 5720 158956 5772
rect 227904 5720 227956 5772
rect 329656 5720 329708 5772
rect 427268 5720 427320 5772
rect 163688 5652 163740 5704
rect 229192 5652 229244 5704
rect 328276 5652 328328 5704
rect 423772 5652 423824 5704
rect 167184 5584 167236 5636
rect 230572 5584 230624 5636
rect 313924 5516 313976 5568
rect 315028 5516 315080 5568
rect 323584 5516 323636 5568
rect 324412 5516 324464 5568
rect 65524 5448 65576 5500
rect 191932 5448 191984 5500
rect 302148 5448 302200 5500
rect 354036 5448 354088 5500
rect 372252 5448 372304 5500
rect 540796 5448 540848 5500
rect 62028 5380 62080 5432
rect 190552 5380 190604 5432
rect 302056 5380 302108 5432
rect 356336 5380 356388 5432
rect 373908 5380 373960 5432
rect 544384 5380 544436 5432
rect 58440 5312 58492 5364
rect 189172 5312 189224 5364
rect 303528 5312 303580 5364
rect 357532 5312 357584 5364
rect 375288 5312 375340 5364
rect 547880 5312 547932 5364
rect 54944 5244 54996 5296
rect 187792 5244 187844 5296
rect 303436 5244 303488 5296
rect 359924 5244 359976 5296
rect 376668 5244 376720 5296
rect 551468 5244 551520 5296
rect 51356 5176 51408 5228
rect 186320 5176 186372 5228
rect 211068 5176 211120 5228
rect 247132 5176 247184 5228
rect 304816 5176 304868 5228
rect 363512 5176 363564 5228
rect 378048 5176 378100 5228
rect 554964 5176 555016 5228
rect 47860 5108 47912 5160
rect 185124 5108 185176 5160
rect 207388 5108 207440 5160
rect 245844 5108 245896 5160
rect 306196 5108 306248 5160
rect 367008 5108 367060 5160
rect 379428 5108 379480 5160
rect 558552 5108 558604 5160
rect 12348 5040 12400 5092
rect 172704 5040 172756 5092
rect 203892 5040 203944 5092
rect 244372 5040 244424 5092
rect 307576 5040 307628 5092
rect 370596 5040 370648 5092
rect 380808 5040 380860 5092
rect 562048 5040 562100 5092
rect 7656 4972 7708 5024
rect 169852 4972 169904 5024
rect 200304 4972 200356 5024
rect 243084 4972 243136 5024
rect 308956 4972 309008 5024
rect 374092 4972 374144 5024
rect 382096 4972 382148 5024
rect 565636 4972 565688 5024
rect 2872 4904 2924 4956
rect 168380 4904 168432 4956
rect 196808 4904 196860 4956
rect 241704 4904 241756 4956
rect 310336 4904 310388 4956
rect 377680 4904 377732 4956
rect 383476 4904 383528 4956
rect 569132 4904 569184 4956
rect 572 4836 624 4888
rect 167000 4836 167052 4888
rect 193220 4836 193272 4888
rect 240140 4836 240192 4888
rect 311716 4836 311768 4888
rect 381176 4836 381228 4888
rect 384856 4836 384908 4888
rect 572720 4836 572772 4888
rect 1676 4768 1728 4820
rect 168472 4768 168524 4820
rect 189724 4768 189776 4820
rect 238944 4768 238996 4820
rect 277124 4768 277176 4820
rect 288992 4768 289044 4820
rect 313096 4768 313148 4820
rect 384764 4768 384816 4820
rect 386144 4768 386196 4820
rect 576308 4768 576360 4820
rect 69112 4700 69164 4752
rect 193312 4700 193364 4752
rect 301964 4700 302016 4752
rect 352840 4700 352892 4752
rect 371148 4700 371200 4752
rect 537208 4700 537260 4752
rect 72608 4632 72660 4684
rect 194692 4632 194744 4684
rect 300676 4632 300728 4684
rect 349252 4632 349304 4684
rect 369768 4632 369820 4684
rect 533712 4632 533764 4684
rect 126980 4564 127032 4616
rect 215484 4564 215536 4616
rect 300768 4564 300820 4616
rect 350448 4564 350500 4616
rect 368388 4564 368440 4616
rect 530124 4564 530176 4616
rect 150624 4496 150676 4548
rect 223580 4496 223632 4548
rect 299388 4496 299440 4548
rect 154212 4428 154264 4480
rect 224960 4428 225012 4480
rect 298008 4428 298060 4480
rect 343364 4428 343416 4480
rect 157800 4360 157852 4412
rect 226524 4360 226576 4412
rect 296628 4360 296680 4412
rect 339868 4360 339920 4412
rect 366916 4496 366968 4548
rect 526628 4496 526680 4548
rect 365628 4428 365680 4480
rect 523040 4428 523092 4480
rect 346952 4360 347004 4412
rect 364248 4360 364300 4412
rect 519544 4360 519596 4412
rect 162492 4292 162544 4344
rect 229284 4292 229336 4344
rect 295248 4292 295300 4344
rect 336280 4292 336332 4344
rect 362868 4292 362920 4344
rect 515956 4292 516008 4344
rect 166080 4224 166132 4276
rect 230664 4224 230716 4276
rect 361488 4224 361540 4276
rect 512460 4224 512512 4276
rect 135260 4156 135312 4208
rect 136456 4156 136508 4208
rect 143540 4156 143592 4208
rect 144828 4156 144880 4208
rect 151820 4156 151872 4208
rect 153108 4156 153160 4208
rect 178316 4156 178368 4208
rect 291844 4156 291896 4208
rect 292580 4156 292632 4208
rect 314476 4156 314528 4208
rect 385960 4156 386012 4208
rect 6460 4088 6512 4140
rect 7564 4088 7616 4140
rect 78588 4088 78640 4140
rect 197360 4088 197412 4140
rect 233424 4088 233476 4140
rect 254032 4088 254084 4140
rect 279976 4088 280028 4140
rect 297272 4088 297324 4140
rect 332508 4088 332560 4140
rect 436744 4088 436796 4140
rect 75000 4020 75052 4072
rect 195980 4020 196032 4072
rect 231032 4020 231084 4072
rect 254124 4020 254176 4072
rect 288256 4020 288308 4072
rect 316224 4020 316276 4072
rect 335268 4020 335320 4072
rect 443828 4020 443880 4072
rect 71504 3952 71556 4004
rect 194600 3952 194652 4004
rect 229836 3952 229888 4004
rect 252652 3952 252704 4004
rect 277216 3952 277268 4004
rect 287796 3952 287848 4004
rect 288348 3952 288400 4004
rect 319720 3952 319772 4004
rect 328368 3952 328420 4004
rect 338028 3952 338080 4004
rect 340880 3952 340932 4004
rect 342168 3952 342220 4004
rect 450912 3952 450964 4004
rect 14740 3884 14792 3936
rect 17224 3884 17276 3936
rect 67916 3884 67968 3936
rect 193128 3884 193180 3936
rect 228732 3884 228784 3936
rect 231124 3884 231176 3936
rect 252744 3884 252796 3936
rect 281448 3884 281500 3936
rect 300768 3884 300820 3936
rect 304908 3884 304960 3936
rect 357440 3884 357492 3936
rect 358728 3884 358780 3936
rect 362316 3884 362368 3936
rect 382188 3884 382240 3936
rect 568028 3884 568080 3936
rect 45468 3816 45520 3868
rect 47584 3816 47636 3868
rect 64328 3816 64380 3868
rect 60832 3748 60884 3800
rect 190460 3816 190512 3868
rect 227536 3816 227588 3868
rect 57244 3680 57296 3732
rect 191840 3748 191892 3800
rect 223948 3748 224000 3800
rect 251272 3748 251324 3800
rect 226340 3680 226392 3732
rect 251364 3680 251416 3732
rect 53748 3612 53800 3664
rect 187700 3612 187752 3664
rect 219256 3612 219308 3664
rect 247592 3612 247644 3664
rect 248328 3612 248380 3664
rect 25320 3544 25372 3596
rect 32404 3544 32456 3596
rect 34796 3544 34848 3596
rect 39304 3544 39356 3596
rect 43076 3544 43128 3596
rect 183560 3544 183612 3596
rect 216864 3544 216916 3596
rect 13544 3476 13596 3528
rect 14464 3476 14516 3528
rect 18236 3476 18288 3528
rect 21364 3476 21416 3528
rect 24216 3476 24268 3528
rect 15936 3408 15988 3460
rect 22744 3408 22796 3460
rect 27712 3476 27764 3528
rect 28908 3476 28960 3528
rect 39580 3476 39632 3528
rect 43444 3476 43496 3528
rect 35164 3408 35216 3460
rect 35992 3340 36044 3392
rect 9956 3272 10008 3324
rect 15844 3272 15896 3324
rect 28908 3272 28960 3324
rect 171968 3476 172020 3528
rect 172428 3476 172480 3528
rect 173164 3476 173216 3528
rect 173808 3476 173860 3528
rect 175464 3476 175516 3528
rect 176568 3476 176620 3528
rect 176660 3476 176712 3528
rect 177948 3476 178000 3528
rect 180248 3476 180300 3528
rect 180708 3476 180760 3528
rect 182548 3476 182600 3528
rect 183468 3476 183520 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 190828 3476 190880 3528
rect 191748 3476 191800 3528
rect 199108 3476 199160 3528
rect 200028 3476 200080 3528
rect 201500 3476 201552 3528
rect 202788 3476 202840 3528
rect 205088 3476 205140 3528
rect 205548 3476 205600 3528
rect 206192 3476 206244 3528
rect 206928 3476 206980 3528
rect 208584 3476 208636 3528
rect 209688 3476 209740 3528
rect 209780 3476 209832 3528
rect 210976 3476 211028 3528
rect 213368 3476 213420 3528
rect 213828 3476 213880 3528
rect 214472 3476 214524 3528
rect 215208 3476 215260 3528
rect 215668 3476 215720 3528
rect 242900 3544 242952 3596
rect 250536 3612 250588 3664
rect 259644 3816 259696 3868
rect 282828 3816 282880 3868
rect 301964 3816 302016 3868
rect 306288 3816 306340 3868
rect 365812 3816 365864 3868
rect 383568 3816 383620 3868
rect 571524 3816 571576 3868
rect 255872 3748 255924 3800
rect 263784 3748 263836 3800
rect 284208 3748 284260 3800
rect 305552 3748 305604 3800
rect 257068 3680 257120 3732
rect 258724 3680 258776 3732
rect 254676 3612 254728 3664
rect 263692 3680 263744 3732
rect 285588 3680 285640 3732
rect 309048 3680 309100 3732
rect 248512 3476 248564 3528
rect 181076 3408 181128 3460
rect 189080 3408 189132 3460
rect 202696 3408 202748 3460
rect 244188 3408 244240 3460
rect 245200 3408 245252 3460
rect 252376 3544 252428 3596
rect 262312 3612 262364 3664
rect 282736 3612 282788 3664
rect 304356 3612 304408 3664
rect 307668 3612 307720 3664
rect 369400 3748 369452 3800
rect 384948 3748 385000 3800
rect 575112 3748 575164 3800
rect 259460 3544 259512 3596
rect 260656 3544 260708 3596
rect 261760 3544 261812 3596
rect 265624 3544 265676 3596
rect 269120 3544 269172 3596
rect 270040 3544 270092 3596
rect 274364 3544 274416 3596
rect 280712 3544 280764 3596
rect 284116 3544 284168 3596
rect 307944 3544 307996 3596
rect 308956 3544 309008 3596
rect 372896 3680 372948 3732
rect 386328 3680 386380 3732
rect 578608 3680 578660 3732
rect 310428 3612 310480 3664
rect 376484 3612 376536 3664
rect 387616 3612 387668 3664
rect 582196 3612 582248 3664
rect 311808 3544 311860 3596
rect 379980 3544 380032 3596
rect 387524 3544 387576 3596
rect 248788 3476 248840 3528
rect 255504 3408 255556 3460
rect 258264 3476 258316 3528
rect 259368 3476 259420 3528
rect 265348 3476 265400 3528
rect 267004 3476 267056 3528
rect 271696 3476 271748 3528
rect 274824 3476 274876 3528
rect 278596 3476 278648 3528
rect 286968 3476 287020 3528
rect 312636 3476 312688 3528
rect 313188 3476 313240 3528
rect 383568 3476 383620 3528
rect 386236 3476 386288 3528
rect 390652 3476 390704 3528
rect 391848 3476 391900 3528
rect 579804 3544 579856 3596
rect 581000 3476 581052 3528
rect 261024 3408 261076 3460
rect 262956 3408 263008 3460
rect 265716 3408 265768 3460
rect 274456 3408 274508 3460
rect 281908 3408 281960 3460
rect 285496 3408 285548 3460
rect 311440 3408 311492 3460
rect 314568 3408 314620 3460
rect 387156 3408 387208 3460
rect 387708 3408 387760 3460
rect 583392 3408 583444 3460
rect 50160 3340 50212 3392
rect 51724 3340 51776 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 82084 3340 82136 3392
rect 198924 3340 198976 3392
rect 218060 3340 218112 3392
rect 219348 3340 219400 3392
rect 225144 3340 225196 3392
rect 226984 3340 227036 3392
rect 91560 3272 91612 3324
rect 92388 3272 92440 3324
rect 200396 3272 200448 3324
rect 222752 3272 222804 3324
rect 234620 3340 234672 3392
rect 255412 3340 255464 3392
rect 281356 3340 281408 3392
rect 298468 3340 298520 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 238116 3272 238168 3324
rect 248420 3272 248472 3324
rect 253204 3272 253256 3324
rect 282184 3272 282236 3324
rect 285404 3272 285456 3324
rect 89168 3204 89220 3256
rect 201684 3204 201736 3256
rect 241704 3204 241756 3256
rect 258172 3204 258224 3256
rect 280068 3204 280120 3256
rect 294880 3272 294932 3324
rect 329748 3272 329800 3324
rect 429660 3340 429712 3392
rect 431960 3340 432012 3392
rect 433248 3340 433300 3392
rect 473360 3340 473412 3392
rect 474556 3340 474608 3392
rect 481640 3340 481692 3392
rect 482836 3340 482888 3392
rect 489920 3340 489972 3392
rect 491116 3340 491168 3392
rect 531320 3340 531372 3392
rect 532516 3340 532568 3392
rect 556160 3340 556212 3392
rect 557356 3340 557408 3392
rect 422576 3272 422628 3324
rect 23020 3136 23072 3188
rect 25504 3136 25556 3188
rect 31300 3136 31352 3188
rect 33784 3136 33836 3188
rect 38384 3136 38436 3188
rect 40684 3136 40736 3188
rect 46664 3136 46716 3188
rect 50344 3136 50396 3188
rect 85672 3136 85724 3188
rect 92756 3136 92808 3188
rect 203156 3136 203208 3188
rect 248696 3136 248748 3188
rect 251180 3136 251232 3188
rect 262404 3136 262456 3188
rect 264152 3136 264204 3188
rect 266452 3136 266504 3188
rect 278688 3136 278740 3188
rect 293684 3204 293736 3256
rect 325516 3204 325568 3256
rect 415400 3204 415452 3256
rect 415492 3204 415544 3256
rect 416688 3204 416740 3256
rect 291384 3136 291436 3188
rect 322848 3136 322900 3188
rect 408408 3136 408460 3188
rect 98644 3068 98696 3120
rect 99288 3068 99340 3120
rect 102232 3068 102284 3120
rect 103244 3068 103296 3120
rect 105728 3068 105780 3120
rect 106188 3068 106240 3120
rect 109316 3068 109368 3120
rect 110328 3068 110380 3120
rect 41880 3000 41932 3052
rect 46204 3000 46256 3052
rect 96252 3000 96304 3052
rect 204536 3068 204588 3120
rect 240508 3068 240560 3120
rect 251916 3068 251968 3120
rect 266544 3068 266596 3120
rect 268016 3068 268068 3120
rect 274548 3068 274600 3120
rect 32404 2932 32456 2984
rect 36544 2932 36596 2984
rect 99840 2932 99892 2984
rect 204352 3000 204404 3052
rect 232228 3000 232280 3052
rect 242164 3000 242216 3052
rect 244096 3000 244148 3052
rect 251824 3000 251876 3052
rect 275284 3000 275336 3052
rect 277124 3000 277176 3052
rect 277308 3068 277360 3120
rect 290188 3068 290240 3120
rect 321468 3068 321520 3120
rect 404820 3068 404872 3120
rect 279516 3000 279568 3052
rect 320088 3000 320140 3052
rect 110512 2864 110564 2916
rect 111708 2864 111760 2916
rect 106924 2796 106976 2848
rect 207296 2932 207348 2984
rect 249892 2932 249944 2984
rect 271788 2932 271840 2984
rect 273628 2932 273680 2984
rect 318616 2932 318668 2984
rect 397736 2932 397788 2984
rect 398840 3000 398892 3052
rect 400128 3000 400180 3052
rect 401324 2932 401376 2984
rect 116400 2864 116452 2916
rect 117228 2864 117280 2916
rect 117596 2864 117648 2916
rect 118608 2864 118660 2916
rect 123484 2864 123536 2916
rect 124128 2864 124180 2916
rect 124680 2864 124732 2916
rect 125968 2864 126020 2916
rect 126888 2864 126940 2916
rect 114008 2796 114060 2848
rect 130568 2864 130620 2916
rect 131028 2864 131080 2916
rect 131764 2864 131816 2916
rect 132224 2864 132276 2916
rect 210056 2864 210108 2916
rect 237012 2864 237064 2916
rect 214196 2796 214248 2848
rect 239312 2796 239364 2848
rect 246396 2796 246448 2848
rect 249064 2796 249116 2848
rect 249984 2864 250036 2916
rect 253296 2864 253348 2916
rect 317236 2864 317288 2916
rect 394240 2864 394292 2916
rect 250444 2796 250496 2848
rect 248604 2728 248656 2780
rect 256884 2796 256936 2848
rect 315948 2796 316000 2848
rect 390652 2796 390704 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 696998 3464 697303
rect 3424 696992 3476 696998
rect 3424 696934 3476 696940
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2778 645144 2834 645153
rect 2778 645079 2780 645088
rect 2832 645079 2834 645088
rect 2780 645050 2832 645056
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3238 540832 3294 540841
rect 3238 540767 3294 540776
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 3054 514856 3110 514865
rect 3054 514791 3110 514800
rect 2962 501800 3018 501809
rect 2962 501735 3018 501744
rect 2870 488744 2926 488753
rect 2870 488679 2926 488688
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 433294 2820 475623
rect 2884 436082 2912 488679
rect 2976 438870 3004 501735
rect 3068 441590 3096 514791
rect 3160 442950 3188 527847
rect 3252 445738 3280 540767
rect 3344 448526 3372 553823
rect 3436 471986 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3424 471980 3476 471986
rect 3424 471922 3476 471928
rect 3528 469198 3556 658135
rect 4804 645108 4856 645114
rect 4804 645050 4856 645056
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3516 469192 3568 469198
rect 3516 469134 3568 469140
rect 3620 463690 3648 632023
rect 3698 619168 3754 619177
rect 3698 619103 3754 619112
rect 3608 463684 3660 463690
rect 3608 463626 3660 463632
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3332 448520 3384 448526
rect 3332 448462 3384 448468
rect 3240 445732 3292 445738
rect 3240 445674 3292 445680
rect 3148 442944 3200 442950
rect 3148 442886 3200 442892
rect 3056 441584 3108 441590
rect 3056 441526 3108 441532
rect 2964 438864 3016 438870
rect 2964 438806 3016 438812
rect 2872 436076 2924 436082
rect 2872 436018 2924 436024
rect 2780 433288 2832 433294
rect 2780 433230 2832 433236
rect 3436 430574 3464 462567
rect 3712 462330 3740 619103
rect 3790 606112 3846 606121
rect 3790 606047 3846 606056
rect 3700 462324 3752 462330
rect 3700 462266 3752 462272
rect 3804 459542 3832 606047
rect 3882 593056 3938 593065
rect 3882 592991 3938 593000
rect 3792 459536 3844 459542
rect 3792 459478 3844 459484
rect 3896 456754 3924 592991
rect 3974 580000 4030 580009
rect 3974 579935 4030 579944
rect 3884 456748 3936 456754
rect 3884 456690 3936 456696
rect 3988 454034 4016 579935
rect 4066 566944 4122 566953
rect 4066 566879 4122 566888
rect 3976 454028 4028 454034
rect 3976 453970 4028 453976
rect 4080 451246 4108 566879
rect 4816 466410 4844 645050
rect 8220 480962 8248 702406
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 24780 481030 24808 699654
rect 41340 481098 41368 700334
rect 56796 700194 56824 703520
rect 72988 702434 73016 703520
rect 72988 702406 73108 702434
rect 56784 700188 56836 700194
rect 56784 700130 56836 700136
rect 57888 700188 57940 700194
rect 57888 700130 57940 700136
rect 57900 481166 57928 700130
rect 73080 481234 73108 702406
rect 89180 699718 89208 703520
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 106188 700392 106240 700398
rect 106188 700334 106240 700340
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 86224 696992 86276 696998
rect 86224 696934 86276 696940
rect 73068 481228 73120 481234
rect 73068 481170 73120 481176
rect 57888 481160 57940 481166
rect 57888 481102 57940 481108
rect 41328 481092 41380 481098
rect 41328 481034 41380 481040
rect 24768 481024 24820 481030
rect 24768 480966 24820 480972
rect 8208 480956 8260 480962
rect 8208 480898 8260 480904
rect 86236 477494 86264 696934
rect 89640 481302 89668 699654
rect 106200 481370 106228 700334
rect 121656 699718 121684 703520
rect 137848 702434 137876 703520
rect 154132 702434 154160 703520
rect 137848 702406 137968 702434
rect 154132 702406 154528 702434
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 122748 699712 122800 699718
rect 122748 699654 122800 699660
rect 122760 481438 122788 699654
rect 137940 481506 137968 702406
rect 154500 481574 154528 702406
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 171048 700256 171100 700262
rect 171048 700198 171100 700204
rect 171060 489914 171088 700198
rect 186516 700194 186544 703520
rect 186504 700188 186556 700194
rect 186504 700130 186556 700136
rect 187608 700188 187660 700194
rect 187608 700130 187660 700136
rect 170968 489886 171088 489914
rect 154488 481568 154540 481574
rect 154488 481510 154540 481516
rect 137928 481500 137980 481506
rect 137928 481442 137980 481448
rect 122748 481432 122800 481438
rect 122748 481374 122800 481380
rect 106188 481364 106240 481370
rect 106188 481306 106240 481312
rect 89628 481296 89680 481302
rect 89628 481238 89680 481244
rect 170968 480894 170996 489886
rect 183192 481092 183244 481098
rect 183192 481034 183244 481040
rect 177120 481024 177172 481030
rect 177120 480966 177172 480972
rect 171048 480956 171100 480962
rect 171048 480898 171100 480904
rect 170956 480888 171008 480894
rect 170956 480830 171008 480836
rect 171060 477972 171088 480898
rect 177132 477972 177160 480966
rect 183204 477972 183232 481034
rect 187620 481030 187648 700130
rect 201592 481296 201644 481302
rect 201592 481238 201644 481244
rect 195428 481228 195480 481234
rect 195428 481170 195480 481176
rect 189356 481160 189408 481166
rect 189356 481102 189408 481108
rect 187608 481024 187660 481030
rect 187608 480966 187660 480972
rect 189368 477972 189396 481102
rect 195440 477972 195468 481170
rect 201604 477972 201632 481238
rect 202800 481098 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 213736 481432 213788 481438
rect 213736 481374 213788 481380
rect 207664 481364 207716 481370
rect 207664 481306 207716 481312
rect 202788 481092 202840 481098
rect 202788 481034 202840 481040
rect 207676 477972 207704 481306
rect 213748 477972 213776 481374
rect 219360 481166 219388 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 235908 700392 235960 700398
rect 235908 700334 235960 700340
rect 225972 481568 226024 481574
rect 225972 481510 226024 481516
rect 219900 481500 219952 481506
rect 219900 481442 219952 481448
rect 219348 481160 219400 481166
rect 219348 481102 219400 481108
rect 219912 477972 219940 481442
rect 225984 477972 226012 481510
rect 235920 480962 235948 700334
rect 251468 700126 251496 703520
rect 251456 700120 251508 700126
rect 251456 700062 251508 700068
rect 252468 700120 252520 700126
rect 252468 700062 252520 700068
rect 250444 481160 250496 481166
rect 250444 481102 250496 481108
rect 244372 481092 244424 481098
rect 244372 481034 244424 481040
rect 238208 481024 238260 481030
rect 238208 480966 238260 480972
rect 232136 480956 232188 480962
rect 232136 480898 232188 480904
rect 235908 480956 235960 480962
rect 235908 480898 235960 480904
rect 232148 477972 232176 480898
rect 238220 477972 238248 480966
rect 244384 477972 244412 481034
rect 250456 477972 250484 481102
rect 252480 481030 252508 700062
rect 252468 481024 252520 481030
rect 252468 480966 252520 480972
rect 262680 481024 262732 481030
rect 262680 480966 262732 480972
rect 256516 480956 256568 480962
rect 256516 480898 256568 480904
rect 256528 477972 256556 480898
rect 262692 477972 262720 480966
rect 267660 480282 267688 703520
rect 283852 700398 283880 703520
rect 288348 700596 288400 700602
rect 288348 700538 288400 700544
rect 276664 700392 276716 700398
rect 276664 700334 276716 700340
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 276676 481642 276704 700334
rect 281448 700324 281500 700330
rect 281448 700266 281500 700272
rect 274916 481636 274968 481642
rect 274916 481578 274968 481584
rect 276664 481636 276716 481642
rect 276664 481578 276716 481584
rect 267648 480276 267700 480282
rect 267648 480218 267700 480224
rect 268752 480276 268804 480282
rect 268752 480218 268804 480224
rect 268764 477972 268792 480218
rect 274928 477972 274956 481578
rect 281460 480254 281488 700266
rect 288360 481370 288388 700538
rect 293868 700528 293920 700534
rect 293868 700470 293920 700476
rect 287060 481364 287112 481370
rect 287060 481306 287112 481312
rect 288348 481364 288400 481370
rect 288348 481306 288400 481312
rect 281368 480226 281488 480254
rect 281368 477986 281396 480226
rect 281014 477958 281396 477986
rect 287072 477972 287100 481306
rect 293880 480254 293908 700470
rect 299388 700460 299440 700466
rect 299388 700402 299440 700408
rect 293696 480226 293908 480254
rect 293696 477986 293724 480226
rect 299400 477986 299428 700402
rect 300136 700330 300164 703520
rect 316328 700602 316356 703520
rect 324228 701004 324280 701010
rect 324228 700946 324280 700952
rect 316316 700596 316368 700602
rect 316316 700538 316368 700544
rect 306288 700392 306340 700398
rect 306288 700334 306340 700340
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 306300 481642 306328 700334
rect 311808 700324 311860 700330
rect 311808 700266 311860 700272
rect 305460 481636 305512 481642
rect 305460 481578 305512 481584
rect 306288 481636 306340 481642
rect 306288 481578 306340 481584
rect 293250 477958 293724 477986
rect 299322 477958 299428 477986
rect 305472 477972 305500 481578
rect 311820 477986 311848 700266
rect 318708 700256 318760 700262
rect 318708 700198 318760 700204
rect 318720 481234 318748 700198
rect 317696 481228 317748 481234
rect 317696 481170 317748 481176
rect 318708 481228 318760 481234
rect 318708 481170 318760 481176
rect 311558 477958 311848 477986
rect 317708 477972 317736 481170
rect 324240 477986 324268 700946
rect 331128 700936 331180 700942
rect 331128 700878 331180 700884
rect 331140 481642 331168 700878
rect 332520 700534 332548 703520
rect 336648 700868 336700 700874
rect 336648 700810 336700 700816
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 329840 481636 329892 481642
rect 329840 481578 329892 481584
rect 331128 481636 331180 481642
rect 331128 481578 331180 481584
rect 323794 477958 324268 477986
rect 329852 477972 329880 481578
rect 336660 480254 336688 700810
rect 342168 700800 342220 700806
rect 342168 700742 342220 700748
rect 336384 480226 336688 480254
rect 336384 477986 336412 480226
rect 342180 477986 342208 700742
rect 348804 700466 348832 703520
rect 349068 700732 349120 700738
rect 349068 700674 349120 700680
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 349080 481098 349108 700674
rect 354588 700664 354640 700670
rect 354588 700606 354640 700612
rect 348240 481092 348292 481098
rect 348240 481034 348292 481040
rect 349068 481092 349120 481098
rect 349068 481034 349120 481040
rect 336030 477958 336412 477986
rect 342102 477958 342208 477986
rect 348252 477972 348280 481034
rect 354600 477986 354628 700606
rect 361488 700596 361540 700602
rect 361488 700538 361540 700544
rect 361500 481166 361528 700538
rect 364996 700398 365024 703520
rect 367008 700528 367060 700534
rect 367008 700470 367060 700476
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 360384 481160 360436 481166
rect 360384 481102 360436 481108
rect 361488 481160 361540 481166
rect 361488 481102 361540 481108
rect 354338 477958 354628 477986
rect 360396 477972 360424 481102
rect 367020 480254 367048 700470
rect 373908 700460 373960 700466
rect 373908 700402 373960 700408
rect 373920 480826 373948 700402
rect 379428 700392 379480 700398
rect 379428 700334 379480 700340
rect 372620 480820 372672 480826
rect 372620 480762 372672 480768
rect 373908 480820 373960 480826
rect 373908 480762 373960 480768
rect 366928 480226 367048 480254
rect 366928 477986 366956 480226
rect 366574 477958 366956 477986
rect 372632 477972 372660 480762
rect 379440 480254 379468 700334
rect 381188 700330 381216 703520
rect 381176 700324 381228 700330
rect 381176 700266 381228 700272
rect 384948 700324 385000 700330
rect 384948 700266 385000 700272
rect 379256 480226 379468 480254
rect 379256 477986 379284 480226
rect 384960 477986 384988 700266
rect 397472 700262 397500 703520
rect 413664 701010 413692 703520
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 429856 700942 429884 703520
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 446140 700874 446168 703520
rect 446128 700868 446180 700874
rect 446128 700810 446180 700816
rect 462332 700806 462360 703520
rect 462320 700800 462372 700806
rect 462320 700742 462372 700748
rect 478524 700738 478552 703520
rect 478512 700732 478564 700738
rect 478512 700674 478564 700680
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 511000 700602 511028 703520
rect 510988 700596 511040 700602
rect 510988 700538 511040 700544
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 575860 700330 575888 703520
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 389824 696992 389876 696998
rect 389824 696934 389876 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 389732 536852 389784 536858
rect 389732 536794 389784 536800
rect 389640 524476 389692 524482
rect 389640 524418 389692 524424
rect 389548 484424 389600 484430
rect 389548 484366 389600 484372
rect 378810 477958 379284 477986
rect 384882 477958 384988 477986
rect 86224 477488 86276 477494
rect 86224 477430 86276 477436
rect 165620 477488 165672 477494
rect 165620 477430 165672 477436
rect 165632 476513 165660 477430
rect 165618 476504 165674 476513
rect 165618 476439 165674 476448
rect 165620 471980 165672 471986
rect 165620 471922 165672 471928
rect 165632 471345 165660 471922
rect 165618 471336 165674 471345
rect 165618 471271 165674 471280
rect 165620 469192 165672 469198
rect 165620 469134 165672 469140
rect 165632 468761 165660 469134
rect 165618 468752 165674 468761
rect 165618 468687 165674 468696
rect 4804 466404 4856 466410
rect 4804 466346 4856 466352
rect 165620 466404 165672 466410
rect 165620 466346 165672 466352
rect 165632 466177 165660 466346
rect 165618 466168 165674 466177
rect 165618 466103 165674 466112
rect 165620 463684 165672 463690
rect 165620 463626 165672 463632
rect 165632 463593 165660 463626
rect 165618 463584 165674 463593
rect 165618 463519 165674 463528
rect 165620 462324 165672 462330
rect 165620 462266 165672 462272
rect 165632 461009 165660 462266
rect 165618 461000 165674 461009
rect 165618 460935 165674 460944
rect 165620 459536 165672 459542
rect 165620 459478 165672 459484
rect 165632 458425 165660 459478
rect 165618 458416 165674 458425
rect 165618 458351 165674 458360
rect 165620 456748 165672 456754
rect 165620 456690 165672 456696
rect 165632 455841 165660 456690
rect 165618 455832 165674 455841
rect 165618 455767 165674 455776
rect 165620 454028 165672 454034
rect 165620 453970 165672 453976
rect 165632 453257 165660 453970
rect 165618 453248 165674 453257
rect 165618 453183 165674 453192
rect 4068 451240 4120 451246
rect 4068 451182 4120 451188
rect 165620 451240 165672 451246
rect 165620 451182 165672 451188
rect 165632 450673 165660 451182
rect 165618 450664 165674 450673
rect 165618 450599 165674 450608
rect 3514 449576 3570 449585
rect 3514 449511 3570 449520
rect 3424 430568 3476 430574
rect 3424 430510 3476 430516
rect 3528 427786 3556 449511
rect 165620 448520 165672 448526
rect 165620 448462 165672 448468
rect 165632 448089 165660 448462
rect 165618 448080 165674 448089
rect 165618 448015 165674 448024
rect 165620 445732 165672 445738
rect 165620 445674 165672 445680
rect 165632 445505 165660 445674
rect 165618 445496 165674 445505
rect 165618 445431 165674 445440
rect 165620 442944 165672 442950
rect 165618 442912 165620 442921
rect 165672 442912 165674 442921
rect 165618 442847 165674 442856
rect 165620 441584 165672 441590
rect 165620 441526 165672 441532
rect 165632 440337 165660 441526
rect 165618 440328 165674 440337
rect 165618 440263 165674 440272
rect 165620 438864 165672 438870
rect 165620 438806 165672 438812
rect 165632 437753 165660 438806
rect 165618 437744 165674 437753
rect 165618 437679 165674 437688
rect 3606 436656 3662 436665
rect 3606 436591 3662 436600
rect 3516 427780 3568 427786
rect 3516 427722 3568 427728
rect 3620 425066 3648 436591
rect 165620 436076 165672 436082
rect 165620 436018 165672 436024
rect 165632 435169 165660 436018
rect 165618 435160 165674 435169
rect 165618 435095 165674 435104
rect 389560 434217 389588 484366
rect 389652 442241 389680 524418
rect 389744 444825 389772 536794
rect 389836 476513 389864 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 389916 683188 389968 683194
rect 389916 683130 389968 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 389822 476504 389878 476513
rect 389822 476439 389878 476448
rect 389928 473929 389956 683130
rect 390008 670744 390060 670750
rect 580172 670744 580224 670750
rect 390008 670686 390060 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 389914 473920 389970 473929
rect 389914 473855 389970 473864
rect 390020 471209 390048 670686
rect 580170 670647 580226 670656
rect 580262 657384 580318 657393
rect 580262 657319 580318 657328
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 390100 643136 390152 643142
rect 390100 643078 390152 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 390006 471200 390062 471209
rect 390006 471135 390062 471144
rect 389824 470620 389876 470626
rect 390112 470594 390140 643078
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 390192 630692 390244 630698
rect 390192 630634 390244 630640
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 389824 470562 389876 470568
rect 390020 470566 390140 470594
rect 389730 444816 389786 444825
rect 389730 444751 389786 444760
rect 389638 442232 389694 442241
rect 389638 442167 389694 442176
rect 389546 434208 389602 434217
rect 389546 434143 389602 434152
rect 165620 433288 165672 433294
rect 165620 433230 165672 433236
rect 165632 432585 165660 433230
rect 165618 432576 165674 432585
rect 165618 432511 165674 432520
rect 389836 431633 389864 470562
rect 390020 465905 390048 470566
rect 390100 469192 390152 469198
rect 390100 469134 390152 469140
rect 390112 468625 390140 469134
rect 390098 468616 390154 468625
rect 390098 468551 390154 468560
rect 390006 465896 390062 465905
rect 390006 465831 390062 465840
rect 390204 463321 390232 630634
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 390284 616888 390336 616894
rect 390284 616830 390336 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 390190 463312 390246 463321
rect 390190 463247 390246 463256
rect 390296 460737 390324 616830
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 390376 590708 390428 590714
rect 390376 590650 390428 590656
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 390282 460728 390338 460737
rect 390282 460663 390338 460672
rect 390192 458176 390244 458182
rect 390192 458118 390244 458124
rect 390204 458017 390232 458118
rect 390190 458008 390246 458017
rect 390190 457943 390246 457952
rect 389916 456816 389968 456822
rect 389916 456758 389968 456764
rect 389822 431624 389878 431633
rect 389822 431559 389878 431568
rect 389824 430636 389876 430642
rect 389824 430578 389876 430584
rect 165620 430568 165672 430574
rect 165620 430510 165672 430516
rect 165632 429865 165660 430510
rect 165618 429856 165674 429865
rect 165618 429791 165674 429800
rect 165620 427780 165672 427786
rect 165620 427722 165672 427728
rect 165632 427281 165660 427722
rect 165618 427272 165674 427281
rect 165618 427207 165674 427216
rect 3608 425060 3660 425066
rect 3608 425002 3660 425008
rect 165620 425060 165672 425066
rect 165620 425002 165672 425008
rect 165632 424697 165660 425002
rect 165618 424688 165674 424697
rect 165618 424623 165674 424632
rect 389836 423745 389864 430578
rect 389928 429049 389956 456758
rect 390388 455433 390416 590650
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 390468 576904 390520 576910
rect 390468 576846 390520 576852
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 390374 455424 390430 455433
rect 390374 455359 390430 455368
rect 390480 452713 390508 576846
rect 579618 537840 579674 537849
rect 579618 537775 579674 537784
rect 579632 536858 579660 537775
rect 579620 536852 579672 536858
rect 579620 536794 579672 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580276 469198 580304 657319
rect 580354 604208 580410 604217
rect 580354 604143 580410 604152
rect 580264 469192 580316 469198
rect 580264 469134 580316 469140
rect 580368 458182 580396 604143
rect 580446 564360 580502 564369
rect 580446 564295 580502 564304
rect 580356 458176 580408 458182
rect 579802 458144 579858 458153
rect 580356 458118 580408 458124
rect 579802 458079 579858 458088
rect 579816 456822 579844 458079
rect 579804 456816 579856 456822
rect 579804 456758 579856 456764
rect 390466 452704 390522 452713
rect 390466 452639 390522 452648
rect 580460 451246 580488 564295
rect 580538 551168 580594 551177
rect 580538 551103 580594 551112
rect 390192 451240 390244 451246
rect 390192 451182 390244 451188
rect 580448 451240 580500 451246
rect 580448 451182 580500 451188
rect 390204 450129 390232 451182
rect 390190 450120 390246 450129
rect 390190 450055 390246 450064
rect 580552 448526 580580 551103
rect 580630 511320 580686 511329
rect 580630 511255 580686 511264
rect 390192 448520 390244 448526
rect 390192 448462 390244 448468
rect 580540 448520 580592 448526
rect 580540 448462 580592 448468
rect 390204 447545 390232 448462
rect 390190 447536 390246 447545
rect 390190 447471 390246 447480
rect 580170 444816 580226 444825
rect 580170 444751 580226 444760
rect 580184 444446 580212 444751
rect 390008 444440 390060 444446
rect 390008 444382 390060 444388
rect 580172 444440 580224 444446
rect 580172 444382 580224 444388
rect 389914 429040 389970 429049
rect 389914 428975 389970 428984
rect 390020 426329 390048 444382
rect 580644 440230 580672 511255
rect 580722 497992 580778 498001
rect 580722 497927 580778 497936
rect 390192 440224 390244 440230
rect 390192 440166 390244 440172
rect 580632 440224 580684 440230
rect 580632 440166 580684 440172
rect 390204 439521 390232 440166
rect 390190 439512 390246 439521
rect 390190 439447 390246 439456
rect 580736 437442 580764 497927
rect 390284 437436 390336 437442
rect 390284 437378 390336 437384
rect 580724 437436 580776 437442
rect 580724 437378 580776 437384
rect 390296 436937 390324 437378
rect 390282 436928 390338 436937
rect 390282 436863 390338 436872
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 390006 426320 390062 426329
rect 390006 426255 390062 426264
rect 389822 423736 389878 423745
rect 389822 423671 389878 423680
rect 3790 423600 3846 423609
rect 3790 423535 3846 423544
rect 3804 422278 3832 423535
rect 3792 422272 3844 422278
rect 3792 422214 3844 422220
rect 165620 422272 165672 422278
rect 165620 422214 165672 422220
rect 165632 422113 165660 422214
rect 165618 422104 165674 422113
rect 165618 422039 165674 422048
rect 390098 421016 390154 421025
rect 390098 420951 390154 420960
rect 165618 419520 165674 419529
rect 390112 419490 390140 420951
rect 165618 419455 165674 419464
rect 390100 419484 390152 419490
rect 165632 418198 165660 419455
rect 390100 419426 390152 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 390190 418432 390246 418441
rect 390190 418367 390246 418376
rect 3424 418192 3476 418198
rect 3424 418134 3476 418140
rect 165620 418192 165672 418198
rect 165620 418134 165672 418140
rect 3436 410553 3464 418134
rect 165618 416936 165674 416945
rect 165618 416871 165674 416880
rect 165632 416838 165660 416871
rect 3792 416832 3844 416838
rect 3792 416774 3844 416780
rect 165620 416832 165672 416838
rect 165620 416774 165672 416780
rect 3700 414044 3752 414050
rect 3700 413986 3752 413992
rect 3608 411324 3660 411330
rect 3608 411266 3660 411272
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3516 408536 3568 408542
rect 3516 408478 3568 408484
rect 3424 405748 3476 405754
rect 3424 405690 3476 405696
rect 3148 398880 3200 398886
rect 3148 398822 3200 398828
rect 3056 332580 3108 332586
rect 3056 332522 3108 332528
rect 3068 332353 3096 332522
rect 3054 332344 3110 332353
rect 3054 332279 3110 332288
rect 3056 320136 3108 320142
rect 3056 320078 3108 320084
rect 3068 319297 3096 320078
rect 3054 319288 3110 319297
rect 3054 319223 3110 319232
rect 3160 306241 3188 398822
rect 3240 385076 3292 385082
rect 3240 385018 3292 385024
rect 3146 306232 3202 306241
rect 3146 306167 3202 306176
rect 2780 293616 2832 293622
rect 2780 293558 2832 293564
rect 2792 293185 2820 293558
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3252 241097 3280 385018
rect 3332 376780 3384 376786
rect 3332 376722 3384 376728
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3240 229084 3292 229090
rect 3240 229026 3292 229032
rect 3252 228041 3280 229026
rect 3238 228032 3294 228041
rect 3238 227967 3294 227976
rect 3240 215280 3292 215286
rect 3240 215222 3292 215228
rect 3252 214985 3280 215222
rect 3238 214976 3294 214985
rect 3238 214911 3294 214920
rect 3344 201929 3372 376722
rect 3436 345409 3464 405690
rect 3528 358465 3556 408478
rect 3620 371385 3648 411266
rect 3712 384441 3740 413986
rect 3804 397497 3832 416774
rect 390098 415848 390154 415857
rect 390098 415783 390154 415792
rect 165618 414352 165674 414361
rect 165618 414287 165674 414296
rect 165632 414050 165660 414287
rect 165620 414044 165672 414050
rect 165620 413986 165672 413992
rect 390006 413128 390062 413137
rect 390006 413063 390062 413072
rect 165618 411768 165674 411777
rect 165618 411703 165674 411712
rect 165632 411330 165660 411703
rect 165620 411324 165672 411330
rect 165620 411266 165672 411272
rect 389914 410544 389970 410553
rect 389914 410479 389970 410488
rect 165618 409184 165674 409193
rect 165618 409119 165674 409128
rect 165632 408542 165660 409119
rect 165620 408536 165672 408542
rect 165620 408478 165672 408484
rect 389822 407824 389878 407833
rect 389822 407759 389878 407768
rect 165618 406600 165674 406609
rect 165618 406535 165674 406544
rect 165632 405754 165660 406535
rect 165620 405748 165672 405754
rect 165620 405690 165672 405696
rect 389178 405240 389234 405249
rect 389178 405175 389234 405184
rect 389192 404530 389220 405175
rect 389180 404524 389232 404530
rect 389180 404466 389232 404472
rect 166906 404016 166962 404025
rect 166906 403951 166962 403960
rect 166814 401432 166870 401441
rect 166814 401367 166870 401376
rect 165620 398880 165672 398886
rect 165618 398848 165620 398857
rect 165672 398848 165674 398857
rect 165618 398783 165674 398792
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 165618 396264 165674 396273
rect 165618 396199 165674 396208
rect 165632 396098 165660 396199
rect 4804 396092 4856 396098
rect 4804 396034 4856 396040
rect 165620 396092 165672 396098
rect 165620 396034 165672 396040
rect 3698 384432 3754 384441
rect 3698 384367 3754 384376
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 4068 369912 4120 369918
rect 4068 369854 4120 369860
rect 3976 364404 4028 364410
rect 3976 364346 4028 364352
rect 3884 358828 3936 358834
rect 3884 358770 3936 358776
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 3792 356108 3844 356114
rect 3792 356050 3844 356056
rect 3700 351960 3752 351966
rect 3700 351902 3752 351908
rect 3608 346452 3660 346458
rect 3608 346394 3660 346400
rect 3422 345400 3478 345409
rect 3422 345335 3478 345344
rect 3516 343664 3568 343670
rect 3516 343606 3568 343612
rect 3424 340944 3476 340950
rect 3424 340886 3476 340892
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3332 176656 3384 176662
rect 3332 176598 3384 176604
rect 3344 175953 3372 176598
rect 3330 175944 3386 175953
rect 3330 175879 3386 175888
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3148 124160 3200 124166
rect 3148 124102 3200 124108
rect 3160 123729 3188 124102
rect 3146 123720 3202 123729
rect 3146 123655 3202 123664
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 2872 59356 2924 59362
rect 2872 59298 2924 59304
rect 2884 58585 2912 59298
rect 2870 58576 2926 58585
rect 2870 58511 2926 58520
rect 3436 19417 3464 340886
rect 3528 32473 3556 343606
rect 3620 45529 3648 346394
rect 3712 71641 3740 351902
rect 3804 97617 3832 356050
rect 3896 110673 3924 358770
rect 3988 136785 4016 364346
rect 4080 162897 4108 369854
rect 4816 293622 4844 396034
rect 166722 393680 166778 393689
rect 166722 393615 166778 393624
rect 166630 391096 166686 391105
rect 166630 391031 166686 391040
rect 165618 388512 165674 388521
rect 165618 388447 165674 388456
rect 165632 387870 165660 388447
rect 21456 387864 21508 387870
rect 21456 387806 21508 387812
rect 165620 387864 165672 387870
rect 165620 387806 165672 387812
rect 10324 375420 10376 375426
rect 10324 375362 10376 375368
rect 7564 336048 7616 336054
rect 7564 335990 7616 335996
rect 4804 293616 4856 293622
rect 4804 293558 4856 293564
rect 4066 162888 4122 162897
rect 4066 162823 4122 162832
rect 3974 136776 4030 136785
rect 3974 136711 4030 136720
rect 3882 110664 3938 110673
rect 3882 110599 3938 110608
rect 3790 97608 3846 97617
rect 3790 97543 3846 97552
rect 3698 71632 3754 71641
rect 3698 71567 3754 71576
rect 3606 45520 3662 45529
rect 3606 45455 3662 45464
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 7576 4146 7604 335990
rect 10336 189038 10364 375362
rect 11704 354748 11756 354754
rect 11704 354690 11756 354696
rect 10324 189032 10376 189038
rect 10324 188974 10376 188980
rect 11716 85542 11744 354690
rect 18604 338156 18656 338162
rect 18604 338098 18656 338104
rect 17224 336116 17276 336122
rect 17224 336058 17276 336064
rect 15844 330540 15896 330546
rect 15844 330482 15896 330488
rect 14464 320884 14516 320890
rect 14464 320826 14516 320832
rect 11704 85536 11756 85542
rect 11704 85478 11756 85484
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 4082
rect 7668 480 7696 4966
rect 8772 480 8800 6190
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11150 3496 11206 3505
rect 11150 3431 11206 3440
rect 9956 3324 10008 3330
rect 9956 3266 10008 3272
rect 9968 480 9996 3266
rect 11164 480 11192 3431
rect 12360 480 12388 5034
rect 14476 3534 14504 320826
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 13556 480 13584 3470
rect 14752 480 14780 3878
rect 15856 3330 15884 330482
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15844 3324 15896 3330
rect 15844 3266 15896 3272
rect 15948 480 15976 3402
rect 17052 480 17080 6258
rect 17236 3942 17264 336058
rect 18616 6866 18644 338098
rect 21468 255270 21496 387806
rect 165618 385928 165674 385937
rect 165618 385863 165674 385872
rect 165632 385082 165660 385863
rect 165620 385076 165672 385082
rect 165620 385018 165672 385024
rect 166538 383208 166594 383217
rect 166538 383143 166594 383152
rect 166446 380624 166502 380633
rect 166446 380559 166502 380568
rect 165618 378040 165674 378049
rect 165618 377975 165674 377984
rect 165632 376786 165660 377975
rect 165620 376780 165672 376786
rect 165620 376722 165672 376728
rect 165618 375456 165674 375465
rect 165618 375391 165620 375400
rect 165672 375391 165674 375400
rect 165620 375362 165672 375368
rect 166354 372872 166410 372881
rect 166354 372807 166410 372816
rect 165618 370288 165674 370297
rect 165618 370223 165674 370232
rect 165632 369918 165660 370223
rect 165620 369912 165672 369918
rect 165620 369854 165672 369860
rect 165618 367704 165674 367713
rect 165618 367639 165674 367648
rect 165632 367130 165660 367639
rect 28264 367124 28316 367130
rect 28264 367066 28316 367072
rect 165620 367124 165672 367130
rect 165620 367066 165672 367072
rect 22744 336184 22796 336190
rect 22744 336126 22796 336132
rect 21456 255264 21508 255270
rect 21456 255206 21508 255212
rect 21364 254584 21416 254590
rect 21364 254526 21416 254532
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 20626 3768 20682 3777
rect 20626 3703 20682 3712
rect 19430 3632 19486 3641
rect 19430 3567 19486 3576
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 480 18276 3470
rect 19444 480 19472 3567
rect 20640 480 20668 3703
rect 21376 3534 21404 254526
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21836 480 21864 6326
rect 22756 3466 22784 336126
rect 25504 334620 25556 334626
rect 25504 334562 25556 334568
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23032 480 23060 3130
rect 24228 480 24256 3470
rect 25332 480 25360 3538
rect 25516 3194 25544 334562
rect 28276 150414 28304 367066
rect 165618 365120 165674 365129
rect 165618 365055 165674 365064
rect 165632 364410 165660 365055
rect 165620 364404 165672 364410
rect 165620 364346 165672 364352
rect 166262 362536 166318 362545
rect 166262 362471 166318 362480
rect 165618 359952 165674 359961
rect 165618 359887 165674 359896
rect 165632 358834 165660 359887
rect 165620 358828 165672 358834
rect 165620 358770 165672 358776
rect 165618 357368 165674 357377
rect 165618 357303 165674 357312
rect 165632 356114 165660 357303
rect 165620 356108 165672 356114
rect 165620 356050 165672 356056
rect 165618 354784 165674 354793
rect 165618 354719 165620 354728
rect 165672 354719 165674 354728
rect 165620 354690 165672 354696
rect 165618 352200 165674 352209
rect 165618 352135 165674 352144
rect 165632 351966 165660 352135
rect 165620 351960 165672 351966
rect 165620 351902 165672 351908
rect 165618 349616 165674 349625
rect 165618 349551 165674 349560
rect 165632 349178 165660 349551
rect 29644 349172 29696 349178
rect 29644 349114 29696 349120
rect 165620 349172 165672 349178
rect 165620 349114 165672 349120
rect 28908 323604 28960 323610
rect 28908 323546 28960 323552
rect 28264 150408 28316 150414
rect 28264 150350 28316 150356
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 26528 480 26556 6394
rect 28920 3534 28948 323546
rect 29656 59362 29684 349114
rect 165618 347032 165674 347041
rect 165618 346967 165674 346976
rect 165632 346458 165660 346967
rect 165620 346452 165672 346458
rect 165620 346394 165672 346400
rect 165618 344448 165674 344457
rect 165618 344383 165674 344392
rect 165632 343670 165660 344383
rect 165620 343664 165672 343670
rect 165620 343606 165672 343612
rect 165618 341864 165674 341873
rect 165618 341799 165674 341808
rect 165632 340950 165660 341799
rect 165620 340944 165672 340950
rect 165620 340886 165672 340892
rect 165618 339280 165674 339289
rect 165618 339215 165674 339224
rect 165632 338162 165660 339215
rect 165620 338156 165672 338162
rect 165620 338098 165672 338104
rect 118608 336728 118660 336734
rect 118608 336670 118660 336676
rect 111708 336660 111760 336666
rect 111708 336602 111760 336608
rect 103428 336592 103480 336598
rect 103428 336534 103480 336540
rect 50344 336524 50396 336530
rect 50344 336466 50396 336472
rect 43444 336456 43496 336462
rect 43444 336398 43496 336404
rect 35164 336388 35216 336394
rect 35164 336330 35216 336336
rect 32404 336252 32456 336258
rect 32404 336194 32456 336200
rect 29644 59356 29696 59362
rect 29644 59298 29696 59304
rect 30104 6520 30156 6526
rect 30104 6462 30156 6468
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 27724 480 27752 3470
rect 28908 3324 28960 3330
rect 28908 3266 28960 3272
rect 28920 480 28948 3266
rect 30116 480 30144 6462
rect 32416 3602 32444 336194
rect 33784 324964 33836 324970
rect 33784 324906 33836 324912
rect 33600 6588 33652 6594
rect 33600 6530 33652 6536
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31312 480 31340 3130
rect 32404 2984 32456 2990
rect 32404 2926 32456 2932
rect 32416 480 32444 2926
rect 33612 480 33640 6530
rect 33796 3194 33824 324906
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 34808 480 34836 3538
rect 35176 3466 35204 336330
rect 36544 336320 36596 336326
rect 36544 336262 36596 336268
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 36004 480 36032 3334
rect 36556 2990 36584 336262
rect 39304 326392 39356 326398
rect 39304 326334 39356 326340
rect 37188 6656 37240 6662
rect 37188 6598 37240 6604
rect 36544 2984 36596 2990
rect 36544 2926 36596 2932
rect 37200 480 37228 6598
rect 39316 3602 39344 326334
rect 40684 301504 40736 301510
rect 40684 301446 40736 301452
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 39580 3528 39632 3534
rect 39580 3470 39632 3476
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 39592 480 39620 3470
rect 40696 3194 40724 301446
rect 40776 6724 40828 6730
rect 40776 6666 40828 6672
rect 40684 3188 40736 3194
rect 40684 3130 40736 3136
rect 40788 3074 40816 6666
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 40696 3046 40816 3074
rect 41880 3052 41932 3058
rect 40696 480 40724 3046
rect 41880 2994 41932 3000
rect 41892 480 41920 2994
rect 43088 480 43116 3538
rect 43456 3534 43484 336398
rect 46204 327752 46256 327758
rect 46204 327694 46256 327700
rect 44272 6792 44324 6798
rect 44272 6734 44324 6740
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 44284 480 44312 6734
rect 45468 3868 45520 3874
rect 45468 3810 45520 3816
rect 45480 480 45508 3810
rect 46216 3058 46244 327694
rect 47584 302932 47636 302938
rect 47584 302874 47636 302880
rect 47596 3874 47624 302874
rect 48964 6860 49016 6866
rect 48964 6802 49016 6808
rect 47860 5160 47912 5166
rect 47860 5102 47912 5108
rect 47584 3868 47636 3874
rect 47584 3810 47636 3816
rect 46664 3188 46716 3194
rect 46664 3130 46716 3136
rect 46204 3052 46256 3058
rect 46204 2994 46256 3000
rect 46676 480 46704 3130
rect 47872 480 47900 5102
rect 48976 480 49004 6802
rect 50160 3392 50212 3398
rect 50160 3334 50212 3340
rect 50172 480 50200 3334
rect 50356 3194 50384 336466
rect 51724 322244 51776 322250
rect 51724 322186 51776 322192
rect 51356 5228 51408 5234
rect 51356 5170 51408 5176
rect 50344 3188 50396 3194
rect 50344 3130 50396 3136
rect 51368 480 51396 5170
rect 51736 3398 51764 322186
rect 88248 312588 88300 312594
rect 88248 312530 88300 312536
rect 81348 28280 81400 28286
rect 81348 28222 81400 28228
rect 79692 7948 79744 7954
rect 79692 7890 79744 7896
rect 77392 7880 77444 7886
rect 77392 7822 77444 7828
rect 73804 7812 73856 7818
rect 73804 7754 73856 7760
rect 70308 7744 70360 7750
rect 70308 7686 70360 7692
rect 66720 7676 66772 7682
rect 66720 7618 66772 7624
rect 63224 7608 63276 7614
rect 63224 7550 63276 7556
rect 52552 6112 52604 6118
rect 52552 6054 52604 6060
rect 51724 3392 51776 3398
rect 51724 3334 51776 3340
rect 52564 480 52592 6054
rect 56048 6044 56100 6050
rect 56048 5986 56100 5992
rect 54944 5296 54996 5302
rect 54944 5238 54996 5244
rect 53748 3664 53800 3670
rect 53748 3606 53800 3612
rect 53760 480 53788 3606
rect 54956 480 54984 5238
rect 56060 480 56088 5986
rect 59636 5976 59688 5982
rect 59636 5918 59688 5924
rect 58440 5364 58492 5370
rect 58440 5306 58492 5312
rect 57244 3732 57296 3738
rect 57244 3674 57296 3680
rect 57256 480 57284 3674
rect 58452 480 58480 5306
rect 59648 480 59676 5918
rect 62028 5432 62080 5438
rect 62028 5374 62080 5380
rect 60832 3800 60884 3806
rect 60832 3742 60884 3748
rect 60844 480 60872 3742
rect 62040 480 62068 5374
rect 63236 480 63264 7550
rect 65524 5500 65576 5506
rect 65524 5442 65576 5448
rect 64328 3868 64380 3874
rect 64328 3810 64380 3816
rect 64340 480 64368 3810
rect 65536 480 65564 5442
rect 66732 480 66760 7618
rect 69112 4752 69164 4758
rect 69112 4694 69164 4700
rect 67916 3936 67968 3942
rect 67916 3878 67968 3884
rect 67928 480 67956 3878
rect 69124 480 69152 4694
rect 70320 480 70348 7686
rect 72608 4684 72660 4690
rect 72608 4626 72660 4632
rect 71504 4004 71556 4010
rect 71504 3946 71556 3952
rect 71516 480 71544 3946
rect 72620 480 72648 4626
rect 73816 480 73844 7754
rect 76196 5908 76248 5914
rect 76196 5850 76248 5856
rect 75000 4072 75052 4078
rect 75000 4014 75052 4020
rect 75012 480 75040 4014
rect 76208 480 76236 5850
rect 77404 480 77432 7822
rect 78588 4140 78640 4146
rect 78588 4082 78640 4088
rect 78600 480 78628 4082
rect 79704 480 79732 7890
rect 81360 3398 81388 28222
rect 84476 8968 84528 8974
rect 84476 8910 84528 8916
rect 83280 8016 83332 8022
rect 83280 7958 83332 7964
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 82084 3392 82136 3398
rect 82084 3334 82136 3340
rect 80900 480 80928 3334
rect 82096 480 82124 3334
rect 83292 480 83320 7958
rect 84488 480 84516 8910
rect 86868 8084 86920 8090
rect 86868 8026 86920 8032
rect 85672 3188 85724 3194
rect 85672 3130 85724 3136
rect 85684 480 85712 3130
rect 86880 480 86908 8026
rect 88260 6914 88288 312530
rect 95148 311160 95200 311166
rect 95148 311102 95200 311108
rect 92388 10328 92440 10334
rect 92388 10270 92440 10276
rect 90364 8152 90416 8158
rect 90364 8094 90416 8100
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 8094
rect 92400 3330 92428 10270
rect 93952 8220 94004 8226
rect 93952 8162 94004 8168
rect 91560 3324 91612 3330
rect 91560 3266 91612 3272
rect 92388 3324 92440 3330
rect 92388 3266 92440 3272
rect 91572 480 91600 3266
rect 92756 3188 92808 3194
rect 92756 3130 92808 3136
rect 92768 480 92796 3130
rect 93964 480 93992 8162
rect 95160 480 95188 311102
rect 99288 307080 99340 307086
rect 99288 307022 99340 307028
rect 97448 8288 97500 8294
rect 97448 8230 97500 8236
rect 96252 3052 96304 3058
rect 96252 2994 96304 3000
rect 96264 480 96292 2994
rect 97460 480 97488 8230
rect 99300 3126 99328 307022
rect 103244 11756 103296 11762
rect 103244 11698 103296 11704
rect 101036 7540 101088 7546
rect 101036 7482 101088 7488
rect 98644 3120 98696 3126
rect 98644 3062 98696 3068
rect 99288 3120 99340 3126
rect 99288 3062 99340 3068
rect 98656 480 98684 3062
rect 99840 2984 99892 2990
rect 99840 2926 99892 2932
rect 99852 480 99880 2926
rect 101048 480 101076 7482
rect 103256 3126 103284 11698
rect 103440 3482 103468 336534
rect 106188 309800 106240 309806
rect 106188 309742 106240 309748
rect 104532 7472 104584 7478
rect 104532 7414 104584 7420
rect 103348 3454 103468 3482
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 103244 3120 103296 3126
rect 103244 3062 103296 3068
rect 102244 480 102272 3062
rect 103348 480 103376 3454
rect 104544 480 104572 7414
rect 106200 3126 106228 309742
rect 110328 21412 110380 21418
rect 110328 21354 110380 21360
rect 108120 7404 108172 7410
rect 108120 7346 108172 7352
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 105740 480 105768 3062
rect 106924 2848 106976 2854
rect 106924 2790 106976 2796
rect 106936 480 106964 2790
rect 108132 480 108160 7346
rect 110340 3126 110368 21354
rect 111616 7336 111668 7342
rect 111616 7278 111668 7284
rect 109316 3120 109368 3126
rect 109316 3062 109368 3068
rect 110328 3120 110380 3126
rect 110328 3062 110380 3068
rect 109328 480 109356 3062
rect 110512 2916 110564 2922
rect 110512 2858 110564 2864
rect 110524 480 110552 2858
rect 111628 480 111656 7278
rect 111720 2922 111748 336602
rect 113088 329112 113140 329118
rect 113088 329054 113140 329060
rect 113100 6914 113128 329054
rect 117228 308440 117280 308446
rect 117228 308382 117280 308388
rect 115204 7268 115256 7274
rect 115204 7210 115256 7216
rect 112824 6886 113128 6914
rect 111708 2916 111760 2922
rect 111708 2858 111760 2864
rect 112824 480 112852 6886
rect 114008 2848 114060 2854
rect 114008 2790 114060 2796
rect 114020 480 114048 2790
rect 115216 480 115244 7210
rect 117240 2922 117268 308382
rect 118620 2922 118648 336670
rect 121368 335980 121420 335986
rect 121368 335922 121420 335928
rect 119988 305652 120040 305658
rect 119988 305594 120040 305600
rect 118792 7200 118844 7206
rect 118792 7142 118844 7148
rect 116400 2916 116452 2922
rect 116400 2858 116452 2864
rect 117228 2916 117280 2922
rect 117228 2858 117280 2864
rect 117596 2916 117648 2922
rect 117596 2858 117648 2864
rect 118608 2916 118660 2922
rect 118608 2858 118660 2864
rect 116412 480 116440 2858
rect 117608 480 117636 2858
rect 118804 480 118832 7142
rect 120000 6914 120028 305594
rect 121380 6914 121408 335922
rect 126888 334688 126940 334694
rect 126888 334630 126940 334636
rect 124128 304292 124180 304298
rect 124128 304234 124180 304240
rect 122288 7132 122340 7138
rect 122288 7074 122340 7080
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122300 480 122328 7074
rect 124140 2922 124168 304234
rect 126900 2922 126928 334630
rect 161388 333328 161440 333334
rect 161388 333270 161440 333276
rect 135168 333260 135220 333266
rect 135168 333202 135220 333208
rect 133788 329180 133840 329186
rect 133788 329122 133840 329128
rect 129648 327820 129700 327826
rect 129648 327762 129700 327768
rect 129660 6914 129688 327762
rect 131028 322312 131080 322318
rect 131028 322254 131080 322260
rect 129384 6886 129688 6914
rect 128176 5840 128228 5846
rect 128176 5782 128228 5788
rect 126980 4616 127032 4622
rect 126980 4558 127032 4564
rect 123484 2916 123536 2922
rect 123484 2858 123536 2864
rect 124128 2916 124180 2922
rect 124128 2858 124180 2864
rect 124680 2916 124732 2922
rect 124680 2858 124732 2864
rect 125968 2916 126020 2922
rect 125968 2858 126020 2864
rect 126888 2916 126940 2922
rect 126888 2858 126940 2864
rect 123496 480 123524 2858
rect 124692 480 124720 2858
rect 125980 2802 126008 2858
rect 125888 2774 126008 2802
rect 125888 480 125916 2774
rect 126992 480 127020 4558
rect 128188 480 128216 5782
rect 129384 480 129412 6886
rect 131040 2922 131068 322254
rect 132224 14476 132276 14482
rect 132224 14418 132276 14424
rect 132236 2922 132264 14418
rect 133800 6914 133828 329122
rect 135180 6914 135208 333202
rect 136548 331900 136600 331906
rect 136548 331842 136600 331848
rect 136456 22772 136508 22778
rect 136456 22714 136508 22720
rect 132972 6886 133828 6914
rect 134168 6886 135208 6914
rect 130568 2916 130620 2922
rect 130568 2858 130620 2864
rect 131028 2916 131080 2922
rect 131028 2858 131080 2864
rect 131764 2916 131816 2922
rect 131764 2858 131816 2864
rect 132224 2916 132276 2922
rect 132224 2858 132276 2864
rect 130580 480 130608 2858
rect 131776 480 131804 2858
rect 132972 480 133000 6886
rect 134168 480 134196 6886
rect 136468 4214 136496 22714
rect 135260 4208 135312 4214
rect 135260 4150 135312 4156
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 135272 480 135300 4150
rect 136560 1442 136588 331842
rect 155868 330608 155920 330614
rect 155868 330550 155920 330556
rect 140688 326460 140740 326466
rect 140688 326402 140740 326408
rect 137928 316736 137980 316742
rect 137928 316678 137980 316684
rect 137940 6914 137968 316678
rect 138848 13116 138900 13122
rect 138848 13058 138900 13064
rect 136468 1414 136588 1442
rect 137664 6886 137968 6914
rect 136468 480 136496 1414
rect 137664 480 137692 6886
rect 138860 480 138888 13058
rect 140700 6914 140728 326402
rect 144828 325032 144880 325038
rect 144828 324974 144880 324980
rect 142068 318096 142120 318102
rect 142068 318038 142120 318044
rect 142080 6914 142108 318038
rect 144736 315308 144788 315314
rect 144736 315250 144788 315256
rect 143448 220108 143500 220114
rect 143448 220050 143500 220056
rect 143460 6914 143488 220050
rect 140056 6886 140728 6914
rect 141252 6886 142108 6914
rect 142448 6886 143488 6914
rect 140056 480 140084 6886
rect 141252 480 141280 6886
rect 142448 480 142476 6886
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 144748 480 144776 315250
rect 144840 4214 144868 324974
rect 147588 323672 147640 323678
rect 147588 323614 147640 323620
rect 146208 24132 146260 24138
rect 146208 24074 146260 24080
rect 146220 6914 146248 24074
rect 147600 6914 147628 323614
rect 153108 319456 153160 319462
rect 153108 319398 153160 319404
rect 148968 313948 149020 313954
rect 148968 313890 149020 313896
rect 148980 6914 149008 313890
rect 153016 221468 153068 221474
rect 153016 221410 153068 221416
rect 150348 25560 150400 25566
rect 150348 25502 150400 25508
rect 150360 6914 150388 25502
rect 145944 6886 146248 6914
rect 147140 6886 147628 6914
rect 148336 6886 149008 6914
rect 149532 6886 150388 6914
rect 144828 4208 144880 4214
rect 144828 4150 144880 4156
rect 145944 480 145972 6886
rect 147140 480 147168 6886
rect 148336 480 148364 6886
rect 149532 480 149560 6886
rect 150624 4548 150676 4554
rect 150624 4490 150676 4496
rect 150636 480 150664 4490
rect 151820 4208 151872 4214
rect 151820 4150 151872 4156
rect 151832 480 151860 4150
rect 153028 480 153056 221410
rect 153120 4214 153148 319398
rect 155880 6914 155908 330550
rect 157248 26920 157300 26926
rect 157248 26862 157300 26868
rect 157260 6914 157288 26862
rect 160100 7064 160152 7070
rect 160100 7006 160152 7012
rect 155420 6886 155908 6914
rect 156616 6886 157288 6914
rect 154212 4480 154264 4486
rect 154212 4422 154264 4428
rect 153108 4208 153160 4214
rect 153108 4150 153160 4156
rect 154224 480 154252 4422
rect 155420 480 155448 6886
rect 156616 480 156644 6886
rect 158904 5772 158956 5778
rect 158904 5714 158956 5720
rect 157800 4412 157852 4418
rect 157800 4354 157852 4360
rect 157812 480 157840 4354
rect 158916 480 158944 5714
rect 160112 480 160140 7006
rect 161400 6914 161428 333270
rect 165528 330676 165580 330682
rect 165528 330618 165580 330624
rect 165540 6914 165568 330618
rect 166276 124166 166304 362471
rect 166368 176662 166396 372807
rect 166460 215286 166488 380559
rect 166552 229090 166580 383143
rect 166644 267714 166672 391031
rect 166736 280158 166764 393615
rect 166828 320142 166856 401367
rect 166920 332586 166948 403951
rect 389178 402520 389234 402529
rect 389178 402455 389234 402464
rect 389086 341320 389142 341329
rect 389086 341255 389142 341264
rect 389100 340950 389128 341255
rect 389088 340944 389140 340950
rect 389088 340886 389140 340892
rect 389086 338736 389142 338745
rect 389086 338671 389142 338680
rect 389100 338162 389128 338671
rect 389088 338156 389140 338162
rect 389088 338098 389140 338104
rect 167748 338014 168222 338042
rect 168484 338014 168590 338042
rect 168760 338014 169050 338042
rect 169128 338014 169510 338042
rect 166908 332580 166960 332586
rect 166908 332522 166960 332528
rect 166816 320136 166868 320142
rect 166816 320078 166868 320084
rect 167748 316034 167776 338014
rect 168380 336796 168432 336802
rect 168380 336738 168432 336744
rect 167012 316006 167776 316034
rect 166724 280152 166776 280158
rect 166724 280094 166776 280100
rect 166632 267708 166684 267714
rect 166632 267650 166684 267656
rect 166540 229084 166592 229090
rect 166540 229026 166592 229032
rect 166448 215280 166500 215286
rect 166448 215222 166500 215228
rect 166356 176656 166408 176662
rect 166356 176598 166408 176604
rect 166264 124160 166316 124166
rect 166264 124102 166316 124108
rect 161308 6886 161428 6914
rect 164896 6886 165568 6914
rect 161308 480 161336 6886
rect 163688 5704 163740 5710
rect 163688 5646 163740 5652
rect 162492 4344 162544 4350
rect 162492 4286 162544 4292
rect 162504 480 162532 4286
rect 163700 480 163728 5646
rect 164896 480 164924 6886
rect 167012 4894 167040 316006
rect 167184 5636 167236 5642
rect 167184 5578 167236 5584
rect 167000 4888 167052 4894
rect 167000 4830 167052 4836
rect 166080 4276 166132 4282
rect 166080 4218 166132 4224
rect 166092 480 166120 4218
rect 167196 480 167224 5578
rect 168392 4962 168420 336738
rect 168380 4956 168432 4962
rect 168380 4898 168432 4904
rect 168484 4826 168512 338014
rect 168760 336802 168788 338014
rect 168748 336796 168800 336802
rect 168748 336738 168800 336744
rect 169128 316034 169156 338014
rect 169852 330472 169904 330478
rect 169852 330414 169904 330420
rect 168576 316006 169156 316034
rect 168576 6186 168604 316006
rect 169576 15904 169628 15910
rect 169576 15846 169628 15852
rect 168656 9036 168708 9042
rect 168656 8978 168708 8984
rect 168564 6180 168616 6186
rect 168564 6122 168616 6128
rect 168472 4820 168524 4826
rect 168472 4762 168524 4768
rect 168668 3482 168696 8978
rect 168392 3454 168696 3482
rect 168392 480 168420 3454
rect 169588 480 169616 15846
rect 169864 5030 169892 330414
rect 169852 5024 169904 5030
rect 169852 4966 169904 4972
rect 169956 3369 169984 338028
rect 170416 336054 170444 338028
rect 170600 338014 170890 338042
rect 170404 336048 170456 336054
rect 170404 335990 170456 335996
rect 170600 330478 170628 338014
rect 170588 330472 170640 330478
rect 170588 330414 170640 330420
rect 171244 6254 171272 338028
rect 171704 330546 171732 338028
rect 171796 338014 172178 338042
rect 172638 338014 172744 338042
rect 171692 330540 171744 330546
rect 171692 330482 171744 330488
rect 171796 316034 171824 338014
rect 172612 330540 172664 330546
rect 172612 330482 172664 330488
rect 172624 320890 172652 330482
rect 172612 320884 172664 320890
rect 172612 320826 172664 320832
rect 171336 316006 171824 316034
rect 171232 6248 171284 6254
rect 171232 6190 171284 6196
rect 170772 6180 170824 6186
rect 170772 6122 170824 6128
rect 169942 3360 169998 3369
rect 169942 3295 169998 3304
rect 170784 480 170812 6122
rect 171336 3505 171364 316006
rect 172428 10396 172480 10402
rect 172428 10338 172480 10344
rect 172440 3534 172468 10338
rect 172716 5098 172744 338014
rect 172808 338014 173098 338042
rect 172808 330546 172836 338014
rect 173544 336122 173572 338028
rect 173912 336190 173940 338028
rect 174096 338014 174386 338042
rect 174464 338014 174846 338042
rect 175306 338014 175412 338042
rect 173900 336184 173952 336190
rect 173900 336126 173952 336132
rect 173532 336116 173584 336122
rect 173532 336058 173584 336064
rect 173164 336048 173216 336054
rect 173164 335990 173216 335996
rect 172796 330540 172848 330546
rect 172796 330482 172848 330488
rect 173176 8974 173204 335990
rect 173992 330540 174044 330546
rect 173992 330482 174044 330488
rect 174004 254590 174032 330482
rect 173992 254584 174044 254590
rect 173992 254526 174044 254532
rect 173808 17264 173860 17270
rect 173808 17206 173860 17212
rect 173164 8968 173216 8974
rect 173164 8910 173216 8916
rect 172704 5092 172756 5098
rect 172704 5034 172756 5040
rect 173820 3534 173848 17206
rect 174096 6322 174124 338014
rect 174464 330546 174492 338014
rect 174452 330540 174504 330546
rect 174452 330482 174504 330488
rect 174084 6316 174136 6322
rect 174084 6258 174136 6264
rect 174268 6248 174320 6254
rect 174268 6190 174320 6196
rect 171968 3528 172020 3534
rect 171322 3496 171378 3505
rect 171968 3470 172020 3476
rect 172428 3528 172480 3534
rect 172428 3470 172480 3476
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 173808 3528 173860 3534
rect 173808 3470 173860 3476
rect 171322 3431 171378 3440
rect 171980 480 172008 3470
rect 173176 480 173204 3470
rect 174280 480 174308 6190
rect 175384 3641 175412 338014
rect 175568 338014 175766 338042
rect 175936 338014 176226 338042
rect 175464 330540 175516 330546
rect 175464 330482 175516 330488
rect 175476 6390 175504 330482
rect 175464 6384 175516 6390
rect 175464 6326 175516 6332
rect 175568 3777 175596 338014
rect 175936 330546 175964 338014
rect 176580 334626 176608 338028
rect 177040 336394 177068 338028
rect 177132 338014 177514 338042
rect 177592 338014 177974 338042
rect 178236 338014 178434 338042
rect 178512 338014 178894 338042
rect 179064 338014 179354 338042
rect 179524 338014 179722 338042
rect 177028 336388 177080 336394
rect 177028 336330 177080 336336
rect 177132 336258 177160 338014
rect 177592 336682 177620 338014
rect 177224 336654 177620 336682
rect 177120 336252 177172 336258
rect 177120 336194 177172 336200
rect 176568 334620 176620 334626
rect 176568 334562 176620 334568
rect 175924 330540 175976 330546
rect 175924 330482 175976 330488
rect 177224 316034 177252 336654
rect 177304 336116 177356 336122
rect 177304 336058 177356 336064
rect 176764 316006 177252 316034
rect 176568 11824 176620 11830
rect 176568 11766 176620 11772
rect 175554 3768 175610 3777
rect 175554 3703 175610 3712
rect 175370 3632 175426 3641
rect 175370 3567 175426 3576
rect 176580 3534 176608 11766
rect 176764 6458 176792 316006
rect 177316 10334 177344 336058
rect 178132 330540 178184 330546
rect 178132 330482 178184 330488
rect 177948 320884 178000 320890
rect 177948 320826 178000 320832
rect 177304 10328 177356 10334
rect 177304 10270 177356 10276
rect 176752 6452 176804 6458
rect 176752 6394 176804 6400
rect 177856 6316 177908 6322
rect 177856 6258 177908 6264
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 176568 3528 176620 3534
rect 176568 3470 176620 3476
rect 176660 3528 176712 3534
rect 176660 3470 176712 3476
rect 175476 480 175504 3470
rect 176672 480 176700 3470
rect 177868 480 177896 6258
rect 177960 3534 177988 320826
rect 178144 6526 178172 330482
rect 178236 323610 178264 338014
rect 178224 323604 178276 323610
rect 178224 323546 178276 323552
rect 178512 316034 178540 338014
rect 179064 330546 179092 338014
rect 179052 330540 179104 330546
rect 179052 330482 179104 330488
rect 179524 324970 179552 338014
rect 180168 336326 180196 338028
rect 180260 338014 180642 338042
rect 180996 338014 181102 338042
rect 181180 338014 181562 338042
rect 181640 338014 182022 338042
rect 182284 338014 182390 338042
rect 180156 336320 180208 336326
rect 180156 336262 180208 336268
rect 179512 324964 179564 324970
rect 179512 324906 179564 324912
rect 180260 316034 180288 338014
rect 180708 334620 180760 334626
rect 180708 334562 180760 334568
rect 178328 316006 178540 316034
rect 179616 316006 180288 316034
rect 178132 6520 178184 6526
rect 178132 6462 178184 6468
rect 178328 4214 178356 316006
rect 179052 13184 179104 13190
rect 179052 13126 179104 13132
rect 178316 4208 178368 4214
rect 178316 4150 178368 4156
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 179064 480 179092 13126
rect 179616 6594 179644 316006
rect 179604 6588 179656 6594
rect 179604 6530 179656 6536
rect 180720 3534 180748 334562
rect 180892 328976 180944 328982
rect 180892 328918 180944 328924
rect 180904 6662 180932 328918
rect 180996 326398 181024 338014
rect 180984 326392 181036 326398
rect 180984 326334 181036 326340
rect 181180 316034 181208 338014
rect 181640 328982 181668 338014
rect 181628 328976 181680 328982
rect 181628 328918 181680 328924
rect 181088 316006 181208 316034
rect 180892 6656 180944 6662
rect 180892 6598 180944 6604
rect 180248 3528 180300 3534
rect 180248 3470 180300 3476
rect 180708 3528 180760 3534
rect 180708 3470 180760 3476
rect 180260 480 180288 3470
rect 181088 3466 181116 316006
rect 182284 301510 182312 338014
rect 182836 336462 182864 338028
rect 182928 338014 183310 338042
rect 182824 336456 182876 336462
rect 182824 336398 182876 336404
rect 182928 316034 182956 338014
rect 183560 336252 183612 336258
rect 183560 336194 183612 336200
rect 182376 316006 182956 316034
rect 182272 301504 182324 301510
rect 182272 301446 182324 301452
rect 182376 6730 182404 316006
rect 183468 217320 183520 217326
rect 183468 217262 183520 217268
rect 182364 6724 182416 6730
rect 182364 6666 182416 6672
rect 181444 6384 181496 6390
rect 181444 6326 181496 6332
rect 181076 3460 181128 3466
rect 181076 3402 181128 3408
rect 181456 480 181484 6326
rect 183480 3534 183508 217262
rect 183572 3602 183600 336194
rect 183756 327758 183784 338028
rect 183848 338014 184230 338042
rect 184400 338014 184690 338042
rect 183848 336258 183876 338014
rect 183836 336252 183888 336258
rect 183836 336194 183888 336200
rect 183744 327752 183796 327758
rect 183744 327694 183796 327700
rect 184400 316034 184428 338014
rect 183664 316006 184428 316034
rect 183664 6798 183692 316006
rect 185044 302938 185072 338028
rect 185504 336530 185532 338028
rect 185596 338014 185978 338042
rect 185492 336524 185544 336530
rect 185492 336466 185544 336472
rect 185596 316034 185624 338014
rect 186320 326392 186372 326398
rect 186320 326334 186372 326340
rect 185136 316006 185624 316034
rect 185032 302932 185084 302938
rect 185032 302874 185084 302880
rect 184848 18624 184900 18630
rect 184848 18566 184900 18572
rect 183652 6792 183704 6798
rect 183652 6734 183704 6740
rect 183560 3596 183612 3602
rect 183560 3538 183612 3544
rect 184860 3534 184888 18566
rect 184940 6452 184992 6458
rect 184940 6394 184992 6400
rect 182548 3528 182600 3534
rect 182548 3470 182600 3476
rect 183468 3528 183520 3534
rect 183468 3470 183520 3476
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 182560 480 182588 3470
rect 183756 480 183784 3470
rect 184952 480 184980 6394
rect 185136 5166 185164 316006
rect 186136 8968 186188 8974
rect 186136 8910 186188 8916
rect 185124 5160 185176 5166
rect 185124 5102 185176 5108
rect 186148 480 186176 8910
rect 186332 5234 186360 326334
rect 186424 6866 186452 338028
rect 186516 338014 186898 338042
rect 186976 338014 187358 338042
rect 187726 338014 187924 338042
rect 186516 322250 186544 338014
rect 186976 326398 187004 338014
rect 187896 331226 187924 338014
rect 187988 338014 188186 338042
rect 188264 338014 188646 338042
rect 189106 338014 189304 338042
rect 187884 331220 187936 331226
rect 187884 331162 187936 331168
rect 187988 326618 188016 338014
rect 188068 331220 188120 331226
rect 188068 331162 188120 331168
rect 187712 326590 188016 326618
rect 186964 326392 187016 326398
rect 186964 326334 187016 326340
rect 186504 322244 186556 322250
rect 186504 322186 186556 322192
rect 187608 19984 187660 19990
rect 187608 19926 187660 19932
rect 187620 6914 187648 19926
rect 187344 6886 187648 6914
rect 186412 6860 186464 6866
rect 186412 6802 186464 6808
rect 186320 5228 186372 5234
rect 186320 5170 186372 5176
rect 187344 480 187372 6886
rect 187712 3670 187740 326590
rect 187792 326392 187844 326398
rect 187792 326334 187844 326340
rect 187804 5302 187832 326334
rect 188080 316034 188108 331162
rect 188264 326398 188292 338014
rect 189080 336796 189132 336802
rect 189080 336738 189132 336744
rect 188252 326392 188304 326398
rect 188252 326334 188304 326340
rect 187896 316006 188108 316034
rect 187896 6118 187924 316006
rect 188528 6520 188580 6526
rect 188528 6462 188580 6468
rect 187884 6112 187936 6118
rect 187884 6054 187936 6060
rect 187792 5296 187844 5302
rect 187792 5238 187844 5244
rect 187700 3664 187752 3670
rect 187700 3606 187752 3612
rect 188540 480 188568 6462
rect 189092 3466 189120 336738
rect 189172 326392 189224 326398
rect 189172 326334 189224 326340
rect 189184 5370 189212 326334
rect 189276 6050 189304 338014
rect 189368 338014 189566 338042
rect 189736 338014 190026 338042
rect 190486 338014 190592 338042
rect 189368 336802 189396 338014
rect 189356 336796 189408 336802
rect 189356 336738 189408 336744
rect 189736 326398 189764 338014
rect 189724 326392 189776 326398
rect 189724 326334 189776 326340
rect 190460 326392 190512 326398
rect 190460 326334 190512 326340
rect 190564 326346 190592 338014
rect 190748 338014 190854 338042
rect 191024 338014 191314 338042
rect 191392 338014 191774 338042
rect 191852 338014 192234 338042
rect 192312 338014 192694 338042
rect 192864 338014 193154 338042
rect 193232 338014 193522 338042
rect 193600 338014 193982 338042
rect 194152 338014 194442 338042
rect 194612 338014 194902 338042
rect 195072 338014 195362 338042
rect 195440 338014 195822 338042
rect 195992 338014 196190 338042
rect 196360 338014 196650 338042
rect 196728 338014 197110 338042
rect 197372 338014 197570 338042
rect 197648 338014 198030 338042
rect 198200 338014 198490 338042
rect 198858 338014 198964 338042
rect 190748 326398 190776 338014
rect 190736 326392 190788 326398
rect 189264 6044 189316 6050
rect 189264 5986 189316 5992
rect 189172 5364 189224 5370
rect 189172 5306 189224 5312
rect 189724 4820 189776 4826
rect 189724 4762 189776 4768
rect 189080 3460 189132 3466
rect 189080 3402 189132 3408
rect 189736 480 189764 4762
rect 190472 3874 190500 326334
rect 190564 326318 190684 326346
rect 190736 326334 190788 326340
rect 190552 326256 190604 326262
rect 190552 326198 190604 326204
rect 190564 5438 190592 326198
rect 190656 5982 190684 326318
rect 191024 326262 191052 338014
rect 191012 326256 191064 326262
rect 191012 326198 191064 326204
rect 191392 316034 191420 338014
rect 190748 316006 191420 316034
rect 190748 7614 190776 316006
rect 191748 14544 191800 14550
rect 191748 14486 191800 14492
rect 190736 7608 190788 7614
rect 190736 7550 190788 7556
rect 190644 5976 190696 5982
rect 190644 5918 190696 5924
rect 190552 5432 190604 5438
rect 190552 5374 190604 5380
rect 190460 3868 190512 3874
rect 190460 3810 190512 3816
rect 191760 3534 191788 14486
rect 191852 3806 191880 338014
rect 192312 335354 192340 338014
rect 191944 335326 192340 335354
rect 191944 5506 191972 335326
rect 192864 316034 192892 338014
rect 192036 316006 192892 316034
rect 192036 7682 192064 316006
rect 192024 7676 192076 7682
rect 192024 7618 192076 7624
rect 192024 6588 192076 6594
rect 192024 6530 192076 6536
rect 191932 5500 191984 5506
rect 191932 5442 191984 5448
rect 191840 3800 191892 3806
rect 191840 3742 191892 3748
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 191748 3528 191800 3534
rect 191748 3470 191800 3476
rect 190840 480 190868 3470
rect 192036 480 192064 6530
rect 193232 4978 193260 338014
rect 193600 335354 193628 338014
rect 193140 4950 193260 4978
rect 193324 335326 193628 335354
rect 193140 3942 193168 4950
rect 193220 4888 193272 4894
rect 193220 4830 193272 4836
rect 193128 3936 193180 3942
rect 193128 3878 193180 3884
rect 193232 480 193260 4830
rect 193324 4758 193352 335326
rect 194152 316034 194180 338014
rect 193416 316006 194180 316034
rect 193416 7750 193444 316006
rect 194416 21480 194468 21486
rect 194416 21422 194468 21428
rect 193404 7744 193456 7750
rect 193404 7686 193456 7692
rect 193312 4752 193364 4758
rect 193312 4694 193364 4700
rect 194428 480 194456 21422
rect 194612 4010 194640 338014
rect 195072 335354 195100 338014
rect 194704 335326 195100 335354
rect 194704 4690 194732 335326
rect 195440 316034 195468 338014
rect 194796 316006 195468 316034
rect 194796 7818 194824 316006
rect 195888 215960 195940 215966
rect 195888 215902 195940 215908
rect 194784 7812 194836 7818
rect 194784 7754 194836 7760
rect 195900 6914 195928 215902
rect 195624 6886 195928 6914
rect 194692 4684 194744 4690
rect 194692 4626 194744 4632
rect 194600 4004 194652 4010
rect 194600 3946 194652 3952
rect 195624 480 195652 6886
rect 195992 4078 196020 338014
rect 196360 335354 196388 338014
rect 196084 335326 196388 335354
rect 196084 5914 196112 335326
rect 196728 311894 196756 338014
rect 196176 311866 196756 311894
rect 196176 7886 196204 311866
rect 196164 7880 196216 7886
rect 196164 7822 196216 7828
rect 196072 5908 196124 5914
rect 196072 5850 196124 5856
rect 196808 4956 196860 4962
rect 196808 4898 196860 4904
rect 195980 4072 196032 4078
rect 195980 4014 196032 4020
rect 196820 480 196848 4898
rect 197372 4146 197400 338014
rect 197648 335354 197676 338014
rect 197464 335326 197676 335354
rect 197464 7954 197492 335326
rect 198200 311894 198228 338014
rect 198936 318794 198964 338014
rect 198844 318766 198964 318794
rect 199028 338014 199318 338042
rect 198844 314106 198872 318766
rect 198844 314078 198964 314106
rect 198832 314016 198884 314022
rect 198832 313958 198884 313964
rect 197556 311866 198228 311894
rect 197556 28286 197584 311866
rect 197544 28280 197596 28286
rect 197544 28222 197596 28228
rect 198844 8022 198872 313958
rect 198832 8016 198884 8022
rect 198832 7958 198884 7964
rect 197452 7948 197504 7954
rect 197452 7890 197504 7896
rect 197912 6656 197964 6662
rect 197912 6598 197964 6604
rect 197360 4140 197412 4146
rect 197360 4082 197412 4088
rect 197924 480 197952 6598
rect 198936 3398 198964 314078
rect 199028 314022 199056 338014
rect 199764 336054 199792 338028
rect 200238 338014 200436 338042
rect 199752 336048 199804 336054
rect 199752 335990 199804 335996
rect 200408 331226 200436 338014
rect 200500 338014 200698 338042
rect 200776 338014 201158 338042
rect 201618 338014 201724 338042
rect 200396 331220 200448 331226
rect 200396 331162 200448 331168
rect 200500 326618 200528 338014
rect 200580 331220 200632 331226
rect 200580 331162 200632 331168
rect 200224 326590 200528 326618
rect 199016 314016 199068 314022
rect 199016 313958 199068 313964
rect 200028 11892 200080 11898
rect 200028 11834 200080 11840
rect 200040 3534 200068 11834
rect 200224 8090 200252 326590
rect 200304 326392 200356 326398
rect 200304 326334 200356 326340
rect 200316 312594 200344 326334
rect 200304 312588 200356 312594
rect 200304 312530 200356 312536
rect 200592 311894 200620 331162
rect 200776 326398 200804 338014
rect 200764 326392 200816 326398
rect 200764 326334 200816 326340
rect 201696 318794 201724 338014
rect 201604 318766 201724 318794
rect 201788 338014 201986 338042
rect 201604 313970 201632 318766
rect 201604 313942 201724 313970
rect 201592 313880 201644 313886
rect 201592 313822 201644 313828
rect 200408 311866 200620 311894
rect 200212 8084 200264 8090
rect 200212 8026 200264 8032
rect 200304 5024 200356 5030
rect 200304 4966 200356 4972
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 200028 3528 200080 3534
rect 200028 3470 200080 3476
rect 198924 3392 198976 3398
rect 198924 3334 198976 3340
rect 199120 480 199148 3470
rect 200316 480 200344 4966
rect 200408 3330 200436 311866
rect 201604 8158 201632 313822
rect 201592 8152 201644 8158
rect 201592 8094 201644 8100
rect 201500 3528 201552 3534
rect 201500 3470 201552 3476
rect 200396 3324 200448 3330
rect 200396 3266 200448 3272
rect 201512 480 201540 3470
rect 201696 3262 201724 313942
rect 201788 313886 201816 338014
rect 202144 336592 202196 336598
rect 202144 336534 202196 336540
rect 201776 313880 201828 313886
rect 201776 313822 201828 313828
rect 202156 307086 202184 336534
rect 202432 336122 202460 338028
rect 202906 338014 203196 338042
rect 202420 336116 202472 336122
rect 202420 336058 202472 336064
rect 203168 331226 203196 338014
rect 203260 338014 203366 338042
rect 203536 338014 203826 338042
rect 204286 338014 204392 338042
rect 203156 331220 203208 331226
rect 203156 331162 203208 331168
rect 203260 326618 203288 338014
rect 203340 331220 203392 331226
rect 203340 331162 203392 331168
rect 202984 326590 203288 326618
rect 202144 307080 202196 307086
rect 202144 307022 202196 307028
rect 202788 218748 202840 218754
rect 202788 218690 202840 218696
rect 202800 3534 202828 218690
rect 202984 8226 203012 326590
rect 203064 326392 203116 326398
rect 203064 326334 203116 326340
rect 203076 311166 203104 326334
rect 203352 311894 203380 331162
rect 203536 326398 203564 338014
rect 204364 326482 204392 338014
rect 204456 338014 204654 338042
rect 204456 326618 204484 338014
rect 205100 336598 205128 338028
rect 205192 338014 205574 338042
rect 205836 338014 206034 338042
rect 206112 338014 206494 338042
rect 205088 336592 205140 336598
rect 205088 336534 205140 336540
rect 204456 326590 204668 326618
rect 204364 326454 204576 326482
rect 203524 326392 203576 326398
rect 203524 326334 203576 326340
rect 204352 326392 204404 326398
rect 204352 326334 204404 326340
rect 203168 311866 203380 311894
rect 203064 311160 203116 311166
rect 203064 311102 203116 311108
rect 202972 8220 203024 8226
rect 202972 8162 203024 8168
rect 202788 3528 202840 3534
rect 202788 3470 202840 3476
rect 202696 3460 202748 3466
rect 202696 3402 202748 3408
rect 201684 3256 201736 3262
rect 201684 3198 201736 3204
rect 202708 480 202736 3402
rect 203168 3194 203196 311866
rect 203892 5092 203944 5098
rect 203892 5034 203944 5040
rect 203156 3188 203208 3194
rect 203156 3130 203208 3136
rect 203904 480 203932 5034
rect 204364 3058 204392 326334
rect 204444 326324 204496 326330
rect 204444 326266 204496 326272
rect 204456 8294 204484 326266
rect 204444 8288 204496 8294
rect 204444 8230 204496 8236
rect 204548 3126 204576 326454
rect 204640 326330 204668 326590
rect 205192 326398 205220 338014
rect 205180 326392 205232 326398
rect 205180 326334 205232 326340
rect 205732 326392 205784 326398
rect 205732 326334 205784 326340
rect 204628 326324 204680 326330
rect 204628 326266 204680 326272
rect 205744 11762 205772 326334
rect 205732 11756 205784 11762
rect 205732 11698 205784 11704
rect 205548 10328 205600 10334
rect 205548 10270 205600 10276
rect 205560 3534 205588 10270
rect 205836 7546 205864 338014
rect 206112 326398 206140 338014
rect 206940 336530 206968 338028
rect 207124 338014 207322 338042
rect 207400 338014 207782 338042
rect 207952 338014 208242 338042
rect 208596 338014 208702 338042
rect 208780 338014 209162 338042
rect 206928 336524 206980 336530
rect 206928 336466 206980 336472
rect 206928 336048 206980 336054
rect 206928 335990 206980 335996
rect 206100 326392 206152 326398
rect 206100 326334 206152 326340
rect 205824 7540 205876 7546
rect 205824 7482 205876 7488
rect 206940 3534 206968 335990
rect 207124 7478 207152 338014
rect 207400 335354 207428 338014
rect 207216 335326 207428 335354
rect 207216 309806 207244 335326
rect 207952 316034 207980 338014
rect 208492 324420 208544 324426
rect 208492 324362 208544 324368
rect 207308 316006 207980 316034
rect 207204 309800 207256 309806
rect 207204 309742 207256 309748
rect 207112 7472 207164 7478
rect 207112 7414 207164 7420
rect 205088 3528 205140 3534
rect 205088 3470 205140 3476
rect 205548 3528 205600 3534
rect 205548 3470 205600 3476
rect 206192 3528 206244 3534
rect 206192 3470 206244 3476
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 204536 3120 204588 3126
rect 204536 3062 204588 3068
rect 204352 3052 204404 3058
rect 204352 2994 204404 3000
rect 205100 480 205128 3470
rect 206204 480 206232 3470
rect 207308 2990 207336 316006
rect 208504 21418 208532 324362
rect 208492 21412 208544 21418
rect 208492 21354 208544 21360
rect 208596 7410 208624 338014
rect 208780 324426 208808 338014
rect 209608 336666 209636 338028
rect 209884 338014 209990 338042
rect 209596 336660 209648 336666
rect 209596 336602 209648 336608
rect 209688 336116 209740 336122
rect 209688 336058 209740 336064
rect 208768 324420 208820 324426
rect 208768 324362 208820 324368
rect 208584 7404 208636 7410
rect 208584 7346 208636 7352
rect 207388 5160 207440 5166
rect 207388 5102 207440 5108
rect 207296 2984 207348 2990
rect 207296 2926 207348 2932
rect 207400 480 207428 5102
rect 209700 3534 209728 336058
rect 209884 7342 209912 338014
rect 210436 329118 210464 338028
rect 210528 338014 210910 338042
rect 210424 329112 210476 329118
rect 210424 329054 210476 329060
rect 210528 316034 210556 338014
rect 210976 336184 211028 336190
rect 210976 336126 211028 336132
rect 210068 316006 210556 316034
rect 209872 7336 209924 7342
rect 209872 7278 209924 7284
rect 208584 3528 208636 3534
rect 208584 3470 208636 3476
rect 209688 3528 209740 3534
rect 209688 3470 209740 3476
rect 209780 3528 209832 3534
rect 209780 3470 209832 3476
rect 208596 480 208624 3470
rect 209792 480 209820 3470
rect 210068 2922 210096 316006
rect 210988 3534 211016 336126
rect 211252 326392 211304 326398
rect 211252 326334 211304 326340
rect 211264 308446 211292 326334
rect 211252 308440 211304 308446
rect 211252 308382 211304 308388
rect 211356 7274 211384 338028
rect 211448 338014 211830 338042
rect 211448 326398 211476 338014
rect 212276 336734 212304 338028
rect 212264 336728 212316 336734
rect 212264 336670 212316 336676
rect 212448 336252 212500 336258
rect 212448 336194 212500 336200
rect 211436 326392 211488 326398
rect 211436 326334 211488 326340
rect 211344 7268 211396 7274
rect 211344 7210 211396 7216
rect 212460 6914 212488 336194
rect 212736 326534 212764 338028
rect 212828 338014 213118 338042
rect 212724 326528 212776 326534
rect 212724 326470 212776 326476
rect 212828 323762 212856 338014
rect 213564 335986 213592 338028
rect 213828 336388 213880 336394
rect 213828 336330 213880 336336
rect 213552 335980 213604 335986
rect 213552 335922 213604 335928
rect 212644 323734 212856 323762
rect 212644 305658 212672 323734
rect 212724 323604 212776 323610
rect 212724 323546 212776 323552
rect 212632 305652 212684 305658
rect 212632 305594 212684 305600
rect 212736 7206 212764 323546
rect 212724 7200 212776 7206
rect 212724 7142 212776 7148
rect 212184 6886 212488 6914
rect 211068 5228 211120 5234
rect 211068 5170 211120 5176
rect 210976 3528 211028 3534
rect 210976 3470 211028 3476
rect 210056 2916 210108 2922
rect 210056 2858 210108 2864
rect 211080 2666 211108 5170
rect 210988 2638 211108 2666
rect 210988 480 211016 2638
rect 212184 480 212212 6886
rect 213840 3534 213868 336330
rect 214024 7138 214052 338028
rect 214116 338014 214498 338042
rect 214576 338014 214958 338042
rect 214116 304298 214144 338014
rect 214576 316034 214604 338014
rect 215404 334694 215432 338028
rect 215496 338014 215786 338042
rect 215864 338014 216246 338042
rect 215392 334688 215444 334694
rect 215392 334630 215444 334636
rect 215392 326392 215444 326398
rect 215392 326334 215444 326340
rect 214208 316006 214604 316034
rect 214104 304292 214156 304298
rect 214104 304234 214156 304240
rect 214012 7132 214064 7138
rect 214012 7074 214064 7080
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 213828 3528 213880 3534
rect 213828 3470 213880 3476
rect 213380 480 213408 3470
rect 214208 2854 214236 316006
rect 215208 14612 215260 14618
rect 215208 14554 215260 14560
rect 215220 3534 215248 14554
rect 215404 5846 215432 326334
rect 215392 5840 215444 5846
rect 215392 5782 215444 5788
rect 215496 4622 215524 338014
rect 215864 326398 215892 338014
rect 216692 327826 216720 338028
rect 216784 338014 217166 338042
rect 217336 338014 217626 338042
rect 216680 327820 216732 327826
rect 216680 327762 216732 327768
rect 215852 326392 215904 326398
rect 215852 326334 215904 326340
rect 216784 322318 216812 338014
rect 216772 322312 216824 322318
rect 216772 322254 216824 322260
rect 217336 321554 217364 338014
rect 218072 329186 218100 338028
rect 218440 333266 218468 338028
rect 218532 338014 218914 338042
rect 218992 338014 219374 338042
rect 219544 338014 219834 338042
rect 219912 338014 220294 338042
rect 220372 338014 220754 338042
rect 220924 338014 221122 338042
rect 221200 338014 221582 338042
rect 221660 338014 222042 338042
rect 222304 338014 222502 338042
rect 222672 338014 222962 338042
rect 223040 338014 223422 338042
rect 223776 338014 223882 338042
rect 223960 338014 224250 338042
rect 224328 338014 224710 338042
rect 218428 333260 218480 333266
rect 218428 333202 218480 333208
rect 218060 329180 218112 329186
rect 218060 329122 218112 329128
rect 216692 321526 217364 321554
rect 216692 14482 216720 321526
rect 218532 316034 218560 338014
rect 218992 331906 219020 338014
rect 219348 336320 219400 336326
rect 219348 336262 219400 336268
rect 218980 331900 219032 331906
rect 218980 331842 219032 331848
rect 218348 316006 218560 316034
rect 218348 22778 218376 316006
rect 218336 22772 218388 22778
rect 218336 22714 218388 22720
rect 216680 14476 216732 14482
rect 216680 14418 216732 14424
rect 215484 4616 215536 4622
rect 215484 4558 215536 4564
rect 219256 3664 219308 3670
rect 219256 3606 219308 3612
rect 216864 3596 216916 3602
rect 216864 3538 216916 3544
rect 214472 3528 214524 3534
rect 214472 3470 214524 3476
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215668 3528 215720 3534
rect 215668 3470 215720 3476
rect 214196 2848 214248 2854
rect 214196 2790 214248 2796
rect 214484 480 214512 3470
rect 215680 480 215708 3470
rect 216876 480 216904 3538
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218072 480 218100 3334
rect 219268 480 219296 3606
rect 219360 3398 219388 336262
rect 219440 326392 219492 326398
rect 219440 326334 219492 326340
rect 219452 13122 219480 326334
rect 219544 316742 219572 338014
rect 219912 326398 219940 338014
rect 220372 326466 220400 338014
rect 220820 336728 220872 336734
rect 220820 336670 220872 336676
rect 220728 336456 220780 336462
rect 220728 336398 220780 336404
rect 220360 326460 220412 326466
rect 220360 326402 220412 326408
rect 219900 326392 219952 326398
rect 219900 326334 219952 326340
rect 219532 316736 219584 316742
rect 219532 316678 219584 316684
rect 219440 13116 219492 13122
rect 219440 13058 219492 13064
rect 220740 6914 220768 336398
rect 220832 220114 220860 336670
rect 220924 318102 220952 338014
rect 221200 336734 221228 338014
rect 221188 336728 221240 336734
rect 221188 336670 221240 336676
rect 221660 325038 221688 338014
rect 221648 325032 221700 325038
rect 221648 324974 221700 324980
rect 222200 324284 222252 324290
rect 222200 324226 222252 324232
rect 220912 318096 220964 318102
rect 220912 318038 220964 318044
rect 220820 220108 220872 220114
rect 220820 220050 220872 220056
rect 222212 24138 222240 324226
rect 222304 315314 222332 338014
rect 222672 324290 222700 338014
rect 223040 336682 223068 338014
rect 222764 336654 223068 336682
rect 222660 324284 222712 324290
rect 222660 324226 222712 324232
rect 222764 323678 222792 336654
rect 222844 336592 222896 336598
rect 222844 336534 222896 336540
rect 222752 323672 222804 323678
rect 222752 323614 222804 323620
rect 222292 315308 222344 315314
rect 222292 315250 222344 315256
rect 222200 24132 222252 24138
rect 222200 24074 222252 24080
rect 222856 15910 222884 336534
rect 223776 326534 223804 338014
rect 223960 335354 223988 338014
rect 223868 335326 223988 335354
rect 223764 326528 223816 326534
rect 223764 326470 223816 326476
rect 223580 326392 223632 326398
rect 223580 326334 223632 326340
rect 222844 15904 222896 15910
rect 222844 15846 222896 15852
rect 221556 7608 221608 7614
rect 221556 7550 221608 7556
rect 220464 6886 220768 6914
rect 219348 3392 219400 3398
rect 219348 3334 219400 3340
rect 220464 480 220492 6886
rect 221568 480 221596 7550
rect 223592 4554 223620 326334
rect 223868 323626 223896 335326
rect 224328 326398 224356 338014
rect 224960 326460 225012 326466
rect 224960 326402 225012 326408
rect 224316 326392 224368 326398
rect 224316 326334 224368 326340
rect 223684 323598 223896 323626
rect 223684 25566 223712 323598
rect 223764 321972 223816 321978
rect 223764 321914 223816 321920
rect 223776 313954 223804 321914
rect 223764 313948 223816 313954
rect 223764 313890 223816 313896
rect 223672 25560 223724 25566
rect 223672 25502 223724 25508
rect 223580 4548 223632 4554
rect 223580 4490 223632 4496
rect 224972 4486 225000 326402
rect 225052 326392 225104 326398
rect 225052 326334 225104 326340
rect 225064 221474 225092 326334
rect 225156 319462 225184 338028
rect 225248 338014 225630 338042
rect 225800 338014 226090 338042
rect 226352 338014 226550 338042
rect 226628 338014 226918 338042
rect 226996 338014 227378 338042
rect 227838 338014 227944 338042
rect 225248 326398 225276 338014
rect 225800 326466 225828 338014
rect 226352 330614 226380 338014
rect 226340 330608 226392 330614
rect 226340 330550 226392 330556
rect 225788 326460 225840 326466
rect 225788 326402 225840 326408
rect 225236 326392 225288 326398
rect 225236 326334 225288 326340
rect 226628 321554 226656 338014
rect 226996 336682 227024 338014
rect 226444 321526 226656 321554
rect 226812 336654 227024 336682
rect 225144 319456 225196 319462
rect 225144 319398 225196 319404
rect 225052 221468 225104 221474
rect 225052 221410 225104 221416
rect 226444 26926 226472 321526
rect 226812 316034 226840 336654
rect 226984 336524 227036 336530
rect 226984 336466 227036 336472
rect 226536 316006 226840 316034
rect 226432 26920 226484 26926
rect 226432 26862 226484 26868
rect 224960 4480 225012 4486
rect 224960 4422 225012 4428
rect 226536 4418 226564 316006
rect 226524 4412 226576 4418
rect 226524 4354 226576 4360
rect 223948 3800 224000 3806
rect 223948 3742 224000 3748
rect 222752 3324 222804 3330
rect 222752 3266 222804 3272
rect 222764 480 222792 3266
rect 223960 480 223988 3742
rect 226340 3732 226392 3738
rect 226340 3674 226392 3680
rect 225144 3392 225196 3398
rect 225144 3334 225196 3340
rect 225156 480 225184 3334
rect 226352 480 226380 3674
rect 226996 3398 227024 336466
rect 227812 326392 227864 326398
rect 227812 326334 227864 326340
rect 227824 7070 227852 326334
rect 227812 7064 227864 7070
rect 227812 7006 227864 7012
rect 227916 5778 227944 338014
rect 228008 338014 228298 338042
rect 228008 326398 228036 338014
rect 228744 333334 228772 338028
rect 229218 338014 229324 338042
rect 228732 333328 228784 333334
rect 228732 333270 228784 333276
rect 229296 326466 229324 338014
rect 229388 338014 229586 338042
rect 229284 326460 229336 326466
rect 229284 326402 229336 326408
rect 227996 326392 228048 326398
rect 227996 326334 228048 326340
rect 229284 326256 229336 326262
rect 229284 326198 229336 326204
rect 229192 323604 229244 323610
rect 229192 323546 229244 323552
rect 227904 5772 227956 5778
rect 227904 5714 227956 5720
rect 229204 5710 229232 323546
rect 229192 5704 229244 5710
rect 229192 5646 229244 5652
rect 229296 4350 229324 326198
rect 229388 323610 229416 338014
rect 229744 335980 229796 335986
rect 229744 335922 229796 335928
rect 229376 323604 229428 323610
rect 229376 323546 229428 323552
rect 229756 9042 229784 335922
rect 230032 330682 230060 338028
rect 230506 338014 230704 338042
rect 230020 330676 230072 330682
rect 230020 330618 230072 330624
rect 230572 326392 230624 326398
rect 230572 326334 230624 326340
rect 229744 9036 229796 9042
rect 229744 8978 229796 8984
rect 230584 5642 230612 326334
rect 230572 5636 230624 5642
rect 230572 5578 230624 5584
rect 229284 4344 229336 4350
rect 229284 4286 229336 4292
rect 230676 4282 230704 338014
rect 230768 338014 230966 338042
rect 230768 326398 230796 338014
rect 231124 336592 231176 336598
rect 231124 336534 231176 336540
rect 230756 326392 230808 326398
rect 230756 326334 230808 326340
rect 230664 4276 230716 4282
rect 230664 4218 230716 4224
rect 231032 4072 231084 4078
rect 231032 4014 231084 4020
rect 229836 4004 229888 4010
rect 229836 3946 229888 3952
rect 228732 3936 228784 3942
rect 228732 3878 228784 3884
rect 227536 3868 227588 3874
rect 227536 3810 227588 3816
rect 226984 3392 227036 3398
rect 226984 3334 227036 3340
rect 227548 480 227576 3810
rect 228744 480 228772 3878
rect 229848 480 229876 3946
rect 231044 480 231072 4014
rect 231136 3942 231164 336534
rect 231412 335986 231440 338028
rect 231872 336666 231900 338028
rect 232148 338014 232254 338042
rect 232424 338014 232714 338042
rect 232792 338014 233174 338042
rect 233252 338014 233634 338042
rect 233712 338014 234094 338042
rect 234264 338014 234554 338042
rect 234816 338014 235014 338042
rect 235092 338014 235382 338042
rect 231860 336660 231912 336666
rect 231860 336602 231912 336608
rect 231400 335980 231452 335986
rect 231400 335922 231452 335928
rect 231952 326392 232004 326398
rect 231952 326334 232004 326340
rect 231964 10402 231992 326334
rect 232044 325916 232096 325922
rect 232044 325858 232096 325864
rect 232056 17270 232084 325858
rect 232044 17264 232096 17270
rect 232044 17206 232096 17212
rect 231952 10396 232004 10402
rect 231952 10338 232004 10344
rect 232148 6186 232176 338014
rect 232424 326398 232452 338014
rect 232412 326392 232464 326398
rect 232412 326334 232464 326340
rect 232792 325922 232820 338014
rect 232780 325916 232832 325922
rect 232780 325858 232832 325864
rect 233252 6254 233280 338014
rect 233712 335354 233740 338014
rect 233884 336728 233936 336734
rect 233884 336670 233936 336676
rect 233344 335326 233740 335354
rect 233344 11830 233372 335326
rect 233424 326392 233476 326398
rect 233424 326334 233476 326340
rect 233436 320890 233464 326334
rect 233424 320884 233476 320890
rect 233424 320826 233476 320832
rect 233896 18630 233924 336670
rect 234264 326398 234292 338014
rect 234816 328454 234844 338014
rect 235092 335354 235120 338014
rect 234724 328426 234844 328454
rect 234908 335326 235120 335354
rect 234252 326392 234304 326398
rect 234252 326334 234304 326340
rect 234724 323728 234752 328426
rect 234724 323700 234844 323728
rect 234712 323604 234764 323610
rect 234712 323546 234764 323552
rect 233884 18624 233936 18630
rect 233884 18566 233936 18572
rect 234724 13190 234752 323546
rect 234712 13184 234764 13190
rect 234712 13126 234764 13132
rect 233332 11824 233384 11830
rect 233332 11766 233384 11772
rect 234816 6322 234844 323700
rect 234908 323610 234936 335326
rect 235828 334626 235856 338028
rect 236196 338014 236302 338042
rect 236380 338014 236762 338042
rect 235908 336660 235960 336666
rect 235908 336602 235960 336608
rect 235816 334620 235868 334626
rect 235816 334562 235868 334568
rect 234896 323604 234948 323610
rect 234896 323546 234948 323552
rect 234804 6316 234856 6322
rect 234804 6258 234856 6264
rect 233240 6248 233292 6254
rect 233240 6190 233292 6196
rect 232136 6180 232188 6186
rect 232136 6122 232188 6128
rect 233424 4140 233476 4146
rect 233424 4082 233476 4088
rect 231124 3936 231176 3942
rect 231124 3878 231176 3884
rect 232228 3052 232280 3058
rect 232228 2994 232280 3000
rect 232240 480 232268 2994
rect 233436 480 233464 4082
rect 234620 3392 234672 3398
rect 234620 3334 234672 3340
rect 234632 480 234660 3334
rect 235920 2774 235948 336602
rect 236092 323740 236144 323746
rect 236092 323682 236144 323688
rect 236104 217326 236132 323682
rect 236092 217320 236144 217326
rect 236092 217262 236144 217268
rect 236196 6390 236224 338014
rect 236380 323746 236408 338014
rect 237208 336734 237236 338028
rect 237392 338014 237682 338042
rect 237760 338014 238050 338042
rect 238128 338014 238510 338042
rect 238864 338014 238970 338042
rect 239048 338014 239430 338042
rect 237196 336728 237248 336734
rect 237196 336670 237248 336676
rect 236644 335436 236696 335442
rect 236644 335378 236696 335384
rect 236368 323740 236420 323746
rect 236368 323682 236420 323688
rect 236656 14550 236684 335378
rect 236644 14544 236696 14550
rect 236644 14486 236696 14492
rect 237392 6458 237420 338014
rect 237760 335354 237788 338014
rect 237484 335326 237788 335354
rect 237484 8974 237512 335326
rect 238128 316034 238156 338014
rect 237576 316006 238156 316034
rect 237576 19990 237604 316006
rect 237564 19984 237616 19990
rect 237564 19926 237616 19932
rect 237472 8968 237524 8974
rect 237472 8910 237524 8916
rect 238864 6526 238892 338014
rect 239048 316034 239076 338014
rect 239404 336728 239456 336734
rect 239404 336670 239456 336676
rect 238956 316006 239076 316034
rect 238852 6520 238904 6526
rect 238852 6462 238904 6468
rect 237380 6452 237432 6458
rect 237380 6394 237432 6400
rect 236184 6384 236236 6390
rect 236184 6326 236236 6332
rect 238956 4826 238984 316006
rect 239416 215966 239444 336670
rect 239876 335442 239904 338028
rect 240244 338014 240350 338042
rect 240428 338014 240718 338042
rect 240796 338014 241178 338042
rect 240140 336796 240192 336802
rect 240140 336738 240192 336744
rect 239864 335436 239916 335442
rect 239864 335378 239916 335384
rect 239404 215960 239456 215966
rect 239404 215902 239456 215908
rect 240152 4894 240180 336738
rect 240244 6594 240272 338014
rect 240428 336802 240456 338014
rect 240416 336796 240468 336802
rect 240416 336738 240468 336744
rect 240796 316034 240824 338014
rect 241624 336734 241652 338028
rect 241716 338014 242098 338042
rect 242176 338014 242558 338042
rect 241612 336728 241664 336734
rect 241612 336670 241664 336676
rect 241612 326392 241664 326398
rect 241612 326334 241664 326340
rect 240336 316006 240824 316034
rect 240336 21486 240364 316006
rect 240324 21480 240376 21486
rect 240324 21422 240376 21428
rect 241624 6662 241652 326334
rect 241612 6656 241664 6662
rect 241612 6598 241664 6604
rect 240232 6588 240284 6594
rect 240232 6530 240284 6536
rect 241716 4962 241744 338014
rect 242072 336728 242124 336734
rect 242072 336670 242124 336676
rect 242084 321554 242112 336670
rect 242176 326398 242204 338014
rect 243004 335646 243032 338028
rect 243096 338014 243386 338042
rect 243464 338014 243846 338042
rect 242256 335640 242308 335646
rect 242256 335582 242308 335588
rect 242992 335640 243044 335646
rect 242992 335582 243044 335588
rect 242164 326392 242216 326398
rect 242164 326334 242216 326340
rect 242084 321526 242204 321554
rect 241704 4956 241756 4962
rect 241704 4898 241756 4904
rect 240140 4888 240192 4894
rect 240140 4830 240192 4836
rect 238944 4820 238996 4826
rect 238944 4762 238996 4768
rect 238116 3324 238168 3330
rect 238116 3266 238168 3272
rect 237012 2916 237064 2922
rect 237012 2858 237064 2864
rect 235828 2746 235948 2774
rect 235828 480 235856 2746
rect 237024 480 237052 2858
rect 238128 480 238156 3266
rect 241704 3256 241756 3262
rect 241704 3198 241756 3204
rect 240508 3120 240560 3126
rect 240508 3062 240560 3068
rect 239312 2848 239364 2854
rect 239312 2790 239364 2796
rect 239324 480 239352 2790
rect 240520 480 240548 3062
rect 241716 480 241744 3198
rect 242176 3058 242204 321526
rect 242268 11898 242296 335582
rect 242992 326392 243044 326398
rect 242992 326334 243044 326340
rect 243004 218754 243032 326334
rect 242992 218748 243044 218754
rect 242992 218690 243044 218696
rect 242256 11892 242308 11898
rect 242256 11834 242308 11840
rect 243096 5030 243124 338014
rect 243464 326398 243492 338014
rect 243452 326392 243504 326398
rect 243452 326334 243504 326340
rect 243084 5024 243136 5030
rect 243084 4966 243136 4972
rect 242900 3596 242952 3602
rect 242900 3538 242952 3544
rect 242164 3052 242216 3058
rect 242164 2994 242216 3000
rect 242912 480 242940 3538
rect 244188 3460 244240 3466
rect 244188 3402 244240 3408
rect 244200 3176 244228 3402
rect 244292 3176 244320 338028
rect 244384 338014 244766 338042
rect 244844 338014 245226 338042
rect 244384 5098 244412 338014
rect 244844 316034 244872 338014
rect 245672 336054 245700 338028
rect 245856 338014 246146 338042
rect 245660 336048 245712 336054
rect 245660 335990 245712 335996
rect 244476 316006 244872 316034
rect 244476 10334 244504 316006
rect 244464 10328 244516 10334
rect 244464 10270 244516 10276
rect 245856 5166 245884 338014
rect 246500 336122 246528 338028
rect 246960 336190 246988 338028
rect 247144 338014 247434 338042
rect 247512 338014 247894 338042
rect 246948 336184 247000 336190
rect 246948 336126 247000 336132
rect 246488 336116 246540 336122
rect 246488 336058 246540 336064
rect 246304 335368 246356 335374
rect 246304 335310 246356 335316
rect 246316 14618 246344 335310
rect 246304 14612 246356 14618
rect 246304 14554 246356 14560
rect 247144 5234 247172 338014
rect 247512 336258 247540 338014
rect 248340 336394 248368 338028
rect 248328 336388 248380 336394
rect 248328 336330 248380 336336
rect 247500 336252 247552 336258
rect 247500 336194 247552 336200
rect 247684 336252 247736 336258
rect 247684 336194 247736 336200
rect 247696 7614 247724 336194
rect 248328 336048 248380 336054
rect 248328 335990 248380 335996
rect 247684 7608 247736 7614
rect 247684 7550 247736 7556
rect 247132 5228 247184 5234
rect 247132 5170 247184 5176
rect 245844 5160 245896 5166
rect 245844 5102 245896 5108
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 248340 3670 248368 335990
rect 248800 335374 248828 338028
rect 248892 338014 249182 338042
rect 249352 338014 249642 338042
rect 248788 335368 248840 335374
rect 248788 335310 248840 335316
rect 248512 330540 248564 330546
rect 248512 330482 248564 330488
rect 247592 3664 247644 3670
rect 247592 3606 247644 3612
rect 248328 3664 248380 3670
rect 248328 3606 248380 3612
rect 245200 3460 245252 3466
rect 245200 3402 245252 3408
rect 244200 3148 244320 3176
rect 244096 3052 244148 3058
rect 244096 2994 244148 3000
rect 244108 480 244136 2994
rect 245212 480 245240 3402
rect 246396 2848 246448 2854
rect 246396 2790 246448 2796
rect 246408 480 246436 2790
rect 247604 480 247632 3606
rect 248524 3534 248552 330482
rect 248892 316034 248920 338014
rect 249064 336116 249116 336122
rect 249064 336058 249116 336064
rect 248708 316006 248920 316034
rect 248512 3528 248564 3534
rect 248512 3470 248564 3476
rect 248420 3324 248472 3330
rect 248420 3266 248472 3272
rect 248432 3074 248460 3266
rect 248708 3194 248736 316006
rect 248788 3528 248840 3534
rect 248788 3470 248840 3476
rect 248696 3188 248748 3194
rect 248696 3130 248748 3136
rect 248432 3046 248644 3074
rect 248616 2786 248644 3046
rect 248604 2780 248656 2786
rect 248604 2722 248656 2728
rect 248800 480 248828 3470
rect 249076 2854 249104 336058
rect 249352 330546 249380 338014
rect 250088 336326 250116 338028
rect 250180 338014 250562 338042
rect 250076 336320 250128 336326
rect 250076 336262 250128 336268
rect 249340 330540 249392 330546
rect 249340 330482 249392 330488
rect 250180 316034 250208 338014
rect 251008 336462 251036 338028
rect 250996 336456 251048 336462
rect 250996 336398 251048 336404
rect 251468 336258 251496 338028
rect 251560 338014 251850 338042
rect 251928 338014 252310 338042
rect 251456 336252 251508 336258
rect 251456 336194 251508 336200
rect 250536 336184 250588 336190
rect 250536 336126 250588 336132
rect 250444 335980 250496 335986
rect 250444 335922 250496 335928
rect 249904 316006 250208 316034
rect 249904 2990 249932 316006
rect 249892 2984 249944 2990
rect 249892 2926 249944 2932
rect 249984 2916 250036 2922
rect 249984 2858 250036 2864
rect 249064 2848 249116 2854
rect 249064 2790 249116 2796
rect 249996 480 250024 2858
rect 250456 2854 250484 335922
rect 250548 3670 250576 336126
rect 251272 330540 251324 330546
rect 251272 330482 251324 330488
rect 251284 3806 251312 330482
rect 251560 316034 251588 338014
rect 251824 336320 251876 336326
rect 251824 336262 251876 336268
rect 251376 316006 251588 316034
rect 251272 3800 251324 3806
rect 251272 3742 251324 3748
rect 251376 3738 251404 316006
rect 251364 3732 251416 3738
rect 251364 3674 251416 3680
rect 250536 3664 250588 3670
rect 250536 3606 250588 3612
rect 251180 3188 251232 3194
rect 251180 3130 251232 3136
rect 250444 2848 250496 2854
rect 250444 2790 250496 2796
rect 251192 480 251220 3130
rect 251836 3058 251864 336262
rect 251928 330546 251956 338014
rect 252756 336530 252784 338028
rect 252848 338014 253230 338042
rect 253400 338014 253690 338042
rect 252744 336524 252796 336530
rect 252744 336466 252796 336472
rect 252008 335640 252060 335646
rect 252008 335582 252060 335588
rect 251916 330540 251968 330546
rect 251916 330482 251968 330488
rect 252020 316034 252048 335582
rect 252652 330540 252704 330546
rect 252652 330482 252704 330488
rect 251928 316006 252048 316034
rect 251928 3126 251956 316006
rect 252664 4010 252692 330482
rect 252848 316034 252876 338014
rect 253296 336388 253348 336394
rect 253296 336330 253348 336336
rect 253204 335368 253256 335374
rect 253204 335310 253256 335316
rect 252756 316006 252876 316034
rect 252652 4004 252704 4010
rect 252652 3946 252704 3952
rect 252756 3942 252784 316006
rect 252744 3936 252796 3942
rect 252744 3878 252796 3884
rect 252376 3596 252428 3602
rect 252376 3538 252428 3544
rect 251916 3120 251968 3126
rect 251916 3062 251968 3068
rect 251824 3052 251876 3058
rect 251824 2994 251876 3000
rect 252388 480 252416 3538
rect 253216 3330 253244 335310
rect 253204 3324 253256 3330
rect 253204 3266 253256 3272
rect 253308 2922 253336 336330
rect 253400 330546 253428 338014
rect 254136 336598 254164 338028
rect 254228 338014 254518 338042
rect 254596 338014 254978 338042
rect 254124 336592 254176 336598
rect 254124 336534 254176 336540
rect 253848 336252 253900 336258
rect 253848 336194 253900 336200
rect 253388 330540 253440 330546
rect 253388 330482 253440 330488
rect 253860 6914 253888 336194
rect 254228 335354 254256 338014
rect 253492 6886 253888 6914
rect 254044 335326 254256 335354
rect 253296 2916 253348 2922
rect 253296 2858 253348 2864
rect 253492 480 253520 6886
rect 254044 4146 254072 335326
rect 254596 316034 254624 338014
rect 255424 336734 255452 338028
rect 255516 338014 255898 338042
rect 255976 338014 256358 338042
rect 255412 336728 255464 336734
rect 255412 336670 255464 336676
rect 255412 326392 255464 326398
rect 255412 326334 255464 326340
rect 254136 316006 254624 316034
rect 254032 4140 254084 4146
rect 254032 4082 254084 4088
rect 254136 4078 254164 316006
rect 254124 4072 254176 4078
rect 254124 4014 254176 4020
rect 254676 3664 254728 3670
rect 254676 3606 254728 3612
rect 254688 480 254716 3606
rect 255424 3398 255452 326334
rect 255516 3466 255544 338014
rect 255976 326398 256004 338014
rect 256804 336666 256832 338028
rect 256792 336660 256844 336666
rect 256792 336602 256844 336608
rect 257264 335986 257292 338028
rect 257356 338014 257646 338042
rect 257252 335980 257304 335986
rect 257252 335922 257304 335928
rect 255964 326392 256016 326398
rect 255964 326334 256016 326340
rect 257356 316034 257384 338014
rect 258092 336122 258120 338028
rect 258080 336116 258132 336122
rect 258080 336058 258132 336064
rect 258552 335646 258580 338028
rect 258644 338014 259026 338042
rect 258540 335640 258592 335646
rect 258540 335582 258592 335588
rect 258644 316034 258672 338014
rect 258724 336660 258776 336666
rect 258724 336602 258776 336608
rect 256896 316006 257384 316034
rect 258184 316006 258672 316034
rect 255872 3800 255924 3806
rect 255872 3742 255924 3748
rect 255504 3460 255556 3466
rect 255504 3402 255556 3408
rect 255412 3392 255464 3398
rect 255412 3334 255464 3340
rect 255884 480 255912 3742
rect 256896 2854 256924 316006
rect 257068 3732 257120 3738
rect 257068 3674 257120 3680
rect 256884 2848 256936 2854
rect 256884 2790 256936 2796
rect 257080 480 257108 3674
rect 258184 3262 258212 316006
rect 258736 3738 258764 336602
rect 259472 336190 259500 338028
rect 259460 336184 259512 336190
rect 259460 336126 259512 336132
rect 259368 335640 259420 335646
rect 259368 335582 259420 335588
rect 258724 3732 258776 3738
rect 258724 3674 258776 3680
rect 259380 3534 259408 335582
rect 259932 335374 259960 338028
rect 260024 338014 260314 338042
rect 259920 335368 259972 335374
rect 259920 335310 259972 335316
rect 260024 316034 260052 338014
rect 260656 336728 260708 336734
rect 260656 336670 260708 336676
rect 259656 316006 260052 316034
rect 259656 3874 259684 316006
rect 259644 3868 259696 3874
rect 259644 3810 259696 3816
rect 260668 3602 260696 336670
rect 260760 336326 260788 338028
rect 260748 336320 260800 336326
rect 260748 336262 260800 336268
rect 260748 336184 260800 336190
rect 260748 336126 260800 336132
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 258172 3256 258224 3262
rect 258172 3198 258224 3204
rect 258276 480 258304 3470
rect 259472 480 259500 3538
rect 260760 3482 260788 336126
rect 261220 336054 261248 338028
rect 261312 338014 261694 338042
rect 261208 336048 261260 336054
rect 261208 335990 261260 335996
rect 261312 316034 261340 338014
rect 262140 336394 262168 338028
rect 262416 338014 262614 338042
rect 262692 338014 262982 338042
rect 262128 336388 262180 336394
rect 262128 336330 262180 336336
rect 262416 326466 262444 338014
rect 262692 335354 262720 338014
rect 263428 336258 263456 338028
rect 263704 338014 263902 338042
rect 263980 338014 264362 338042
rect 263416 336252 263468 336258
rect 263416 336194 263468 336200
rect 262508 335326 262720 335354
rect 262404 326460 262456 326466
rect 262404 326402 262456 326408
rect 262404 326256 262456 326262
rect 262404 326198 262456 326204
rect 262312 319388 262364 319394
rect 262312 319330 262364 319336
rect 260668 3454 260788 3482
rect 261036 316006 261340 316034
rect 261036 3466 261064 316006
rect 262324 3670 262352 319330
rect 262312 3664 262364 3670
rect 262312 3606 262364 3612
rect 261760 3596 261812 3602
rect 261760 3538 261812 3544
rect 261024 3460 261076 3466
rect 260668 480 260696 3454
rect 261024 3402 261076 3408
rect 261772 480 261800 3538
rect 262416 3194 262444 326198
rect 262508 319394 262536 335326
rect 262496 319388 262548 319394
rect 262496 319330 262548 319336
rect 263704 3738 263732 338014
rect 263980 316034 264008 338014
rect 264808 336666 264836 338028
rect 264796 336660 264848 336666
rect 264796 336602 264848 336608
rect 265268 335646 265296 338028
rect 265636 336734 265664 338028
rect 265624 336728 265676 336734
rect 265624 336670 265676 336676
rect 266096 336190 266124 338028
rect 266084 336184 266136 336190
rect 266084 336126 266136 336132
rect 265716 335980 265768 335986
rect 265716 335922 265768 335928
rect 265624 335844 265676 335850
rect 265624 335786 265676 335792
rect 265256 335640 265308 335646
rect 265256 335582 265308 335588
rect 263796 316006 264008 316034
rect 263796 3806 263824 316006
rect 263784 3800 263836 3806
rect 263784 3742 263836 3748
rect 263692 3732 263744 3738
rect 263692 3674 263744 3680
rect 265636 3602 265664 335786
rect 265624 3596 265676 3602
rect 265624 3538 265676 3544
rect 265348 3528 265400 3534
rect 265348 3470 265400 3476
rect 262956 3460 263008 3466
rect 262956 3402 263008 3408
rect 262404 3188 262456 3194
rect 262404 3130 262456 3136
rect 262968 480 262996 3402
rect 264152 3188 264204 3194
rect 264152 3130 264204 3136
rect 264164 480 264192 3130
rect 265360 480 265388 3470
rect 265728 3466 265756 335922
rect 266556 335850 266584 338028
rect 266648 338014 267030 338042
rect 267108 338014 267490 338042
rect 266648 335986 266676 338014
rect 267108 336682 267136 338014
rect 266924 336654 267136 336682
rect 266636 335980 266688 335986
rect 266636 335922 266688 335928
rect 266544 335844 266596 335850
rect 266544 335786 266596 335792
rect 266924 316034 266952 336654
rect 267936 335782 267964 338028
rect 268028 338014 268410 338042
rect 268488 338014 268778 338042
rect 267004 335776 267056 335782
rect 267004 335718 267056 335724
rect 267924 335776 267976 335782
rect 267924 335718 267976 335724
rect 266464 316006 266952 316034
rect 265716 3460 265768 3466
rect 265716 3402 265768 3408
rect 266464 3194 266492 316006
rect 267016 3534 267044 335718
rect 267832 326392 267884 326398
rect 267832 326334 267884 326340
rect 267844 6914 267872 326334
rect 267752 6886 267872 6914
rect 267004 3528 267056 3534
rect 267004 3470 267056 3476
rect 266452 3188 266504 3194
rect 266452 3130 266504 3136
rect 266544 3120 266596 3126
rect 266544 3062 266596 3068
rect 266556 480 266584 3062
rect 267752 480 267780 6886
rect 268028 3126 268056 338014
rect 268488 326398 268516 338014
rect 269224 326466 269252 338028
rect 269316 338014 269698 338042
rect 270158 338014 270448 338042
rect 269212 326460 269264 326466
rect 269212 326402 269264 326408
rect 268476 326392 268528 326398
rect 268476 326334 268528 326340
rect 269212 326256 269264 326262
rect 269212 326198 269264 326204
rect 269120 319388 269172 319394
rect 269120 319330 269172 319336
rect 269132 3602 269160 319330
rect 269120 3596 269172 3602
rect 269120 3538 269172 3544
rect 269224 3482 269252 326198
rect 269316 319394 269344 338014
rect 270420 335354 270448 338014
rect 270604 336666 270632 338028
rect 271064 336734 271092 338028
rect 271446 338014 271736 338042
rect 271906 338014 272288 338042
rect 271052 336728 271104 336734
rect 271052 336670 271104 336676
rect 270592 336660 270644 336666
rect 270592 336602 270644 336608
rect 270420 335326 270816 335354
rect 269304 319388 269356 319394
rect 269304 319330 269356 319336
rect 270788 16574 270816 335326
rect 270788 16546 271276 16574
rect 270040 3596 270092 3602
rect 270040 3538 270092 3544
rect 268856 3454 269252 3482
rect 268016 3120 268068 3126
rect 268016 3062 268068 3068
rect 268856 480 268884 3454
rect 270052 480 270080 3538
rect 271248 480 271276 16546
rect 271708 3534 271736 338014
rect 272260 336734 272288 338014
rect 271788 336728 271840 336734
rect 271788 336670 271840 336676
rect 272248 336728 272300 336734
rect 272248 336670 272300 336676
rect 271696 3528 271748 3534
rect 271696 3470 271748 3476
rect 271800 2990 271828 336670
rect 271880 336660 271932 336666
rect 271880 336602 271932 336608
rect 271892 16574 271920 336602
rect 272352 335714 272380 338028
rect 272340 335708 272392 335714
rect 272340 335650 272392 335656
rect 272812 335578 272840 338028
rect 272800 335572 272852 335578
rect 272800 335514 272852 335520
rect 273272 335510 273300 338028
rect 273746 338014 274036 338042
rect 274114 338014 274496 338042
rect 273260 335504 273312 335510
rect 273260 335446 273312 335452
rect 274008 335354 274036 338014
rect 274008 335326 274404 335354
rect 271892 16546 272472 16574
rect 271788 2984 271840 2990
rect 271788 2926 271840 2932
rect 272444 480 272472 16546
rect 274376 3602 274404 335326
rect 274364 3596 274416 3602
rect 274364 3538 274416 3544
rect 274468 3466 274496 338014
rect 274560 336190 274588 338028
rect 274548 336184 274600 336190
rect 274548 336126 274600 336132
rect 275020 336122 275048 338028
rect 275480 336258 275508 338028
rect 275468 336252 275520 336258
rect 275468 336194 275520 336200
rect 275008 336116 275060 336122
rect 275008 336058 275060 336064
rect 275940 336054 275968 338028
rect 276400 336734 276428 338028
rect 276782 338014 277164 338042
rect 277242 338014 277348 338042
rect 276204 336728 276256 336734
rect 276204 336670 276256 336676
rect 276388 336728 276440 336734
rect 276388 336670 276440 336676
rect 275928 336048 275980 336054
rect 275928 335990 275980 335996
rect 275284 335708 275336 335714
rect 275284 335650 275336 335656
rect 274548 335504 274600 335510
rect 274548 335446 274600 335452
rect 274456 3460 274508 3466
rect 274456 3402 274508 3408
rect 274560 3126 274588 335446
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 274548 3120 274600 3126
rect 274548 3062 274600 3068
rect 273628 2984 273680 2990
rect 273628 2926 273680 2932
rect 273640 480 273668 2926
rect 274836 480 274864 3470
rect 275296 3058 275324 335650
rect 276216 6914 276244 336670
rect 276032 6886 276244 6914
rect 275284 3052 275336 3058
rect 275284 2994 275336 3000
rect 276032 480 276060 6886
rect 277136 4826 277164 338014
rect 277216 336728 277268 336734
rect 277216 336670 277268 336676
rect 277124 4820 277176 4826
rect 277124 4762 277176 4768
rect 277228 4010 277256 336670
rect 277216 4004 277268 4010
rect 277216 3946 277268 3952
rect 277320 3126 277348 338014
rect 277688 336666 277716 338028
rect 277676 336660 277728 336666
rect 277676 336602 277728 336608
rect 278148 336326 278176 338028
rect 278622 338014 278728 338042
rect 278596 336660 278648 336666
rect 278596 336602 278648 336608
rect 278136 336320 278188 336326
rect 278136 336262 278188 336268
rect 277584 335572 277636 335578
rect 277584 335514 277636 335520
rect 277596 325694 277624 335514
rect 277596 325666 277716 325694
rect 277688 16574 277716 325666
rect 277688 16546 278360 16574
rect 277308 3120 277360 3126
rect 277308 3062 277360 3068
rect 277124 3052 277176 3058
rect 277124 2994 277176 3000
rect 277136 480 277164 2994
rect 278332 480 278360 16546
rect 278608 3534 278636 336602
rect 278596 3528 278648 3534
rect 278596 3470 278648 3476
rect 278700 3194 278728 338014
rect 279068 336734 279096 338028
rect 279542 338014 279832 338042
rect 279910 338014 280016 338042
rect 279056 336728 279108 336734
rect 279056 336670 279108 336676
rect 279804 335354 279832 338014
rect 279804 335326 279924 335354
rect 279896 217394 279924 335326
rect 279884 217388 279936 217394
rect 279884 217330 279936 217336
rect 279988 4146 280016 338014
rect 280356 336734 280384 338028
rect 280830 338014 281120 338042
rect 281290 338014 281488 338042
rect 280068 336728 280120 336734
rect 280068 336670 280120 336676
rect 280344 336728 280396 336734
rect 280344 336670 280396 336676
rect 279976 4140 280028 4146
rect 279976 4082 280028 4088
rect 280080 3262 280108 336670
rect 281092 335354 281120 338014
rect 281356 336728 281408 336734
rect 281356 336670 281408 336676
rect 281092 335326 281304 335354
rect 281276 6254 281304 335326
rect 281264 6248 281316 6254
rect 281264 6190 281316 6196
rect 280712 3596 280764 3602
rect 280712 3538 280764 3544
rect 280068 3256 280120 3262
rect 280068 3198 280120 3204
rect 278688 3188 278740 3194
rect 278688 3130 278740 3136
rect 279516 3052 279568 3058
rect 279516 2994 279568 3000
rect 279528 480 279556 2994
rect 280724 480 280752 3538
rect 281368 3398 281396 336670
rect 281460 3942 281488 338014
rect 281736 336734 281764 338028
rect 282210 338014 282500 338042
rect 282578 338014 282776 338042
rect 281724 336728 281776 336734
rect 281724 336670 281776 336676
rect 282184 336252 282236 336258
rect 282184 336194 282236 336200
rect 281448 3936 281500 3942
rect 281448 3878 281500 3884
rect 281908 3460 281960 3466
rect 281908 3402 281960 3408
rect 281356 3392 281408 3398
rect 281356 3334 281408 3340
rect 281920 480 281948 3402
rect 282196 3330 282224 336194
rect 282472 335354 282500 338014
rect 282472 335326 282684 335354
rect 282656 215966 282684 335326
rect 282644 215960 282696 215966
rect 282644 215902 282696 215908
rect 282748 3670 282776 338014
rect 282828 336728 282880 336734
rect 282828 336670 282880 336676
rect 282840 3874 282868 336670
rect 283024 335442 283052 338028
rect 283498 338014 283880 338042
rect 283958 338014 284156 338042
rect 283196 336184 283248 336190
rect 283196 336126 283248 336132
rect 283012 335436 283064 335442
rect 283012 335378 283064 335384
rect 283208 6914 283236 336126
rect 283852 335354 283880 338014
rect 283852 335326 284064 335354
rect 284036 218754 284064 335326
rect 284024 218748 284076 218754
rect 284024 218690 284076 218696
rect 283116 6886 283236 6914
rect 282828 3868 282880 3874
rect 282828 3810 282880 3816
rect 282736 3664 282788 3670
rect 282736 3606 282788 3612
rect 282184 3324 282236 3330
rect 282184 3266 282236 3272
rect 283116 480 283144 6886
rect 284128 3602 284156 338014
rect 284404 335578 284432 338028
rect 284878 338014 285168 338042
rect 285246 338014 285536 338042
rect 284484 336116 284536 336122
rect 284484 336058 284536 336064
rect 284392 335572 284444 335578
rect 284392 335514 284444 335520
rect 284208 335436 284260 335442
rect 284208 335378 284260 335384
rect 284220 3806 284248 335378
rect 284496 6914 284524 336058
rect 285140 335354 285168 338014
rect 285140 335326 285444 335354
rect 285416 8974 285444 335326
rect 285404 8968 285456 8974
rect 285404 8910 285456 8916
rect 284312 6886 284524 6914
rect 284208 3800 284260 3806
rect 284208 3742 284260 3748
rect 284116 3596 284168 3602
rect 284116 3538 284168 3544
rect 284312 480 284340 6886
rect 285508 3466 285536 338014
rect 285692 336054 285720 338028
rect 286152 336734 286180 338028
rect 286140 336728 286192 336734
rect 286140 336670 286192 336676
rect 286612 336258 286640 338028
rect 286876 336728 286928 336734
rect 286876 336670 286928 336676
rect 286600 336252 286652 336258
rect 286600 336194 286652 336200
rect 285680 336048 285732 336054
rect 285680 335990 285732 335996
rect 285772 335980 285824 335986
rect 285772 335922 285824 335928
rect 285588 335572 285640 335578
rect 285588 335514 285640 335520
rect 285600 3738 285628 335514
rect 285784 16574 285812 335922
rect 286888 18698 286916 336670
rect 287072 336394 287100 338028
rect 287546 338014 287836 338042
rect 287060 336388 287112 336394
rect 287060 336330 287112 336336
rect 286968 336048 287020 336054
rect 286968 335990 287020 335996
rect 286876 18692 286928 18698
rect 286876 18634 286928 18640
rect 285784 16546 286640 16574
rect 285588 3732 285640 3738
rect 285588 3674 285640 3680
rect 285496 3460 285548 3466
rect 285496 3402 285548 3408
rect 285404 3324 285456 3330
rect 285404 3266 285456 3272
rect 285416 480 285444 3266
rect 286612 480 286640 16546
rect 286980 3534 287008 335990
rect 287808 335354 287836 338014
rect 287900 336190 287928 338028
rect 288256 336388 288308 336394
rect 288256 336330 288308 336336
rect 287888 336184 287940 336190
rect 287888 336126 287940 336132
rect 287808 335326 288204 335354
rect 288176 6186 288204 335326
rect 288164 6180 288216 6186
rect 288164 6122 288216 6128
rect 288268 4078 288296 336330
rect 288256 4072 288308 4078
rect 288256 4014 288308 4020
rect 288360 4010 288388 338028
rect 288820 335918 288848 338028
rect 289294 338014 289676 338042
rect 288808 335912 288860 335918
rect 288808 335854 288860 335860
rect 289648 15910 289676 338014
rect 289740 336734 289768 338028
rect 289728 336728 289780 336734
rect 289728 336670 289780 336676
rect 290200 336122 290228 338028
rect 290464 336728 290516 336734
rect 290464 336670 290516 336676
rect 290188 336116 290240 336122
rect 290188 336058 290240 336064
rect 289728 335912 289780 335918
rect 289728 335854 289780 335860
rect 289636 15904 289688 15910
rect 289636 15846 289688 15852
rect 289740 10470 289768 335854
rect 290476 224262 290504 336670
rect 290660 336394 290688 338028
rect 291042 338014 291148 338042
rect 290648 336388 290700 336394
rect 290648 336330 290700 336336
rect 290464 224256 290516 224262
rect 290464 224198 290516 224204
rect 289728 10464 289780 10470
rect 289728 10406 289780 10412
rect 291120 10402 291148 338014
rect 291488 336734 291516 338028
rect 291476 336728 291528 336734
rect 291476 336670 291528 336676
rect 291844 336320 291896 336326
rect 291844 336262 291896 336268
rect 291108 10396 291160 10402
rect 291108 10338 291160 10344
rect 288992 4820 289044 4826
rect 288992 4762 289044 4768
rect 287796 4004 287848 4010
rect 287796 3946 287848 3952
rect 288348 4004 288400 4010
rect 288348 3946 288400 3952
rect 286968 3528 287020 3534
rect 286968 3470 287020 3476
rect 287808 480 287836 3946
rect 289004 480 289032 4762
rect 291856 4214 291884 336262
rect 291948 336054 291976 338028
rect 291936 336048 291988 336054
rect 291936 335990 291988 335996
rect 292408 19990 292436 338028
rect 292868 336734 292896 338028
rect 292488 336728 292540 336734
rect 292488 336670 292540 336676
rect 292856 336728 292908 336734
rect 292856 336670 292908 336676
rect 292396 19984 292448 19990
rect 292396 19926 292448 19932
rect 292500 11830 292528 336670
rect 293328 336326 293356 338028
rect 293710 338014 293908 338042
rect 293776 336728 293828 336734
rect 293776 336670 293828 336676
rect 293316 336320 293368 336326
rect 293316 336262 293368 336268
rect 293788 217326 293816 336670
rect 293776 217320 293828 217326
rect 293776 217262 293828 217268
rect 292488 11824 292540 11830
rect 292488 11766 292540 11772
rect 293880 11762 293908 338014
rect 294156 335986 294184 338028
rect 294616 336734 294644 338028
rect 295090 338014 295196 338042
rect 294604 336728 294656 336734
rect 294604 336670 294656 336676
rect 294144 335980 294196 335986
rect 294144 335922 294196 335928
rect 295064 335980 295116 335986
rect 295064 335922 295116 335928
rect 295076 13122 295104 335922
rect 295064 13116 295116 13122
rect 295064 13058 295116 13064
rect 293868 11756 293920 11762
rect 293868 11698 293920 11704
rect 295168 10334 295196 338014
rect 295248 336728 295300 336734
rect 295248 336670 295300 336676
rect 295156 10328 295208 10334
rect 295156 10270 295208 10276
rect 295260 4350 295288 336670
rect 295536 335578 295564 338028
rect 295996 336734 296024 338028
rect 296378 338014 296576 338042
rect 295984 336728 296036 336734
rect 295984 336670 296036 336676
rect 295524 335572 295576 335578
rect 295524 335514 295576 335520
rect 296444 335572 296496 335578
rect 296444 335514 296496 335520
rect 296456 220114 296484 335514
rect 296444 220108 296496 220114
rect 296444 220050 296496 220056
rect 295340 217388 295392 217394
rect 295340 217330 295392 217336
rect 295352 16574 295380 217330
rect 296548 21418 296576 338014
rect 296628 336728 296680 336734
rect 296628 336670 296680 336676
rect 296536 21412 296588 21418
rect 296536 21354 296588 21360
rect 295352 16546 296116 16574
rect 295248 4344 295300 4350
rect 295248 4286 295300 4292
rect 291844 4208 291896 4214
rect 291844 4150 291896 4156
rect 292580 4208 292632 4214
rect 292580 4150 292632 4156
rect 291384 3188 291436 3194
rect 291384 3130 291436 3136
rect 290188 3120 290240 3126
rect 290188 3062 290240 3068
rect 290200 480 290228 3062
rect 291396 480 291424 3130
rect 292592 480 292620 4150
rect 294880 3324 294932 3330
rect 294880 3266 294932 3272
rect 293684 3256 293736 3262
rect 293684 3198 293736 3204
rect 293696 480 293724 3198
rect 294892 480 294920 3266
rect 296088 480 296116 16546
rect 296640 4418 296668 336670
rect 296824 336598 296852 338028
rect 297298 338014 297680 338042
rect 297758 338014 298048 338042
rect 297652 336682 297680 338014
rect 298020 336818 298048 338014
rect 298020 336790 298140 336818
rect 297652 336654 298048 336682
rect 296812 336592 296864 336598
rect 296812 336534 296864 336540
rect 297916 336592 297968 336598
rect 297916 336534 297968 336540
rect 297928 221474 297956 336534
rect 297916 221468 297968 221474
rect 297916 221410 297968 221416
rect 298020 4486 298048 336654
rect 298112 336462 298140 336790
rect 298100 336456 298152 336462
rect 298100 336398 298152 336404
rect 298204 335578 298232 338028
rect 298664 336734 298692 338028
rect 299046 338014 299244 338042
rect 298652 336728 298704 336734
rect 298652 336670 298704 336676
rect 298192 335572 298244 335578
rect 298192 335514 298244 335520
rect 299216 22778 299244 338014
rect 299388 336728 299440 336734
rect 299388 336670 299440 336676
rect 299296 335572 299348 335578
rect 299296 335514 299348 335520
rect 299204 22772 299256 22778
rect 299204 22714 299256 22720
rect 299308 14482 299336 335514
rect 299296 14476 299348 14482
rect 299296 14418 299348 14424
rect 299400 4554 299428 336670
rect 299492 336666 299520 338028
rect 299952 336734 299980 338028
rect 300426 338014 300624 338042
rect 299940 336728 299992 336734
rect 299940 336670 299992 336676
rect 299480 336660 299532 336666
rect 299480 336602 299532 336608
rect 300596 18630 300624 338014
rect 300872 336734 300900 338028
rect 300768 336728 300820 336734
rect 300768 336670 300820 336676
rect 300860 336728 300912 336734
rect 300860 336670 300912 336676
rect 300676 336660 300728 336666
rect 300676 336602 300728 336608
rect 300584 18624 300636 18630
rect 300584 18566 300636 18572
rect 299664 6248 299716 6254
rect 299664 6190 299716 6196
rect 299388 4548 299440 4554
rect 299388 4490 299440 4496
rect 298008 4480 298060 4486
rect 298008 4422 298060 4428
rect 296628 4412 296680 4418
rect 296628 4354 296680 4360
rect 297272 4140 297324 4146
rect 297272 4082 297324 4088
rect 297284 480 297312 4082
rect 298468 3392 298520 3398
rect 298468 3334 298520 3340
rect 298480 480 298508 3334
rect 299676 480 299704 6190
rect 300688 4690 300716 336602
rect 300676 4684 300728 4690
rect 300676 4626 300728 4632
rect 300780 4622 300808 336670
rect 301332 336666 301360 338028
rect 301320 336660 301372 336666
rect 301320 336602 301372 336608
rect 301792 330546 301820 338028
rect 302068 338014 302174 338042
rect 301964 336728 302016 336734
rect 301964 336670 302016 336676
rect 301780 330540 301832 330546
rect 301780 330482 301832 330488
rect 301976 4758 302004 336670
rect 302068 5438 302096 338014
rect 302148 336660 302200 336666
rect 302148 336602 302200 336608
rect 302160 5506 302188 336602
rect 302620 335714 302648 338028
rect 303094 338014 303384 338042
rect 302608 335708 302660 335714
rect 302608 335650 302660 335656
rect 303356 305658 303384 338014
rect 303448 338014 303554 338042
rect 303344 305652 303396 305658
rect 303344 305594 303396 305600
rect 302240 215960 302292 215966
rect 302240 215902 302292 215908
rect 302252 16574 302280 215902
rect 302252 16546 303200 16574
rect 302148 5500 302200 5506
rect 302148 5442 302200 5448
rect 302056 5432 302108 5438
rect 302056 5374 302108 5380
rect 301964 4752 302016 4758
rect 301964 4694 302016 4700
rect 300768 4616 300820 4622
rect 300768 4558 300820 4564
rect 300768 3936 300820 3942
rect 300768 3878 300820 3884
rect 300780 480 300808 3878
rect 301964 3868 302016 3874
rect 301964 3810 302016 3816
rect 301976 480 302004 3810
rect 303172 480 303200 16546
rect 303448 5302 303476 338014
rect 304000 336734 304028 338028
rect 303988 336728 304040 336734
rect 303988 336670 304040 336676
rect 304460 336666 304488 338028
rect 304724 336728 304776 336734
rect 304724 336670 304776 336676
rect 304448 336660 304500 336666
rect 304448 336602 304500 336608
rect 303528 335708 303580 335714
rect 303528 335650 303580 335656
rect 303540 5370 303568 335650
rect 304736 8022 304764 336670
rect 304724 8016 304776 8022
rect 304724 7958 304776 7964
rect 303528 5364 303580 5370
rect 303528 5306 303580 5312
rect 303436 5296 303488 5302
rect 303436 5238 303488 5244
rect 304828 5234 304856 338028
rect 305288 336734 305316 338028
rect 305276 336728 305328 336734
rect 305276 336670 305328 336676
rect 305748 336666 305776 338028
rect 306104 336728 306156 336734
rect 306104 336670 306156 336676
rect 304908 336660 304960 336666
rect 304908 336602 304960 336608
rect 305736 336660 305788 336666
rect 305736 336602 305788 336608
rect 304816 5228 304868 5234
rect 304816 5170 304868 5176
rect 304920 3942 304948 336602
rect 306116 7954 306144 336670
rect 306104 7948 306156 7954
rect 306104 7890 306156 7896
rect 306208 5166 306236 338028
rect 306668 336734 306696 338028
rect 306656 336728 306708 336734
rect 306656 336670 306708 336676
rect 307128 336666 307156 338028
rect 307510 338014 307616 338042
rect 307484 336728 307536 336734
rect 307484 336670 307536 336676
rect 306288 336660 306340 336666
rect 306288 336602 306340 336608
rect 307116 336660 307168 336666
rect 307116 336602 307168 336608
rect 306196 5160 306248 5166
rect 306196 5102 306248 5108
rect 304908 3936 304960 3942
rect 304908 3878 304960 3884
rect 306300 3874 306328 336602
rect 306380 218748 306432 218754
rect 306380 218690 306432 218696
rect 306392 16574 306420 218690
rect 306392 16546 306788 16574
rect 306288 3868 306340 3874
rect 306288 3810 306340 3816
rect 305552 3800 305604 3806
rect 305552 3742 305604 3748
rect 304356 3664 304408 3670
rect 304356 3606 304408 3612
rect 304368 480 304396 3606
rect 305564 480 305592 3742
rect 306760 480 306788 16546
rect 307496 7886 307524 336670
rect 307484 7880 307536 7886
rect 307484 7822 307536 7828
rect 307588 5098 307616 338014
rect 307956 336734 307984 338028
rect 307944 336728 307996 336734
rect 307944 336670 307996 336676
rect 308416 336666 308444 338028
rect 308890 338014 308996 338042
rect 308864 336728 308916 336734
rect 308864 336670 308916 336676
rect 307668 336660 307720 336666
rect 307668 336602 307720 336608
rect 308404 336660 308456 336666
rect 308404 336602 308456 336608
rect 307576 5092 307628 5098
rect 307576 5034 307628 5040
rect 307680 3670 307708 336602
rect 308876 7818 308904 336670
rect 308864 7812 308916 7818
rect 308864 7754 308916 7760
rect 308968 5030 308996 338014
rect 309336 336734 309364 338028
rect 309324 336728 309376 336734
rect 309324 336670 309376 336676
rect 309796 336666 309824 338028
rect 310178 338014 310376 338042
rect 310244 336728 310296 336734
rect 310244 336670 310296 336676
rect 309048 336660 309100 336666
rect 309048 336602 309100 336608
rect 309784 336660 309836 336666
rect 309784 336602 309836 336608
rect 308956 5024 309008 5030
rect 308956 4966 309008 4972
rect 309060 4842 309088 336602
rect 310256 16574 310284 336670
rect 310164 16546 310284 16574
rect 310164 7750 310192 16546
rect 310244 8968 310296 8974
rect 310244 8910 310296 8916
rect 310152 7744 310204 7750
rect 310152 7686 310204 7692
rect 308968 4814 309088 4842
rect 307668 3664 307720 3670
rect 307668 3606 307720 3612
rect 308968 3602 308996 4814
rect 309048 3732 309100 3738
rect 309048 3674 309100 3680
rect 307944 3596 307996 3602
rect 307944 3538 307996 3544
rect 308956 3596 309008 3602
rect 308956 3538 309008 3544
rect 307956 480 307984 3538
rect 309060 480 309088 3674
rect 310256 480 310284 8910
rect 310348 4962 310376 338014
rect 310624 336734 310652 338028
rect 310612 336728 310664 336734
rect 310612 336670 310664 336676
rect 311084 336666 311112 338028
rect 311558 338014 311756 338042
rect 311624 336728 311676 336734
rect 311624 336670 311676 336676
rect 310428 336660 310480 336666
rect 310428 336602 310480 336608
rect 311072 336660 311124 336666
rect 311072 336602 311124 336608
rect 310336 4956 310388 4962
rect 310336 4898 310388 4904
rect 310440 3670 310468 336602
rect 311636 7682 311664 336670
rect 311624 7676 311676 7682
rect 311624 7618 311676 7624
rect 311728 4894 311756 338014
rect 311808 336660 311860 336666
rect 311808 336602 311860 336608
rect 311716 4888 311768 4894
rect 311716 4830 311768 4836
rect 310428 3664 310480 3670
rect 310428 3606 310480 3612
rect 311820 3602 311848 336602
rect 312004 335918 312032 338028
rect 312464 336734 312492 338028
rect 312938 338014 313136 338042
rect 312452 336728 312504 336734
rect 312452 336670 312504 336676
rect 311992 335912 312044 335918
rect 311992 335854 312044 335860
rect 313004 335912 313056 335918
rect 313004 335854 313056 335860
rect 313016 7614 313044 335854
rect 313004 7608 313056 7614
rect 313004 7550 313056 7556
rect 313108 4826 313136 338014
rect 313292 336734 313320 338028
rect 313188 336728 313240 336734
rect 313188 336670 313240 336676
rect 313280 336728 313332 336734
rect 313280 336670 313332 336676
rect 313096 4820 313148 4826
rect 313096 4762 313148 4768
rect 311808 3596 311860 3602
rect 311808 3538 311860 3544
rect 313200 3534 313228 336670
rect 313752 336598 313780 338028
rect 313740 336592 313792 336598
rect 313740 336534 313792 336540
rect 313924 336252 313976 336258
rect 313924 336194 313976 336200
rect 313280 18692 313332 18698
rect 313280 18634 313332 18640
rect 313292 16574 313320 18634
rect 313292 16546 313872 16574
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 313188 3528 313240 3534
rect 313188 3470 313240 3476
rect 311440 3460 311492 3466
rect 311440 3402 311492 3408
rect 311452 480 311480 3402
rect 312648 480 312676 3470
rect 313844 480 313872 16546
rect 313936 5574 313964 336194
rect 314212 329186 314240 338028
rect 314672 336734 314700 338028
rect 314476 336728 314528 336734
rect 314476 336670 314528 336676
rect 314660 336728 314712 336734
rect 314660 336670 314712 336676
rect 314200 329180 314252 329186
rect 314200 329122 314252 329128
rect 313924 5568 313976 5574
rect 313924 5510 313976 5516
rect 314488 4214 314516 336670
rect 315132 336666 315160 338028
rect 315120 336660 315172 336666
rect 315120 336602 315172 336608
rect 314568 336592 314620 336598
rect 314568 336534 314620 336540
rect 314476 4208 314528 4214
rect 314476 4150 314528 4156
rect 314580 3466 314608 336534
rect 315592 336258 315620 338028
rect 315776 338014 315974 338042
rect 315580 336252 315632 336258
rect 315580 336194 315632 336200
rect 315776 7138 315804 338014
rect 316420 336734 316448 338028
rect 316894 338014 317184 338042
rect 315856 336728 315908 336734
rect 315856 336670 315908 336676
rect 316408 336728 316460 336734
rect 316408 336670 316460 336676
rect 315764 7132 315816 7138
rect 315764 7074 315816 7080
rect 315868 7070 315896 336670
rect 315948 336660 316000 336666
rect 315948 336602 316000 336608
rect 315856 7064 315908 7070
rect 315856 7006 315908 7012
rect 315028 5568 315080 5574
rect 315028 5510 315080 5516
rect 314568 3460 314620 3466
rect 314568 3402 314620 3408
rect 315040 480 315068 5510
rect 315960 2854 315988 336602
rect 316684 336388 316736 336394
rect 316684 336330 316736 336336
rect 316696 17950 316724 336330
rect 317156 327826 317184 338014
rect 317248 338014 317354 338042
rect 317814 338014 318196 338042
rect 318274 338014 318564 338042
rect 317144 327820 317196 327826
rect 317144 327762 317196 327768
rect 317248 324970 317276 338014
rect 317328 336728 317380 336734
rect 317328 336670 317380 336676
rect 317236 324964 317288 324970
rect 317236 324906 317288 324912
rect 316684 17944 316736 17950
rect 316684 17886 316736 17892
rect 317340 6914 317368 336670
rect 318064 336456 318116 336462
rect 318064 336398 318116 336404
rect 317696 336184 317748 336190
rect 317696 336126 317748 336132
rect 317248 6886 317368 6914
rect 317708 6914 317736 336126
rect 318076 10538 318104 336398
rect 318168 325694 318196 338014
rect 318536 326466 318564 338014
rect 318628 334694 318656 338028
rect 319088 336734 319116 338028
rect 319562 338014 319944 338042
rect 319076 336728 319128 336734
rect 319076 336670 319128 336676
rect 318616 334688 318668 334694
rect 318616 334630 318668 334636
rect 318524 326460 318576 326466
rect 318524 326402 318576 326408
rect 318168 325666 318564 325694
rect 318536 16574 318564 325666
rect 319916 322318 319944 338014
rect 319904 322312 319956 322318
rect 319904 322254 319956 322260
rect 320008 222902 320036 338028
rect 320468 336734 320496 338028
rect 320942 338014 321232 338042
rect 321310 338014 321416 338042
rect 320088 336728 320140 336734
rect 320088 336670 320140 336676
rect 320456 336728 320508 336734
rect 320456 336670 320508 336676
rect 319996 222896 320048 222902
rect 319996 222838 320048 222844
rect 318536 16546 318656 16574
rect 318064 10532 318116 10538
rect 318064 10474 318116 10480
rect 317708 6886 318472 6914
rect 316224 4072 316276 4078
rect 316224 4014 316276 4020
rect 315948 2848 316000 2854
rect 315948 2790 316000 2796
rect 316236 480 316264 4014
rect 317248 2922 317276 6886
rect 317328 6180 317380 6186
rect 317328 6122 317380 6128
rect 317236 2916 317288 2922
rect 317236 2858 317288 2864
rect 317340 480 317368 6122
rect 318444 3482 318472 6886
rect 318444 3454 318564 3482
rect 318536 480 318564 3454
rect 318628 2990 318656 16546
rect 319720 4004 319772 4010
rect 319720 3946 319772 3952
rect 318616 2984 318668 2990
rect 318616 2926 318668 2932
rect 319732 480 319760 3946
rect 320100 3058 320128 336670
rect 320824 336320 320876 336326
rect 320824 336262 320876 336268
rect 320732 10464 320784 10470
rect 320732 10406 320784 10412
rect 320744 3482 320772 10406
rect 320836 6186 320864 336262
rect 321204 335354 321232 338014
rect 321204 335326 321324 335354
rect 321296 320958 321324 335326
rect 321284 320952 321336 320958
rect 321284 320894 321336 320900
rect 321388 8430 321416 338014
rect 321468 336728 321520 336734
rect 321468 336670 321520 336676
rect 321376 8424 321428 8430
rect 321376 8366 321428 8372
rect 320824 6180 320876 6186
rect 320824 6122 320876 6128
rect 320744 3454 320956 3482
rect 320088 3052 320140 3058
rect 320088 2994 320140 3000
rect 320928 480 320956 3454
rect 321480 3126 321508 336670
rect 321756 336122 321784 338028
rect 322230 338014 322520 338042
rect 322690 338014 322796 338042
rect 321744 336116 321796 336122
rect 321744 336058 321796 336064
rect 322492 335354 322520 338014
rect 322492 335326 322704 335354
rect 322676 15910 322704 335326
rect 322112 15904 322164 15910
rect 322112 15846 322164 15852
rect 322664 15904 322716 15910
rect 322664 15846 322716 15852
rect 321468 3120 321520 3126
rect 321468 3062 321520 3068
rect 322124 480 322152 15846
rect 322768 8498 322796 338014
rect 323136 336666 323164 338028
rect 323610 338014 323992 338042
rect 324070 338014 324268 338042
rect 323124 336660 323176 336666
rect 323124 336602 323176 336608
rect 323584 336184 323636 336190
rect 323584 336126 323636 336132
rect 322848 336116 322900 336122
rect 322848 336058 322900 336064
rect 322756 8492 322808 8498
rect 322756 8434 322808 8440
rect 322860 3194 322888 336058
rect 322940 224256 322992 224262
rect 322940 224198 322992 224204
rect 322952 16574 322980 224198
rect 322952 16546 323348 16574
rect 322848 3188 322900 3194
rect 322848 3130 322900 3136
rect 323320 480 323348 16546
rect 323596 5574 323624 336126
rect 323964 335354 323992 338014
rect 323964 335326 324176 335354
rect 324148 323678 324176 335326
rect 324136 323672 324188 323678
rect 324136 323614 324188 323620
rect 324240 8566 324268 338014
rect 324424 336734 324452 338028
rect 324898 338014 325280 338042
rect 325358 338014 325556 338042
rect 324412 336728 324464 336734
rect 324412 336670 324464 336676
rect 325252 335354 325280 338014
rect 325252 335326 325464 335354
rect 324320 17944 324372 17950
rect 324320 17886 324372 17892
rect 324228 8560 324280 8566
rect 324228 8502 324280 8508
rect 323584 5568 323636 5574
rect 323584 5510 323636 5516
rect 324332 3398 324360 17886
rect 325436 17270 325464 335326
rect 325424 17264 325476 17270
rect 325424 17206 325476 17212
rect 325528 8634 325556 338014
rect 325608 336728 325660 336734
rect 325608 336670 325660 336676
rect 325516 8628 325568 8634
rect 325516 8570 325568 8576
rect 325620 6914 325648 336670
rect 325804 336462 325832 338028
rect 326278 338014 326568 338042
rect 326738 338014 327028 338042
rect 325792 336456 325844 336462
rect 325792 336398 325844 336404
rect 326540 335354 326568 338014
rect 326540 335326 326936 335354
rect 326908 319530 326936 335326
rect 326896 319524 326948 319530
rect 326896 319466 326948 319472
rect 326804 10396 326856 10402
rect 326804 10338 326856 10344
rect 325528 6886 325648 6914
rect 324412 5568 324464 5574
rect 324412 5510 324464 5516
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 5510
rect 325528 3262 325556 6886
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325516 3256 325568 3262
rect 325516 3198 325568 3204
rect 325620 480 325648 3334
rect 326816 480 326844 10338
rect 327000 8702 327028 338014
rect 327092 335850 327120 338028
rect 327552 336734 327580 338028
rect 328026 338014 328224 338042
rect 327540 336728 327592 336734
rect 327540 336670 327592 336676
rect 327080 335844 327132 335850
rect 327080 335786 327132 335792
rect 328000 11824 328052 11830
rect 328000 11766 328052 11772
rect 326988 8696 327040 8702
rect 326988 8638 327040 8644
rect 328012 480 328040 11766
rect 328196 8770 328224 338014
rect 328276 336728 328328 336734
rect 328276 336670 328328 336676
rect 328184 8764 328236 8770
rect 328184 8706 328236 8712
rect 328288 5710 328316 336670
rect 328472 336598 328500 338028
rect 328932 336734 328960 338028
rect 329406 338014 329604 338042
rect 328920 336728 328972 336734
rect 328920 336670 328972 336676
rect 328460 336592 328512 336598
rect 328460 336534 328512 336540
rect 328552 336048 328604 336054
rect 328552 335990 328604 335996
rect 328368 335844 328420 335850
rect 328368 335786 328420 335792
rect 328276 5704 328328 5710
rect 328276 5646 328328 5652
rect 328380 4010 328408 335786
rect 328564 16574 328592 335990
rect 328564 16546 329236 16574
rect 328368 4004 328420 4010
rect 328368 3946 328420 3952
rect 329208 480 329236 16546
rect 329576 8838 329604 338014
rect 329656 336728 329708 336734
rect 329656 336670 329708 336676
rect 329564 8832 329616 8838
rect 329564 8774 329616 8780
rect 329668 5778 329696 336670
rect 329656 5772 329708 5778
rect 329656 5714 329708 5720
rect 329760 3330 329788 338028
rect 330220 336734 330248 338028
rect 330694 338014 331076 338042
rect 330208 336728 330260 336734
rect 330208 336670 330260 336676
rect 329840 19984 329892 19990
rect 329840 19926 329892 19932
rect 329852 16574 329880 19926
rect 329852 16546 330432 16574
rect 329748 3324 329800 3330
rect 329748 3266 329800 3272
rect 330404 480 330432 16546
rect 331048 8906 331076 338014
rect 331140 336818 331168 338028
rect 331140 336790 331260 336818
rect 331128 336728 331180 336734
rect 331128 336670 331180 336676
rect 331036 8900 331088 8906
rect 331036 8842 331088 8848
rect 331140 5846 331168 336670
rect 331232 336530 331260 336790
rect 331600 336734 331628 338028
rect 332074 338014 332364 338042
rect 332442 338014 332548 338042
rect 331588 336728 331640 336734
rect 331588 336670 331640 336676
rect 331220 336524 331272 336530
rect 331220 336466 331272 336472
rect 331220 217320 331272 217326
rect 331220 217262 331272 217268
rect 331232 16574 331260 217262
rect 331232 16546 331628 16574
rect 331128 5840 331180 5846
rect 331128 5782 331180 5788
rect 331600 480 331628 16546
rect 332336 9654 332364 338014
rect 332416 336728 332468 336734
rect 332416 336670 332468 336676
rect 332324 9648 332376 9654
rect 332324 9590 332376 9596
rect 332428 5914 332456 336670
rect 332416 5908 332468 5914
rect 332416 5850 332468 5856
rect 332520 4146 332548 338014
rect 332888 336734 332916 338028
rect 333362 338014 333744 338042
rect 332876 336728 332928 336734
rect 332876 336670 332928 336676
rect 333716 335354 333744 338014
rect 333808 336394 333836 338028
rect 334268 336734 334296 338028
rect 334742 338014 335124 338042
rect 335202 338014 335308 338042
rect 333888 336728 333940 336734
rect 333888 336670 333940 336676
rect 334256 336728 334308 336734
rect 334256 336670 334308 336676
rect 333796 336388 333848 336394
rect 333796 336330 333848 336336
rect 333716 335326 333836 335354
rect 332600 11756 332652 11762
rect 332600 11698 332652 11704
rect 332508 4140 332560 4146
rect 332508 4082 332560 4088
rect 332612 3398 332640 11698
rect 333808 9586 333836 335326
rect 333796 9580 333848 9586
rect 333796 9522 333848 9528
rect 332692 6180 332744 6186
rect 332692 6122 332744 6128
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 6122
rect 333900 5982 333928 336670
rect 334992 13116 335044 13122
rect 334992 13058 335044 13064
rect 335004 6914 335032 13058
rect 335096 9518 335124 338014
rect 335176 336728 335228 336734
rect 335176 336670 335228 336676
rect 335084 9512 335136 9518
rect 335084 9454 335136 9460
rect 335004 6886 335124 6914
rect 333888 5976 333940 5982
rect 333888 5918 333940 5924
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 335096 480 335124 6886
rect 335188 6050 335216 336670
rect 335176 6044 335228 6050
rect 335176 5986 335228 5992
rect 335280 4078 335308 338014
rect 335556 336734 335584 338028
rect 336030 338014 336320 338042
rect 335544 336728 335596 336734
rect 335544 336670 335596 336676
rect 336004 336252 336056 336258
rect 336004 336194 336056 336200
rect 336016 13190 336044 336194
rect 336292 335354 336320 338014
rect 336476 336054 336504 338028
rect 336936 336734 336964 338028
rect 337410 338014 337792 338042
rect 337870 338014 338068 338042
rect 336648 336728 336700 336734
rect 336648 336670 336700 336676
rect 336924 336728 336976 336734
rect 336924 336670 336976 336676
rect 336464 336048 336516 336054
rect 336464 335990 336516 335996
rect 336292 335326 336596 335354
rect 336004 13184 336056 13190
rect 336004 13126 336056 13132
rect 336568 9450 336596 335326
rect 336556 9444 336608 9450
rect 336556 9386 336608 9392
rect 336660 6118 336688 336670
rect 337764 335354 337792 338014
rect 337936 336728 337988 336734
rect 337936 336670 337988 336676
rect 337764 335326 337884 335354
rect 337476 10328 337528 10334
rect 337476 10270 337528 10276
rect 336648 6112 336700 6118
rect 336648 6054 336700 6060
rect 336280 4344 336332 4350
rect 336280 4286 336332 4292
rect 335268 4072 335320 4078
rect 335268 4014 335320 4020
rect 336292 480 336320 4286
rect 337488 480 337516 10270
rect 337856 9382 337884 335326
rect 337844 9376 337896 9382
rect 337844 9318 337896 9324
rect 337948 6866 337976 336670
rect 337936 6860 337988 6866
rect 337936 6802 337988 6808
rect 338040 4010 338068 338014
rect 338224 336734 338252 338028
rect 338698 338014 339080 338042
rect 338212 336728 338264 336734
rect 338212 336670 338264 336676
rect 339052 335354 339080 338014
rect 339144 336122 339172 338028
rect 339604 336734 339632 338028
rect 340078 338014 340368 338042
rect 340538 338014 340828 338042
rect 339408 336728 339460 336734
rect 339408 336670 339460 336676
rect 339592 336728 339644 336734
rect 339592 336670 339644 336676
rect 339132 336116 339184 336122
rect 339132 336058 339184 336064
rect 339052 335326 339356 335354
rect 338120 220108 338172 220114
rect 338120 220050 338172 220056
rect 338132 16574 338160 220050
rect 338132 16546 338712 16574
rect 338028 4004 338080 4010
rect 338028 3946 338080 3952
rect 338684 480 338712 16546
rect 339328 9314 339356 335326
rect 339316 9308 339368 9314
rect 339316 9250 339368 9256
rect 339420 6798 339448 336670
rect 340340 335354 340368 338014
rect 340696 336728 340748 336734
rect 340696 336670 340748 336676
rect 340340 335326 340644 335354
rect 340616 9246 340644 335326
rect 340604 9240 340656 9246
rect 340604 9182 340656 9188
rect 339408 6792 339460 6798
rect 339408 6734 339460 6740
rect 340708 6730 340736 336670
rect 340696 6724 340748 6730
rect 340696 6666 340748 6672
rect 339868 4412 339920 4418
rect 339868 4354 339920 4360
rect 339880 480 339908 4354
rect 340800 3777 340828 338014
rect 340892 336734 340920 338028
rect 340880 336728 340932 336734
rect 340880 336670 340932 336676
rect 341352 336258 341380 338028
rect 341340 336252 341392 336258
rect 341340 336194 341392 336200
rect 341812 335986 341840 338028
rect 342168 336728 342220 336734
rect 342168 336670 342220 336676
rect 342076 336252 342128 336258
rect 342076 336194 342128 336200
rect 341800 335980 341852 335986
rect 341800 335922 341852 335928
rect 340880 221468 340932 221474
rect 340880 221410 340932 221416
rect 340892 4010 340920 221410
rect 340972 21412 341024 21418
rect 340972 21354 341024 21360
rect 340880 4004 340932 4010
rect 340880 3946 340932 3952
rect 340786 3768 340842 3777
rect 340786 3703 340842 3712
rect 340984 480 341012 21354
rect 342088 9178 342116 336194
rect 342076 9172 342128 9178
rect 342076 9114 342128 9120
rect 342180 6662 342208 336670
rect 342272 336530 342300 338028
rect 342746 338014 343128 338042
rect 342260 336524 342312 336530
rect 342260 336466 342312 336472
rect 343100 325694 343128 338014
rect 343192 336734 343220 338028
rect 343376 338014 343574 338042
rect 343180 336728 343232 336734
rect 343180 336670 343232 336676
rect 343100 325666 343312 325694
rect 343284 9110 343312 325666
rect 343272 9104 343324 9110
rect 343272 9046 343324 9052
rect 342168 6656 342220 6662
rect 342168 6598 342220 6604
rect 343376 6526 343404 338014
rect 343548 336728 343600 336734
rect 343548 336670 343600 336676
rect 343456 336524 343508 336530
rect 343456 336466 343508 336472
rect 343468 6594 343496 336466
rect 343456 6588 343508 6594
rect 343456 6530 343508 6536
rect 343364 6520 343416 6526
rect 343364 6462 343416 6468
rect 343364 4480 343416 4486
rect 343364 4422 343416 4428
rect 342168 4004 342220 4010
rect 342168 3946 342220 3952
rect 342180 480 342208 3946
rect 343376 480 343404 4422
rect 343560 3641 343588 336670
rect 344020 335918 344048 338028
rect 344480 336122 344508 338028
rect 344468 336116 344520 336122
rect 344468 336058 344520 336064
rect 344008 335912 344060 335918
rect 344008 335854 344060 335860
rect 344836 335912 344888 335918
rect 344836 335854 344888 335860
rect 344560 10532 344612 10538
rect 344560 10474 344612 10480
rect 343546 3632 343602 3641
rect 343546 3567 343602 3576
rect 344572 480 344600 10474
rect 344848 9042 344876 335854
rect 344836 9036 344888 9042
rect 344836 8978 344888 8984
rect 344940 6458 344968 338028
rect 345400 336734 345428 338028
rect 345388 336728 345440 336734
rect 345388 336670 345440 336676
rect 345860 336054 345888 338028
rect 346228 338014 346334 338042
rect 346124 336728 346176 336734
rect 346124 336670 346176 336676
rect 345848 336048 345900 336054
rect 345848 335990 345900 335996
rect 345756 14476 345808 14482
rect 345756 14418 345808 14424
rect 344928 6452 344980 6458
rect 344928 6394 344980 6400
rect 345768 480 345796 14418
rect 346136 8974 346164 336670
rect 346124 8968 346176 8974
rect 346124 8910 346176 8916
rect 346228 6390 346256 338014
rect 346308 336048 346360 336054
rect 346308 335990 346360 335996
rect 346216 6384 346268 6390
rect 346216 6326 346268 6332
rect 346320 3505 346348 335990
rect 346688 335442 346716 338028
rect 347148 335986 347176 338028
rect 347622 338014 347728 338042
rect 347136 335980 347188 335986
rect 347136 335922 347188 335928
rect 346676 335436 346728 335442
rect 346676 335378 346728 335384
rect 347596 335436 347648 335442
rect 347596 335378 347648 335384
rect 347608 21418 347636 335378
rect 347596 21412 347648 21418
rect 347596 21354 347648 21360
rect 347700 6322 347728 338014
rect 348068 336734 348096 338028
rect 348056 336728 348108 336734
rect 348056 336670 348108 336676
rect 348528 336054 348556 338028
rect 348884 336728 348936 336734
rect 348884 336670 348936 336676
rect 348516 336048 348568 336054
rect 348516 335990 348568 335996
rect 348896 311166 348924 336670
rect 348884 311160 348936 311166
rect 348884 311102 348936 311108
rect 347780 22772 347832 22778
rect 347780 22714 347832 22720
rect 347792 16574 347820 22714
rect 347792 16546 348096 16574
rect 347688 6316 347740 6322
rect 347688 6258 347740 6264
rect 346952 4412 347004 4418
rect 346952 4354 347004 4360
rect 346306 3496 346362 3505
rect 346306 3431 346362 3440
rect 346964 480 346992 4354
rect 348068 480 348096 16546
rect 348988 11762 349016 338028
rect 349068 336048 349120 336054
rect 349068 335990 349120 335996
rect 348976 11756 349028 11762
rect 348976 11698 349028 11704
rect 349080 3369 349108 335990
rect 349356 335442 349384 338028
rect 349830 338014 350212 338042
rect 350290 338014 350488 338042
rect 350184 336682 350212 338014
rect 350184 336654 350396 336682
rect 349344 335436 349396 335442
rect 349344 335378 349396 335384
rect 350264 335436 350316 335442
rect 350264 335378 350316 335384
rect 350276 6254 350304 335378
rect 350368 308446 350396 336654
rect 350460 334626 350488 338014
rect 350736 336734 350764 338028
rect 351210 338014 351592 338042
rect 351670 338014 351776 338042
rect 350724 336728 350776 336734
rect 350724 336670 350776 336676
rect 350448 334620 350500 334626
rect 350448 334562 350500 334568
rect 351564 327758 351592 338014
rect 351552 327752 351604 327758
rect 351552 327694 351604 327700
rect 350356 308440 350408 308446
rect 350356 308382 350408 308388
rect 351748 217326 351776 338014
rect 352024 336734 352052 338028
rect 352498 338014 352880 338042
rect 351828 336728 351880 336734
rect 351828 336670 351880 336676
rect 352012 336728 352064 336734
rect 352012 336670 352064 336676
rect 351736 217320 351788 217326
rect 351736 217262 351788 217268
rect 350540 18624 350592 18630
rect 350540 18566 350592 18572
rect 350552 16574 350580 18566
rect 350552 16546 351684 16574
rect 350264 6248 350316 6254
rect 350264 6190 350316 6196
rect 349252 4684 349304 4690
rect 349252 4626 349304 4632
rect 349066 3360 349122 3369
rect 349066 3295 349122 3304
rect 349264 480 349292 4626
rect 350448 4616 350500 4622
rect 350448 4558 350500 4564
rect 350460 480 350488 4558
rect 351656 480 351684 16546
rect 351840 6186 351868 336670
rect 352852 325694 352880 338014
rect 352944 333334 352972 338028
rect 353116 336728 353168 336734
rect 353116 336670 353168 336676
rect 352932 333328 352984 333334
rect 352932 333270 352984 333276
rect 352852 325666 353064 325694
rect 353036 22778 353064 325666
rect 353128 318102 353156 336670
rect 353404 336054 353432 338028
rect 353878 338014 354260 338042
rect 354338 338014 354628 338042
rect 353392 336048 353444 336054
rect 353392 335990 353444 335996
rect 354232 326398 354260 338014
rect 354496 336048 354548 336054
rect 354496 335990 354548 335996
rect 354220 326392 354272 326398
rect 354220 326334 354272 326340
rect 353116 318096 353168 318102
rect 353116 318038 353168 318044
rect 353024 22772 353076 22778
rect 353024 22714 353076 22720
rect 354508 14482 354536 335990
rect 354496 14476 354548 14482
rect 354496 14418 354548 14424
rect 354600 10334 354628 338014
rect 354692 335918 354720 338028
rect 355152 336734 355180 338028
rect 355626 338014 356008 338042
rect 355140 336728 355192 336734
rect 355140 336670 355192 336676
rect 355876 336728 355928 336734
rect 355876 336670 355928 336676
rect 354680 335912 354732 335918
rect 354680 335854 354732 335860
rect 355784 335912 355836 335918
rect 355784 335854 355836 335860
rect 354680 330540 354732 330546
rect 354680 330482 354732 330488
rect 354692 16574 354720 330482
rect 355796 316742 355824 335854
rect 355784 316736 355836 316742
rect 355784 316678 355836 316684
rect 355888 309806 355916 336670
rect 355876 309800 355928 309806
rect 355876 309742 355928 309748
rect 355980 215966 356008 338014
rect 356072 336734 356100 338028
rect 356546 338014 356928 338042
rect 356060 336728 356112 336734
rect 356060 336670 356112 336676
rect 356900 325694 356928 338014
rect 356992 331974 357020 338028
rect 357348 336728 357400 336734
rect 357348 336670 357400 336676
rect 356980 331968 357032 331974
rect 356980 331910 357032 331916
rect 356900 325666 357296 325694
rect 357268 307086 357296 325666
rect 357256 307080 357308 307086
rect 357256 307022 357308 307028
rect 355968 215960 356020 215966
rect 355968 215902 356020 215908
rect 354692 16546 355272 16574
rect 354588 10328 354640 10334
rect 354588 10270 354640 10276
rect 351828 6180 351880 6186
rect 351828 6122 351880 6128
rect 354036 5500 354088 5506
rect 354036 5442 354088 5448
rect 352840 4752 352892 4758
rect 352840 4694 352892 4700
rect 352852 480 352880 4694
rect 354048 480 354076 5442
rect 355244 480 355272 16546
rect 357360 13122 357388 336670
rect 357452 329118 357480 338028
rect 357820 336734 357848 338028
rect 357808 336728 357860 336734
rect 357808 336670 357860 336676
rect 358280 335918 358308 338028
rect 358556 338014 358754 338042
rect 358268 335912 358320 335918
rect 358268 335854 358320 335860
rect 357440 329112 357492 329118
rect 357440 329054 357492 329060
rect 358556 315314 358584 338014
rect 359200 336734 359228 338028
rect 358636 336728 358688 336734
rect 358636 336670 358688 336676
rect 359188 336728 359240 336734
rect 359188 336670 359240 336676
rect 358544 315308 358596 315314
rect 358544 315250 358596 315256
rect 358648 305658 358676 336670
rect 358728 335912 358780 335918
rect 358728 335854 358780 335860
rect 357440 305652 357492 305658
rect 357440 305594 357492 305600
rect 358636 305652 358688 305658
rect 358636 305594 358688 305600
rect 357348 13116 357400 13122
rect 357348 13058 357400 13064
rect 356336 5432 356388 5438
rect 356336 5374 356388 5380
rect 356348 480 356376 5374
rect 357452 3942 357480 305594
rect 358740 42090 358768 335854
rect 359660 330546 359688 338028
rect 360016 336728 360068 336734
rect 360016 336670 360068 336676
rect 359648 330540 359700 330546
rect 359648 330482 359700 330488
rect 358728 42084 358780 42090
rect 358728 42026 358780 42032
rect 360028 24138 360056 336670
rect 360016 24132 360068 24138
rect 360016 24074 360068 24080
rect 360120 18630 360148 338028
rect 360488 336734 360516 338028
rect 360476 336728 360528 336734
rect 360476 336670 360528 336676
rect 360948 335986 360976 338028
rect 361316 338014 361422 338042
rect 360936 335980 360988 335986
rect 360936 335922 360988 335928
rect 361316 313954 361344 338014
rect 361868 336734 361896 338028
rect 361396 336728 361448 336734
rect 361396 336670 361448 336676
rect 361856 336728 361908 336734
rect 361856 336670 361908 336676
rect 361304 313948 361356 313954
rect 361304 313890 361356 313896
rect 361408 302938 361436 336670
rect 361488 335980 361540 335986
rect 361488 335922 361540 335928
rect 361396 302932 361448 302938
rect 361396 302874 361448 302880
rect 360108 18624 360160 18630
rect 360108 18566 360160 18572
rect 361120 8016 361172 8022
rect 361120 7958 361172 7964
rect 357532 5364 357584 5370
rect 357532 5306 357584 5312
rect 357440 3936 357492 3942
rect 357440 3878 357492 3884
rect 357544 480 357572 5306
rect 359924 5296 359976 5302
rect 359924 5238 359976 5244
rect 358728 3936 358780 3942
rect 358728 3878 358780 3884
rect 358740 480 358768 3878
rect 359936 480 359964 5238
rect 361132 480 361160 7958
rect 361500 4282 361528 335922
rect 362328 335646 362356 338028
rect 362684 336728 362736 336734
rect 362684 336670 362736 336676
rect 362316 335640 362368 335646
rect 362316 335582 362368 335588
rect 362696 322250 362724 336670
rect 362684 322244 362736 322250
rect 362684 322186 362736 322192
rect 362788 220114 362816 338028
rect 363156 336734 363184 338028
rect 363144 336728 363196 336734
rect 363144 336670 363196 336676
rect 363616 335986 363644 338028
rect 364090 338014 364196 338042
rect 364064 336728 364116 336734
rect 364064 336670 364116 336676
rect 363604 335980 363656 335986
rect 363604 335922 363656 335928
rect 362868 335640 362920 335646
rect 362868 335582 362920 335588
rect 362776 220108 362828 220114
rect 362776 220050 362828 220056
rect 362880 4350 362908 335582
rect 364076 320890 364104 336670
rect 364064 320884 364116 320890
rect 364064 320826 364116 320832
rect 364168 7206 364196 338014
rect 364536 336734 364564 338028
rect 364524 336728 364576 336734
rect 364524 336670 364576 336676
rect 364996 335986 365024 338028
rect 365470 338014 365576 338042
rect 365444 336728 365496 336734
rect 365444 336670 365496 336676
rect 364248 335980 364300 335986
rect 364248 335922 364300 335928
rect 364984 335980 365036 335986
rect 364984 335922 365036 335928
rect 364156 7200 364208 7206
rect 364156 7142 364208 7148
rect 363512 5228 363564 5234
rect 363512 5170 363564 5176
rect 362868 4344 362920 4350
rect 362868 4286 362920 4292
rect 361488 4276 361540 4282
rect 361488 4218 361540 4224
rect 362316 3936 362368 3942
rect 362316 3878 362368 3884
rect 362328 480 362356 3878
rect 363524 480 363552 5170
rect 364260 4418 364288 335922
rect 365456 323610 365484 336670
rect 365444 323604 365496 323610
rect 365444 323546 365496 323552
rect 364616 7948 364668 7954
rect 364616 7890 364668 7896
rect 364248 4412 364300 4418
rect 364248 4354 364300 4360
rect 364628 480 364656 7890
rect 365548 7274 365576 338014
rect 365824 336734 365852 338028
rect 365812 336728 365864 336734
rect 365812 336670 365864 336676
rect 366284 335986 366312 338028
rect 366758 338014 366956 338042
rect 366824 336728 366876 336734
rect 366824 336670 366876 336676
rect 365628 335980 365680 335986
rect 365628 335922 365680 335928
rect 366272 335980 366324 335986
rect 366272 335922 366324 335928
rect 365536 7268 365588 7274
rect 365536 7210 365588 7216
rect 365640 4486 365668 335922
rect 366836 304298 366864 336670
rect 366824 304292 366876 304298
rect 366824 304234 366876 304240
rect 366928 7342 366956 338014
rect 367204 336734 367232 338028
rect 367192 336728 367244 336734
rect 367192 336670 367244 336676
rect 367664 335986 367692 338028
rect 368138 338014 368336 338042
rect 368204 336728 368256 336734
rect 368204 336670 368256 336676
rect 367008 335980 367060 335986
rect 367008 335922 367060 335928
rect 367652 335980 367704 335986
rect 367652 335922 367704 335928
rect 366916 7336 366968 7342
rect 366916 7278 366968 7284
rect 367020 6914 367048 335922
rect 368216 301510 368244 336670
rect 368204 301504 368256 301510
rect 368204 301446 368256 301452
rect 368204 7880 368256 7886
rect 368204 7822 368256 7828
rect 366928 6886 367048 6914
rect 366928 4554 366956 6886
rect 367008 5160 367060 5166
rect 367008 5102 367060 5108
rect 366916 4548 366968 4554
rect 366916 4490 366968 4496
rect 365628 4480 365680 4486
rect 365628 4422 365680 4428
rect 365812 3868 365864 3874
rect 365812 3810 365864 3816
rect 365824 480 365852 3810
rect 367020 480 367048 5102
rect 368216 480 368244 7822
rect 368308 7410 368336 338014
rect 368584 335986 368612 338028
rect 368952 336734 368980 338028
rect 369426 338014 369716 338042
rect 368940 336728 368992 336734
rect 368940 336670 368992 336676
rect 368388 335980 368440 335986
rect 368388 335922 368440 335928
rect 368572 335980 368624 335986
rect 368572 335922 368624 335928
rect 369584 335980 369636 335986
rect 369584 335922 369636 335928
rect 368296 7404 368348 7410
rect 368296 7346 368348 7352
rect 368400 4622 368428 335922
rect 369596 297430 369624 335922
rect 369584 297424 369636 297430
rect 369584 297366 369636 297372
rect 369688 7478 369716 338014
rect 369872 336734 369900 338028
rect 369768 336728 369820 336734
rect 369768 336670 369820 336676
rect 369860 336728 369912 336734
rect 369860 336670 369912 336676
rect 369676 7472 369728 7478
rect 369676 7414 369728 7420
rect 369780 4690 369808 336670
rect 370332 335986 370360 338028
rect 370806 338014 371096 338042
rect 370964 336728 371016 336734
rect 370964 336670 371016 336676
rect 370320 335980 370372 335986
rect 370320 335922 370372 335928
rect 370976 319462 371004 336670
rect 370964 319456 371016 319462
rect 370964 319398 371016 319404
rect 371068 7546 371096 338014
rect 371148 335980 371200 335986
rect 371148 335922 371200 335928
rect 371056 7540 371108 7546
rect 371056 7482 371108 7488
rect 370596 5092 370648 5098
rect 370596 5034 370648 5040
rect 369768 4684 369820 4690
rect 369768 4626 369820 4632
rect 368388 4616 368440 4622
rect 368388 4558 368440 4564
rect 369400 3800 369452 3806
rect 369400 3742 369452 3748
rect 369412 480 369440 3742
rect 370608 480 370636 5034
rect 371160 4758 371188 335922
rect 371252 333198 371280 338028
rect 371634 338014 372016 338042
rect 371240 333192 371292 333198
rect 371240 333134 371292 333140
rect 371988 325694 372016 338014
rect 372080 336734 372108 338028
rect 372356 338014 372554 338042
rect 373014 338014 373304 338042
rect 372068 336728 372120 336734
rect 372068 336670 372120 336676
rect 371988 325666 372292 325694
rect 371700 7812 371752 7818
rect 371700 7754 371752 7760
rect 371148 4752 371200 4758
rect 371148 4694 371200 4700
rect 371712 480 371740 7754
rect 372264 5506 372292 325666
rect 372356 300150 372384 338014
rect 372436 336728 372488 336734
rect 372436 336670 372488 336676
rect 372344 300144 372396 300150
rect 372344 300086 372396 300092
rect 372448 8294 372476 336670
rect 373276 330750 373304 338014
rect 373460 336734 373488 338028
rect 373736 338014 373934 338042
rect 373448 336728 373500 336734
rect 373448 336670 373500 336676
rect 373264 330744 373316 330750
rect 373264 330686 373316 330692
rect 373736 296002 373764 338014
rect 373816 336728 373868 336734
rect 373816 336670 373868 336676
rect 373724 295996 373776 296002
rect 373724 295938 373776 295944
rect 372436 8288 372488 8294
rect 372436 8230 372488 8236
rect 373828 8226 373856 336670
rect 374288 335578 374316 338028
rect 374748 336734 374776 338028
rect 375116 338014 375222 338042
rect 374736 336728 374788 336734
rect 374736 336670 374788 336676
rect 374276 335572 374328 335578
rect 374276 335514 374328 335520
rect 373908 330744 373960 330750
rect 373908 330686 373960 330692
rect 373816 8220 373868 8226
rect 373816 8162 373868 8168
rect 372252 5500 372304 5506
rect 372252 5442 372304 5448
rect 373920 5438 373948 330686
rect 375116 293282 375144 338014
rect 375668 336734 375696 338028
rect 375196 336728 375248 336734
rect 375196 336670 375248 336676
rect 375656 336728 375708 336734
rect 375656 336670 375708 336676
rect 375104 293276 375156 293282
rect 375104 293218 375156 293224
rect 375208 8158 375236 336670
rect 376128 335646 376156 338028
rect 376496 338014 376602 338042
rect 376116 335640 376168 335646
rect 376116 335582 376168 335588
rect 375288 335572 375340 335578
rect 375288 335514 375340 335520
rect 375196 8152 375248 8158
rect 375196 8094 375248 8100
rect 375196 7744 375248 7750
rect 375196 7686 375248 7692
rect 373908 5432 373960 5438
rect 373908 5374 373960 5380
rect 374092 5024 374144 5030
rect 374092 4966 374144 4972
rect 372896 3732 372948 3738
rect 372896 3674 372948 3680
rect 372908 480 372936 3674
rect 374104 480 374132 4966
rect 375208 3482 375236 7686
rect 375300 5370 375328 335514
rect 376496 294642 376524 338014
rect 376956 336734 376984 338028
rect 377430 338014 377812 338042
rect 376668 336728 376720 336734
rect 376668 336670 376720 336676
rect 376944 336728 376996 336734
rect 376944 336670 376996 336676
rect 376576 335640 376628 335646
rect 376576 335582 376628 335588
rect 376484 294636 376536 294642
rect 376484 294578 376536 294584
rect 376588 8090 376616 335582
rect 376576 8084 376628 8090
rect 376576 8026 376628 8032
rect 375288 5364 375340 5370
rect 375288 5306 375340 5312
rect 376680 5302 376708 336670
rect 377784 325694 377812 338014
rect 377876 331906 377904 338028
rect 378048 336728 378100 336734
rect 378048 336670 378100 336676
rect 377864 331900 377916 331906
rect 377864 331842 377916 331848
rect 377784 325666 377996 325694
rect 377968 8022 377996 325666
rect 377956 8016 378008 8022
rect 377956 7958 378008 7964
rect 376668 5296 376720 5302
rect 376668 5238 376720 5244
rect 378060 5234 378088 336670
rect 378336 335986 378364 338028
rect 378796 336734 378824 338028
rect 378784 336728 378836 336734
rect 378784 336670 378836 336676
rect 378324 335980 378376 335986
rect 378324 335922 378376 335928
rect 379256 291854 379284 338028
rect 379336 336728 379388 336734
rect 379336 336670 379388 336676
rect 379244 291848 379296 291854
rect 379244 291790 379296 291796
rect 379348 7954 379376 336670
rect 379716 335986 379744 338028
rect 380084 336734 380112 338028
rect 380558 338014 380664 338042
rect 380072 336728 380124 336734
rect 380072 336670 380124 336676
rect 379428 335980 379480 335986
rect 379428 335922 379480 335928
rect 379704 335980 379756 335986
rect 379704 335922 379756 335928
rect 379336 7948 379388 7954
rect 379336 7890 379388 7896
rect 378876 7676 378928 7682
rect 378876 7618 378928 7624
rect 378048 5228 378100 5234
rect 378048 5170 378100 5176
rect 377680 4956 377732 4962
rect 377680 4898 377732 4904
rect 376484 3664 376536 3670
rect 376484 3606 376536 3612
rect 375208 3454 375328 3482
rect 375300 480 375328 3454
rect 376496 480 376524 3606
rect 377692 480 377720 4898
rect 378888 480 378916 7618
rect 379440 5166 379468 335922
rect 380636 290494 380664 338014
rect 381004 336734 381032 338028
rect 381478 338014 381768 338042
rect 381938 338014 382228 338042
rect 380716 336728 380768 336734
rect 380716 336670 380768 336676
rect 380992 336728 381044 336734
rect 380992 336670 381044 336676
rect 380624 290488 380676 290494
rect 380624 290430 380676 290436
rect 380728 7886 380756 336670
rect 380808 335980 380860 335986
rect 380808 335922 380860 335928
rect 380716 7880 380768 7886
rect 380716 7822 380768 7828
rect 379428 5160 379480 5166
rect 379428 5102 379480 5108
rect 380820 5098 380848 335922
rect 381740 335354 381768 338014
rect 382096 336728 382148 336734
rect 382096 336670 382148 336676
rect 381740 335326 382044 335354
rect 382016 7818 382044 335326
rect 382004 7812 382056 7818
rect 382004 7754 382056 7760
rect 380808 5092 380860 5098
rect 380808 5034 380860 5040
rect 382108 5030 382136 336670
rect 382096 5024 382148 5030
rect 382096 4966 382148 4972
rect 381176 4888 381228 4894
rect 381176 4830 381228 4836
rect 379980 3596 380032 3602
rect 379980 3538 380032 3544
rect 379992 480 380020 3538
rect 381188 480 381216 4830
rect 382200 3942 382228 338014
rect 382384 335918 382412 338028
rect 382766 338014 383056 338042
rect 383226 338014 383608 338042
rect 382372 335912 382424 335918
rect 382372 335854 382424 335860
rect 383028 335354 383056 338014
rect 383476 335912 383528 335918
rect 383476 335854 383528 335860
rect 383028 335326 383424 335354
rect 383396 7750 383424 335326
rect 383384 7744 383436 7750
rect 383384 7686 383436 7692
rect 382372 7608 382424 7614
rect 382372 7550 382424 7556
rect 382188 3936 382240 3942
rect 382188 3878 382240 3884
rect 382384 480 382412 7550
rect 383488 4962 383516 335854
rect 383476 4956 383528 4962
rect 383476 4898 383528 4904
rect 383580 3874 383608 338014
rect 383672 336734 383700 338028
rect 384146 338014 384528 338042
rect 384606 338014 384988 338042
rect 383660 336728 383712 336734
rect 383660 336670 383712 336676
rect 384500 335354 384528 338014
rect 384856 336728 384908 336734
rect 384856 336670 384908 336676
rect 384500 335326 384804 335354
rect 384776 7682 384804 335326
rect 384764 7676 384816 7682
rect 384764 7618 384816 7624
rect 384868 4894 384896 336670
rect 384856 4888 384908 4894
rect 384856 4830 384908 4836
rect 384764 4820 384816 4826
rect 384764 4762 384816 4768
rect 383568 3868 383620 3874
rect 383568 3810 383620 3816
rect 383568 3528 383620 3534
rect 383568 3470 383620 3476
rect 383580 480 383608 3470
rect 384776 480 384804 4762
rect 384960 3806 384988 338014
rect 385052 335986 385080 338028
rect 385434 338014 385816 338042
rect 385040 335980 385092 335986
rect 385040 335922 385092 335928
rect 385788 325694 385816 338014
rect 385880 336734 385908 338028
rect 386248 338014 386354 338042
rect 385868 336728 385920 336734
rect 385868 336670 385920 336676
rect 386144 335980 386196 335986
rect 386144 335922 386196 335928
rect 385788 325666 386092 325694
rect 386064 7614 386092 325666
rect 386052 7608 386104 7614
rect 386052 7550 386104 7556
rect 386156 4826 386184 335922
rect 386144 4820 386196 4826
rect 386144 4762 386196 4768
rect 385960 4208 386012 4214
rect 385960 4150 386012 4156
rect 384948 3800 385000 3806
rect 384948 3742 385000 3748
rect 385972 480 386000 4150
rect 386248 3534 386276 338014
rect 386800 336734 386828 338028
rect 387274 338014 387656 338042
rect 386328 336728 386380 336734
rect 386328 336670 386380 336676
rect 386788 336728 386840 336734
rect 386788 336670 386840 336676
rect 387524 336728 387576 336734
rect 387524 336670 387576 336676
rect 386340 3738 386368 336670
rect 386328 3732 386380 3738
rect 386328 3674 386380 3680
rect 387536 3602 387564 336670
rect 387628 3670 387656 338014
rect 387616 3664 387668 3670
rect 387616 3606 387668 3612
rect 387524 3596 387576 3602
rect 387524 3538 387576 3544
rect 386236 3528 386288 3534
rect 386236 3470 386288 3476
rect 387720 3466 387748 338028
rect 387800 329180 387852 329186
rect 387800 329122 387852 329128
rect 387812 16574 387840 329122
rect 389192 325650 389220 402455
rect 389270 399936 389326 399945
rect 389270 399871 389326 399880
rect 389180 325644 389232 325650
rect 389180 325586 389232 325592
rect 389284 313274 389312 399871
rect 389362 397352 389418 397361
rect 389362 397287 389418 397296
rect 389272 313268 389324 313274
rect 389272 313210 389324 313216
rect 389376 299470 389404 397287
rect 389454 386744 389510 386753
rect 389454 386679 389510 386688
rect 389364 299464 389416 299470
rect 389364 299406 389416 299412
rect 389468 245614 389496 386679
rect 389546 384160 389602 384169
rect 389546 384095 389602 384104
rect 389456 245608 389508 245614
rect 389456 245550 389508 245556
rect 389560 233238 389588 384095
rect 389638 381440 389694 381449
rect 389638 381375 389694 381384
rect 389548 233232 389600 233238
rect 389548 233174 389600 233180
rect 389652 219434 389680 381375
rect 389730 378856 389786 378865
rect 389730 378791 389786 378800
rect 389640 219428 389692 219434
rect 389640 219370 389692 219376
rect 389744 206990 389772 378791
rect 389836 353258 389864 407759
rect 389928 365702 389956 410479
rect 390020 379506 390048 413063
rect 390112 391950 390140 415783
rect 390204 405686 390232 418367
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 390192 405680 390244 405686
rect 390192 405622 390244 405628
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 391204 404524 391256 404530
rect 391204 404466 391256 404472
rect 390190 394632 390246 394641
rect 390190 394567 390246 394576
rect 390204 393378 390232 394567
rect 390192 393372 390244 393378
rect 390192 393314 390244 393320
rect 390190 392048 390246 392057
rect 390190 391983 390192 391992
rect 390244 391983 390246 391992
rect 390192 391954 390244 391960
rect 390100 391944 390152 391950
rect 390100 391886 390152 391892
rect 390190 389328 390246 389337
rect 390190 389263 390246 389272
rect 390204 389230 390232 389263
rect 390192 389224 390244 389230
rect 390192 389166 390244 389172
rect 390008 379500 390060 379506
rect 390008 379442 390060 379448
rect 390466 376136 390522 376145
rect 390466 376071 390522 376080
rect 390098 373552 390154 373561
rect 390098 373487 390154 373496
rect 390112 372638 390140 373487
rect 390100 372632 390152 372638
rect 390100 372574 390152 372580
rect 390374 370832 390430 370841
rect 390374 370767 390430 370776
rect 390282 368248 390338 368257
rect 390282 368183 390338 368192
rect 389916 365696 389968 365702
rect 389916 365638 389968 365644
rect 390190 365664 390246 365673
rect 390190 365599 390246 365608
rect 389914 362944 389970 362953
rect 389914 362879 389970 362888
rect 389928 357338 389956 362879
rect 390006 360360 390062 360369
rect 390006 360295 390062 360304
rect 389916 357332 389968 357338
rect 389916 357274 389968 357280
rect 389914 355056 389970 355065
rect 389914 354991 389970 355000
rect 389928 354754 389956 354991
rect 389916 354748 389968 354754
rect 389916 354690 389968 354696
rect 389824 353252 389876 353258
rect 389824 353194 389876 353200
rect 389914 352472 389970 352481
rect 389914 352407 389970 352416
rect 389822 349752 389878 349761
rect 389822 349687 389878 349696
rect 389732 206984 389784 206990
rect 389732 206926 389784 206932
rect 389836 60722 389864 349687
rect 389928 347274 389956 352407
rect 389916 347268 389968 347274
rect 389916 347210 389968 347216
rect 389914 347168 389970 347177
rect 389914 347103 389970 347112
rect 389928 346458 389956 347103
rect 389916 346452 389968 346458
rect 389916 346394 389968 346400
rect 389916 346316 389968 346322
rect 389916 346258 389968 346264
rect 389928 73166 389956 346258
rect 390020 113150 390048 360295
rect 390098 357640 390154 357649
rect 390098 357575 390154 357584
rect 390112 357474 390140 357575
rect 390100 357468 390152 357474
rect 390100 357410 390152 357416
rect 390100 357332 390152 357338
rect 390100 357274 390152 357280
rect 390112 126954 390140 357274
rect 390204 139398 390232 365599
rect 390296 153202 390324 368183
rect 390388 167006 390416 370767
rect 390480 193186 390508 376071
rect 391216 340202 391244 404466
rect 396816 393372 396868 393378
rect 396816 393314 396868 393320
rect 393964 392012 394016 392018
rect 393964 391954 394016 391960
rect 391204 340196 391256 340202
rect 391204 340138 391256 340144
rect 393976 273222 394004 391954
rect 396828 341562 396856 393314
rect 580172 391944 580224 391950
rect 580172 391886 580224 391892
rect 580184 391785 580212 391886
rect 580170 391776 580226 391785
rect 580170 391711 580226 391720
rect 406384 389224 406436 389230
rect 406384 389166 406436 389172
rect 403624 372632 403676 372638
rect 403624 372574 403676 372580
rect 400864 357468 400916 357474
rect 400864 357410 400916 357416
rect 396816 341556 396868 341562
rect 396816 341498 396868 341504
rect 396724 340944 396776 340950
rect 396724 340886 396776 340892
rect 394700 327820 394752 327826
rect 394700 327762 394752 327768
rect 393964 273216 394016 273222
rect 393964 273158 394016 273164
rect 390468 193180 390520 193186
rect 390468 193122 390520 193128
rect 390376 167000 390428 167006
rect 390376 166942 390428 166948
rect 390284 153196 390336 153202
rect 390284 153138 390336 153144
rect 390192 139392 390244 139398
rect 390192 139334 390244 139340
rect 390100 126948 390152 126954
rect 390100 126890 390152 126896
rect 390008 113144 390060 113150
rect 390008 113086 390060 113092
rect 389916 73160 389968 73166
rect 389916 73102 389968 73108
rect 389824 60716 389876 60722
rect 389824 60658 389876 60664
rect 394712 16574 394740 327762
rect 396080 324964 396132 324970
rect 396080 324906 396132 324912
rect 396092 16574 396120 324906
rect 396736 20670 396764 340886
rect 398840 334688 398892 334694
rect 398840 334630 398892 334636
rect 396724 20664 396776 20670
rect 396724 20606 396776 20612
rect 387812 16546 388300 16574
rect 394712 16546 395384 16574
rect 396092 16546 396580 16574
rect 387156 3460 387208 3466
rect 387156 3402 387208 3408
rect 387708 3460 387760 3466
rect 387708 3402 387760 3408
rect 387168 480 387196 3402
rect 388272 480 388300 16546
rect 390652 13184 390704 13190
rect 390652 13126 390704 13132
rect 389456 7064 389508 7070
rect 389456 7006 389508 7012
rect 389468 480 389496 7006
rect 390664 3534 390692 13126
rect 393044 7132 393096 7138
rect 393044 7074 393096 7080
rect 390652 3528 390704 3534
rect 390652 3470 390704 3476
rect 391848 3528 391900 3534
rect 391848 3470 391900 3476
rect 390652 2848 390704 2854
rect 390652 2790 390704 2796
rect 390664 480 390692 2790
rect 391860 480 391888 3470
rect 393056 480 393084 7074
rect 394240 2916 394292 2922
rect 394240 2858 394292 2864
rect 394252 480 394280 2858
rect 395356 480 395384 16546
rect 396552 480 396580 16546
rect 398852 3058 398880 334630
rect 398932 326460 398984 326466
rect 398932 326402 398984 326408
rect 398840 3052 398892 3058
rect 398840 2994 398892 3000
rect 397736 2984 397788 2990
rect 397736 2926 397788 2932
rect 397748 480 397776 2926
rect 398944 480 398972 326402
rect 400876 100706 400904 357410
rect 401600 322312 401652 322318
rect 401600 322254 401652 322260
rect 400864 100700 400916 100706
rect 400864 100642 400916 100648
rect 401612 16574 401640 322254
rect 402980 222896 403032 222902
rect 402980 222838 403032 222844
rect 402992 16574 403020 222838
rect 403636 179382 403664 372574
rect 405740 320952 405792 320958
rect 405740 320894 405792 320900
rect 403624 179376 403676 179382
rect 403624 179318 403676 179324
rect 405752 16574 405780 320894
rect 406396 259418 406424 389166
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 547144 354748 547196 354754
rect 547144 354690 547196 354696
rect 543004 346452 543056 346458
rect 543004 346394 543056 346400
rect 519544 338156 519596 338162
rect 519544 338098 519596 338104
rect 411260 336660 411312 336666
rect 411260 336602 411312 336608
rect 406384 259412 406436 259418
rect 406384 259354 406436 259360
rect 411272 16574 411300 336602
rect 418160 336592 418212 336598
rect 418160 336534 418212 336540
rect 412640 323672 412692 323678
rect 412640 323614 412692 323620
rect 412652 16574 412680 323614
rect 415492 17264 415544 17270
rect 415492 17206 415544 17212
rect 401612 16546 402560 16574
rect 402992 16546 403664 16574
rect 405752 16546 406056 16574
rect 411272 16546 411944 16574
rect 412652 16546 413140 16574
rect 400128 3052 400180 3058
rect 400128 2994 400180 3000
rect 400140 480 400168 2994
rect 401324 2984 401376 2990
rect 401324 2926 401376 2932
rect 401336 480 401364 2926
rect 402532 480 402560 16546
rect 403636 480 403664 16546
rect 404820 3120 404872 3126
rect 404820 3062 404872 3068
rect 404832 480 404860 3062
rect 406028 480 406056 16546
rect 409604 15904 409656 15910
rect 409604 15846 409656 15852
rect 407212 8424 407264 8430
rect 407212 8366 407264 8372
rect 407224 480 407252 8366
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 408420 480 408448 3130
rect 409616 480 409644 15846
rect 410800 8492 410852 8498
rect 410800 8434 410852 8440
rect 410812 480 410840 8434
rect 411916 480 411944 16546
rect 413112 480 413140 16546
rect 414296 8560 414348 8566
rect 414296 8502 414348 8508
rect 414308 480 414336 8502
rect 415504 3262 415532 17206
rect 418172 16574 418200 336534
rect 425060 336524 425112 336530
rect 425060 336466 425112 336472
rect 419540 319524 419592 319530
rect 419540 319466 419592 319472
rect 419552 16574 419580 319466
rect 425072 16574 425100 336466
rect 431960 336456 432012 336462
rect 431960 336398 432012 336404
rect 418172 16546 419028 16574
rect 419552 16546 420224 16574
rect 425072 16546 426204 16574
rect 417884 8628 417936 8634
rect 417884 8570 417936 8576
rect 415400 3256 415452 3262
rect 415400 3198 415452 3204
rect 415492 3256 415544 3262
rect 415492 3198 415544 3204
rect 416688 3256 416740 3262
rect 416688 3198 416740 3204
rect 415412 1714 415440 3198
rect 415412 1686 415532 1714
rect 415504 480 415532 1686
rect 416700 480 416728 3198
rect 417896 480 417924 8570
rect 419000 480 419028 16546
rect 420196 480 420224 16546
rect 424968 8764 425020 8770
rect 424968 8706 425020 8712
rect 421380 8696 421432 8702
rect 421380 8638 421432 8644
rect 421392 480 421420 8638
rect 423772 5704 423824 5710
rect 423772 5646 423824 5652
rect 422576 3324 422628 3330
rect 422576 3266 422628 3272
rect 422588 480 422616 3266
rect 423784 480 423812 5646
rect 424980 480 425008 8706
rect 426176 480 426204 16546
rect 428464 8832 428516 8838
rect 428464 8774 428516 8780
rect 427268 5772 427320 5778
rect 427268 5714 427320 5720
rect 427280 480 427308 5714
rect 428476 480 428504 8774
rect 430856 5840 430908 5846
rect 430856 5782 430908 5788
rect 429660 3392 429712 3398
rect 429660 3334 429712 3340
rect 429672 480 429700 3334
rect 430868 480 430896 5782
rect 431972 3398 432000 336398
rect 440240 336388 440292 336394
rect 440240 336330 440292 336336
rect 440252 16574 440280 336330
rect 447140 336320 447192 336326
rect 447140 336262 447192 336268
rect 447152 16574 447180 336262
rect 454040 336252 454092 336258
rect 454040 336194 454092 336200
rect 454052 16574 454080 336194
rect 460940 336184 460992 336190
rect 460940 336126 460992 336132
rect 460952 16574 460980 336126
rect 467840 336116 467892 336122
rect 467840 336058 467892 336064
rect 467852 16574 467880 336058
rect 474740 336048 474792 336054
rect 474740 335990 474792 335996
rect 473360 21412 473412 21418
rect 473360 21354 473412 21360
rect 440252 16546 440372 16574
rect 447152 16546 447456 16574
rect 454052 16546 454540 16574
rect 460952 16546 461624 16574
rect 467852 16546 468708 16574
rect 435548 9648 435600 9654
rect 435548 9590 435600 9596
rect 432052 8900 432104 8906
rect 432052 8842 432104 8848
rect 431960 3392 432012 3398
rect 431960 3334 432012 3340
rect 432064 480 432092 8842
rect 434444 5908 434496 5914
rect 434444 5850 434496 5856
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 434456 480 434484 5850
rect 435560 480 435588 9590
rect 439136 9580 439188 9586
rect 439136 9522 439188 9528
rect 437940 5976 437992 5982
rect 437940 5918 437992 5924
rect 436744 4140 436796 4146
rect 436744 4082 436796 4088
rect 436756 480 436784 4082
rect 437952 480 437980 5918
rect 439148 480 439176 9522
rect 440344 480 440372 16546
rect 442632 9512 442684 9518
rect 442632 9454 442684 9460
rect 441528 6044 441580 6050
rect 441528 5986 441580 5992
rect 441540 480 441568 5986
rect 442644 480 442672 9454
rect 446220 9444 446272 9450
rect 446220 9386 446272 9392
rect 445024 6112 445076 6118
rect 445024 6054 445076 6060
rect 443828 4072 443880 4078
rect 443828 4014 443880 4020
rect 443840 480 443868 4014
rect 445036 480 445064 6054
rect 446232 480 446260 9386
rect 447428 480 447456 16546
rect 449808 9376 449860 9382
rect 449808 9318 449860 9324
rect 448612 6860 448664 6866
rect 448612 6802 448664 6808
rect 448624 480 448652 6802
rect 449820 480 449848 9318
rect 453304 9308 453356 9314
rect 453304 9250 453356 9256
rect 452108 6792 452160 6798
rect 452108 6734 452160 6740
rect 450912 4004 450964 4010
rect 450912 3946 450964 3952
rect 450924 480 450952 3946
rect 452120 480 452148 6734
rect 453316 480 453344 9250
rect 454512 480 454540 16546
rect 456892 9240 456944 9246
rect 456892 9182 456944 9188
rect 455696 6724 455748 6730
rect 455696 6666 455748 6672
rect 455708 480 455736 6666
rect 456904 480 456932 9182
rect 460388 9172 460440 9178
rect 460388 9114 460440 9120
rect 459192 6656 459244 6662
rect 459192 6598 459244 6604
rect 458086 3768 458142 3777
rect 458086 3703 458142 3712
rect 458100 480 458128 3703
rect 459204 480 459232 6598
rect 460400 480 460428 9114
rect 461596 480 461624 16546
rect 463976 9104 464028 9110
rect 463976 9046 464028 9052
rect 462780 6588 462832 6594
rect 462780 6530 462832 6536
rect 462792 480 462820 6530
rect 463988 480 464016 9046
rect 467472 9036 467524 9042
rect 467472 8978 467524 8984
rect 466276 6520 466328 6526
rect 466276 6462 466328 6468
rect 465170 3632 465226 3641
rect 465170 3567 465226 3576
rect 465184 480 465212 3567
rect 466288 480 466316 6462
rect 467484 480 467512 8978
rect 468680 480 468708 16546
rect 471060 8968 471112 8974
rect 471060 8910 471112 8916
rect 469864 6452 469916 6458
rect 469864 6394 469916 6400
rect 469876 480 469904 6394
rect 471072 480 471100 8910
rect 472254 3496 472310 3505
rect 472254 3431 472310 3440
rect 472268 480 472296 3431
rect 473372 3398 473400 21354
rect 474752 16574 474780 335990
rect 483020 334620 483072 334626
rect 483020 334562 483072 334568
rect 477500 311160 477552 311166
rect 477500 311102 477552 311108
rect 477512 16574 477540 311102
rect 481640 308440 481692 308446
rect 481640 308382 481692 308388
rect 474752 16546 475792 16574
rect 477512 16546 478184 16574
rect 473452 6384 473504 6390
rect 473452 6326 473504 6332
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 6326
rect 474556 3392 474608 3398
rect 474556 3334 474608 3340
rect 474568 480 474596 3334
rect 475764 480 475792 16546
rect 476948 6316 477000 6322
rect 476948 6258 477000 6264
rect 476960 480 476988 6258
rect 478156 480 478184 16546
rect 480536 11756 480588 11762
rect 480536 11698 480588 11704
rect 479338 3360 479394 3369
rect 479338 3295 479394 3304
rect 479352 480 479380 3295
rect 480548 480 480576 11698
rect 481652 3398 481680 308382
rect 483032 16574 483060 334562
rect 489920 333328 489972 333334
rect 489920 333270 489972 333276
rect 485780 327752 485832 327758
rect 485780 327694 485832 327700
rect 485792 16574 485820 327694
rect 488540 318096 488592 318102
rect 488540 318038 488592 318044
rect 487160 217320 487212 217326
rect 487160 217262 487212 217268
rect 487172 16574 487200 217262
rect 488552 16574 488580 318038
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 487172 16546 487660 16574
rect 488552 16546 488856 16574
rect 481732 6248 481784 6254
rect 481732 6190 481784 6196
rect 481640 3392 481692 3398
rect 481640 3334 481692 3340
rect 481744 480 481772 6190
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482848 480 482876 3334
rect 484044 480 484072 16546
rect 485228 6180 485280 6186
rect 485228 6122 485280 6128
rect 485240 480 485268 6122
rect 486436 480 486464 16546
rect 487632 480 487660 16546
rect 488828 480 488856 16546
rect 489932 3398 489960 333270
rect 500960 331968 501012 331974
rect 500960 331910 501012 331916
rect 492680 326392 492732 326398
rect 492680 326334 492732 326340
rect 490012 22772 490064 22778
rect 490012 22714 490064 22720
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 490024 1442 490052 22714
rect 492692 16574 492720 326334
rect 495440 316736 495492 316742
rect 495440 316678 495492 316684
rect 495452 16574 495480 316678
rect 496820 309800 496872 309806
rect 496820 309742 496872 309748
rect 496832 16574 496860 309742
rect 499580 307080 499632 307086
rect 499580 307022 499632 307028
rect 498200 215960 498252 215966
rect 498200 215902 498252 215908
rect 492692 16546 493548 16574
rect 495452 16546 495940 16574
rect 496832 16546 497136 16574
rect 492312 14476 492364 14482
rect 492312 14418 492364 14424
rect 491116 3392 491168 3398
rect 491116 3334 491168 3340
rect 489932 1414 490052 1442
rect 489932 480 489960 1414
rect 491128 480 491156 3334
rect 492324 480 492352 14418
rect 493520 480 493548 16546
rect 494704 10328 494756 10334
rect 494704 10270 494756 10276
rect 494716 480 494744 10270
rect 495912 480 495940 16546
rect 497108 480 497136 16546
rect 498212 480 498240 215902
rect 499592 16574 499620 307022
rect 500972 16574 501000 331910
rect 507860 330540 507912 330546
rect 507860 330482 507912 330488
rect 502340 329112 502392 329118
rect 502340 329054 502392 329060
rect 502352 16574 502380 329054
rect 506480 315308 506532 315314
rect 506480 315250 506532 315256
rect 503720 305652 503772 305658
rect 503720 305594 503772 305600
rect 503732 16574 503760 305594
rect 505100 42084 505152 42090
rect 505100 42026 505152 42032
rect 505112 16574 505140 42026
rect 499592 16546 500632 16574
rect 500972 16546 501828 16574
rect 502352 16546 503024 16574
rect 503732 16546 504220 16574
rect 505112 16546 505416 16574
rect 499396 13116 499448 13122
rect 499396 13058 499448 13064
rect 499408 480 499436 13058
rect 500604 480 500632 16546
rect 501800 480 501828 16546
rect 502996 480 503024 16546
rect 504192 480 504220 16546
rect 505388 480 505416 16546
rect 506492 480 506520 315250
rect 506572 24132 506624 24138
rect 506572 24074 506624 24080
rect 506584 16574 506612 24074
rect 507872 16574 507900 330482
rect 514760 322244 514812 322250
rect 514760 322186 514812 322192
rect 513380 313948 513432 313954
rect 513380 313890 513432 313896
rect 510620 302932 510672 302938
rect 510620 302874 510672 302880
rect 509240 18624 509292 18630
rect 509240 18566 509292 18572
rect 509252 16574 509280 18566
rect 510632 16574 510660 302874
rect 513392 16574 513420 313890
rect 506584 16546 507716 16574
rect 507872 16546 508912 16574
rect 509252 16546 510108 16574
rect 510632 16546 511304 16574
rect 513392 16546 513604 16574
rect 507688 480 507716 16546
rect 508884 480 508912 16546
rect 510080 480 510108 16546
rect 511276 480 511304 16546
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 513576 480 513604 16546
rect 514772 480 514800 322186
rect 517520 320884 517572 320890
rect 517520 320826 517572 320832
rect 516140 220108 516192 220114
rect 516140 220050 516192 220056
rect 516152 16574 516180 220050
rect 517532 16574 517560 320826
rect 516152 16546 517192 16574
rect 517532 16546 518388 16574
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517164 480 517192 16546
rect 518360 480 518388 16546
rect 519556 6866 519584 338098
rect 539600 333260 539652 333266
rect 539600 333202 539652 333208
rect 521660 323604 521712 323610
rect 521660 323546 521712 323552
rect 521672 16574 521700 323546
rect 535460 319456 535512 319462
rect 535460 319398 535512 319404
rect 524420 304292 524472 304298
rect 524420 304234 524472 304240
rect 524432 16574 524460 304234
rect 528560 301504 528612 301510
rect 528560 301446 528612 301452
rect 528572 16574 528600 301446
rect 531320 297424 531372 297430
rect 531320 297366 531372 297372
rect 521672 16546 521884 16574
rect 524432 16546 525472 16574
rect 528572 16546 529060 16574
rect 520740 7200 520792 7206
rect 520740 7142 520792 7148
rect 519544 6860 519596 6866
rect 519544 6802 519596 6808
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 519556 480 519584 4354
rect 520752 480 520780 7142
rect 521856 480 521884 16546
rect 524236 7268 524288 7274
rect 524236 7210 524288 7216
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 523052 480 523080 4422
rect 524248 480 524276 7210
rect 525444 480 525472 16546
rect 527824 7336 527876 7342
rect 527824 7278 527876 7284
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526640 480 526668 4490
rect 527836 480 527864 7278
rect 529032 480 529060 16546
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 530136 480 530164 4558
rect 531332 3398 531360 297366
rect 535472 16574 535500 319398
rect 535472 16546 536144 16574
rect 534908 7472 534960 7478
rect 534908 7414 534960 7420
rect 531412 7404 531464 7410
rect 531412 7346 531464 7352
rect 531320 3392 531372 3398
rect 531320 3334 531372 3340
rect 531424 1442 531452 7346
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 532516 3392 532568 3398
rect 532516 3334 532568 3340
rect 531332 1414 531452 1442
rect 531332 480 531360 1414
rect 532528 480 532556 3334
rect 533724 480 533752 4626
rect 534920 480 534948 7414
rect 536116 480 536144 16546
rect 538404 7540 538456 7546
rect 538404 7482 538456 7488
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 538416 480 538444 7482
rect 539612 480 539640 333202
rect 542360 300144 542412 300150
rect 542360 300086 542412 300092
rect 542372 16574 542400 300086
rect 543016 46918 543044 346394
rect 546500 295996 546552 296002
rect 546500 295938 546552 295944
rect 543004 46912 543056 46918
rect 543004 46854 543056 46860
rect 546512 16574 546540 295938
rect 547156 86970 547184 354690
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580264 341556 580316 341562
rect 580264 341498 580316 341504
rect 580172 340196 580224 340202
rect 580172 340138 580224 340144
rect 580184 338609 580212 340138
rect 580170 338600 580226 338609
rect 580170 338535 580226 338544
rect 556160 331900 556212 331906
rect 556160 331842 556212 331848
rect 553400 294636 553452 294642
rect 553400 294578 553452 294584
rect 549260 293276 549312 293282
rect 549260 293218 549312 293224
rect 547144 86964 547196 86970
rect 547144 86906 547196 86912
rect 549272 16574 549300 293218
rect 553412 16574 553440 294578
rect 542372 16546 543228 16574
rect 546512 16546 546724 16574
rect 549272 16546 550312 16574
rect 553412 16546 553808 16574
rect 541992 8288 542044 8294
rect 541992 8230 542044 8236
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 540808 480 540836 5442
rect 542004 480 542032 8230
rect 543200 480 543228 16546
rect 545488 8220 545540 8226
rect 545488 8162 545540 8168
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 544396 480 544424 5374
rect 545500 480 545528 8162
rect 546696 480 546724 16546
rect 549076 8152 549128 8158
rect 549076 8094 549128 8100
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 547892 480 547920 5306
rect 549088 480 549116 8094
rect 550284 480 550312 16546
rect 552664 8084 552716 8090
rect 552664 8026 552716 8032
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 551480 480 551508 5238
rect 552676 480 552704 8026
rect 553780 480 553808 16546
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 554976 480 555004 5170
rect 556172 3398 556200 331842
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 560300 291848 560352 291854
rect 560300 291790 560352 291796
rect 560312 16574 560340 291790
rect 564440 290488 564492 290494
rect 564440 290430 564492 290436
rect 560312 16546 560892 16574
rect 556252 8016 556304 8022
rect 556252 7958 556304 7964
rect 556160 3392 556212 3398
rect 556160 3334 556212 3340
rect 556264 1442 556292 7958
rect 559748 7948 559800 7954
rect 559748 7890 559800 7896
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3392 557408 3398
rect 557356 3334 557408 3340
rect 556172 1414 556292 1442
rect 556172 480 556200 1414
rect 557368 480 557396 3334
rect 558564 480 558592 5102
rect 559760 480 559788 7890
rect 560864 480 560892 16546
rect 563244 7880 563296 7886
rect 563244 7822 563296 7828
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 562060 480 562088 5034
rect 563256 480 563284 7822
rect 564452 480 564480 290430
rect 580276 285433 580304 341498
rect 580262 285424 580318 285433
rect 580262 285359 580318 285368
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 566832 7812 566884 7818
rect 566832 7754 566884 7760
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 565648 480 565676 4966
rect 566844 480 566872 7754
rect 570328 7744 570380 7750
rect 570328 7686 570380 7692
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3936 568080 3942
rect 568028 3878 568080 3884
rect 568040 480 568068 3878
rect 569144 480 569172 4898
rect 570340 480 570368 7686
rect 573916 7676 573968 7682
rect 573916 7618 573968 7624
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 571524 3868 571576 3874
rect 571524 3810 571576 3816
rect 571536 480 571564 3810
rect 572732 480 572760 4830
rect 573928 480 573956 7618
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 575112 3800 575164 3806
rect 575112 3742 575164 3748
rect 575124 480 575152 3742
rect 576320 480 576348 4762
rect 577424 480 577452 7550
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 578608 3732 578660 3738
rect 578608 3674 578660 3680
rect 578620 480 578648 3674
rect 582196 3664 582248 3670
rect 582196 3606 582248 3612
rect 579804 3596 579856 3602
rect 579804 3538 579856 3544
rect 579816 480 579844 3538
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 582208 480 582236 3606
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3422 671200 3478 671256
rect 2778 645108 2834 645144
rect 2778 645088 2780 645108
rect 2780 645088 2832 645108
rect 2832 645088 2834 645108
rect 3330 553832 3386 553888
rect 3238 540776 3294 540832
rect 3146 527856 3202 527912
rect 3054 514800 3110 514856
rect 2962 501744 3018 501800
rect 2870 488688 2926 488744
rect 2778 475632 2834 475688
rect 3514 658144 3570 658200
rect 3606 632032 3662 632088
rect 3698 619112 3754 619168
rect 3422 462576 3478 462632
rect 3790 606056 3846 606112
rect 3882 593000 3938 593056
rect 3974 579944 4030 580000
rect 4066 566888 4122 566944
rect 580170 697176 580226 697232
rect 165618 476448 165674 476504
rect 165618 471280 165674 471336
rect 165618 468696 165674 468752
rect 165618 466112 165674 466168
rect 165618 463528 165674 463584
rect 165618 460944 165674 461000
rect 165618 458360 165674 458416
rect 165618 455776 165674 455832
rect 165618 453192 165674 453248
rect 165618 450608 165674 450664
rect 3514 449520 3570 449576
rect 165618 448024 165674 448080
rect 165618 445440 165674 445496
rect 165618 442892 165620 442912
rect 165620 442892 165672 442912
rect 165672 442892 165674 442912
rect 165618 442856 165674 442892
rect 165618 440272 165674 440328
rect 165618 437688 165674 437744
rect 3606 436600 3662 436656
rect 165618 435104 165674 435160
rect 580170 683848 580226 683904
rect 389822 476448 389878 476504
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 389914 473864 389970 473920
rect 580170 670656 580226 670692
rect 580262 657328 580318 657384
rect 580170 644000 580226 644056
rect 390006 471144 390062 471200
rect 579986 630808 580042 630864
rect 389730 444760 389786 444816
rect 389638 442176 389694 442232
rect 389546 434152 389602 434208
rect 165618 432520 165674 432576
rect 390098 468560 390154 468616
rect 390006 465840 390062 465896
rect 580170 617480 580226 617536
rect 390190 463256 390246 463312
rect 579618 590960 579674 591016
rect 390282 460672 390338 460728
rect 390190 457952 390246 458008
rect 389822 431568 389878 431624
rect 165618 429800 165674 429856
rect 165618 427216 165674 427272
rect 165618 424632 165674 424688
rect 579618 577632 579674 577688
rect 390374 455368 390430 455424
rect 579618 537784 579674 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580354 604152 580410 604208
rect 580446 564304 580502 564360
rect 579802 458088 579858 458144
rect 390466 452648 390522 452704
rect 580538 551112 580594 551168
rect 390190 450064 390246 450120
rect 580630 511264 580686 511320
rect 390190 447480 390246 447536
rect 580170 444760 580226 444816
rect 389914 428984 389970 429040
rect 580722 497936 580778 497992
rect 390190 439456 390246 439512
rect 390282 436872 390338 436928
rect 580170 431568 580226 431624
rect 390006 426264 390062 426320
rect 389822 423680 389878 423736
rect 3790 423544 3846 423600
rect 165618 422048 165674 422104
rect 390098 420960 390154 421016
rect 165618 419464 165674 419520
rect 390190 418376 390246 418432
rect 165618 416880 165674 416936
rect 3422 410488 3478 410544
rect 3054 332288 3110 332344
rect 3054 319232 3110 319288
rect 3146 306176 3202 306232
rect 2778 293120 2834 293176
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3238 227976 3294 228032
rect 3238 214920 3294 214976
rect 390098 415792 390154 415848
rect 165618 414296 165674 414352
rect 390006 413072 390062 413128
rect 165618 411712 165674 411768
rect 389914 410488 389970 410544
rect 165618 409128 165674 409184
rect 389822 407768 389878 407824
rect 165618 406544 165674 406600
rect 389178 405184 389234 405240
rect 166906 403960 166962 404016
rect 166814 401376 166870 401432
rect 165618 398828 165620 398848
rect 165620 398828 165672 398848
rect 165672 398828 165674 398848
rect 165618 398792 165674 398828
rect 3790 397432 3846 397488
rect 165618 396208 165674 396264
rect 3698 384376 3754 384432
rect 3606 371320 3662 371376
rect 3514 358400 3570 358456
rect 3422 345344 3478 345400
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3330 175888 3386 175944
rect 3330 149776 3386 149832
rect 3146 123664 3202 123720
rect 3146 84632 3202 84688
rect 2870 58520 2926 58576
rect 166722 393624 166778 393680
rect 166630 391040 166686 391096
rect 165618 388456 165674 388512
rect 4066 162832 4122 162888
rect 3974 136720 4030 136776
rect 3882 110608 3938 110664
rect 3790 97552 3846 97608
rect 3698 71576 3754 71632
rect 3606 45464 3662 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 11150 3440 11206 3496
rect 165618 385872 165674 385928
rect 166538 383152 166594 383208
rect 166446 380568 166502 380624
rect 165618 377984 165674 378040
rect 165618 375420 165674 375456
rect 165618 375400 165620 375420
rect 165620 375400 165672 375420
rect 165672 375400 165674 375420
rect 166354 372816 166410 372872
rect 165618 370232 165674 370288
rect 165618 367648 165674 367704
rect 20626 3712 20682 3768
rect 19430 3576 19486 3632
rect 165618 365064 165674 365120
rect 166262 362480 166318 362536
rect 165618 359896 165674 359952
rect 165618 357312 165674 357368
rect 165618 354748 165674 354784
rect 165618 354728 165620 354748
rect 165620 354728 165672 354748
rect 165672 354728 165674 354748
rect 165618 352144 165674 352200
rect 165618 349560 165674 349616
rect 165618 346976 165674 347032
rect 165618 344392 165674 344448
rect 165618 341808 165674 341864
rect 165618 339224 165674 339280
rect 389178 402464 389234 402520
rect 389086 341264 389142 341320
rect 389086 338680 389142 338736
rect 169942 3304 169998 3360
rect 171322 3440 171378 3496
rect 175554 3712 175610 3768
rect 175370 3576 175426 3632
rect 340786 3712 340842 3768
rect 343546 3576 343602 3632
rect 346306 3440 346362 3496
rect 349066 3304 349122 3360
rect 389270 399880 389326 399936
rect 389362 397296 389418 397352
rect 389454 386688 389510 386744
rect 389546 384104 389602 384160
rect 389638 381384 389694 381440
rect 389730 378800 389786 378856
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 390190 394576 390246 394632
rect 390190 392012 390246 392048
rect 390190 391992 390192 392012
rect 390192 391992 390244 392012
rect 390244 391992 390246 392012
rect 390190 389272 390246 389328
rect 390466 376080 390522 376136
rect 390098 373496 390154 373552
rect 390374 370776 390430 370832
rect 390282 368192 390338 368248
rect 390190 365608 390246 365664
rect 389914 362888 389970 362944
rect 390006 360304 390062 360360
rect 389914 355000 389970 355056
rect 389914 352416 389970 352472
rect 389822 349696 389878 349752
rect 389914 347112 389970 347168
rect 390098 357584 390154 357640
rect 580170 391720 580226 391776
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 458086 3712 458142 3768
rect 465170 3576 465226 3632
rect 472254 3440 472310 3496
rect 479338 3304 479394 3360
rect 580170 351872 580226 351928
rect 580170 338544 580226 338600
rect 579894 325216 579950 325272
rect 580170 312024 580226 312080
rect 579618 298696 579674 298752
rect 580262 285368 580318 285424
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3366 684314 3372 684316
rect -960 684254 3372 684314
rect -960 684164 480 684254
rect 3366 684252 3372 684254
rect 3436 684252 3442 684316
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 580257 657386 580323 657389
rect 583520 657386 584960 657476
rect 580257 657384 584960 657386
rect 580257 657328 580262 657384
rect 580318 657328 584960 657384
rect 580257 657326 584960 657328
rect 580257 657323 580323 657326
rect 583520 657236 584960 657326
rect -960 645146 480 645236
rect 2773 645146 2839 645149
rect -960 645144 2839 645146
rect -960 645088 2778 645144
rect 2834 645088 2839 645144
rect -960 645086 2839 645088
rect -960 644996 480 645086
rect 2773 645083 2839 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3693 619170 3759 619173
rect -960 619168 3759 619170
rect -960 619112 3698 619168
rect 3754 619112 3759 619168
rect -960 619110 3759 619112
rect -960 619020 480 619110
rect 3693 619107 3759 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3785 606114 3851 606117
rect -960 606112 3851 606114
rect -960 606056 3790 606112
rect 3846 606056 3851 606112
rect -960 606054 3851 606056
rect -960 605964 480 606054
rect 3785 606051 3851 606054
rect 580349 604210 580415 604213
rect 583520 604210 584960 604300
rect 580349 604208 584960 604210
rect 580349 604152 580354 604208
rect 580410 604152 584960 604208
rect 580349 604150 584960 604152
rect 580349 604147 580415 604150
rect 583520 604060 584960 604150
rect -960 593058 480 593148
rect 3877 593058 3943 593061
rect -960 593056 3943 593058
rect -960 593000 3882 593056
rect 3938 593000 3943 593056
rect -960 592998 3943 593000
rect -960 592908 480 592998
rect 3877 592995 3943 592998
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3969 580002 4035 580005
rect -960 580000 4035 580002
rect -960 579944 3974 580000
rect 4030 579944 4035 580000
rect -960 579942 4035 579944
rect -960 579852 480 579942
rect 3969 579939 4035 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 4061 566946 4127 566949
rect -960 566944 4127 566946
rect -960 566888 4066 566944
rect 4122 566888 4127 566944
rect -960 566886 4127 566888
rect -960 566796 480 566886
rect 4061 566883 4127 566886
rect 580441 564362 580507 564365
rect 583520 564362 584960 564452
rect 580441 564360 584960 564362
rect 580441 564304 580446 564360
rect 580502 564304 584960 564360
rect 580441 564302 584960 564304
rect 580441 564299 580507 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 580533 551170 580599 551173
rect 583520 551170 584960 551260
rect 580533 551168 584960 551170
rect 580533 551112 580538 551168
rect 580594 551112 584960 551168
rect 580533 551110 584960 551112
rect 580533 551107 580599 551110
rect 583520 551020 584960 551110
rect -960 540834 480 540924
rect 3233 540834 3299 540837
rect -960 540832 3299 540834
rect -960 540776 3238 540832
rect 3294 540776 3299 540832
rect -960 540774 3299 540776
rect -960 540684 480 540774
rect 3233 540771 3299 540774
rect 579613 537842 579679 537845
rect 583520 537842 584960 537932
rect 579613 537840 584960 537842
rect 579613 537784 579618 537840
rect 579674 537784 584960 537840
rect 579613 537782 584960 537784
rect 579613 537779 579679 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3049 514858 3115 514861
rect -960 514856 3115 514858
rect -960 514800 3054 514856
rect 3110 514800 3115 514856
rect -960 514798 3115 514800
rect -960 514708 480 514798
rect 3049 514795 3115 514798
rect 580625 511322 580691 511325
rect 583520 511322 584960 511412
rect 580625 511320 584960 511322
rect 580625 511264 580630 511320
rect 580686 511264 584960 511320
rect 580625 511262 584960 511264
rect 580625 511259 580691 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 2957 501802 3023 501805
rect -960 501800 3023 501802
rect -960 501744 2962 501800
rect 3018 501744 3023 501800
rect -960 501742 3023 501744
rect -960 501652 480 501742
rect 2957 501739 3023 501742
rect 580717 497994 580783 497997
rect 583520 497994 584960 498084
rect 580717 497992 584960 497994
rect 580717 497936 580722 497992
rect 580778 497936 584960 497992
rect 580717 497934 584960 497936
rect 580717 497931 580783 497934
rect 583520 497844 584960 497934
rect -960 488746 480 488836
rect 2865 488746 2931 488749
rect -960 488744 2931 488746
rect -960 488688 2870 488744
rect 2926 488688 2931 488744
rect -960 488686 2931 488688
rect -960 488596 480 488686
rect 2865 488683 2931 488686
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 165613 476506 165679 476509
rect 389817 476506 389883 476509
rect 165613 476504 168084 476506
rect 165613 476448 165618 476504
rect 165674 476448 168084 476504
rect 165613 476446 168084 476448
rect 387964 476504 389883 476506
rect 387964 476448 389822 476504
rect 389878 476448 389883 476504
rect 387964 476446 389883 476448
rect 165613 476443 165679 476446
rect 389817 476443 389883 476446
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 389909 473922 389975 473925
rect 387964 473920 389975 473922
rect 3366 473316 3372 473380
rect 3436 473378 3442 473380
rect 168054 473378 168114 473892
rect 387964 473864 389914 473920
rect 389970 473864 389975 473920
rect 387964 473862 389975 473864
rect 389909 473859 389975 473862
rect 3436 473318 168114 473378
rect 3436 473316 3442 473318
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 165613 471338 165679 471341
rect 165613 471336 168084 471338
rect 165613 471280 165618 471336
rect 165674 471280 168084 471336
rect 583520 471324 584960 471414
rect 165613 471278 168084 471280
rect 165613 471275 165679 471278
rect 390001 471202 390067 471205
rect 387964 471200 390067 471202
rect 387964 471144 390006 471200
rect 390062 471144 390067 471200
rect 387964 471142 390067 471144
rect 390001 471139 390067 471142
rect 165613 468754 165679 468757
rect 165613 468752 168084 468754
rect 165613 468696 165618 468752
rect 165674 468696 168084 468752
rect 165613 468694 168084 468696
rect 165613 468691 165679 468694
rect 390093 468618 390159 468621
rect 387964 468616 390159 468618
rect 387964 468560 390098 468616
rect 390154 468560 390159 468616
rect 387964 468558 390159 468560
rect 390093 468555 390159 468558
rect 165613 466170 165679 466173
rect 165613 466168 168084 466170
rect 165613 466112 165618 466168
rect 165674 466112 168084 466168
rect 165613 466110 168084 466112
rect 165613 466107 165679 466110
rect 390001 465898 390067 465901
rect 387964 465896 390067 465898
rect 387964 465840 390006 465896
rect 390062 465840 390067 465896
rect 387964 465838 390067 465840
rect 390001 465835 390067 465838
rect 165613 463586 165679 463589
rect 165613 463584 168084 463586
rect 165613 463528 165618 463584
rect 165674 463528 168084 463584
rect 165613 463526 168084 463528
rect 165613 463523 165679 463526
rect 390185 463314 390251 463317
rect 387964 463312 390251 463314
rect 387964 463256 390190 463312
rect 390246 463256 390251 463312
rect 387964 463254 390251 463256
rect 390185 463251 390251 463254
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 165613 461002 165679 461005
rect 165613 461000 168084 461002
rect 165613 460944 165618 461000
rect 165674 460944 168084 461000
rect 165613 460942 168084 460944
rect 165613 460939 165679 460942
rect 390277 460730 390343 460733
rect 387964 460728 390343 460730
rect 387964 460672 390282 460728
rect 390338 460672 390343 460728
rect 387964 460670 390343 460672
rect 390277 460667 390343 460670
rect 165613 458418 165679 458421
rect 165613 458416 168084 458418
rect 165613 458360 165618 458416
rect 165674 458360 168084 458416
rect 165613 458358 168084 458360
rect 165613 458355 165679 458358
rect 579797 458146 579863 458149
rect 583520 458146 584960 458236
rect 579797 458144 584960 458146
rect 579797 458088 579802 458144
rect 579858 458088 584960 458144
rect 579797 458086 584960 458088
rect 579797 458083 579863 458086
rect 390185 458010 390251 458013
rect 387964 458008 390251 458010
rect 387964 457952 390190 458008
rect 390246 457952 390251 458008
rect 583520 457996 584960 458086
rect 387964 457950 390251 457952
rect 390185 457947 390251 457950
rect 165613 455834 165679 455837
rect 165613 455832 168084 455834
rect 165613 455776 165618 455832
rect 165674 455776 168084 455832
rect 165613 455774 168084 455776
rect 165613 455771 165679 455774
rect 390369 455426 390435 455429
rect 387964 455424 390435 455426
rect 387964 455368 390374 455424
rect 390430 455368 390435 455424
rect 387964 455366 390435 455368
rect 390369 455363 390435 455366
rect 165613 453250 165679 453253
rect 165613 453248 168084 453250
rect 165613 453192 165618 453248
rect 165674 453192 168084 453248
rect 165613 453190 168084 453192
rect 165613 453187 165679 453190
rect 390461 452706 390527 452709
rect 387964 452704 390527 452706
rect 387964 452648 390466 452704
rect 390522 452648 390527 452704
rect 387964 452646 390527 452648
rect 390461 452643 390527 452646
rect 165613 450666 165679 450669
rect 165613 450664 168084 450666
rect 165613 450608 165618 450664
rect 165674 450608 168084 450664
rect 165613 450606 168084 450608
rect 165613 450603 165679 450606
rect 390185 450122 390251 450125
rect 387964 450120 390251 450122
rect 387964 450064 390190 450120
rect 390246 450064 390251 450120
rect 387964 450062 390251 450064
rect 390185 450059 390251 450062
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 165613 448082 165679 448085
rect 165613 448080 168084 448082
rect 165613 448024 165618 448080
rect 165674 448024 168084 448080
rect 165613 448022 168084 448024
rect 165613 448019 165679 448022
rect 390185 447538 390251 447541
rect 387964 447536 390251 447538
rect 387964 447480 390190 447536
rect 390246 447480 390251 447536
rect 387964 447478 390251 447480
rect 390185 447475 390251 447478
rect 165613 445498 165679 445501
rect 165613 445496 168084 445498
rect 165613 445440 165618 445496
rect 165674 445440 168084 445496
rect 165613 445438 168084 445440
rect 165613 445435 165679 445438
rect 389725 444818 389791 444821
rect 387964 444816 389791 444818
rect 387964 444760 389730 444816
rect 389786 444760 389791 444816
rect 387964 444758 389791 444760
rect 389725 444755 389791 444758
rect 580165 444818 580231 444821
rect 583520 444818 584960 444908
rect 580165 444816 584960 444818
rect 580165 444760 580170 444816
rect 580226 444760 584960 444816
rect 580165 444758 584960 444760
rect 580165 444755 580231 444758
rect 583520 444668 584960 444758
rect 165613 442914 165679 442917
rect 165613 442912 168084 442914
rect 165613 442856 165618 442912
rect 165674 442856 168084 442912
rect 165613 442854 168084 442856
rect 165613 442851 165679 442854
rect 389633 442234 389699 442237
rect 387964 442232 389699 442234
rect 387964 442176 389638 442232
rect 389694 442176 389699 442232
rect 387964 442174 389699 442176
rect 389633 442171 389699 442174
rect 165613 440330 165679 440333
rect 165613 440328 168084 440330
rect 165613 440272 165618 440328
rect 165674 440272 168084 440328
rect 165613 440270 168084 440272
rect 165613 440267 165679 440270
rect 390185 439514 390251 439517
rect 387964 439512 390251 439514
rect 387964 439456 390190 439512
rect 390246 439456 390251 439512
rect 387964 439454 390251 439456
rect 390185 439451 390251 439454
rect 165613 437746 165679 437749
rect 165613 437744 168084 437746
rect 165613 437688 165618 437744
rect 165674 437688 168084 437744
rect 165613 437686 168084 437688
rect 165613 437683 165679 437686
rect 390277 436930 390343 436933
rect 387964 436928 390343 436930
rect 387964 436872 390282 436928
rect 390338 436872 390343 436928
rect 387964 436870 390343 436872
rect 390277 436867 390343 436870
rect -960 436658 480 436748
rect 3601 436658 3667 436661
rect -960 436656 3667 436658
rect -960 436600 3606 436656
rect 3662 436600 3667 436656
rect -960 436598 3667 436600
rect -960 436508 480 436598
rect 3601 436595 3667 436598
rect 165613 435162 165679 435165
rect 165613 435160 168084 435162
rect 165613 435104 165618 435160
rect 165674 435104 168084 435160
rect 165613 435102 168084 435104
rect 165613 435099 165679 435102
rect 389541 434210 389607 434213
rect 387964 434208 389607 434210
rect 387964 434152 389546 434208
rect 389602 434152 389607 434208
rect 387964 434150 389607 434152
rect 389541 434147 389607 434150
rect 165613 432578 165679 432581
rect 165613 432576 168084 432578
rect 165613 432520 165618 432576
rect 165674 432520 168084 432576
rect 165613 432518 168084 432520
rect 165613 432515 165679 432518
rect 389817 431626 389883 431629
rect 387964 431624 389883 431626
rect 387964 431568 389822 431624
rect 389878 431568 389883 431624
rect 387964 431566 389883 431568
rect 389817 431563 389883 431566
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 165613 429858 165679 429861
rect 165613 429856 168084 429858
rect 165613 429800 165618 429856
rect 165674 429800 168084 429856
rect 165613 429798 168084 429800
rect 165613 429795 165679 429798
rect 389909 429042 389975 429045
rect 387964 429040 389975 429042
rect 387964 428984 389914 429040
rect 389970 428984 389975 429040
rect 387964 428982 389975 428984
rect 389909 428979 389975 428982
rect 165613 427274 165679 427277
rect 165613 427272 168084 427274
rect 165613 427216 165618 427272
rect 165674 427216 168084 427272
rect 165613 427214 168084 427216
rect 165613 427211 165679 427214
rect 390001 426322 390067 426325
rect 387964 426320 390067 426322
rect 387964 426264 390006 426320
rect 390062 426264 390067 426320
rect 387964 426262 390067 426264
rect 390001 426259 390067 426262
rect 165613 424690 165679 424693
rect 165613 424688 168084 424690
rect 165613 424632 165618 424688
rect 165674 424632 168084 424688
rect 165613 424630 168084 424632
rect 165613 424627 165679 424630
rect 389817 423738 389883 423741
rect 387964 423736 389883 423738
rect -960 423602 480 423692
rect 387964 423680 389822 423736
rect 389878 423680 389883 423736
rect 387964 423678 389883 423680
rect 389817 423675 389883 423678
rect 3785 423602 3851 423605
rect -960 423600 3851 423602
rect -960 423544 3790 423600
rect 3846 423544 3851 423600
rect -960 423542 3851 423544
rect -960 423452 480 423542
rect 3785 423539 3851 423542
rect 165613 422106 165679 422109
rect 165613 422104 168084 422106
rect 165613 422048 165618 422104
rect 165674 422048 168084 422104
rect 165613 422046 168084 422048
rect 165613 422043 165679 422046
rect 390093 421018 390159 421021
rect 387964 421016 390159 421018
rect 387964 420960 390098 421016
rect 390154 420960 390159 421016
rect 387964 420958 390159 420960
rect 390093 420955 390159 420958
rect 165613 419522 165679 419525
rect 165613 419520 168084 419522
rect 165613 419464 165618 419520
rect 165674 419464 168084 419520
rect 165613 419462 168084 419464
rect 165613 419459 165679 419462
rect 390185 418434 390251 418437
rect 387964 418432 390251 418434
rect 387964 418376 390190 418432
rect 390246 418376 390251 418432
rect 387964 418374 390251 418376
rect 390185 418371 390251 418374
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 165613 416938 165679 416941
rect 165613 416936 168084 416938
rect 165613 416880 165618 416936
rect 165674 416880 168084 416936
rect 165613 416878 168084 416880
rect 165613 416875 165679 416878
rect 390093 415850 390159 415853
rect 387964 415848 390159 415850
rect 387964 415792 390098 415848
rect 390154 415792 390159 415848
rect 387964 415790 390159 415792
rect 390093 415787 390159 415790
rect 165613 414354 165679 414357
rect 165613 414352 168084 414354
rect 165613 414296 165618 414352
rect 165674 414296 168084 414352
rect 165613 414294 168084 414296
rect 165613 414291 165679 414294
rect 390001 413130 390067 413133
rect 387964 413128 390067 413130
rect 387964 413072 390006 413128
rect 390062 413072 390067 413128
rect 387964 413070 390067 413072
rect 390001 413067 390067 413070
rect 165613 411770 165679 411773
rect 165613 411768 168084 411770
rect 165613 411712 165618 411768
rect 165674 411712 168084 411768
rect 165613 411710 168084 411712
rect 165613 411707 165679 411710
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect 389909 410546 389975 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect 387964 410544 389975 410546
rect 387964 410488 389914 410544
rect 389970 410488 389975 410544
rect 387964 410486 389975 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 389909 410483 389975 410486
rect 165613 409186 165679 409189
rect 165613 409184 168084 409186
rect 165613 409128 165618 409184
rect 165674 409128 168084 409184
rect 165613 409126 168084 409128
rect 165613 409123 165679 409126
rect 389817 407826 389883 407829
rect 387964 407824 389883 407826
rect 387964 407768 389822 407824
rect 389878 407768 389883 407824
rect 387964 407766 389883 407768
rect 389817 407763 389883 407766
rect 165613 406602 165679 406605
rect 165613 406600 168084 406602
rect 165613 406544 165618 406600
rect 165674 406544 168084 406600
rect 165613 406542 168084 406544
rect 165613 406539 165679 406542
rect 389173 405242 389239 405245
rect 387964 405240 389239 405242
rect 387964 405184 389178 405240
rect 389234 405184 389239 405240
rect 387964 405182 389239 405184
rect 389173 405179 389239 405182
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 166901 404018 166967 404021
rect 166901 404016 168084 404018
rect 166901 403960 166906 404016
rect 166962 403960 168084 404016
rect 166901 403958 168084 403960
rect 166901 403955 166967 403958
rect 389173 402522 389239 402525
rect 387964 402520 389239 402522
rect 387964 402464 389178 402520
rect 389234 402464 389239 402520
rect 387964 402462 389239 402464
rect 389173 402459 389239 402462
rect 166809 401434 166875 401437
rect 166809 401432 168084 401434
rect 166809 401376 166814 401432
rect 166870 401376 168084 401432
rect 166809 401374 168084 401376
rect 166809 401371 166875 401374
rect 389265 399938 389331 399941
rect 387964 399936 389331 399938
rect 387964 399880 389270 399936
rect 389326 399880 389331 399936
rect 387964 399878 389331 399880
rect 389265 399875 389331 399878
rect 165613 398850 165679 398853
rect 165613 398848 168084 398850
rect 165613 398792 165618 398848
rect 165674 398792 168084 398848
rect 165613 398790 168084 398792
rect 165613 398787 165679 398790
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 389357 397354 389423 397357
rect 387964 397352 389423 397354
rect 387964 397296 389362 397352
rect 389418 397296 389423 397352
rect 387964 397294 389423 397296
rect 389357 397291 389423 397294
rect 165613 396266 165679 396269
rect 165613 396264 168084 396266
rect 165613 396208 165618 396264
rect 165674 396208 168084 396264
rect 165613 396206 168084 396208
rect 165613 396203 165679 396206
rect 390185 394634 390251 394637
rect 387964 394632 390251 394634
rect 387964 394576 390190 394632
rect 390246 394576 390251 394632
rect 387964 394574 390251 394576
rect 390185 394571 390251 394574
rect 166717 393682 166783 393685
rect 166717 393680 168084 393682
rect 166717 393624 166722 393680
rect 166778 393624 168084 393680
rect 166717 393622 168084 393624
rect 166717 393619 166783 393622
rect 390185 392050 390251 392053
rect 387964 392048 390251 392050
rect 387964 391992 390190 392048
rect 390246 391992 390251 392048
rect 387964 391990 390251 391992
rect 390185 391987 390251 391990
rect 580165 391778 580231 391781
rect 583520 391778 584960 391868
rect 580165 391776 584960 391778
rect 580165 391720 580170 391776
rect 580226 391720 584960 391776
rect 580165 391718 584960 391720
rect 580165 391715 580231 391718
rect 583520 391628 584960 391718
rect 166625 391098 166691 391101
rect 166625 391096 168084 391098
rect 166625 391040 166630 391096
rect 166686 391040 168084 391096
rect 166625 391038 168084 391040
rect 166625 391035 166691 391038
rect 390185 389330 390251 389333
rect 387964 389328 390251 389330
rect 387964 389272 390190 389328
rect 390246 389272 390251 389328
rect 387964 389270 390251 389272
rect 390185 389267 390251 389270
rect 165613 388514 165679 388517
rect 165613 388512 168084 388514
rect 165613 388456 165618 388512
rect 165674 388456 168084 388512
rect 165613 388454 168084 388456
rect 165613 388451 165679 388454
rect 389449 386746 389515 386749
rect 387964 386744 389515 386746
rect 387964 386688 389454 386744
rect 389510 386688 389515 386744
rect 387964 386686 389515 386688
rect 389449 386683 389515 386686
rect 165613 385930 165679 385933
rect 165613 385928 168084 385930
rect 165613 385872 165618 385928
rect 165674 385872 168084 385928
rect 165613 385870 168084 385872
rect 165613 385867 165679 385870
rect -960 384434 480 384524
rect 3693 384434 3759 384437
rect -960 384432 3759 384434
rect -960 384376 3698 384432
rect 3754 384376 3759 384432
rect -960 384374 3759 384376
rect -960 384284 480 384374
rect 3693 384371 3759 384374
rect 389541 384162 389607 384165
rect 387964 384160 389607 384162
rect 387964 384104 389546 384160
rect 389602 384104 389607 384160
rect 387964 384102 389607 384104
rect 389541 384099 389607 384102
rect 166533 383210 166599 383213
rect 166533 383208 168084 383210
rect 166533 383152 166538 383208
rect 166594 383152 168084 383208
rect 166533 383150 168084 383152
rect 166533 383147 166599 383150
rect 389633 381442 389699 381445
rect 387964 381440 389699 381442
rect 387964 381384 389638 381440
rect 389694 381384 389699 381440
rect 387964 381382 389699 381384
rect 389633 381379 389699 381382
rect 166441 380626 166507 380629
rect 166441 380624 168084 380626
rect 166441 380568 166446 380624
rect 166502 380568 168084 380624
rect 166441 380566 168084 380568
rect 166441 380563 166507 380566
rect 389725 378858 389791 378861
rect 387964 378856 389791 378858
rect 387964 378800 389730 378856
rect 389786 378800 389791 378856
rect 387964 378798 389791 378800
rect 389725 378795 389791 378798
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 165613 378042 165679 378045
rect 165613 378040 168084 378042
rect 165613 377984 165618 378040
rect 165674 377984 168084 378040
rect 165613 377982 168084 377984
rect 165613 377979 165679 377982
rect 390461 376138 390527 376141
rect 387964 376136 390527 376138
rect 387964 376080 390466 376136
rect 390522 376080 390527 376136
rect 387964 376078 390527 376080
rect 390461 376075 390527 376078
rect 165613 375458 165679 375461
rect 165613 375456 168084 375458
rect 165613 375400 165618 375456
rect 165674 375400 168084 375456
rect 165613 375398 168084 375400
rect 165613 375395 165679 375398
rect 390093 373554 390159 373557
rect 387964 373552 390159 373554
rect 387964 373496 390098 373552
rect 390154 373496 390159 373552
rect 387964 373494 390159 373496
rect 390093 373491 390159 373494
rect 166349 372874 166415 372877
rect 166349 372872 168084 372874
rect 166349 372816 166354 372872
rect 166410 372816 168084 372872
rect 166349 372814 168084 372816
rect 166349 372811 166415 372814
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 390369 370834 390435 370837
rect 387964 370832 390435 370834
rect 387964 370776 390374 370832
rect 390430 370776 390435 370832
rect 387964 370774 390435 370776
rect 390369 370771 390435 370774
rect 165613 370290 165679 370293
rect 165613 370288 168084 370290
rect 165613 370232 165618 370288
rect 165674 370232 168084 370288
rect 165613 370230 168084 370232
rect 165613 370227 165679 370230
rect 390277 368250 390343 368253
rect 387964 368248 390343 368250
rect 387964 368192 390282 368248
rect 390338 368192 390343 368248
rect 387964 368190 390343 368192
rect 390277 368187 390343 368190
rect 165613 367706 165679 367709
rect 165613 367704 168084 367706
rect 165613 367648 165618 367704
rect 165674 367648 168084 367704
rect 165613 367646 168084 367648
rect 165613 367643 165679 367646
rect 390185 365666 390251 365669
rect 387964 365664 390251 365666
rect 387964 365608 390190 365664
rect 390246 365608 390251 365664
rect 387964 365606 390251 365608
rect 390185 365603 390251 365606
rect 165613 365122 165679 365125
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 165613 365120 168084 365122
rect 165613 365064 165618 365120
rect 165674 365064 168084 365120
rect 165613 365062 168084 365064
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 165613 365059 165679 365062
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 389909 362946 389975 362949
rect 387964 362944 389975 362946
rect 387964 362888 389914 362944
rect 389970 362888 389975 362944
rect 387964 362886 389975 362888
rect 389909 362883 389975 362886
rect 166257 362538 166323 362541
rect 166257 362536 168084 362538
rect 166257 362480 166262 362536
rect 166318 362480 168084 362536
rect 166257 362478 168084 362480
rect 166257 362475 166323 362478
rect 390001 360362 390067 360365
rect 387964 360360 390067 360362
rect 387964 360304 390006 360360
rect 390062 360304 390067 360360
rect 387964 360302 390067 360304
rect 390001 360299 390067 360302
rect 165613 359954 165679 359957
rect 165613 359952 168084 359954
rect 165613 359896 165618 359952
rect 165674 359896 168084 359952
rect 165613 359894 168084 359896
rect 165613 359891 165679 359894
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 390093 357642 390159 357645
rect 387964 357640 390159 357642
rect 387964 357584 390098 357640
rect 390154 357584 390159 357640
rect 387964 357582 390159 357584
rect 390093 357579 390159 357582
rect 165613 357370 165679 357373
rect 165613 357368 168084 357370
rect 165613 357312 165618 357368
rect 165674 357312 168084 357368
rect 165613 357310 168084 357312
rect 165613 357307 165679 357310
rect 389909 355058 389975 355061
rect 387964 355056 389975 355058
rect 387964 355000 389914 355056
rect 389970 355000 389975 355056
rect 387964 354998 389975 355000
rect 389909 354995 389975 354998
rect 165613 354786 165679 354789
rect 165613 354784 168084 354786
rect 165613 354728 165618 354784
rect 165674 354728 168084 354784
rect 165613 354726 168084 354728
rect 165613 354723 165679 354726
rect 389909 352474 389975 352477
rect 387964 352472 389975 352474
rect 387964 352416 389914 352472
rect 389970 352416 389975 352472
rect 387964 352414 389975 352416
rect 389909 352411 389975 352414
rect 165613 352202 165679 352205
rect 165613 352200 168084 352202
rect 165613 352144 165618 352200
rect 165674 352144 168084 352200
rect 165613 352142 168084 352144
rect 165613 352139 165679 352142
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 389817 349754 389883 349757
rect 387964 349752 389883 349754
rect 387964 349696 389822 349752
rect 389878 349696 389883 349752
rect 387964 349694 389883 349696
rect 389817 349691 389883 349694
rect 165613 349618 165679 349621
rect 165613 349616 168084 349618
rect 165613 349560 165618 349616
rect 165674 349560 168084 349616
rect 165613 349558 168084 349560
rect 165613 349555 165679 349558
rect 389909 347170 389975 347173
rect 387964 347168 389975 347170
rect 387964 347112 389914 347168
rect 389970 347112 389975 347168
rect 387964 347110 389975 347112
rect 389909 347107 389975 347110
rect 165613 347034 165679 347037
rect 165613 347032 168084 347034
rect 165613 346976 165618 347032
rect 165674 346976 168084 347032
rect 165613 346974 168084 346976
rect 165613 346971 165679 346974
rect -960 345402 480 345492
rect 3417 345402 3483 345405
rect -960 345400 3483 345402
rect -960 345344 3422 345400
rect 3478 345344 3483 345400
rect -960 345342 3483 345344
rect -960 345252 480 345342
rect 3417 345339 3483 345342
rect 165613 344450 165679 344453
rect 389766 344450 389772 344452
rect 165613 344448 168084 344450
rect 165613 344392 165618 344448
rect 165674 344392 168084 344448
rect 165613 344390 168084 344392
rect 387964 344390 389772 344450
rect 165613 344387 165679 344390
rect 389766 344388 389772 344390
rect 389836 344388 389842 344452
rect 165613 341866 165679 341869
rect 165613 341864 168084 341866
rect 165613 341808 165618 341864
rect 165674 341808 168084 341864
rect 165613 341806 168084 341808
rect 165613 341803 165679 341806
rect 387934 341322 387994 341836
rect 389081 341322 389147 341325
rect 387934 341320 389147 341322
rect 387934 341264 389086 341320
rect 389142 341264 389147 341320
rect 387934 341262 389147 341264
rect 389081 341259 389147 341262
rect 165613 339282 165679 339285
rect 165613 339280 168084 339282
rect 165613 339224 165618 339280
rect 165674 339224 168084 339280
rect 165613 339222 168084 339224
rect 165613 339219 165679 339222
rect 387934 338738 387994 339252
rect 389081 338738 389147 338741
rect 387934 338736 389147 338738
rect 387934 338680 389086 338736
rect 389142 338680 389147 338736
rect 387934 338678 389147 338680
rect 389081 338675 389147 338678
rect 580165 338602 580231 338605
rect 583520 338602 584960 338692
rect 580165 338600 584960 338602
rect 580165 338544 580170 338600
rect 580226 338544 584960 338600
rect 580165 338542 584960 338544
rect 580165 338539 580231 338542
rect 583520 338452 584960 338542
rect -960 332346 480 332436
rect 3049 332346 3115 332349
rect -960 332344 3115 332346
rect -960 332288 3054 332344
rect 3110 332288 3115 332344
rect -960 332286 3115 332288
rect -960 332196 480 332286
rect 3049 332283 3115 332286
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3049 319290 3115 319293
rect -960 319288 3115 319290
rect -960 319232 3054 319288
rect 3110 319232 3115 319288
rect -960 319230 3115 319232
rect -960 319140 480 319230
rect 3049 319227 3115 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3141 306234 3207 306237
rect -960 306232 3207 306234
rect -960 306176 3146 306232
rect 3202 306176 3207 306232
rect -960 306174 3207 306176
rect -960 306084 480 306174
rect 3141 306171 3207 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 580257 285426 580323 285429
rect 583520 285426 584960 285516
rect 580257 285424 584960 285426
rect 580257 285368 580262 285424
rect 580318 285368 584960 285424
rect 580257 285366 584960 285368
rect 580257 285363 580323 285366
rect 583520 285276 584960 285366
rect -960 280122 480 280212
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 228034 480 228124
rect 3233 228034 3299 228037
rect -960 228032 3299 228034
rect -960 227976 3238 228032
rect 3294 227976 3299 228032
rect -960 227974 3299 227976
rect -960 227884 480 227974
rect 3233 227971 3299 227974
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3233 214978 3299 214981
rect -960 214976 3299 214978
rect -960 214920 3238 214976
rect 3294 214920 3299 214976
rect -960 214918 3299 214920
rect -960 214828 480 214918
rect 3233 214915 3299 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 3325 175946 3391 175949
rect -960 175944 3391 175946
rect -960 175888 3330 175944
rect 3386 175888 3391 175944
rect -960 175886 3391 175888
rect -960 175796 480 175886
rect 3325 175883 3391 175886
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 4061 162890 4127 162893
rect -960 162888 4127 162890
rect -960 162832 4066 162888
rect 4122 162832 4127 162888
rect -960 162830 4127 162832
rect -960 162740 480 162830
rect 4061 162827 4127 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3969 136778 4035 136781
rect -960 136776 4035 136778
rect -960 136720 3974 136776
rect 4030 136720 4035 136776
rect -960 136718 4035 136720
rect -960 136628 480 136718
rect 3969 136715 4035 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 3141 123722 3207 123725
rect -960 123720 3207 123722
rect -960 123664 3146 123720
rect 3202 123664 3207 123720
rect -960 123662 3207 123664
rect -960 123572 480 123662
rect 3141 123659 3207 123662
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3877 110666 3943 110669
rect -960 110664 3943 110666
rect -960 110608 3882 110664
rect 3938 110608 3943 110664
rect -960 110606 3943 110608
rect -960 110516 480 110606
rect 3877 110603 3943 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3785 97610 3851 97613
rect -960 97608 3851 97610
rect -960 97552 3790 97608
rect 3846 97552 3851 97608
rect -960 97550 3851 97552
rect -960 97460 480 97550
rect 3785 97547 3851 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3693 71634 3759 71637
rect -960 71632 3759 71634
rect -960 71576 3698 71632
rect 3754 71576 3759 71632
rect -960 71574 3759 71576
rect -960 71484 480 71574
rect 3693 71571 3759 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2865 58578 2931 58581
rect -960 58576 2931 58578
rect -960 58520 2870 58576
rect 2926 58520 2931 58576
rect -960 58518 2931 58520
rect -960 58428 480 58518
rect 2865 58515 2931 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3601 45522 3667 45525
rect -960 45520 3667 45522
rect -960 45464 3606 45520
rect 3662 45464 3667 45520
rect -960 45462 3667 45464
rect -960 45372 480 45462
rect 3601 45459 3667 45462
rect 583520 33146 584960 33236
rect 567150 33086 584960 33146
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 389766 31724 389772 31788
rect 389836 31786 389842 31788
rect 567150 31786 567210 33086
rect 583520 32996 584960 33086
rect 389836 31726 567210 31786
rect 389836 31724 389842 31726
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 20621 3770 20687 3773
rect 175549 3770 175615 3773
rect 20621 3768 175615 3770
rect 20621 3712 20626 3768
rect 20682 3712 175554 3768
rect 175610 3712 175615 3768
rect 20621 3710 175615 3712
rect 20621 3707 20687 3710
rect 175549 3707 175615 3710
rect 340781 3770 340847 3773
rect 458081 3770 458147 3773
rect 340781 3768 458147 3770
rect 340781 3712 340786 3768
rect 340842 3712 458086 3768
rect 458142 3712 458147 3768
rect 340781 3710 458147 3712
rect 340781 3707 340847 3710
rect 458081 3707 458147 3710
rect 19425 3634 19491 3637
rect 175365 3634 175431 3637
rect 19425 3632 175431 3634
rect 19425 3576 19430 3632
rect 19486 3576 175370 3632
rect 175426 3576 175431 3632
rect 19425 3574 175431 3576
rect 19425 3571 19491 3574
rect 175365 3571 175431 3574
rect 343541 3634 343607 3637
rect 465165 3634 465231 3637
rect 343541 3632 465231 3634
rect 343541 3576 343546 3632
rect 343602 3576 465170 3632
rect 465226 3576 465231 3632
rect 343541 3574 465231 3576
rect 343541 3571 343607 3574
rect 465165 3571 465231 3574
rect 11145 3498 11211 3501
rect 171317 3498 171383 3501
rect 11145 3496 171383 3498
rect 11145 3440 11150 3496
rect 11206 3440 171322 3496
rect 171378 3440 171383 3496
rect 11145 3438 171383 3440
rect 11145 3435 11211 3438
rect 171317 3435 171383 3438
rect 346301 3498 346367 3501
rect 472249 3498 472315 3501
rect 346301 3496 472315 3498
rect 346301 3440 346306 3496
rect 346362 3440 472254 3496
rect 472310 3440 472315 3496
rect 346301 3438 472315 3440
rect 346301 3435 346367 3438
rect 472249 3435 472315 3438
rect 5257 3362 5323 3365
rect 169937 3362 170003 3365
rect 5257 3360 170003 3362
rect 5257 3304 5262 3360
rect 5318 3304 169942 3360
rect 169998 3304 170003 3360
rect 5257 3302 170003 3304
rect 5257 3299 5323 3302
rect 169937 3299 170003 3302
rect 349061 3362 349127 3365
rect 479333 3362 479399 3365
rect 349061 3360 479399 3362
rect 349061 3304 349066 3360
rect 349122 3304 479338 3360
rect 479394 3304 479399 3360
rect 349061 3302 479399 3304
rect 349061 3299 349127 3302
rect 479333 3299 479399 3302
<< via3 >>
rect 3372 684252 3436 684316
rect 3372 473316 3436 473380
rect 389772 344388 389836 344452
rect 389772 31724 389836 31788
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 680254 -7976 710862
rect -8576 680018 -8394 680254
rect -8158 680018 -7976 680254
rect -8576 679934 -7976 680018
rect -8576 679698 -8394 679934
rect -8158 679698 -7976 679934
rect -8576 644254 -7976 679698
rect -8576 644018 -8394 644254
rect -8158 644018 -7976 644254
rect -8576 643934 -7976 644018
rect -8576 643698 -8394 643934
rect -8158 643698 -7976 643934
rect -8576 608254 -7976 643698
rect -8576 608018 -8394 608254
rect -8158 608018 -7976 608254
rect -8576 607934 -7976 608018
rect -8576 607698 -8394 607934
rect -8158 607698 -7976 607934
rect -8576 572254 -7976 607698
rect -8576 572018 -8394 572254
rect -8158 572018 -7976 572254
rect -8576 571934 -7976 572018
rect -8576 571698 -8394 571934
rect -8158 571698 -7976 571934
rect -8576 536254 -7976 571698
rect -8576 536018 -8394 536254
rect -8158 536018 -7976 536254
rect -8576 535934 -7976 536018
rect -8576 535698 -8394 535934
rect -8158 535698 -7976 535934
rect -8576 500254 -7976 535698
rect -8576 500018 -8394 500254
rect -8158 500018 -7976 500254
rect -8576 499934 -7976 500018
rect -8576 499698 -8394 499934
rect -8158 499698 -7976 499934
rect -8576 464254 -7976 499698
rect -8576 464018 -8394 464254
rect -8158 464018 -7976 464254
rect -8576 463934 -7976 464018
rect -8576 463698 -8394 463934
rect -8158 463698 -7976 463934
rect -8576 428254 -7976 463698
rect -8576 428018 -8394 428254
rect -8158 428018 -7976 428254
rect -8576 427934 -7976 428018
rect -8576 427698 -8394 427934
rect -8158 427698 -7976 427934
rect -8576 392254 -7976 427698
rect -8576 392018 -8394 392254
rect -8158 392018 -7976 392254
rect -8576 391934 -7976 392018
rect -8576 391698 -8394 391934
rect -8158 391698 -7976 391934
rect -8576 356254 -7976 391698
rect -8576 356018 -8394 356254
rect -8158 356018 -7976 356254
rect -8576 355934 -7976 356018
rect -8576 355698 -8394 355934
rect -8158 355698 -7976 355934
rect -8576 320254 -7976 355698
rect -8576 320018 -8394 320254
rect -8158 320018 -7976 320254
rect -8576 319934 -7976 320018
rect -8576 319698 -8394 319934
rect -8158 319698 -7976 319934
rect -8576 284254 -7976 319698
rect -8576 284018 -8394 284254
rect -8158 284018 -7976 284254
rect -8576 283934 -7976 284018
rect -8576 283698 -8394 283934
rect -8158 283698 -7976 283934
rect -8576 248254 -7976 283698
rect -8576 248018 -8394 248254
rect -8158 248018 -7976 248254
rect -8576 247934 -7976 248018
rect -8576 247698 -8394 247934
rect -8158 247698 -7976 247934
rect -8576 212254 -7976 247698
rect -8576 212018 -8394 212254
rect -8158 212018 -7976 212254
rect -8576 211934 -7976 212018
rect -8576 211698 -8394 211934
rect -8158 211698 -7976 211934
rect -8576 176254 -7976 211698
rect -8576 176018 -8394 176254
rect -8158 176018 -7976 176254
rect -8576 175934 -7976 176018
rect -8576 175698 -8394 175934
rect -8158 175698 -7976 175934
rect -8576 140254 -7976 175698
rect -8576 140018 -8394 140254
rect -8158 140018 -7976 140254
rect -8576 139934 -7976 140018
rect -8576 139698 -8394 139934
rect -8158 139698 -7976 139934
rect -8576 104254 -7976 139698
rect -8576 104018 -8394 104254
rect -8158 104018 -7976 104254
rect -8576 103934 -7976 104018
rect -8576 103698 -8394 103934
rect -8158 103698 -7976 103934
rect -8576 68254 -7976 103698
rect -8576 68018 -8394 68254
rect -8158 68018 -7976 68254
rect -8576 67934 -7976 68018
rect -8576 67698 -8394 67934
rect -8158 67698 -7976 67934
rect -8576 32254 -7976 67698
rect -8576 32018 -8394 32254
rect -8158 32018 -7976 32254
rect -8576 31934 -7976 32018
rect -8576 31698 -8394 31934
rect -8158 31698 -7976 31934
rect -8576 -6926 -7976 31698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 698254 -7036 709922
rect 12604 710478 13204 711440
rect 12604 710242 12786 710478
rect 13022 710242 13204 710478
rect 12604 710158 13204 710242
rect 12604 709922 12786 710158
rect 13022 709922 13204 710158
rect -7636 698018 -7454 698254
rect -7218 698018 -7036 698254
rect -7636 697934 -7036 698018
rect -7636 697698 -7454 697934
rect -7218 697698 -7036 697934
rect -7636 662254 -7036 697698
rect -7636 662018 -7454 662254
rect -7218 662018 -7036 662254
rect -7636 661934 -7036 662018
rect -7636 661698 -7454 661934
rect -7218 661698 -7036 661934
rect -7636 626254 -7036 661698
rect -7636 626018 -7454 626254
rect -7218 626018 -7036 626254
rect -7636 625934 -7036 626018
rect -7636 625698 -7454 625934
rect -7218 625698 -7036 625934
rect -7636 590254 -7036 625698
rect -7636 590018 -7454 590254
rect -7218 590018 -7036 590254
rect -7636 589934 -7036 590018
rect -7636 589698 -7454 589934
rect -7218 589698 -7036 589934
rect -7636 554254 -7036 589698
rect -7636 554018 -7454 554254
rect -7218 554018 -7036 554254
rect -7636 553934 -7036 554018
rect -7636 553698 -7454 553934
rect -7218 553698 -7036 553934
rect -7636 518254 -7036 553698
rect -7636 518018 -7454 518254
rect -7218 518018 -7036 518254
rect -7636 517934 -7036 518018
rect -7636 517698 -7454 517934
rect -7218 517698 -7036 517934
rect -7636 482254 -7036 517698
rect -7636 482018 -7454 482254
rect -7218 482018 -7036 482254
rect -7636 481934 -7036 482018
rect -7636 481698 -7454 481934
rect -7218 481698 -7036 481934
rect -7636 446254 -7036 481698
rect -7636 446018 -7454 446254
rect -7218 446018 -7036 446254
rect -7636 445934 -7036 446018
rect -7636 445698 -7454 445934
rect -7218 445698 -7036 445934
rect -7636 410254 -7036 445698
rect -7636 410018 -7454 410254
rect -7218 410018 -7036 410254
rect -7636 409934 -7036 410018
rect -7636 409698 -7454 409934
rect -7218 409698 -7036 409934
rect -7636 374254 -7036 409698
rect -7636 374018 -7454 374254
rect -7218 374018 -7036 374254
rect -7636 373934 -7036 374018
rect -7636 373698 -7454 373934
rect -7218 373698 -7036 373934
rect -7636 338254 -7036 373698
rect -7636 338018 -7454 338254
rect -7218 338018 -7036 338254
rect -7636 337934 -7036 338018
rect -7636 337698 -7454 337934
rect -7218 337698 -7036 337934
rect -7636 302254 -7036 337698
rect -7636 302018 -7454 302254
rect -7218 302018 -7036 302254
rect -7636 301934 -7036 302018
rect -7636 301698 -7454 301934
rect -7218 301698 -7036 301934
rect -7636 266254 -7036 301698
rect -7636 266018 -7454 266254
rect -7218 266018 -7036 266254
rect -7636 265934 -7036 266018
rect -7636 265698 -7454 265934
rect -7218 265698 -7036 265934
rect -7636 230254 -7036 265698
rect -7636 230018 -7454 230254
rect -7218 230018 -7036 230254
rect -7636 229934 -7036 230018
rect -7636 229698 -7454 229934
rect -7218 229698 -7036 229934
rect -7636 194254 -7036 229698
rect -7636 194018 -7454 194254
rect -7218 194018 -7036 194254
rect -7636 193934 -7036 194018
rect -7636 193698 -7454 193934
rect -7218 193698 -7036 193934
rect -7636 158254 -7036 193698
rect -7636 158018 -7454 158254
rect -7218 158018 -7036 158254
rect -7636 157934 -7036 158018
rect -7636 157698 -7454 157934
rect -7218 157698 -7036 157934
rect -7636 122254 -7036 157698
rect -7636 122018 -7454 122254
rect -7218 122018 -7036 122254
rect -7636 121934 -7036 122018
rect -7636 121698 -7454 121934
rect -7218 121698 -7036 121934
rect -7636 86254 -7036 121698
rect -7636 86018 -7454 86254
rect -7218 86018 -7036 86254
rect -7636 85934 -7036 86018
rect -7636 85698 -7454 85934
rect -7218 85698 -7036 85934
rect -7636 50254 -7036 85698
rect -7636 50018 -7454 50254
rect -7218 50018 -7036 50254
rect -7636 49934 -7036 50018
rect -7636 49698 -7454 49934
rect -7218 49698 -7036 49934
rect -7636 14254 -7036 49698
rect -7636 14018 -7454 14254
rect -7218 14018 -7036 14254
rect -7636 13934 -7036 14018
rect -7636 13698 -7454 13934
rect -7218 13698 -7036 13934
rect -7636 -5986 -7036 13698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 676654 -6096 708982
rect -6696 676418 -6514 676654
rect -6278 676418 -6096 676654
rect -6696 676334 -6096 676418
rect -6696 676098 -6514 676334
rect -6278 676098 -6096 676334
rect -6696 640654 -6096 676098
rect -6696 640418 -6514 640654
rect -6278 640418 -6096 640654
rect -6696 640334 -6096 640418
rect -6696 640098 -6514 640334
rect -6278 640098 -6096 640334
rect -6696 604654 -6096 640098
rect -6696 604418 -6514 604654
rect -6278 604418 -6096 604654
rect -6696 604334 -6096 604418
rect -6696 604098 -6514 604334
rect -6278 604098 -6096 604334
rect -6696 568654 -6096 604098
rect -6696 568418 -6514 568654
rect -6278 568418 -6096 568654
rect -6696 568334 -6096 568418
rect -6696 568098 -6514 568334
rect -6278 568098 -6096 568334
rect -6696 532654 -6096 568098
rect -6696 532418 -6514 532654
rect -6278 532418 -6096 532654
rect -6696 532334 -6096 532418
rect -6696 532098 -6514 532334
rect -6278 532098 -6096 532334
rect -6696 496654 -6096 532098
rect -6696 496418 -6514 496654
rect -6278 496418 -6096 496654
rect -6696 496334 -6096 496418
rect -6696 496098 -6514 496334
rect -6278 496098 -6096 496334
rect -6696 460654 -6096 496098
rect -6696 460418 -6514 460654
rect -6278 460418 -6096 460654
rect -6696 460334 -6096 460418
rect -6696 460098 -6514 460334
rect -6278 460098 -6096 460334
rect -6696 424654 -6096 460098
rect -6696 424418 -6514 424654
rect -6278 424418 -6096 424654
rect -6696 424334 -6096 424418
rect -6696 424098 -6514 424334
rect -6278 424098 -6096 424334
rect -6696 388654 -6096 424098
rect -6696 388418 -6514 388654
rect -6278 388418 -6096 388654
rect -6696 388334 -6096 388418
rect -6696 388098 -6514 388334
rect -6278 388098 -6096 388334
rect -6696 352654 -6096 388098
rect -6696 352418 -6514 352654
rect -6278 352418 -6096 352654
rect -6696 352334 -6096 352418
rect -6696 352098 -6514 352334
rect -6278 352098 -6096 352334
rect -6696 316654 -6096 352098
rect -6696 316418 -6514 316654
rect -6278 316418 -6096 316654
rect -6696 316334 -6096 316418
rect -6696 316098 -6514 316334
rect -6278 316098 -6096 316334
rect -6696 280654 -6096 316098
rect -6696 280418 -6514 280654
rect -6278 280418 -6096 280654
rect -6696 280334 -6096 280418
rect -6696 280098 -6514 280334
rect -6278 280098 -6096 280334
rect -6696 244654 -6096 280098
rect -6696 244418 -6514 244654
rect -6278 244418 -6096 244654
rect -6696 244334 -6096 244418
rect -6696 244098 -6514 244334
rect -6278 244098 -6096 244334
rect -6696 208654 -6096 244098
rect -6696 208418 -6514 208654
rect -6278 208418 -6096 208654
rect -6696 208334 -6096 208418
rect -6696 208098 -6514 208334
rect -6278 208098 -6096 208334
rect -6696 172654 -6096 208098
rect -6696 172418 -6514 172654
rect -6278 172418 -6096 172654
rect -6696 172334 -6096 172418
rect -6696 172098 -6514 172334
rect -6278 172098 -6096 172334
rect -6696 136654 -6096 172098
rect -6696 136418 -6514 136654
rect -6278 136418 -6096 136654
rect -6696 136334 -6096 136418
rect -6696 136098 -6514 136334
rect -6278 136098 -6096 136334
rect -6696 100654 -6096 136098
rect -6696 100418 -6514 100654
rect -6278 100418 -6096 100654
rect -6696 100334 -6096 100418
rect -6696 100098 -6514 100334
rect -6278 100098 -6096 100334
rect -6696 64654 -6096 100098
rect -6696 64418 -6514 64654
rect -6278 64418 -6096 64654
rect -6696 64334 -6096 64418
rect -6696 64098 -6514 64334
rect -6278 64098 -6096 64334
rect -6696 28654 -6096 64098
rect -6696 28418 -6514 28654
rect -6278 28418 -6096 28654
rect -6696 28334 -6096 28418
rect -6696 28098 -6514 28334
rect -6278 28098 -6096 28334
rect -6696 -5046 -6096 28098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 694654 -5156 708042
rect 9004 708598 9604 709560
rect 9004 708362 9186 708598
rect 9422 708362 9604 708598
rect 9004 708278 9604 708362
rect 9004 708042 9186 708278
rect 9422 708042 9604 708278
rect -5756 694418 -5574 694654
rect -5338 694418 -5156 694654
rect -5756 694334 -5156 694418
rect -5756 694098 -5574 694334
rect -5338 694098 -5156 694334
rect -5756 658654 -5156 694098
rect -5756 658418 -5574 658654
rect -5338 658418 -5156 658654
rect -5756 658334 -5156 658418
rect -5756 658098 -5574 658334
rect -5338 658098 -5156 658334
rect -5756 622654 -5156 658098
rect -5756 622418 -5574 622654
rect -5338 622418 -5156 622654
rect -5756 622334 -5156 622418
rect -5756 622098 -5574 622334
rect -5338 622098 -5156 622334
rect -5756 586654 -5156 622098
rect -5756 586418 -5574 586654
rect -5338 586418 -5156 586654
rect -5756 586334 -5156 586418
rect -5756 586098 -5574 586334
rect -5338 586098 -5156 586334
rect -5756 550654 -5156 586098
rect -5756 550418 -5574 550654
rect -5338 550418 -5156 550654
rect -5756 550334 -5156 550418
rect -5756 550098 -5574 550334
rect -5338 550098 -5156 550334
rect -5756 514654 -5156 550098
rect -5756 514418 -5574 514654
rect -5338 514418 -5156 514654
rect -5756 514334 -5156 514418
rect -5756 514098 -5574 514334
rect -5338 514098 -5156 514334
rect -5756 478654 -5156 514098
rect -5756 478418 -5574 478654
rect -5338 478418 -5156 478654
rect -5756 478334 -5156 478418
rect -5756 478098 -5574 478334
rect -5338 478098 -5156 478334
rect -5756 442654 -5156 478098
rect -5756 442418 -5574 442654
rect -5338 442418 -5156 442654
rect -5756 442334 -5156 442418
rect -5756 442098 -5574 442334
rect -5338 442098 -5156 442334
rect -5756 406654 -5156 442098
rect -5756 406418 -5574 406654
rect -5338 406418 -5156 406654
rect -5756 406334 -5156 406418
rect -5756 406098 -5574 406334
rect -5338 406098 -5156 406334
rect -5756 370654 -5156 406098
rect -5756 370418 -5574 370654
rect -5338 370418 -5156 370654
rect -5756 370334 -5156 370418
rect -5756 370098 -5574 370334
rect -5338 370098 -5156 370334
rect -5756 334654 -5156 370098
rect -5756 334418 -5574 334654
rect -5338 334418 -5156 334654
rect -5756 334334 -5156 334418
rect -5756 334098 -5574 334334
rect -5338 334098 -5156 334334
rect -5756 298654 -5156 334098
rect -5756 298418 -5574 298654
rect -5338 298418 -5156 298654
rect -5756 298334 -5156 298418
rect -5756 298098 -5574 298334
rect -5338 298098 -5156 298334
rect -5756 262654 -5156 298098
rect -5756 262418 -5574 262654
rect -5338 262418 -5156 262654
rect -5756 262334 -5156 262418
rect -5756 262098 -5574 262334
rect -5338 262098 -5156 262334
rect -5756 226654 -5156 262098
rect -5756 226418 -5574 226654
rect -5338 226418 -5156 226654
rect -5756 226334 -5156 226418
rect -5756 226098 -5574 226334
rect -5338 226098 -5156 226334
rect -5756 190654 -5156 226098
rect -5756 190418 -5574 190654
rect -5338 190418 -5156 190654
rect -5756 190334 -5156 190418
rect -5756 190098 -5574 190334
rect -5338 190098 -5156 190334
rect -5756 154654 -5156 190098
rect -5756 154418 -5574 154654
rect -5338 154418 -5156 154654
rect -5756 154334 -5156 154418
rect -5756 154098 -5574 154334
rect -5338 154098 -5156 154334
rect -5756 118654 -5156 154098
rect -5756 118418 -5574 118654
rect -5338 118418 -5156 118654
rect -5756 118334 -5156 118418
rect -5756 118098 -5574 118334
rect -5338 118098 -5156 118334
rect -5756 82654 -5156 118098
rect -5756 82418 -5574 82654
rect -5338 82418 -5156 82654
rect -5756 82334 -5156 82418
rect -5756 82098 -5574 82334
rect -5338 82098 -5156 82334
rect -5756 46654 -5156 82098
rect -5756 46418 -5574 46654
rect -5338 46418 -5156 46654
rect -5756 46334 -5156 46418
rect -5756 46098 -5574 46334
rect -5338 46098 -5156 46334
rect -5756 10654 -5156 46098
rect -5756 10418 -5574 10654
rect -5338 10418 -5156 10654
rect -5756 10334 -5156 10418
rect -5756 10098 -5574 10334
rect -5338 10098 -5156 10334
rect -5756 -4106 -5156 10098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 673054 -4216 707102
rect -4816 672818 -4634 673054
rect -4398 672818 -4216 673054
rect -4816 672734 -4216 672818
rect -4816 672498 -4634 672734
rect -4398 672498 -4216 672734
rect -4816 637054 -4216 672498
rect -4816 636818 -4634 637054
rect -4398 636818 -4216 637054
rect -4816 636734 -4216 636818
rect -4816 636498 -4634 636734
rect -4398 636498 -4216 636734
rect -4816 601054 -4216 636498
rect -4816 600818 -4634 601054
rect -4398 600818 -4216 601054
rect -4816 600734 -4216 600818
rect -4816 600498 -4634 600734
rect -4398 600498 -4216 600734
rect -4816 565054 -4216 600498
rect -4816 564818 -4634 565054
rect -4398 564818 -4216 565054
rect -4816 564734 -4216 564818
rect -4816 564498 -4634 564734
rect -4398 564498 -4216 564734
rect -4816 529054 -4216 564498
rect -4816 528818 -4634 529054
rect -4398 528818 -4216 529054
rect -4816 528734 -4216 528818
rect -4816 528498 -4634 528734
rect -4398 528498 -4216 528734
rect -4816 493054 -4216 528498
rect -4816 492818 -4634 493054
rect -4398 492818 -4216 493054
rect -4816 492734 -4216 492818
rect -4816 492498 -4634 492734
rect -4398 492498 -4216 492734
rect -4816 457054 -4216 492498
rect -4816 456818 -4634 457054
rect -4398 456818 -4216 457054
rect -4816 456734 -4216 456818
rect -4816 456498 -4634 456734
rect -4398 456498 -4216 456734
rect -4816 421054 -4216 456498
rect -4816 420818 -4634 421054
rect -4398 420818 -4216 421054
rect -4816 420734 -4216 420818
rect -4816 420498 -4634 420734
rect -4398 420498 -4216 420734
rect -4816 385054 -4216 420498
rect -4816 384818 -4634 385054
rect -4398 384818 -4216 385054
rect -4816 384734 -4216 384818
rect -4816 384498 -4634 384734
rect -4398 384498 -4216 384734
rect -4816 349054 -4216 384498
rect -4816 348818 -4634 349054
rect -4398 348818 -4216 349054
rect -4816 348734 -4216 348818
rect -4816 348498 -4634 348734
rect -4398 348498 -4216 348734
rect -4816 313054 -4216 348498
rect -4816 312818 -4634 313054
rect -4398 312818 -4216 313054
rect -4816 312734 -4216 312818
rect -4816 312498 -4634 312734
rect -4398 312498 -4216 312734
rect -4816 277054 -4216 312498
rect -4816 276818 -4634 277054
rect -4398 276818 -4216 277054
rect -4816 276734 -4216 276818
rect -4816 276498 -4634 276734
rect -4398 276498 -4216 276734
rect -4816 241054 -4216 276498
rect -4816 240818 -4634 241054
rect -4398 240818 -4216 241054
rect -4816 240734 -4216 240818
rect -4816 240498 -4634 240734
rect -4398 240498 -4216 240734
rect -4816 205054 -4216 240498
rect -4816 204818 -4634 205054
rect -4398 204818 -4216 205054
rect -4816 204734 -4216 204818
rect -4816 204498 -4634 204734
rect -4398 204498 -4216 204734
rect -4816 169054 -4216 204498
rect -4816 168818 -4634 169054
rect -4398 168818 -4216 169054
rect -4816 168734 -4216 168818
rect -4816 168498 -4634 168734
rect -4398 168498 -4216 168734
rect -4816 133054 -4216 168498
rect -4816 132818 -4634 133054
rect -4398 132818 -4216 133054
rect -4816 132734 -4216 132818
rect -4816 132498 -4634 132734
rect -4398 132498 -4216 132734
rect -4816 97054 -4216 132498
rect -4816 96818 -4634 97054
rect -4398 96818 -4216 97054
rect -4816 96734 -4216 96818
rect -4816 96498 -4634 96734
rect -4398 96498 -4216 96734
rect -4816 61054 -4216 96498
rect -4816 60818 -4634 61054
rect -4398 60818 -4216 61054
rect -4816 60734 -4216 60818
rect -4816 60498 -4634 60734
rect -4398 60498 -4216 60734
rect -4816 25054 -4216 60498
rect -4816 24818 -4634 25054
rect -4398 24818 -4216 25054
rect -4816 24734 -4216 24818
rect -4816 24498 -4634 24734
rect -4398 24498 -4216 24734
rect -4816 -3166 -4216 24498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 691054 -3276 706162
rect 5404 706718 6004 707680
rect 5404 706482 5586 706718
rect 5822 706482 6004 706718
rect 5404 706398 6004 706482
rect 5404 706162 5586 706398
rect 5822 706162 6004 706398
rect -3876 690818 -3694 691054
rect -3458 690818 -3276 691054
rect -3876 690734 -3276 690818
rect -3876 690498 -3694 690734
rect -3458 690498 -3276 690734
rect -3876 655054 -3276 690498
rect -3876 654818 -3694 655054
rect -3458 654818 -3276 655054
rect -3876 654734 -3276 654818
rect -3876 654498 -3694 654734
rect -3458 654498 -3276 654734
rect -3876 619054 -3276 654498
rect -3876 618818 -3694 619054
rect -3458 618818 -3276 619054
rect -3876 618734 -3276 618818
rect -3876 618498 -3694 618734
rect -3458 618498 -3276 618734
rect -3876 583054 -3276 618498
rect -3876 582818 -3694 583054
rect -3458 582818 -3276 583054
rect -3876 582734 -3276 582818
rect -3876 582498 -3694 582734
rect -3458 582498 -3276 582734
rect -3876 547054 -3276 582498
rect -3876 546818 -3694 547054
rect -3458 546818 -3276 547054
rect -3876 546734 -3276 546818
rect -3876 546498 -3694 546734
rect -3458 546498 -3276 546734
rect -3876 511054 -3276 546498
rect -3876 510818 -3694 511054
rect -3458 510818 -3276 511054
rect -3876 510734 -3276 510818
rect -3876 510498 -3694 510734
rect -3458 510498 -3276 510734
rect -3876 475054 -3276 510498
rect -3876 474818 -3694 475054
rect -3458 474818 -3276 475054
rect -3876 474734 -3276 474818
rect -3876 474498 -3694 474734
rect -3458 474498 -3276 474734
rect -3876 439054 -3276 474498
rect -3876 438818 -3694 439054
rect -3458 438818 -3276 439054
rect -3876 438734 -3276 438818
rect -3876 438498 -3694 438734
rect -3458 438498 -3276 438734
rect -3876 403054 -3276 438498
rect -3876 402818 -3694 403054
rect -3458 402818 -3276 403054
rect -3876 402734 -3276 402818
rect -3876 402498 -3694 402734
rect -3458 402498 -3276 402734
rect -3876 367054 -3276 402498
rect -3876 366818 -3694 367054
rect -3458 366818 -3276 367054
rect -3876 366734 -3276 366818
rect -3876 366498 -3694 366734
rect -3458 366498 -3276 366734
rect -3876 331054 -3276 366498
rect -3876 330818 -3694 331054
rect -3458 330818 -3276 331054
rect -3876 330734 -3276 330818
rect -3876 330498 -3694 330734
rect -3458 330498 -3276 330734
rect -3876 295054 -3276 330498
rect -3876 294818 -3694 295054
rect -3458 294818 -3276 295054
rect -3876 294734 -3276 294818
rect -3876 294498 -3694 294734
rect -3458 294498 -3276 294734
rect -3876 259054 -3276 294498
rect -3876 258818 -3694 259054
rect -3458 258818 -3276 259054
rect -3876 258734 -3276 258818
rect -3876 258498 -3694 258734
rect -3458 258498 -3276 258734
rect -3876 223054 -3276 258498
rect -3876 222818 -3694 223054
rect -3458 222818 -3276 223054
rect -3876 222734 -3276 222818
rect -3876 222498 -3694 222734
rect -3458 222498 -3276 222734
rect -3876 187054 -3276 222498
rect -3876 186818 -3694 187054
rect -3458 186818 -3276 187054
rect -3876 186734 -3276 186818
rect -3876 186498 -3694 186734
rect -3458 186498 -3276 186734
rect -3876 151054 -3276 186498
rect -3876 150818 -3694 151054
rect -3458 150818 -3276 151054
rect -3876 150734 -3276 150818
rect -3876 150498 -3694 150734
rect -3458 150498 -3276 150734
rect -3876 115054 -3276 150498
rect -3876 114818 -3694 115054
rect -3458 114818 -3276 115054
rect -3876 114734 -3276 114818
rect -3876 114498 -3694 114734
rect -3458 114498 -3276 114734
rect -3876 79054 -3276 114498
rect -3876 78818 -3694 79054
rect -3458 78818 -3276 79054
rect -3876 78734 -3276 78818
rect -3876 78498 -3694 78734
rect -3458 78498 -3276 78734
rect -3876 43054 -3276 78498
rect -3876 42818 -3694 43054
rect -3458 42818 -3276 43054
rect -3876 42734 -3276 42818
rect -3876 42498 -3694 42734
rect -3458 42498 -3276 42734
rect -3876 7054 -3276 42498
rect -3876 6818 -3694 7054
rect -3458 6818 -3276 7054
rect -3876 6734 -3276 6818
rect -3876 6498 -3694 6734
rect -3458 6498 -3276 6734
rect -3876 -2226 -3276 6498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 669454 -2336 705222
rect -2936 669218 -2754 669454
rect -2518 669218 -2336 669454
rect -2936 669134 -2336 669218
rect -2936 668898 -2754 669134
rect -2518 668898 -2336 669134
rect -2936 633454 -2336 668898
rect -2936 633218 -2754 633454
rect -2518 633218 -2336 633454
rect -2936 633134 -2336 633218
rect -2936 632898 -2754 633134
rect -2518 632898 -2336 633134
rect -2936 597454 -2336 632898
rect -2936 597218 -2754 597454
rect -2518 597218 -2336 597454
rect -2936 597134 -2336 597218
rect -2936 596898 -2754 597134
rect -2518 596898 -2336 597134
rect -2936 561454 -2336 596898
rect -2936 561218 -2754 561454
rect -2518 561218 -2336 561454
rect -2936 561134 -2336 561218
rect -2936 560898 -2754 561134
rect -2518 560898 -2336 561134
rect -2936 525454 -2336 560898
rect -2936 525218 -2754 525454
rect -2518 525218 -2336 525454
rect -2936 525134 -2336 525218
rect -2936 524898 -2754 525134
rect -2518 524898 -2336 525134
rect -2936 489454 -2336 524898
rect -2936 489218 -2754 489454
rect -2518 489218 -2336 489454
rect -2936 489134 -2336 489218
rect -2936 488898 -2754 489134
rect -2518 488898 -2336 489134
rect -2936 453454 -2336 488898
rect -2936 453218 -2754 453454
rect -2518 453218 -2336 453454
rect -2936 453134 -2336 453218
rect -2936 452898 -2754 453134
rect -2518 452898 -2336 453134
rect -2936 417454 -2336 452898
rect -2936 417218 -2754 417454
rect -2518 417218 -2336 417454
rect -2936 417134 -2336 417218
rect -2936 416898 -2754 417134
rect -2518 416898 -2336 417134
rect -2936 381454 -2336 416898
rect -2936 381218 -2754 381454
rect -2518 381218 -2336 381454
rect -2936 381134 -2336 381218
rect -2936 380898 -2754 381134
rect -2518 380898 -2336 381134
rect -2936 345454 -2336 380898
rect -2936 345218 -2754 345454
rect -2518 345218 -2336 345454
rect -2936 345134 -2336 345218
rect -2936 344898 -2754 345134
rect -2518 344898 -2336 345134
rect -2936 309454 -2336 344898
rect -2936 309218 -2754 309454
rect -2518 309218 -2336 309454
rect -2936 309134 -2336 309218
rect -2936 308898 -2754 309134
rect -2518 308898 -2336 309134
rect -2936 273454 -2336 308898
rect -2936 273218 -2754 273454
rect -2518 273218 -2336 273454
rect -2936 273134 -2336 273218
rect -2936 272898 -2754 273134
rect -2518 272898 -2336 273134
rect -2936 237454 -2336 272898
rect -2936 237218 -2754 237454
rect -2518 237218 -2336 237454
rect -2936 237134 -2336 237218
rect -2936 236898 -2754 237134
rect -2518 236898 -2336 237134
rect -2936 201454 -2336 236898
rect -2936 201218 -2754 201454
rect -2518 201218 -2336 201454
rect -2936 201134 -2336 201218
rect -2936 200898 -2754 201134
rect -2518 200898 -2336 201134
rect -2936 165454 -2336 200898
rect -2936 165218 -2754 165454
rect -2518 165218 -2336 165454
rect -2936 165134 -2336 165218
rect -2936 164898 -2754 165134
rect -2518 164898 -2336 165134
rect -2936 129454 -2336 164898
rect -2936 129218 -2754 129454
rect -2518 129218 -2336 129454
rect -2936 129134 -2336 129218
rect -2936 128898 -2754 129134
rect -2518 128898 -2336 129134
rect -2936 93454 -2336 128898
rect -2936 93218 -2754 93454
rect -2518 93218 -2336 93454
rect -2936 93134 -2336 93218
rect -2936 92898 -2754 93134
rect -2518 92898 -2336 93134
rect -2936 57454 -2336 92898
rect -2936 57218 -2754 57454
rect -2518 57218 -2336 57454
rect -2936 57134 -2336 57218
rect -2936 56898 -2754 57134
rect -2518 56898 -2336 57134
rect -2936 21454 -2336 56898
rect -2936 21218 -2754 21454
rect -2518 21218 -2336 21454
rect -2936 21134 -2336 21218
rect -2936 20898 -2754 21134
rect -2518 20898 -2336 21134
rect -2936 -1286 -2336 20898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 687454 -1396 704282
rect -1996 687218 -1814 687454
rect -1578 687218 -1396 687454
rect -1996 687134 -1396 687218
rect -1996 686898 -1814 687134
rect -1578 686898 -1396 687134
rect -1996 651454 -1396 686898
rect -1996 651218 -1814 651454
rect -1578 651218 -1396 651454
rect -1996 651134 -1396 651218
rect -1996 650898 -1814 651134
rect -1578 650898 -1396 651134
rect -1996 615454 -1396 650898
rect -1996 615218 -1814 615454
rect -1578 615218 -1396 615454
rect -1996 615134 -1396 615218
rect -1996 614898 -1814 615134
rect -1578 614898 -1396 615134
rect -1996 579454 -1396 614898
rect -1996 579218 -1814 579454
rect -1578 579218 -1396 579454
rect -1996 579134 -1396 579218
rect -1996 578898 -1814 579134
rect -1578 578898 -1396 579134
rect -1996 543454 -1396 578898
rect -1996 543218 -1814 543454
rect -1578 543218 -1396 543454
rect -1996 543134 -1396 543218
rect -1996 542898 -1814 543134
rect -1578 542898 -1396 543134
rect -1996 507454 -1396 542898
rect -1996 507218 -1814 507454
rect -1578 507218 -1396 507454
rect -1996 507134 -1396 507218
rect -1996 506898 -1814 507134
rect -1578 506898 -1396 507134
rect -1996 471454 -1396 506898
rect -1996 471218 -1814 471454
rect -1578 471218 -1396 471454
rect -1996 471134 -1396 471218
rect -1996 470898 -1814 471134
rect -1578 470898 -1396 471134
rect -1996 435454 -1396 470898
rect -1996 435218 -1814 435454
rect -1578 435218 -1396 435454
rect -1996 435134 -1396 435218
rect -1996 434898 -1814 435134
rect -1578 434898 -1396 435134
rect -1996 399454 -1396 434898
rect -1996 399218 -1814 399454
rect -1578 399218 -1396 399454
rect -1996 399134 -1396 399218
rect -1996 398898 -1814 399134
rect -1578 398898 -1396 399134
rect -1996 363454 -1396 398898
rect -1996 363218 -1814 363454
rect -1578 363218 -1396 363454
rect -1996 363134 -1396 363218
rect -1996 362898 -1814 363134
rect -1578 362898 -1396 363134
rect -1996 327454 -1396 362898
rect -1996 327218 -1814 327454
rect -1578 327218 -1396 327454
rect -1996 327134 -1396 327218
rect -1996 326898 -1814 327134
rect -1578 326898 -1396 327134
rect -1996 291454 -1396 326898
rect -1996 291218 -1814 291454
rect -1578 291218 -1396 291454
rect -1996 291134 -1396 291218
rect -1996 290898 -1814 291134
rect -1578 290898 -1396 291134
rect -1996 255454 -1396 290898
rect -1996 255218 -1814 255454
rect -1578 255218 -1396 255454
rect -1996 255134 -1396 255218
rect -1996 254898 -1814 255134
rect -1578 254898 -1396 255134
rect -1996 219454 -1396 254898
rect -1996 219218 -1814 219454
rect -1578 219218 -1396 219454
rect -1996 219134 -1396 219218
rect -1996 218898 -1814 219134
rect -1578 218898 -1396 219134
rect -1996 183454 -1396 218898
rect -1996 183218 -1814 183454
rect -1578 183218 -1396 183454
rect -1996 183134 -1396 183218
rect -1996 182898 -1814 183134
rect -1578 182898 -1396 183134
rect -1996 147454 -1396 182898
rect -1996 147218 -1814 147454
rect -1578 147218 -1396 147454
rect -1996 147134 -1396 147218
rect -1996 146898 -1814 147134
rect -1578 146898 -1396 147134
rect -1996 111454 -1396 146898
rect -1996 111218 -1814 111454
rect -1578 111218 -1396 111454
rect -1996 111134 -1396 111218
rect -1996 110898 -1814 111134
rect -1578 110898 -1396 111134
rect -1996 75454 -1396 110898
rect -1996 75218 -1814 75454
rect -1578 75218 -1396 75454
rect -1996 75134 -1396 75218
rect -1996 74898 -1814 75134
rect -1578 74898 -1396 75134
rect -1996 39454 -1396 74898
rect -1996 39218 -1814 39454
rect -1578 39218 -1396 39454
rect -1996 39134 -1396 39218
rect -1996 38898 -1814 39134
rect -1578 38898 -1396 39134
rect -1996 3454 -1396 38898
rect -1996 3218 -1814 3454
rect -1578 3218 -1396 3454
rect -1996 3134 -1396 3218
rect -1996 2898 -1814 3134
rect -1578 2898 -1396 3134
rect -1996 -346 -1396 2898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 1804 704838 2404 705800
rect 1804 704602 1986 704838
rect 2222 704602 2404 704838
rect 1804 704518 2404 704602
rect 1804 704282 1986 704518
rect 2222 704282 2404 704518
rect 1804 687454 2404 704282
rect 1804 687218 1986 687454
rect 2222 687218 2404 687454
rect 1804 687134 2404 687218
rect 1804 686898 1986 687134
rect 2222 686898 2404 687134
rect 1804 651454 2404 686898
rect 5404 691054 6004 706162
rect 5404 690818 5586 691054
rect 5822 690818 6004 691054
rect 5404 690734 6004 690818
rect 5404 690498 5586 690734
rect 5822 690498 6004 690734
rect 3371 684316 3437 684317
rect 3371 684252 3372 684316
rect 3436 684252 3437 684316
rect 3371 684251 3437 684252
rect 1804 651218 1986 651454
rect 2222 651218 2404 651454
rect 1804 651134 2404 651218
rect 1804 650898 1986 651134
rect 2222 650898 2404 651134
rect 1804 615454 2404 650898
rect 1804 615218 1986 615454
rect 2222 615218 2404 615454
rect 1804 615134 2404 615218
rect 1804 614898 1986 615134
rect 2222 614898 2404 615134
rect 1804 579454 2404 614898
rect 1804 579218 1986 579454
rect 2222 579218 2404 579454
rect 1804 579134 2404 579218
rect 1804 578898 1986 579134
rect 2222 578898 2404 579134
rect 1804 543454 2404 578898
rect 1804 543218 1986 543454
rect 2222 543218 2404 543454
rect 1804 543134 2404 543218
rect 1804 542898 1986 543134
rect 2222 542898 2404 543134
rect 1804 507454 2404 542898
rect 1804 507218 1986 507454
rect 2222 507218 2404 507454
rect 1804 507134 2404 507218
rect 1804 506898 1986 507134
rect 2222 506898 2404 507134
rect 1804 471454 2404 506898
rect 3374 473381 3434 684251
rect 5404 655054 6004 690498
rect 5404 654818 5586 655054
rect 5822 654818 6004 655054
rect 5404 654734 6004 654818
rect 5404 654498 5586 654734
rect 5822 654498 6004 654734
rect 5404 619054 6004 654498
rect 5404 618818 5586 619054
rect 5822 618818 6004 619054
rect 5404 618734 6004 618818
rect 5404 618498 5586 618734
rect 5822 618498 6004 618734
rect 5404 583054 6004 618498
rect 5404 582818 5586 583054
rect 5822 582818 6004 583054
rect 5404 582734 6004 582818
rect 5404 582498 5586 582734
rect 5822 582498 6004 582734
rect 5404 547054 6004 582498
rect 5404 546818 5586 547054
rect 5822 546818 6004 547054
rect 5404 546734 6004 546818
rect 5404 546498 5586 546734
rect 5822 546498 6004 546734
rect 5404 511054 6004 546498
rect 5404 510818 5586 511054
rect 5822 510818 6004 511054
rect 5404 510734 6004 510818
rect 5404 510498 5586 510734
rect 5822 510498 6004 510734
rect 5404 475054 6004 510498
rect 5404 474818 5586 475054
rect 5822 474818 6004 475054
rect 5404 474734 6004 474818
rect 5404 474498 5586 474734
rect 5822 474498 6004 474734
rect 3371 473380 3437 473381
rect 3371 473316 3372 473380
rect 3436 473316 3437 473380
rect 3371 473315 3437 473316
rect 1804 471218 1986 471454
rect 2222 471218 2404 471454
rect 1804 471134 2404 471218
rect 1804 470898 1986 471134
rect 2222 470898 2404 471134
rect 1804 435454 2404 470898
rect 1804 435218 1986 435454
rect 2222 435218 2404 435454
rect 1804 435134 2404 435218
rect 1804 434898 1986 435134
rect 2222 434898 2404 435134
rect 1804 399454 2404 434898
rect 1804 399218 1986 399454
rect 2222 399218 2404 399454
rect 1804 399134 2404 399218
rect 1804 398898 1986 399134
rect 2222 398898 2404 399134
rect 1804 363454 2404 398898
rect 1804 363218 1986 363454
rect 2222 363218 2404 363454
rect 1804 363134 2404 363218
rect 1804 362898 1986 363134
rect 2222 362898 2404 363134
rect 1804 327454 2404 362898
rect 1804 327218 1986 327454
rect 2222 327218 2404 327454
rect 1804 327134 2404 327218
rect 1804 326898 1986 327134
rect 2222 326898 2404 327134
rect 1804 291454 2404 326898
rect 1804 291218 1986 291454
rect 2222 291218 2404 291454
rect 1804 291134 2404 291218
rect 1804 290898 1986 291134
rect 2222 290898 2404 291134
rect 1804 255454 2404 290898
rect 1804 255218 1986 255454
rect 2222 255218 2404 255454
rect 1804 255134 2404 255218
rect 1804 254898 1986 255134
rect 2222 254898 2404 255134
rect 1804 219454 2404 254898
rect 1804 219218 1986 219454
rect 2222 219218 2404 219454
rect 1804 219134 2404 219218
rect 1804 218898 1986 219134
rect 2222 218898 2404 219134
rect 1804 183454 2404 218898
rect 1804 183218 1986 183454
rect 2222 183218 2404 183454
rect 1804 183134 2404 183218
rect 1804 182898 1986 183134
rect 2222 182898 2404 183134
rect 1804 147454 2404 182898
rect 1804 147218 1986 147454
rect 2222 147218 2404 147454
rect 1804 147134 2404 147218
rect 1804 146898 1986 147134
rect 2222 146898 2404 147134
rect 1804 111454 2404 146898
rect 1804 111218 1986 111454
rect 2222 111218 2404 111454
rect 1804 111134 2404 111218
rect 1804 110898 1986 111134
rect 2222 110898 2404 111134
rect 1804 75454 2404 110898
rect 1804 75218 1986 75454
rect 2222 75218 2404 75454
rect 1804 75134 2404 75218
rect 1804 74898 1986 75134
rect 2222 74898 2404 75134
rect 1804 39454 2404 74898
rect 1804 39218 1986 39454
rect 2222 39218 2404 39454
rect 1804 39134 2404 39218
rect 1804 38898 1986 39134
rect 2222 38898 2404 39134
rect 1804 3454 2404 38898
rect 1804 3218 1986 3454
rect 2222 3218 2404 3454
rect 1804 3134 2404 3218
rect 1804 2898 1986 3134
rect 2222 2898 2404 3134
rect 1804 -346 2404 2898
rect 1804 -582 1986 -346
rect 2222 -582 2404 -346
rect 1804 -666 2404 -582
rect 1804 -902 1986 -666
rect 2222 -902 2404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 1804 -1864 2404 -902
rect 5404 439054 6004 474498
rect 5404 438818 5586 439054
rect 5822 438818 6004 439054
rect 5404 438734 6004 438818
rect 5404 438498 5586 438734
rect 5822 438498 6004 438734
rect 5404 403054 6004 438498
rect 5404 402818 5586 403054
rect 5822 402818 6004 403054
rect 5404 402734 6004 402818
rect 5404 402498 5586 402734
rect 5822 402498 6004 402734
rect 5404 367054 6004 402498
rect 5404 366818 5586 367054
rect 5822 366818 6004 367054
rect 5404 366734 6004 366818
rect 5404 366498 5586 366734
rect 5822 366498 6004 366734
rect 5404 331054 6004 366498
rect 5404 330818 5586 331054
rect 5822 330818 6004 331054
rect 5404 330734 6004 330818
rect 5404 330498 5586 330734
rect 5822 330498 6004 330734
rect 5404 295054 6004 330498
rect 5404 294818 5586 295054
rect 5822 294818 6004 295054
rect 5404 294734 6004 294818
rect 5404 294498 5586 294734
rect 5822 294498 6004 294734
rect 5404 259054 6004 294498
rect 5404 258818 5586 259054
rect 5822 258818 6004 259054
rect 5404 258734 6004 258818
rect 5404 258498 5586 258734
rect 5822 258498 6004 258734
rect 5404 223054 6004 258498
rect 5404 222818 5586 223054
rect 5822 222818 6004 223054
rect 5404 222734 6004 222818
rect 5404 222498 5586 222734
rect 5822 222498 6004 222734
rect 5404 187054 6004 222498
rect 5404 186818 5586 187054
rect 5822 186818 6004 187054
rect 5404 186734 6004 186818
rect 5404 186498 5586 186734
rect 5822 186498 6004 186734
rect 5404 151054 6004 186498
rect 5404 150818 5586 151054
rect 5822 150818 6004 151054
rect 5404 150734 6004 150818
rect 5404 150498 5586 150734
rect 5822 150498 6004 150734
rect 5404 115054 6004 150498
rect 5404 114818 5586 115054
rect 5822 114818 6004 115054
rect 5404 114734 6004 114818
rect 5404 114498 5586 114734
rect 5822 114498 6004 114734
rect 5404 79054 6004 114498
rect 5404 78818 5586 79054
rect 5822 78818 6004 79054
rect 5404 78734 6004 78818
rect 5404 78498 5586 78734
rect 5822 78498 6004 78734
rect 5404 43054 6004 78498
rect 5404 42818 5586 43054
rect 5822 42818 6004 43054
rect 5404 42734 6004 42818
rect 5404 42498 5586 42734
rect 5822 42498 6004 42734
rect 5404 7054 6004 42498
rect 5404 6818 5586 7054
rect 5822 6818 6004 7054
rect 5404 6734 6004 6818
rect 5404 6498 5586 6734
rect 5822 6498 6004 6734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 5404 -2226 6004 6498
rect 5404 -2462 5586 -2226
rect 5822 -2462 6004 -2226
rect 5404 -2546 6004 -2462
rect 5404 -2782 5586 -2546
rect 5822 -2782 6004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 5404 -3744 6004 -2782
rect 9004 694654 9604 708042
rect 9004 694418 9186 694654
rect 9422 694418 9604 694654
rect 9004 694334 9604 694418
rect 9004 694098 9186 694334
rect 9422 694098 9604 694334
rect 9004 658654 9604 694098
rect 9004 658418 9186 658654
rect 9422 658418 9604 658654
rect 9004 658334 9604 658418
rect 9004 658098 9186 658334
rect 9422 658098 9604 658334
rect 9004 622654 9604 658098
rect 9004 622418 9186 622654
rect 9422 622418 9604 622654
rect 9004 622334 9604 622418
rect 9004 622098 9186 622334
rect 9422 622098 9604 622334
rect 9004 586654 9604 622098
rect 9004 586418 9186 586654
rect 9422 586418 9604 586654
rect 9004 586334 9604 586418
rect 9004 586098 9186 586334
rect 9422 586098 9604 586334
rect 9004 550654 9604 586098
rect 9004 550418 9186 550654
rect 9422 550418 9604 550654
rect 9004 550334 9604 550418
rect 9004 550098 9186 550334
rect 9422 550098 9604 550334
rect 9004 514654 9604 550098
rect 9004 514418 9186 514654
rect 9422 514418 9604 514654
rect 9004 514334 9604 514418
rect 9004 514098 9186 514334
rect 9422 514098 9604 514334
rect 9004 478654 9604 514098
rect 9004 478418 9186 478654
rect 9422 478418 9604 478654
rect 9004 478334 9604 478418
rect 9004 478098 9186 478334
rect 9422 478098 9604 478334
rect 9004 442654 9604 478098
rect 9004 442418 9186 442654
rect 9422 442418 9604 442654
rect 9004 442334 9604 442418
rect 9004 442098 9186 442334
rect 9422 442098 9604 442334
rect 9004 406654 9604 442098
rect 9004 406418 9186 406654
rect 9422 406418 9604 406654
rect 9004 406334 9604 406418
rect 9004 406098 9186 406334
rect 9422 406098 9604 406334
rect 9004 370654 9604 406098
rect 9004 370418 9186 370654
rect 9422 370418 9604 370654
rect 9004 370334 9604 370418
rect 9004 370098 9186 370334
rect 9422 370098 9604 370334
rect 9004 334654 9604 370098
rect 9004 334418 9186 334654
rect 9422 334418 9604 334654
rect 9004 334334 9604 334418
rect 9004 334098 9186 334334
rect 9422 334098 9604 334334
rect 9004 298654 9604 334098
rect 9004 298418 9186 298654
rect 9422 298418 9604 298654
rect 9004 298334 9604 298418
rect 9004 298098 9186 298334
rect 9422 298098 9604 298334
rect 9004 262654 9604 298098
rect 9004 262418 9186 262654
rect 9422 262418 9604 262654
rect 9004 262334 9604 262418
rect 9004 262098 9186 262334
rect 9422 262098 9604 262334
rect 9004 226654 9604 262098
rect 9004 226418 9186 226654
rect 9422 226418 9604 226654
rect 9004 226334 9604 226418
rect 9004 226098 9186 226334
rect 9422 226098 9604 226334
rect 9004 190654 9604 226098
rect 9004 190418 9186 190654
rect 9422 190418 9604 190654
rect 9004 190334 9604 190418
rect 9004 190098 9186 190334
rect 9422 190098 9604 190334
rect 9004 154654 9604 190098
rect 9004 154418 9186 154654
rect 9422 154418 9604 154654
rect 9004 154334 9604 154418
rect 9004 154098 9186 154334
rect 9422 154098 9604 154334
rect 9004 118654 9604 154098
rect 9004 118418 9186 118654
rect 9422 118418 9604 118654
rect 9004 118334 9604 118418
rect 9004 118098 9186 118334
rect 9422 118098 9604 118334
rect 9004 82654 9604 118098
rect 9004 82418 9186 82654
rect 9422 82418 9604 82654
rect 9004 82334 9604 82418
rect 9004 82098 9186 82334
rect 9422 82098 9604 82334
rect 9004 46654 9604 82098
rect 9004 46418 9186 46654
rect 9422 46418 9604 46654
rect 9004 46334 9604 46418
rect 9004 46098 9186 46334
rect 9422 46098 9604 46334
rect 9004 10654 9604 46098
rect 9004 10418 9186 10654
rect 9422 10418 9604 10654
rect 9004 10334 9604 10418
rect 9004 10098 9186 10334
rect 9422 10098 9604 10334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 9004 -4106 9604 10098
rect 9004 -4342 9186 -4106
rect 9422 -4342 9604 -4106
rect 9004 -4426 9604 -4342
rect 9004 -4662 9186 -4426
rect 9422 -4662 9604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 9004 -5624 9604 -4662
rect 12604 698254 13204 709922
rect 30604 711418 31204 711440
rect 30604 711182 30786 711418
rect 31022 711182 31204 711418
rect 30604 711098 31204 711182
rect 30604 710862 30786 711098
rect 31022 710862 31204 711098
rect 27004 709538 27604 709560
rect 27004 709302 27186 709538
rect 27422 709302 27604 709538
rect 27004 709218 27604 709302
rect 27004 708982 27186 709218
rect 27422 708982 27604 709218
rect 23404 707658 24004 707680
rect 23404 707422 23586 707658
rect 23822 707422 24004 707658
rect 23404 707338 24004 707422
rect 23404 707102 23586 707338
rect 23822 707102 24004 707338
rect 12604 698018 12786 698254
rect 13022 698018 13204 698254
rect 12604 697934 13204 698018
rect 12604 697698 12786 697934
rect 13022 697698 13204 697934
rect 12604 662254 13204 697698
rect 12604 662018 12786 662254
rect 13022 662018 13204 662254
rect 12604 661934 13204 662018
rect 12604 661698 12786 661934
rect 13022 661698 13204 661934
rect 12604 626254 13204 661698
rect 12604 626018 12786 626254
rect 13022 626018 13204 626254
rect 12604 625934 13204 626018
rect 12604 625698 12786 625934
rect 13022 625698 13204 625934
rect 12604 590254 13204 625698
rect 12604 590018 12786 590254
rect 13022 590018 13204 590254
rect 12604 589934 13204 590018
rect 12604 589698 12786 589934
rect 13022 589698 13204 589934
rect 12604 554254 13204 589698
rect 12604 554018 12786 554254
rect 13022 554018 13204 554254
rect 12604 553934 13204 554018
rect 12604 553698 12786 553934
rect 13022 553698 13204 553934
rect 12604 518254 13204 553698
rect 12604 518018 12786 518254
rect 13022 518018 13204 518254
rect 12604 517934 13204 518018
rect 12604 517698 12786 517934
rect 13022 517698 13204 517934
rect 12604 482254 13204 517698
rect 12604 482018 12786 482254
rect 13022 482018 13204 482254
rect 12604 481934 13204 482018
rect 12604 481698 12786 481934
rect 13022 481698 13204 481934
rect 12604 446254 13204 481698
rect 12604 446018 12786 446254
rect 13022 446018 13204 446254
rect 12604 445934 13204 446018
rect 12604 445698 12786 445934
rect 13022 445698 13204 445934
rect 12604 410254 13204 445698
rect 12604 410018 12786 410254
rect 13022 410018 13204 410254
rect 12604 409934 13204 410018
rect 12604 409698 12786 409934
rect 13022 409698 13204 409934
rect 12604 374254 13204 409698
rect 12604 374018 12786 374254
rect 13022 374018 13204 374254
rect 12604 373934 13204 374018
rect 12604 373698 12786 373934
rect 13022 373698 13204 373934
rect 12604 338254 13204 373698
rect 12604 338018 12786 338254
rect 13022 338018 13204 338254
rect 12604 337934 13204 338018
rect 12604 337698 12786 337934
rect 13022 337698 13204 337934
rect 12604 302254 13204 337698
rect 12604 302018 12786 302254
rect 13022 302018 13204 302254
rect 12604 301934 13204 302018
rect 12604 301698 12786 301934
rect 13022 301698 13204 301934
rect 12604 266254 13204 301698
rect 12604 266018 12786 266254
rect 13022 266018 13204 266254
rect 12604 265934 13204 266018
rect 12604 265698 12786 265934
rect 13022 265698 13204 265934
rect 12604 230254 13204 265698
rect 12604 230018 12786 230254
rect 13022 230018 13204 230254
rect 12604 229934 13204 230018
rect 12604 229698 12786 229934
rect 13022 229698 13204 229934
rect 12604 194254 13204 229698
rect 12604 194018 12786 194254
rect 13022 194018 13204 194254
rect 12604 193934 13204 194018
rect 12604 193698 12786 193934
rect 13022 193698 13204 193934
rect 12604 158254 13204 193698
rect 12604 158018 12786 158254
rect 13022 158018 13204 158254
rect 12604 157934 13204 158018
rect 12604 157698 12786 157934
rect 13022 157698 13204 157934
rect 12604 122254 13204 157698
rect 12604 122018 12786 122254
rect 13022 122018 13204 122254
rect 12604 121934 13204 122018
rect 12604 121698 12786 121934
rect 13022 121698 13204 121934
rect 12604 86254 13204 121698
rect 12604 86018 12786 86254
rect 13022 86018 13204 86254
rect 12604 85934 13204 86018
rect 12604 85698 12786 85934
rect 13022 85698 13204 85934
rect 12604 50254 13204 85698
rect 12604 50018 12786 50254
rect 13022 50018 13204 50254
rect 12604 49934 13204 50018
rect 12604 49698 12786 49934
rect 13022 49698 13204 49934
rect 12604 14254 13204 49698
rect 12604 14018 12786 14254
rect 13022 14018 13204 14254
rect 12604 13934 13204 14018
rect 12604 13698 12786 13934
rect 13022 13698 13204 13934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 12604 -5986 13204 13698
rect 19804 705778 20404 705800
rect 19804 705542 19986 705778
rect 20222 705542 20404 705778
rect 19804 705458 20404 705542
rect 19804 705222 19986 705458
rect 20222 705222 20404 705458
rect 19804 669454 20404 705222
rect 19804 669218 19986 669454
rect 20222 669218 20404 669454
rect 19804 669134 20404 669218
rect 19804 668898 19986 669134
rect 20222 668898 20404 669134
rect 19804 633454 20404 668898
rect 19804 633218 19986 633454
rect 20222 633218 20404 633454
rect 19804 633134 20404 633218
rect 19804 632898 19986 633134
rect 20222 632898 20404 633134
rect 19804 597454 20404 632898
rect 19804 597218 19986 597454
rect 20222 597218 20404 597454
rect 19804 597134 20404 597218
rect 19804 596898 19986 597134
rect 20222 596898 20404 597134
rect 19804 561454 20404 596898
rect 19804 561218 19986 561454
rect 20222 561218 20404 561454
rect 19804 561134 20404 561218
rect 19804 560898 19986 561134
rect 20222 560898 20404 561134
rect 19804 525454 20404 560898
rect 19804 525218 19986 525454
rect 20222 525218 20404 525454
rect 19804 525134 20404 525218
rect 19804 524898 19986 525134
rect 20222 524898 20404 525134
rect 19804 489454 20404 524898
rect 19804 489218 19986 489454
rect 20222 489218 20404 489454
rect 19804 489134 20404 489218
rect 19804 488898 19986 489134
rect 20222 488898 20404 489134
rect 19804 453454 20404 488898
rect 19804 453218 19986 453454
rect 20222 453218 20404 453454
rect 19804 453134 20404 453218
rect 19804 452898 19986 453134
rect 20222 452898 20404 453134
rect 19804 417454 20404 452898
rect 19804 417218 19986 417454
rect 20222 417218 20404 417454
rect 19804 417134 20404 417218
rect 19804 416898 19986 417134
rect 20222 416898 20404 417134
rect 19804 381454 20404 416898
rect 19804 381218 19986 381454
rect 20222 381218 20404 381454
rect 19804 381134 20404 381218
rect 19804 380898 19986 381134
rect 20222 380898 20404 381134
rect 19804 345454 20404 380898
rect 19804 345218 19986 345454
rect 20222 345218 20404 345454
rect 19804 345134 20404 345218
rect 19804 344898 19986 345134
rect 20222 344898 20404 345134
rect 19804 309454 20404 344898
rect 19804 309218 19986 309454
rect 20222 309218 20404 309454
rect 19804 309134 20404 309218
rect 19804 308898 19986 309134
rect 20222 308898 20404 309134
rect 19804 273454 20404 308898
rect 19804 273218 19986 273454
rect 20222 273218 20404 273454
rect 19804 273134 20404 273218
rect 19804 272898 19986 273134
rect 20222 272898 20404 273134
rect 19804 237454 20404 272898
rect 19804 237218 19986 237454
rect 20222 237218 20404 237454
rect 19804 237134 20404 237218
rect 19804 236898 19986 237134
rect 20222 236898 20404 237134
rect 19804 201454 20404 236898
rect 19804 201218 19986 201454
rect 20222 201218 20404 201454
rect 19804 201134 20404 201218
rect 19804 200898 19986 201134
rect 20222 200898 20404 201134
rect 19804 165454 20404 200898
rect 19804 165218 19986 165454
rect 20222 165218 20404 165454
rect 19804 165134 20404 165218
rect 19804 164898 19986 165134
rect 20222 164898 20404 165134
rect 19804 129454 20404 164898
rect 19804 129218 19986 129454
rect 20222 129218 20404 129454
rect 19804 129134 20404 129218
rect 19804 128898 19986 129134
rect 20222 128898 20404 129134
rect 19804 93454 20404 128898
rect 19804 93218 19986 93454
rect 20222 93218 20404 93454
rect 19804 93134 20404 93218
rect 19804 92898 19986 93134
rect 20222 92898 20404 93134
rect 19804 57454 20404 92898
rect 19804 57218 19986 57454
rect 20222 57218 20404 57454
rect 19804 57134 20404 57218
rect 19804 56898 19986 57134
rect 20222 56898 20404 57134
rect 19804 21454 20404 56898
rect 19804 21218 19986 21454
rect 20222 21218 20404 21454
rect 19804 21134 20404 21218
rect 19804 20898 19986 21134
rect 20222 20898 20404 21134
rect 19804 -1286 20404 20898
rect 19804 -1522 19986 -1286
rect 20222 -1522 20404 -1286
rect 19804 -1606 20404 -1522
rect 19804 -1842 19986 -1606
rect 20222 -1842 20404 -1606
rect 19804 -1864 20404 -1842
rect 23404 673054 24004 707102
rect 23404 672818 23586 673054
rect 23822 672818 24004 673054
rect 23404 672734 24004 672818
rect 23404 672498 23586 672734
rect 23822 672498 24004 672734
rect 23404 637054 24004 672498
rect 23404 636818 23586 637054
rect 23822 636818 24004 637054
rect 23404 636734 24004 636818
rect 23404 636498 23586 636734
rect 23822 636498 24004 636734
rect 23404 601054 24004 636498
rect 23404 600818 23586 601054
rect 23822 600818 24004 601054
rect 23404 600734 24004 600818
rect 23404 600498 23586 600734
rect 23822 600498 24004 600734
rect 23404 565054 24004 600498
rect 23404 564818 23586 565054
rect 23822 564818 24004 565054
rect 23404 564734 24004 564818
rect 23404 564498 23586 564734
rect 23822 564498 24004 564734
rect 23404 529054 24004 564498
rect 23404 528818 23586 529054
rect 23822 528818 24004 529054
rect 23404 528734 24004 528818
rect 23404 528498 23586 528734
rect 23822 528498 24004 528734
rect 23404 493054 24004 528498
rect 23404 492818 23586 493054
rect 23822 492818 24004 493054
rect 23404 492734 24004 492818
rect 23404 492498 23586 492734
rect 23822 492498 24004 492734
rect 23404 457054 24004 492498
rect 23404 456818 23586 457054
rect 23822 456818 24004 457054
rect 23404 456734 24004 456818
rect 23404 456498 23586 456734
rect 23822 456498 24004 456734
rect 23404 421054 24004 456498
rect 23404 420818 23586 421054
rect 23822 420818 24004 421054
rect 23404 420734 24004 420818
rect 23404 420498 23586 420734
rect 23822 420498 24004 420734
rect 23404 385054 24004 420498
rect 23404 384818 23586 385054
rect 23822 384818 24004 385054
rect 23404 384734 24004 384818
rect 23404 384498 23586 384734
rect 23822 384498 24004 384734
rect 23404 349054 24004 384498
rect 23404 348818 23586 349054
rect 23822 348818 24004 349054
rect 23404 348734 24004 348818
rect 23404 348498 23586 348734
rect 23822 348498 24004 348734
rect 23404 313054 24004 348498
rect 23404 312818 23586 313054
rect 23822 312818 24004 313054
rect 23404 312734 24004 312818
rect 23404 312498 23586 312734
rect 23822 312498 24004 312734
rect 23404 277054 24004 312498
rect 23404 276818 23586 277054
rect 23822 276818 24004 277054
rect 23404 276734 24004 276818
rect 23404 276498 23586 276734
rect 23822 276498 24004 276734
rect 23404 241054 24004 276498
rect 23404 240818 23586 241054
rect 23822 240818 24004 241054
rect 23404 240734 24004 240818
rect 23404 240498 23586 240734
rect 23822 240498 24004 240734
rect 23404 205054 24004 240498
rect 23404 204818 23586 205054
rect 23822 204818 24004 205054
rect 23404 204734 24004 204818
rect 23404 204498 23586 204734
rect 23822 204498 24004 204734
rect 23404 169054 24004 204498
rect 23404 168818 23586 169054
rect 23822 168818 24004 169054
rect 23404 168734 24004 168818
rect 23404 168498 23586 168734
rect 23822 168498 24004 168734
rect 23404 133054 24004 168498
rect 23404 132818 23586 133054
rect 23822 132818 24004 133054
rect 23404 132734 24004 132818
rect 23404 132498 23586 132734
rect 23822 132498 24004 132734
rect 23404 97054 24004 132498
rect 23404 96818 23586 97054
rect 23822 96818 24004 97054
rect 23404 96734 24004 96818
rect 23404 96498 23586 96734
rect 23822 96498 24004 96734
rect 23404 61054 24004 96498
rect 23404 60818 23586 61054
rect 23822 60818 24004 61054
rect 23404 60734 24004 60818
rect 23404 60498 23586 60734
rect 23822 60498 24004 60734
rect 23404 25054 24004 60498
rect 23404 24818 23586 25054
rect 23822 24818 24004 25054
rect 23404 24734 24004 24818
rect 23404 24498 23586 24734
rect 23822 24498 24004 24734
rect 23404 -3166 24004 24498
rect 23404 -3402 23586 -3166
rect 23822 -3402 24004 -3166
rect 23404 -3486 24004 -3402
rect 23404 -3722 23586 -3486
rect 23822 -3722 24004 -3486
rect 23404 -3744 24004 -3722
rect 27004 676654 27604 708982
rect 27004 676418 27186 676654
rect 27422 676418 27604 676654
rect 27004 676334 27604 676418
rect 27004 676098 27186 676334
rect 27422 676098 27604 676334
rect 27004 640654 27604 676098
rect 27004 640418 27186 640654
rect 27422 640418 27604 640654
rect 27004 640334 27604 640418
rect 27004 640098 27186 640334
rect 27422 640098 27604 640334
rect 27004 604654 27604 640098
rect 27004 604418 27186 604654
rect 27422 604418 27604 604654
rect 27004 604334 27604 604418
rect 27004 604098 27186 604334
rect 27422 604098 27604 604334
rect 27004 568654 27604 604098
rect 27004 568418 27186 568654
rect 27422 568418 27604 568654
rect 27004 568334 27604 568418
rect 27004 568098 27186 568334
rect 27422 568098 27604 568334
rect 27004 532654 27604 568098
rect 27004 532418 27186 532654
rect 27422 532418 27604 532654
rect 27004 532334 27604 532418
rect 27004 532098 27186 532334
rect 27422 532098 27604 532334
rect 27004 496654 27604 532098
rect 27004 496418 27186 496654
rect 27422 496418 27604 496654
rect 27004 496334 27604 496418
rect 27004 496098 27186 496334
rect 27422 496098 27604 496334
rect 27004 460654 27604 496098
rect 27004 460418 27186 460654
rect 27422 460418 27604 460654
rect 27004 460334 27604 460418
rect 27004 460098 27186 460334
rect 27422 460098 27604 460334
rect 27004 424654 27604 460098
rect 27004 424418 27186 424654
rect 27422 424418 27604 424654
rect 27004 424334 27604 424418
rect 27004 424098 27186 424334
rect 27422 424098 27604 424334
rect 27004 388654 27604 424098
rect 27004 388418 27186 388654
rect 27422 388418 27604 388654
rect 27004 388334 27604 388418
rect 27004 388098 27186 388334
rect 27422 388098 27604 388334
rect 27004 352654 27604 388098
rect 27004 352418 27186 352654
rect 27422 352418 27604 352654
rect 27004 352334 27604 352418
rect 27004 352098 27186 352334
rect 27422 352098 27604 352334
rect 27004 316654 27604 352098
rect 27004 316418 27186 316654
rect 27422 316418 27604 316654
rect 27004 316334 27604 316418
rect 27004 316098 27186 316334
rect 27422 316098 27604 316334
rect 27004 280654 27604 316098
rect 27004 280418 27186 280654
rect 27422 280418 27604 280654
rect 27004 280334 27604 280418
rect 27004 280098 27186 280334
rect 27422 280098 27604 280334
rect 27004 244654 27604 280098
rect 27004 244418 27186 244654
rect 27422 244418 27604 244654
rect 27004 244334 27604 244418
rect 27004 244098 27186 244334
rect 27422 244098 27604 244334
rect 27004 208654 27604 244098
rect 27004 208418 27186 208654
rect 27422 208418 27604 208654
rect 27004 208334 27604 208418
rect 27004 208098 27186 208334
rect 27422 208098 27604 208334
rect 27004 172654 27604 208098
rect 27004 172418 27186 172654
rect 27422 172418 27604 172654
rect 27004 172334 27604 172418
rect 27004 172098 27186 172334
rect 27422 172098 27604 172334
rect 27004 136654 27604 172098
rect 27004 136418 27186 136654
rect 27422 136418 27604 136654
rect 27004 136334 27604 136418
rect 27004 136098 27186 136334
rect 27422 136098 27604 136334
rect 27004 100654 27604 136098
rect 27004 100418 27186 100654
rect 27422 100418 27604 100654
rect 27004 100334 27604 100418
rect 27004 100098 27186 100334
rect 27422 100098 27604 100334
rect 27004 64654 27604 100098
rect 27004 64418 27186 64654
rect 27422 64418 27604 64654
rect 27004 64334 27604 64418
rect 27004 64098 27186 64334
rect 27422 64098 27604 64334
rect 27004 28654 27604 64098
rect 27004 28418 27186 28654
rect 27422 28418 27604 28654
rect 27004 28334 27604 28418
rect 27004 28098 27186 28334
rect 27422 28098 27604 28334
rect 27004 -5046 27604 28098
rect 27004 -5282 27186 -5046
rect 27422 -5282 27604 -5046
rect 27004 -5366 27604 -5282
rect 27004 -5602 27186 -5366
rect 27422 -5602 27604 -5366
rect 27004 -5624 27604 -5602
rect 30604 680254 31204 710862
rect 48604 710478 49204 711440
rect 48604 710242 48786 710478
rect 49022 710242 49204 710478
rect 48604 710158 49204 710242
rect 48604 709922 48786 710158
rect 49022 709922 49204 710158
rect 45004 708598 45604 709560
rect 45004 708362 45186 708598
rect 45422 708362 45604 708598
rect 45004 708278 45604 708362
rect 45004 708042 45186 708278
rect 45422 708042 45604 708278
rect 41404 706718 42004 707680
rect 41404 706482 41586 706718
rect 41822 706482 42004 706718
rect 41404 706398 42004 706482
rect 41404 706162 41586 706398
rect 41822 706162 42004 706398
rect 30604 680018 30786 680254
rect 31022 680018 31204 680254
rect 30604 679934 31204 680018
rect 30604 679698 30786 679934
rect 31022 679698 31204 679934
rect 30604 644254 31204 679698
rect 30604 644018 30786 644254
rect 31022 644018 31204 644254
rect 30604 643934 31204 644018
rect 30604 643698 30786 643934
rect 31022 643698 31204 643934
rect 30604 608254 31204 643698
rect 30604 608018 30786 608254
rect 31022 608018 31204 608254
rect 30604 607934 31204 608018
rect 30604 607698 30786 607934
rect 31022 607698 31204 607934
rect 30604 572254 31204 607698
rect 30604 572018 30786 572254
rect 31022 572018 31204 572254
rect 30604 571934 31204 572018
rect 30604 571698 30786 571934
rect 31022 571698 31204 571934
rect 30604 536254 31204 571698
rect 30604 536018 30786 536254
rect 31022 536018 31204 536254
rect 30604 535934 31204 536018
rect 30604 535698 30786 535934
rect 31022 535698 31204 535934
rect 30604 500254 31204 535698
rect 30604 500018 30786 500254
rect 31022 500018 31204 500254
rect 30604 499934 31204 500018
rect 30604 499698 30786 499934
rect 31022 499698 31204 499934
rect 30604 464254 31204 499698
rect 30604 464018 30786 464254
rect 31022 464018 31204 464254
rect 30604 463934 31204 464018
rect 30604 463698 30786 463934
rect 31022 463698 31204 463934
rect 30604 428254 31204 463698
rect 30604 428018 30786 428254
rect 31022 428018 31204 428254
rect 30604 427934 31204 428018
rect 30604 427698 30786 427934
rect 31022 427698 31204 427934
rect 30604 392254 31204 427698
rect 30604 392018 30786 392254
rect 31022 392018 31204 392254
rect 30604 391934 31204 392018
rect 30604 391698 30786 391934
rect 31022 391698 31204 391934
rect 30604 356254 31204 391698
rect 30604 356018 30786 356254
rect 31022 356018 31204 356254
rect 30604 355934 31204 356018
rect 30604 355698 30786 355934
rect 31022 355698 31204 355934
rect 30604 320254 31204 355698
rect 30604 320018 30786 320254
rect 31022 320018 31204 320254
rect 30604 319934 31204 320018
rect 30604 319698 30786 319934
rect 31022 319698 31204 319934
rect 30604 284254 31204 319698
rect 30604 284018 30786 284254
rect 31022 284018 31204 284254
rect 30604 283934 31204 284018
rect 30604 283698 30786 283934
rect 31022 283698 31204 283934
rect 30604 248254 31204 283698
rect 30604 248018 30786 248254
rect 31022 248018 31204 248254
rect 30604 247934 31204 248018
rect 30604 247698 30786 247934
rect 31022 247698 31204 247934
rect 30604 212254 31204 247698
rect 30604 212018 30786 212254
rect 31022 212018 31204 212254
rect 30604 211934 31204 212018
rect 30604 211698 30786 211934
rect 31022 211698 31204 211934
rect 30604 176254 31204 211698
rect 30604 176018 30786 176254
rect 31022 176018 31204 176254
rect 30604 175934 31204 176018
rect 30604 175698 30786 175934
rect 31022 175698 31204 175934
rect 30604 140254 31204 175698
rect 30604 140018 30786 140254
rect 31022 140018 31204 140254
rect 30604 139934 31204 140018
rect 30604 139698 30786 139934
rect 31022 139698 31204 139934
rect 30604 104254 31204 139698
rect 30604 104018 30786 104254
rect 31022 104018 31204 104254
rect 30604 103934 31204 104018
rect 30604 103698 30786 103934
rect 31022 103698 31204 103934
rect 30604 68254 31204 103698
rect 30604 68018 30786 68254
rect 31022 68018 31204 68254
rect 30604 67934 31204 68018
rect 30604 67698 30786 67934
rect 31022 67698 31204 67934
rect 30604 32254 31204 67698
rect 30604 32018 30786 32254
rect 31022 32018 31204 32254
rect 30604 31934 31204 32018
rect 30604 31698 30786 31934
rect 31022 31698 31204 31934
rect 12604 -6222 12786 -5986
rect 13022 -6222 13204 -5986
rect 12604 -6306 13204 -6222
rect 12604 -6542 12786 -6306
rect 13022 -6542 13204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 12604 -7504 13204 -6542
rect 30604 -6926 31204 31698
rect 37804 704838 38404 705800
rect 37804 704602 37986 704838
rect 38222 704602 38404 704838
rect 37804 704518 38404 704602
rect 37804 704282 37986 704518
rect 38222 704282 38404 704518
rect 37804 687454 38404 704282
rect 37804 687218 37986 687454
rect 38222 687218 38404 687454
rect 37804 687134 38404 687218
rect 37804 686898 37986 687134
rect 38222 686898 38404 687134
rect 37804 651454 38404 686898
rect 37804 651218 37986 651454
rect 38222 651218 38404 651454
rect 37804 651134 38404 651218
rect 37804 650898 37986 651134
rect 38222 650898 38404 651134
rect 37804 615454 38404 650898
rect 37804 615218 37986 615454
rect 38222 615218 38404 615454
rect 37804 615134 38404 615218
rect 37804 614898 37986 615134
rect 38222 614898 38404 615134
rect 37804 579454 38404 614898
rect 37804 579218 37986 579454
rect 38222 579218 38404 579454
rect 37804 579134 38404 579218
rect 37804 578898 37986 579134
rect 38222 578898 38404 579134
rect 37804 543454 38404 578898
rect 37804 543218 37986 543454
rect 38222 543218 38404 543454
rect 37804 543134 38404 543218
rect 37804 542898 37986 543134
rect 38222 542898 38404 543134
rect 37804 507454 38404 542898
rect 37804 507218 37986 507454
rect 38222 507218 38404 507454
rect 37804 507134 38404 507218
rect 37804 506898 37986 507134
rect 38222 506898 38404 507134
rect 37804 471454 38404 506898
rect 37804 471218 37986 471454
rect 38222 471218 38404 471454
rect 37804 471134 38404 471218
rect 37804 470898 37986 471134
rect 38222 470898 38404 471134
rect 37804 435454 38404 470898
rect 37804 435218 37986 435454
rect 38222 435218 38404 435454
rect 37804 435134 38404 435218
rect 37804 434898 37986 435134
rect 38222 434898 38404 435134
rect 37804 399454 38404 434898
rect 37804 399218 37986 399454
rect 38222 399218 38404 399454
rect 37804 399134 38404 399218
rect 37804 398898 37986 399134
rect 38222 398898 38404 399134
rect 37804 363454 38404 398898
rect 37804 363218 37986 363454
rect 38222 363218 38404 363454
rect 37804 363134 38404 363218
rect 37804 362898 37986 363134
rect 38222 362898 38404 363134
rect 37804 327454 38404 362898
rect 37804 327218 37986 327454
rect 38222 327218 38404 327454
rect 37804 327134 38404 327218
rect 37804 326898 37986 327134
rect 38222 326898 38404 327134
rect 37804 291454 38404 326898
rect 37804 291218 37986 291454
rect 38222 291218 38404 291454
rect 37804 291134 38404 291218
rect 37804 290898 37986 291134
rect 38222 290898 38404 291134
rect 37804 255454 38404 290898
rect 37804 255218 37986 255454
rect 38222 255218 38404 255454
rect 37804 255134 38404 255218
rect 37804 254898 37986 255134
rect 38222 254898 38404 255134
rect 37804 219454 38404 254898
rect 37804 219218 37986 219454
rect 38222 219218 38404 219454
rect 37804 219134 38404 219218
rect 37804 218898 37986 219134
rect 38222 218898 38404 219134
rect 37804 183454 38404 218898
rect 37804 183218 37986 183454
rect 38222 183218 38404 183454
rect 37804 183134 38404 183218
rect 37804 182898 37986 183134
rect 38222 182898 38404 183134
rect 37804 147454 38404 182898
rect 37804 147218 37986 147454
rect 38222 147218 38404 147454
rect 37804 147134 38404 147218
rect 37804 146898 37986 147134
rect 38222 146898 38404 147134
rect 37804 111454 38404 146898
rect 37804 111218 37986 111454
rect 38222 111218 38404 111454
rect 37804 111134 38404 111218
rect 37804 110898 37986 111134
rect 38222 110898 38404 111134
rect 37804 75454 38404 110898
rect 37804 75218 37986 75454
rect 38222 75218 38404 75454
rect 37804 75134 38404 75218
rect 37804 74898 37986 75134
rect 38222 74898 38404 75134
rect 37804 39454 38404 74898
rect 37804 39218 37986 39454
rect 38222 39218 38404 39454
rect 37804 39134 38404 39218
rect 37804 38898 37986 39134
rect 38222 38898 38404 39134
rect 37804 3454 38404 38898
rect 37804 3218 37986 3454
rect 38222 3218 38404 3454
rect 37804 3134 38404 3218
rect 37804 2898 37986 3134
rect 38222 2898 38404 3134
rect 37804 -346 38404 2898
rect 37804 -582 37986 -346
rect 38222 -582 38404 -346
rect 37804 -666 38404 -582
rect 37804 -902 37986 -666
rect 38222 -902 38404 -666
rect 37804 -1864 38404 -902
rect 41404 691054 42004 706162
rect 41404 690818 41586 691054
rect 41822 690818 42004 691054
rect 41404 690734 42004 690818
rect 41404 690498 41586 690734
rect 41822 690498 42004 690734
rect 41404 655054 42004 690498
rect 41404 654818 41586 655054
rect 41822 654818 42004 655054
rect 41404 654734 42004 654818
rect 41404 654498 41586 654734
rect 41822 654498 42004 654734
rect 41404 619054 42004 654498
rect 41404 618818 41586 619054
rect 41822 618818 42004 619054
rect 41404 618734 42004 618818
rect 41404 618498 41586 618734
rect 41822 618498 42004 618734
rect 41404 583054 42004 618498
rect 41404 582818 41586 583054
rect 41822 582818 42004 583054
rect 41404 582734 42004 582818
rect 41404 582498 41586 582734
rect 41822 582498 42004 582734
rect 41404 547054 42004 582498
rect 41404 546818 41586 547054
rect 41822 546818 42004 547054
rect 41404 546734 42004 546818
rect 41404 546498 41586 546734
rect 41822 546498 42004 546734
rect 41404 511054 42004 546498
rect 41404 510818 41586 511054
rect 41822 510818 42004 511054
rect 41404 510734 42004 510818
rect 41404 510498 41586 510734
rect 41822 510498 42004 510734
rect 41404 475054 42004 510498
rect 41404 474818 41586 475054
rect 41822 474818 42004 475054
rect 41404 474734 42004 474818
rect 41404 474498 41586 474734
rect 41822 474498 42004 474734
rect 41404 439054 42004 474498
rect 41404 438818 41586 439054
rect 41822 438818 42004 439054
rect 41404 438734 42004 438818
rect 41404 438498 41586 438734
rect 41822 438498 42004 438734
rect 41404 403054 42004 438498
rect 41404 402818 41586 403054
rect 41822 402818 42004 403054
rect 41404 402734 42004 402818
rect 41404 402498 41586 402734
rect 41822 402498 42004 402734
rect 41404 367054 42004 402498
rect 41404 366818 41586 367054
rect 41822 366818 42004 367054
rect 41404 366734 42004 366818
rect 41404 366498 41586 366734
rect 41822 366498 42004 366734
rect 41404 331054 42004 366498
rect 41404 330818 41586 331054
rect 41822 330818 42004 331054
rect 41404 330734 42004 330818
rect 41404 330498 41586 330734
rect 41822 330498 42004 330734
rect 41404 295054 42004 330498
rect 41404 294818 41586 295054
rect 41822 294818 42004 295054
rect 41404 294734 42004 294818
rect 41404 294498 41586 294734
rect 41822 294498 42004 294734
rect 41404 259054 42004 294498
rect 41404 258818 41586 259054
rect 41822 258818 42004 259054
rect 41404 258734 42004 258818
rect 41404 258498 41586 258734
rect 41822 258498 42004 258734
rect 41404 223054 42004 258498
rect 41404 222818 41586 223054
rect 41822 222818 42004 223054
rect 41404 222734 42004 222818
rect 41404 222498 41586 222734
rect 41822 222498 42004 222734
rect 41404 187054 42004 222498
rect 41404 186818 41586 187054
rect 41822 186818 42004 187054
rect 41404 186734 42004 186818
rect 41404 186498 41586 186734
rect 41822 186498 42004 186734
rect 41404 151054 42004 186498
rect 41404 150818 41586 151054
rect 41822 150818 42004 151054
rect 41404 150734 42004 150818
rect 41404 150498 41586 150734
rect 41822 150498 42004 150734
rect 41404 115054 42004 150498
rect 41404 114818 41586 115054
rect 41822 114818 42004 115054
rect 41404 114734 42004 114818
rect 41404 114498 41586 114734
rect 41822 114498 42004 114734
rect 41404 79054 42004 114498
rect 41404 78818 41586 79054
rect 41822 78818 42004 79054
rect 41404 78734 42004 78818
rect 41404 78498 41586 78734
rect 41822 78498 42004 78734
rect 41404 43054 42004 78498
rect 41404 42818 41586 43054
rect 41822 42818 42004 43054
rect 41404 42734 42004 42818
rect 41404 42498 41586 42734
rect 41822 42498 42004 42734
rect 41404 7054 42004 42498
rect 41404 6818 41586 7054
rect 41822 6818 42004 7054
rect 41404 6734 42004 6818
rect 41404 6498 41586 6734
rect 41822 6498 42004 6734
rect 41404 -2226 42004 6498
rect 41404 -2462 41586 -2226
rect 41822 -2462 42004 -2226
rect 41404 -2546 42004 -2462
rect 41404 -2782 41586 -2546
rect 41822 -2782 42004 -2546
rect 41404 -3744 42004 -2782
rect 45004 694654 45604 708042
rect 45004 694418 45186 694654
rect 45422 694418 45604 694654
rect 45004 694334 45604 694418
rect 45004 694098 45186 694334
rect 45422 694098 45604 694334
rect 45004 658654 45604 694098
rect 45004 658418 45186 658654
rect 45422 658418 45604 658654
rect 45004 658334 45604 658418
rect 45004 658098 45186 658334
rect 45422 658098 45604 658334
rect 45004 622654 45604 658098
rect 45004 622418 45186 622654
rect 45422 622418 45604 622654
rect 45004 622334 45604 622418
rect 45004 622098 45186 622334
rect 45422 622098 45604 622334
rect 45004 586654 45604 622098
rect 45004 586418 45186 586654
rect 45422 586418 45604 586654
rect 45004 586334 45604 586418
rect 45004 586098 45186 586334
rect 45422 586098 45604 586334
rect 45004 550654 45604 586098
rect 45004 550418 45186 550654
rect 45422 550418 45604 550654
rect 45004 550334 45604 550418
rect 45004 550098 45186 550334
rect 45422 550098 45604 550334
rect 45004 514654 45604 550098
rect 45004 514418 45186 514654
rect 45422 514418 45604 514654
rect 45004 514334 45604 514418
rect 45004 514098 45186 514334
rect 45422 514098 45604 514334
rect 45004 478654 45604 514098
rect 45004 478418 45186 478654
rect 45422 478418 45604 478654
rect 45004 478334 45604 478418
rect 45004 478098 45186 478334
rect 45422 478098 45604 478334
rect 45004 442654 45604 478098
rect 45004 442418 45186 442654
rect 45422 442418 45604 442654
rect 45004 442334 45604 442418
rect 45004 442098 45186 442334
rect 45422 442098 45604 442334
rect 45004 406654 45604 442098
rect 45004 406418 45186 406654
rect 45422 406418 45604 406654
rect 45004 406334 45604 406418
rect 45004 406098 45186 406334
rect 45422 406098 45604 406334
rect 45004 370654 45604 406098
rect 45004 370418 45186 370654
rect 45422 370418 45604 370654
rect 45004 370334 45604 370418
rect 45004 370098 45186 370334
rect 45422 370098 45604 370334
rect 45004 334654 45604 370098
rect 45004 334418 45186 334654
rect 45422 334418 45604 334654
rect 45004 334334 45604 334418
rect 45004 334098 45186 334334
rect 45422 334098 45604 334334
rect 45004 298654 45604 334098
rect 45004 298418 45186 298654
rect 45422 298418 45604 298654
rect 45004 298334 45604 298418
rect 45004 298098 45186 298334
rect 45422 298098 45604 298334
rect 45004 262654 45604 298098
rect 45004 262418 45186 262654
rect 45422 262418 45604 262654
rect 45004 262334 45604 262418
rect 45004 262098 45186 262334
rect 45422 262098 45604 262334
rect 45004 226654 45604 262098
rect 45004 226418 45186 226654
rect 45422 226418 45604 226654
rect 45004 226334 45604 226418
rect 45004 226098 45186 226334
rect 45422 226098 45604 226334
rect 45004 190654 45604 226098
rect 45004 190418 45186 190654
rect 45422 190418 45604 190654
rect 45004 190334 45604 190418
rect 45004 190098 45186 190334
rect 45422 190098 45604 190334
rect 45004 154654 45604 190098
rect 45004 154418 45186 154654
rect 45422 154418 45604 154654
rect 45004 154334 45604 154418
rect 45004 154098 45186 154334
rect 45422 154098 45604 154334
rect 45004 118654 45604 154098
rect 45004 118418 45186 118654
rect 45422 118418 45604 118654
rect 45004 118334 45604 118418
rect 45004 118098 45186 118334
rect 45422 118098 45604 118334
rect 45004 82654 45604 118098
rect 45004 82418 45186 82654
rect 45422 82418 45604 82654
rect 45004 82334 45604 82418
rect 45004 82098 45186 82334
rect 45422 82098 45604 82334
rect 45004 46654 45604 82098
rect 45004 46418 45186 46654
rect 45422 46418 45604 46654
rect 45004 46334 45604 46418
rect 45004 46098 45186 46334
rect 45422 46098 45604 46334
rect 45004 10654 45604 46098
rect 45004 10418 45186 10654
rect 45422 10418 45604 10654
rect 45004 10334 45604 10418
rect 45004 10098 45186 10334
rect 45422 10098 45604 10334
rect 45004 -4106 45604 10098
rect 45004 -4342 45186 -4106
rect 45422 -4342 45604 -4106
rect 45004 -4426 45604 -4342
rect 45004 -4662 45186 -4426
rect 45422 -4662 45604 -4426
rect 45004 -5624 45604 -4662
rect 48604 698254 49204 709922
rect 66604 711418 67204 711440
rect 66604 711182 66786 711418
rect 67022 711182 67204 711418
rect 66604 711098 67204 711182
rect 66604 710862 66786 711098
rect 67022 710862 67204 711098
rect 63004 709538 63604 709560
rect 63004 709302 63186 709538
rect 63422 709302 63604 709538
rect 63004 709218 63604 709302
rect 63004 708982 63186 709218
rect 63422 708982 63604 709218
rect 59404 707658 60004 707680
rect 59404 707422 59586 707658
rect 59822 707422 60004 707658
rect 59404 707338 60004 707422
rect 59404 707102 59586 707338
rect 59822 707102 60004 707338
rect 48604 698018 48786 698254
rect 49022 698018 49204 698254
rect 48604 697934 49204 698018
rect 48604 697698 48786 697934
rect 49022 697698 49204 697934
rect 48604 662254 49204 697698
rect 48604 662018 48786 662254
rect 49022 662018 49204 662254
rect 48604 661934 49204 662018
rect 48604 661698 48786 661934
rect 49022 661698 49204 661934
rect 48604 626254 49204 661698
rect 48604 626018 48786 626254
rect 49022 626018 49204 626254
rect 48604 625934 49204 626018
rect 48604 625698 48786 625934
rect 49022 625698 49204 625934
rect 48604 590254 49204 625698
rect 48604 590018 48786 590254
rect 49022 590018 49204 590254
rect 48604 589934 49204 590018
rect 48604 589698 48786 589934
rect 49022 589698 49204 589934
rect 48604 554254 49204 589698
rect 48604 554018 48786 554254
rect 49022 554018 49204 554254
rect 48604 553934 49204 554018
rect 48604 553698 48786 553934
rect 49022 553698 49204 553934
rect 48604 518254 49204 553698
rect 48604 518018 48786 518254
rect 49022 518018 49204 518254
rect 48604 517934 49204 518018
rect 48604 517698 48786 517934
rect 49022 517698 49204 517934
rect 48604 482254 49204 517698
rect 48604 482018 48786 482254
rect 49022 482018 49204 482254
rect 48604 481934 49204 482018
rect 48604 481698 48786 481934
rect 49022 481698 49204 481934
rect 48604 446254 49204 481698
rect 48604 446018 48786 446254
rect 49022 446018 49204 446254
rect 48604 445934 49204 446018
rect 48604 445698 48786 445934
rect 49022 445698 49204 445934
rect 48604 410254 49204 445698
rect 48604 410018 48786 410254
rect 49022 410018 49204 410254
rect 48604 409934 49204 410018
rect 48604 409698 48786 409934
rect 49022 409698 49204 409934
rect 48604 374254 49204 409698
rect 48604 374018 48786 374254
rect 49022 374018 49204 374254
rect 48604 373934 49204 374018
rect 48604 373698 48786 373934
rect 49022 373698 49204 373934
rect 48604 338254 49204 373698
rect 48604 338018 48786 338254
rect 49022 338018 49204 338254
rect 48604 337934 49204 338018
rect 48604 337698 48786 337934
rect 49022 337698 49204 337934
rect 48604 302254 49204 337698
rect 48604 302018 48786 302254
rect 49022 302018 49204 302254
rect 48604 301934 49204 302018
rect 48604 301698 48786 301934
rect 49022 301698 49204 301934
rect 48604 266254 49204 301698
rect 48604 266018 48786 266254
rect 49022 266018 49204 266254
rect 48604 265934 49204 266018
rect 48604 265698 48786 265934
rect 49022 265698 49204 265934
rect 48604 230254 49204 265698
rect 48604 230018 48786 230254
rect 49022 230018 49204 230254
rect 48604 229934 49204 230018
rect 48604 229698 48786 229934
rect 49022 229698 49204 229934
rect 48604 194254 49204 229698
rect 48604 194018 48786 194254
rect 49022 194018 49204 194254
rect 48604 193934 49204 194018
rect 48604 193698 48786 193934
rect 49022 193698 49204 193934
rect 48604 158254 49204 193698
rect 48604 158018 48786 158254
rect 49022 158018 49204 158254
rect 48604 157934 49204 158018
rect 48604 157698 48786 157934
rect 49022 157698 49204 157934
rect 48604 122254 49204 157698
rect 48604 122018 48786 122254
rect 49022 122018 49204 122254
rect 48604 121934 49204 122018
rect 48604 121698 48786 121934
rect 49022 121698 49204 121934
rect 48604 86254 49204 121698
rect 48604 86018 48786 86254
rect 49022 86018 49204 86254
rect 48604 85934 49204 86018
rect 48604 85698 48786 85934
rect 49022 85698 49204 85934
rect 48604 50254 49204 85698
rect 48604 50018 48786 50254
rect 49022 50018 49204 50254
rect 48604 49934 49204 50018
rect 48604 49698 48786 49934
rect 49022 49698 49204 49934
rect 48604 14254 49204 49698
rect 48604 14018 48786 14254
rect 49022 14018 49204 14254
rect 48604 13934 49204 14018
rect 48604 13698 48786 13934
rect 49022 13698 49204 13934
rect 30604 -7162 30786 -6926
rect 31022 -7162 31204 -6926
rect 30604 -7246 31204 -7162
rect 30604 -7482 30786 -7246
rect 31022 -7482 31204 -7246
rect 30604 -7504 31204 -7482
rect 48604 -5986 49204 13698
rect 55804 705778 56404 705800
rect 55804 705542 55986 705778
rect 56222 705542 56404 705778
rect 55804 705458 56404 705542
rect 55804 705222 55986 705458
rect 56222 705222 56404 705458
rect 55804 669454 56404 705222
rect 55804 669218 55986 669454
rect 56222 669218 56404 669454
rect 55804 669134 56404 669218
rect 55804 668898 55986 669134
rect 56222 668898 56404 669134
rect 55804 633454 56404 668898
rect 55804 633218 55986 633454
rect 56222 633218 56404 633454
rect 55804 633134 56404 633218
rect 55804 632898 55986 633134
rect 56222 632898 56404 633134
rect 55804 597454 56404 632898
rect 55804 597218 55986 597454
rect 56222 597218 56404 597454
rect 55804 597134 56404 597218
rect 55804 596898 55986 597134
rect 56222 596898 56404 597134
rect 55804 561454 56404 596898
rect 55804 561218 55986 561454
rect 56222 561218 56404 561454
rect 55804 561134 56404 561218
rect 55804 560898 55986 561134
rect 56222 560898 56404 561134
rect 55804 525454 56404 560898
rect 55804 525218 55986 525454
rect 56222 525218 56404 525454
rect 55804 525134 56404 525218
rect 55804 524898 55986 525134
rect 56222 524898 56404 525134
rect 55804 489454 56404 524898
rect 55804 489218 55986 489454
rect 56222 489218 56404 489454
rect 55804 489134 56404 489218
rect 55804 488898 55986 489134
rect 56222 488898 56404 489134
rect 55804 453454 56404 488898
rect 55804 453218 55986 453454
rect 56222 453218 56404 453454
rect 55804 453134 56404 453218
rect 55804 452898 55986 453134
rect 56222 452898 56404 453134
rect 55804 417454 56404 452898
rect 55804 417218 55986 417454
rect 56222 417218 56404 417454
rect 55804 417134 56404 417218
rect 55804 416898 55986 417134
rect 56222 416898 56404 417134
rect 55804 381454 56404 416898
rect 55804 381218 55986 381454
rect 56222 381218 56404 381454
rect 55804 381134 56404 381218
rect 55804 380898 55986 381134
rect 56222 380898 56404 381134
rect 55804 345454 56404 380898
rect 55804 345218 55986 345454
rect 56222 345218 56404 345454
rect 55804 345134 56404 345218
rect 55804 344898 55986 345134
rect 56222 344898 56404 345134
rect 55804 309454 56404 344898
rect 55804 309218 55986 309454
rect 56222 309218 56404 309454
rect 55804 309134 56404 309218
rect 55804 308898 55986 309134
rect 56222 308898 56404 309134
rect 55804 273454 56404 308898
rect 55804 273218 55986 273454
rect 56222 273218 56404 273454
rect 55804 273134 56404 273218
rect 55804 272898 55986 273134
rect 56222 272898 56404 273134
rect 55804 237454 56404 272898
rect 55804 237218 55986 237454
rect 56222 237218 56404 237454
rect 55804 237134 56404 237218
rect 55804 236898 55986 237134
rect 56222 236898 56404 237134
rect 55804 201454 56404 236898
rect 55804 201218 55986 201454
rect 56222 201218 56404 201454
rect 55804 201134 56404 201218
rect 55804 200898 55986 201134
rect 56222 200898 56404 201134
rect 55804 165454 56404 200898
rect 55804 165218 55986 165454
rect 56222 165218 56404 165454
rect 55804 165134 56404 165218
rect 55804 164898 55986 165134
rect 56222 164898 56404 165134
rect 55804 129454 56404 164898
rect 55804 129218 55986 129454
rect 56222 129218 56404 129454
rect 55804 129134 56404 129218
rect 55804 128898 55986 129134
rect 56222 128898 56404 129134
rect 55804 93454 56404 128898
rect 55804 93218 55986 93454
rect 56222 93218 56404 93454
rect 55804 93134 56404 93218
rect 55804 92898 55986 93134
rect 56222 92898 56404 93134
rect 55804 57454 56404 92898
rect 55804 57218 55986 57454
rect 56222 57218 56404 57454
rect 55804 57134 56404 57218
rect 55804 56898 55986 57134
rect 56222 56898 56404 57134
rect 55804 21454 56404 56898
rect 55804 21218 55986 21454
rect 56222 21218 56404 21454
rect 55804 21134 56404 21218
rect 55804 20898 55986 21134
rect 56222 20898 56404 21134
rect 55804 -1286 56404 20898
rect 55804 -1522 55986 -1286
rect 56222 -1522 56404 -1286
rect 55804 -1606 56404 -1522
rect 55804 -1842 55986 -1606
rect 56222 -1842 56404 -1606
rect 55804 -1864 56404 -1842
rect 59404 673054 60004 707102
rect 59404 672818 59586 673054
rect 59822 672818 60004 673054
rect 59404 672734 60004 672818
rect 59404 672498 59586 672734
rect 59822 672498 60004 672734
rect 59404 637054 60004 672498
rect 59404 636818 59586 637054
rect 59822 636818 60004 637054
rect 59404 636734 60004 636818
rect 59404 636498 59586 636734
rect 59822 636498 60004 636734
rect 59404 601054 60004 636498
rect 59404 600818 59586 601054
rect 59822 600818 60004 601054
rect 59404 600734 60004 600818
rect 59404 600498 59586 600734
rect 59822 600498 60004 600734
rect 59404 565054 60004 600498
rect 59404 564818 59586 565054
rect 59822 564818 60004 565054
rect 59404 564734 60004 564818
rect 59404 564498 59586 564734
rect 59822 564498 60004 564734
rect 59404 529054 60004 564498
rect 59404 528818 59586 529054
rect 59822 528818 60004 529054
rect 59404 528734 60004 528818
rect 59404 528498 59586 528734
rect 59822 528498 60004 528734
rect 59404 493054 60004 528498
rect 59404 492818 59586 493054
rect 59822 492818 60004 493054
rect 59404 492734 60004 492818
rect 59404 492498 59586 492734
rect 59822 492498 60004 492734
rect 59404 457054 60004 492498
rect 59404 456818 59586 457054
rect 59822 456818 60004 457054
rect 59404 456734 60004 456818
rect 59404 456498 59586 456734
rect 59822 456498 60004 456734
rect 59404 421054 60004 456498
rect 59404 420818 59586 421054
rect 59822 420818 60004 421054
rect 59404 420734 60004 420818
rect 59404 420498 59586 420734
rect 59822 420498 60004 420734
rect 59404 385054 60004 420498
rect 59404 384818 59586 385054
rect 59822 384818 60004 385054
rect 59404 384734 60004 384818
rect 59404 384498 59586 384734
rect 59822 384498 60004 384734
rect 59404 349054 60004 384498
rect 59404 348818 59586 349054
rect 59822 348818 60004 349054
rect 59404 348734 60004 348818
rect 59404 348498 59586 348734
rect 59822 348498 60004 348734
rect 59404 313054 60004 348498
rect 59404 312818 59586 313054
rect 59822 312818 60004 313054
rect 59404 312734 60004 312818
rect 59404 312498 59586 312734
rect 59822 312498 60004 312734
rect 59404 277054 60004 312498
rect 59404 276818 59586 277054
rect 59822 276818 60004 277054
rect 59404 276734 60004 276818
rect 59404 276498 59586 276734
rect 59822 276498 60004 276734
rect 59404 241054 60004 276498
rect 59404 240818 59586 241054
rect 59822 240818 60004 241054
rect 59404 240734 60004 240818
rect 59404 240498 59586 240734
rect 59822 240498 60004 240734
rect 59404 205054 60004 240498
rect 59404 204818 59586 205054
rect 59822 204818 60004 205054
rect 59404 204734 60004 204818
rect 59404 204498 59586 204734
rect 59822 204498 60004 204734
rect 59404 169054 60004 204498
rect 59404 168818 59586 169054
rect 59822 168818 60004 169054
rect 59404 168734 60004 168818
rect 59404 168498 59586 168734
rect 59822 168498 60004 168734
rect 59404 133054 60004 168498
rect 59404 132818 59586 133054
rect 59822 132818 60004 133054
rect 59404 132734 60004 132818
rect 59404 132498 59586 132734
rect 59822 132498 60004 132734
rect 59404 97054 60004 132498
rect 59404 96818 59586 97054
rect 59822 96818 60004 97054
rect 59404 96734 60004 96818
rect 59404 96498 59586 96734
rect 59822 96498 60004 96734
rect 59404 61054 60004 96498
rect 59404 60818 59586 61054
rect 59822 60818 60004 61054
rect 59404 60734 60004 60818
rect 59404 60498 59586 60734
rect 59822 60498 60004 60734
rect 59404 25054 60004 60498
rect 59404 24818 59586 25054
rect 59822 24818 60004 25054
rect 59404 24734 60004 24818
rect 59404 24498 59586 24734
rect 59822 24498 60004 24734
rect 59404 -3166 60004 24498
rect 59404 -3402 59586 -3166
rect 59822 -3402 60004 -3166
rect 59404 -3486 60004 -3402
rect 59404 -3722 59586 -3486
rect 59822 -3722 60004 -3486
rect 59404 -3744 60004 -3722
rect 63004 676654 63604 708982
rect 63004 676418 63186 676654
rect 63422 676418 63604 676654
rect 63004 676334 63604 676418
rect 63004 676098 63186 676334
rect 63422 676098 63604 676334
rect 63004 640654 63604 676098
rect 63004 640418 63186 640654
rect 63422 640418 63604 640654
rect 63004 640334 63604 640418
rect 63004 640098 63186 640334
rect 63422 640098 63604 640334
rect 63004 604654 63604 640098
rect 63004 604418 63186 604654
rect 63422 604418 63604 604654
rect 63004 604334 63604 604418
rect 63004 604098 63186 604334
rect 63422 604098 63604 604334
rect 63004 568654 63604 604098
rect 63004 568418 63186 568654
rect 63422 568418 63604 568654
rect 63004 568334 63604 568418
rect 63004 568098 63186 568334
rect 63422 568098 63604 568334
rect 63004 532654 63604 568098
rect 63004 532418 63186 532654
rect 63422 532418 63604 532654
rect 63004 532334 63604 532418
rect 63004 532098 63186 532334
rect 63422 532098 63604 532334
rect 63004 496654 63604 532098
rect 63004 496418 63186 496654
rect 63422 496418 63604 496654
rect 63004 496334 63604 496418
rect 63004 496098 63186 496334
rect 63422 496098 63604 496334
rect 63004 460654 63604 496098
rect 63004 460418 63186 460654
rect 63422 460418 63604 460654
rect 63004 460334 63604 460418
rect 63004 460098 63186 460334
rect 63422 460098 63604 460334
rect 63004 424654 63604 460098
rect 63004 424418 63186 424654
rect 63422 424418 63604 424654
rect 63004 424334 63604 424418
rect 63004 424098 63186 424334
rect 63422 424098 63604 424334
rect 63004 388654 63604 424098
rect 63004 388418 63186 388654
rect 63422 388418 63604 388654
rect 63004 388334 63604 388418
rect 63004 388098 63186 388334
rect 63422 388098 63604 388334
rect 63004 352654 63604 388098
rect 63004 352418 63186 352654
rect 63422 352418 63604 352654
rect 63004 352334 63604 352418
rect 63004 352098 63186 352334
rect 63422 352098 63604 352334
rect 63004 316654 63604 352098
rect 63004 316418 63186 316654
rect 63422 316418 63604 316654
rect 63004 316334 63604 316418
rect 63004 316098 63186 316334
rect 63422 316098 63604 316334
rect 63004 280654 63604 316098
rect 63004 280418 63186 280654
rect 63422 280418 63604 280654
rect 63004 280334 63604 280418
rect 63004 280098 63186 280334
rect 63422 280098 63604 280334
rect 63004 244654 63604 280098
rect 63004 244418 63186 244654
rect 63422 244418 63604 244654
rect 63004 244334 63604 244418
rect 63004 244098 63186 244334
rect 63422 244098 63604 244334
rect 63004 208654 63604 244098
rect 63004 208418 63186 208654
rect 63422 208418 63604 208654
rect 63004 208334 63604 208418
rect 63004 208098 63186 208334
rect 63422 208098 63604 208334
rect 63004 172654 63604 208098
rect 63004 172418 63186 172654
rect 63422 172418 63604 172654
rect 63004 172334 63604 172418
rect 63004 172098 63186 172334
rect 63422 172098 63604 172334
rect 63004 136654 63604 172098
rect 63004 136418 63186 136654
rect 63422 136418 63604 136654
rect 63004 136334 63604 136418
rect 63004 136098 63186 136334
rect 63422 136098 63604 136334
rect 63004 100654 63604 136098
rect 63004 100418 63186 100654
rect 63422 100418 63604 100654
rect 63004 100334 63604 100418
rect 63004 100098 63186 100334
rect 63422 100098 63604 100334
rect 63004 64654 63604 100098
rect 63004 64418 63186 64654
rect 63422 64418 63604 64654
rect 63004 64334 63604 64418
rect 63004 64098 63186 64334
rect 63422 64098 63604 64334
rect 63004 28654 63604 64098
rect 63004 28418 63186 28654
rect 63422 28418 63604 28654
rect 63004 28334 63604 28418
rect 63004 28098 63186 28334
rect 63422 28098 63604 28334
rect 63004 -5046 63604 28098
rect 63004 -5282 63186 -5046
rect 63422 -5282 63604 -5046
rect 63004 -5366 63604 -5282
rect 63004 -5602 63186 -5366
rect 63422 -5602 63604 -5366
rect 63004 -5624 63604 -5602
rect 66604 680254 67204 710862
rect 84604 710478 85204 711440
rect 84604 710242 84786 710478
rect 85022 710242 85204 710478
rect 84604 710158 85204 710242
rect 84604 709922 84786 710158
rect 85022 709922 85204 710158
rect 81004 708598 81604 709560
rect 81004 708362 81186 708598
rect 81422 708362 81604 708598
rect 81004 708278 81604 708362
rect 81004 708042 81186 708278
rect 81422 708042 81604 708278
rect 77404 706718 78004 707680
rect 77404 706482 77586 706718
rect 77822 706482 78004 706718
rect 77404 706398 78004 706482
rect 77404 706162 77586 706398
rect 77822 706162 78004 706398
rect 66604 680018 66786 680254
rect 67022 680018 67204 680254
rect 66604 679934 67204 680018
rect 66604 679698 66786 679934
rect 67022 679698 67204 679934
rect 66604 644254 67204 679698
rect 66604 644018 66786 644254
rect 67022 644018 67204 644254
rect 66604 643934 67204 644018
rect 66604 643698 66786 643934
rect 67022 643698 67204 643934
rect 66604 608254 67204 643698
rect 66604 608018 66786 608254
rect 67022 608018 67204 608254
rect 66604 607934 67204 608018
rect 66604 607698 66786 607934
rect 67022 607698 67204 607934
rect 66604 572254 67204 607698
rect 66604 572018 66786 572254
rect 67022 572018 67204 572254
rect 66604 571934 67204 572018
rect 66604 571698 66786 571934
rect 67022 571698 67204 571934
rect 66604 536254 67204 571698
rect 66604 536018 66786 536254
rect 67022 536018 67204 536254
rect 66604 535934 67204 536018
rect 66604 535698 66786 535934
rect 67022 535698 67204 535934
rect 66604 500254 67204 535698
rect 66604 500018 66786 500254
rect 67022 500018 67204 500254
rect 66604 499934 67204 500018
rect 66604 499698 66786 499934
rect 67022 499698 67204 499934
rect 66604 464254 67204 499698
rect 66604 464018 66786 464254
rect 67022 464018 67204 464254
rect 66604 463934 67204 464018
rect 66604 463698 66786 463934
rect 67022 463698 67204 463934
rect 66604 428254 67204 463698
rect 66604 428018 66786 428254
rect 67022 428018 67204 428254
rect 66604 427934 67204 428018
rect 66604 427698 66786 427934
rect 67022 427698 67204 427934
rect 66604 392254 67204 427698
rect 66604 392018 66786 392254
rect 67022 392018 67204 392254
rect 66604 391934 67204 392018
rect 66604 391698 66786 391934
rect 67022 391698 67204 391934
rect 66604 356254 67204 391698
rect 66604 356018 66786 356254
rect 67022 356018 67204 356254
rect 66604 355934 67204 356018
rect 66604 355698 66786 355934
rect 67022 355698 67204 355934
rect 66604 320254 67204 355698
rect 66604 320018 66786 320254
rect 67022 320018 67204 320254
rect 66604 319934 67204 320018
rect 66604 319698 66786 319934
rect 67022 319698 67204 319934
rect 66604 284254 67204 319698
rect 66604 284018 66786 284254
rect 67022 284018 67204 284254
rect 66604 283934 67204 284018
rect 66604 283698 66786 283934
rect 67022 283698 67204 283934
rect 66604 248254 67204 283698
rect 66604 248018 66786 248254
rect 67022 248018 67204 248254
rect 66604 247934 67204 248018
rect 66604 247698 66786 247934
rect 67022 247698 67204 247934
rect 66604 212254 67204 247698
rect 66604 212018 66786 212254
rect 67022 212018 67204 212254
rect 66604 211934 67204 212018
rect 66604 211698 66786 211934
rect 67022 211698 67204 211934
rect 66604 176254 67204 211698
rect 66604 176018 66786 176254
rect 67022 176018 67204 176254
rect 66604 175934 67204 176018
rect 66604 175698 66786 175934
rect 67022 175698 67204 175934
rect 66604 140254 67204 175698
rect 66604 140018 66786 140254
rect 67022 140018 67204 140254
rect 66604 139934 67204 140018
rect 66604 139698 66786 139934
rect 67022 139698 67204 139934
rect 66604 104254 67204 139698
rect 66604 104018 66786 104254
rect 67022 104018 67204 104254
rect 66604 103934 67204 104018
rect 66604 103698 66786 103934
rect 67022 103698 67204 103934
rect 66604 68254 67204 103698
rect 66604 68018 66786 68254
rect 67022 68018 67204 68254
rect 66604 67934 67204 68018
rect 66604 67698 66786 67934
rect 67022 67698 67204 67934
rect 66604 32254 67204 67698
rect 66604 32018 66786 32254
rect 67022 32018 67204 32254
rect 66604 31934 67204 32018
rect 66604 31698 66786 31934
rect 67022 31698 67204 31934
rect 48604 -6222 48786 -5986
rect 49022 -6222 49204 -5986
rect 48604 -6306 49204 -6222
rect 48604 -6542 48786 -6306
rect 49022 -6542 49204 -6306
rect 48604 -7504 49204 -6542
rect 66604 -6926 67204 31698
rect 73804 704838 74404 705800
rect 73804 704602 73986 704838
rect 74222 704602 74404 704838
rect 73804 704518 74404 704602
rect 73804 704282 73986 704518
rect 74222 704282 74404 704518
rect 73804 687454 74404 704282
rect 73804 687218 73986 687454
rect 74222 687218 74404 687454
rect 73804 687134 74404 687218
rect 73804 686898 73986 687134
rect 74222 686898 74404 687134
rect 73804 651454 74404 686898
rect 73804 651218 73986 651454
rect 74222 651218 74404 651454
rect 73804 651134 74404 651218
rect 73804 650898 73986 651134
rect 74222 650898 74404 651134
rect 73804 615454 74404 650898
rect 73804 615218 73986 615454
rect 74222 615218 74404 615454
rect 73804 615134 74404 615218
rect 73804 614898 73986 615134
rect 74222 614898 74404 615134
rect 73804 579454 74404 614898
rect 73804 579218 73986 579454
rect 74222 579218 74404 579454
rect 73804 579134 74404 579218
rect 73804 578898 73986 579134
rect 74222 578898 74404 579134
rect 73804 543454 74404 578898
rect 73804 543218 73986 543454
rect 74222 543218 74404 543454
rect 73804 543134 74404 543218
rect 73804 542898 73986 543134
rect 74222 542898 74404 543134
rect 73804 507454 74404 542898
rect 73804 507218 73986 507454
rect 74222 507218 74404 507454
rect 73804 507134 74404 507218
rect 73804 506898 73986 507134
rect 74222 506898 74404 507134
rect 73804 471454 74404 506898
rect 73804 471218 73986 471454
rect 74222 471218 74404 471454
rect 73804 471134 74404 471218
rect 73804 470898 73986 471134
rect 74222 470898 74404 471134
rect 73804 435454 74404 470898
rect 73804 435218 73986 435454
rect 74222 435218 74404 435454
rect 73804 435134 74404 435218
rect 73804 434898 73986 435134
rect 74222 434898 74404 435134
rect 73804 399454 74404 434898
rect 73804 399218 73986 399454
rect 74222 399218 74404 399454
rect 73804 399134 74404 399218
rect 73804 398898 73986 399134
rect 74222 398898 74404 399134
rect 73804 363454 74404 398898
rect 73804 363218 73986 363454
rect 74222 363218 74404 363454
rect 73804 363134 74404 363218
rect 73804 362898 73986 363134
rect 74222 362898 74404 363134
rect 73804 327454 74404 362898
rect 73804 327218 73986 327454
rect 74222 327218 74404 327454
rect 73804 327134 74404 327218
rect 73804 326898 73986 327134
rect 74222 326898 74404 327134
rect 73804 291454 74404 326898
rect 73804 291218 73986 291454
rect 74222 291218 74404 291454
rect 73804 291134 74404 291218
rect 73804 290898 73986 291134
rect 74222 290898 74404 291134
rect 73804 255454 74404 290898
rect 73804 255218 73986 255454
rect 74222 255218 74404 255454
rect 73804 255134 74404 255218
rect 73804 254898 73986 255134
rect 74222 254898 74404 255134
rect 73804 219454 74404 254898
rect 73804 219218 73986 219454
rect 74222 219218 74404 219454
rect 73804 219134 74404 219218
rect 73804 218898 73986 219134
rect 74222 218898 74404 219134
rect 73804 183454 74404 218898
rect 73804 183218 73986 183454
rect 74222 183218 74404 183454
rect 73804 183134 74404 183218
rect 73804 182898 73986 183134
rect 74222 182898 74404 183134
rect 73804 147454 74404 182898
rect 73804 147218 73986 147454
rect 74222 147218 74404 147454
rect 73804 147134 74404 147218
rect 73804 146898 73986 147134
rect 74222 146898 74404 147134
rect 73804 111454 74404 146898
rect 73804 111218 73986 111454
rect 74222 111218 74404 111454
rect 73804 111134 74404 111218
rect 73804 110898 73986 111134
rect 74222 110898 74404 111134
rect 73804 75454 74404 110898
rect 73804 75218 73986 75454
rect 74222 75218 74404 75454
rect 73804 75134 74404 75218
rect 73804 74898 73986 75134
rect 74222 74898 74404 75134
rect 73804 39454 74404 74898
rect 73804 39218 73986 39454
rect 74222 39218 74404 39454
rect 73804 39134 74404 39218
rect 73804 38898 73986 39134
rect 74222 38898 74404 39134
rect 73804 3454 74404 38898
rect 73804 3218 73986 3454
rect 74222 3218 74404 3454
rect 73804 3134 74404 3218
rect 73804 2898 73986 3134
rect 74222 2898 74404 3134
rect 73804 -346 74404 2898
rect 73804 -582 73986 -346
rect 74222 -582 74404 -346
rect 73804 -666 74404 -582
rect 73804 -902 73986 -666
rect 74222 -902 74404 -666
rect 73804 -1864 74404 -902
rect 77404 691054 78004 706162
rect 77404 690818 77586 691054
rect 77822 690818 78004 691054
rect 77404 690734 78004 690818
rect 77404 690498 77586 690734
rect 77822 690498 78004 690734
rect 77404 655054 78004 690498
rect 77404 654818 77586 655054
rect 77822 654818 78004 655054
rect 77404 654734 78004 654818
rect 77404 654498 77586 654734
rect 77822 654498 78004 654734
rect 77404 619054 78004 654498
rect 77404 618818 77586 619054
rect 77822 618818 78004 619054
rect 77404 618734 78004 618818
rect 77404 618498 77586 618734
rect 77822 618498 78004 618734
rect 77404 583054 78004 618498
rect 77404 582818 77586 583054
rect 77822 582818 78004 583054
rect 77404 582734 78004 582818
rect 77404 582498 77586 582734
rect 77822 582498 78004 582734
rect 77404 547054 78004 582498
rect 77404 546818 77586 547054
rect 77822 546818 78004 547054
rect 77404 546734 78004 546818
rect 77404 546498 77586 546734
rect 77822 546498 78004 546734
rect 77404 511054 78004 546498
rect 77404 510818 77586 511054
rect 77822 510818 78004 511054
rect 77404 510734 78004 510818
rect 77404 510498 77586 510734
rect 77822 510498 78004 510734
rect 77404 475054 78004 510498
rect 77404 474818 77586 475054
rect 77822 474818 78004 475054
rect 77404 474734 78004 474818
rect 77404 474498 77586 474734
rect 77822 474498 78004 474734
rect 77404 439054 78004 474498
rect 77404 438818 77586 439054
rect 77822 438818 78004 439054
rect 77404 438734 78004 438818
rect 77404 438498 77586 438734
rect 77822 438498 78004 438734
rect 77404 403054 78004 438498
rect 77404 402818 77586 403054
rect 77822 402818 78004 403054
rect 77404 402734 78004 402818
rect 77404 402498 77586 402734
rect 77822 402498 78004 402734
rect 77404 367054 78004 402498
rect 77404 366818 77586 367054
rect 77822 366818 78004 367054
rect 77404 366734 78004 366818
rect 77404 366498 77586 366734
rect 77822 366498 78004 366734
rect 77404 331054 78004 366498
rect 77404 330818 77586 331054
rect 77822 330818 78004 331054
rect 77404 330734 78004 330818
rect 77404 330498 77586 330734
rect 77822 330498 78004 330734
rect 77404 295054 78004 330498
rect 77404 294818 77586 295054
rect 77822 294818 78004 295054
rect 77404 294734 78004 294818
rect 77404 294498 77586 294734
rect 77822 294498 78004 294734
rect 77404 259054 78004 294498
rect 77404 258818 77586 259054
rect 77822 258818 78004 259054
rect 77404 258734 78004 258818
rect 77404 258498 77586 258734
rect 77822 258498 78004 258734
rect 77404 223054 78004 258498
rect 77404 222818 77586 223054
rect 77822 222818 78004 223054
rect 77404 222734 78004 222818
rect 77404 222498 77586 222734
rect 77822 222498 78004 222734
rect 77404 187054 78004 222498
rect 77404 186818 77586 187054
rect 77822 186818 78004 187054
rect 77404 186734 78004 186818
rect 77404 186498 77586 186734
rect 77822 186498 78004 186734
rect 77404 151054 78004 186498
rect 77404 150818 77586 151054
rect 77822 150818 78004 151054
rect 77404 150734 78004 150818
rect 77404 150498 77586 150734
rect 77822 150498 78004 150734
rect 77404 115054 78004 150498
rect 77404 114818 77586 115054
rect 77822 114818 78004 115054
rect 77404 114734 78004 114818
rect 77404 114498 77586 114734
rect 77822 114498 78004 114734
rect 77404 79054 78004 114498
rect 77404 78818 77586 79054
rect 77822 78818 78004 79054
rect 77404 78734 78004 78818
rect 77404 78498 77586 78734
rect 77822 78498 78004 78734
rect 77404 43054 78004 78498
rect 77404 42818 77586 43054
rect 77822 42818 78004 43054
rect 77404 42734 78004 42818
rect 77404 42498 77586 42734
rect 77822 42498 78004 42734
rect 77404 7054 78004 42498
rect 77404 6818 77586 7054
rect 77822 6818 78004 7054
rect 77404 6734 78004 6818
rect 77404 6498 77586 6734
rect 77822 6498 78004 6734
rect 77404 -2226 78004 6498
rect 77404 -2462 77586 -2226
rect 77822 -2462 78004 -2226
rect 77404 -2546 78004 -2462
rect 77404 -2782 77586 -2546
rect 77822 -2782 78004 -2546
rect 77404 -3744 78004 -2782
rect 81004 694654 81604 708042
rect 81004 694418 81186 694654
rect 81422 694418 81604 694654
rect 81004 694334 81604 694418
rect 81004 694098 81186 694334
rect 81422 694098 81604 694334
rect 81004 658654 81604 694098
rect 81004 658418 81186 658654
rect 81422 658418 81604 658654
rect 81004 658334 81604 658418
rect 81004 658098 81186 658334
rect 81422 658098 81604 658334
rect 81004 622654 81604 658098
rect 81004 622418 81186 622654
rect 81422 622418 81604 622654
rect 81004 622334 81604 622418
rect 81004 622098 81186 622334
rect 81422 622098 81604 622334
rect 81004 586654 81604 622098
rect 81004 586418 81186 586654
rect 81422 586418 81604 586654
rect 81004 586334 81604 586418
rect 81004 586098 81186 586334
rect 81422 586098 81604 586334
rect 81004 550654 81604 586098
rect 81004 550418 81186 550654
rect 81422 550418 81604 550654
rect 81004 550334 81604 550418
rect 81004 550098 81186 550334
rect 81422 550098 81604 550334
rect 81004 514654 81604 550098
rect 81004 514418 81186 514654
rect 81422 514418 81604 514654
rect 81004 514334 81604 514418
rect 81004 514098 81186 514334
rect 81422 514098 81604 514334
rect 81004 478654 81604 514098
rect 81004 478418 81186 478654
rect 81422 478418 81604 478654
rect 81004 478334 81604 478418
rect 81004 478098 81186 478334
rect 81422 478098 81604 478334
rect 81004 442654 81604 478098
rect 81004 442418 81186 442654
rect 81422 442418 81604 442654
rect 81004 442334 81604 442418
rect 81004 442098 81186 442334
rect 81422 442098 81604 442334
rect 81004 406654 81604 442098
rect 81004 406418 81186 406654
rect 81422 406418 81604 406654
rect 81004 406334 81604 406418
rect 81004 406098 81186 406334
rect 81422 406098 81604 406334
rect 81004 370654 81604 406098
rect 81004 370418 81186 370654
rect 81422 370418 81604 370654
rect 81004 370334 81604 370418
rect 81004 370098 81186 370334
rect 81422 370098 81604 370334
rect 81004 334654 81604 370098
rect 81004 334418 81186 334654
rect 81422 334418 81604 334654
rect 81004 334334 81604 334418
rect 81004 334098 81186 334334
rect 81422 334098 81604 334334
rect 81004 298654 81604 334098
rect 81004 298418 81186 298654
rect 81422 298418 81604 298654
rect 81004 298334 81604 298418
rect 81004 298098 81186 298334
rect 81422 298098 81604 298334
rect 81004 262654 81604 298098
rect 81004 262418 81186 262654
rect 81422 262418 81604 262654
rect 81004 262334 81604 262418
rect 81004 262098 81186 262334
rect 81422 262098 81604 262334
rect 81004 226654 81604 262098
rect 81004 226418 81186 226654
rect 81422 226418 81604 226654
rect 81004 226334 81604 226418
rect 81004 226098 81186 226334
rect 81422 226098 81604 226334
rect 81004 190654 81604 226098
rect 81004 190418 81186 190654
rect 81422 190418 81604 190654
rect 81004 190334 81604 190418
rect 81004 190098 81186 190334
rect 81422 190098 81604 190334
rect 81004 154654 81604 190098
rect 81004 154418 81186 154654
rect 81422 154418 81604 154654
rect 81004 154334 81604 154418
rect 81004 154098 81186 154334
rect 81422 154098 81604 154334
rect 81004 118654 81604 154098
rect 81004 118418 81186 118654
rect 81422 118418 81604 118654
rect 81004 118334 81604 118418
rect 81004 118098 81186 118334
rect 81422 118098 81604 118334
rect 81004 82654 81604 118098
rect 81004 82418 81186 82654
rect 81422 82418 81604 82654
rect 81004 82334 81604 82418
rect 81004 82098 81186 82334
rect 81422 82098 81604 82334
rect 81004 46654 81604 82098
rect 81004 46418 81186 46654
rect 81422 46418 81604 46654
rect 81004 46334 81604 46418
rect 81004 46098 81186 46334
rect 81422 46098 81604 46334
rect 81004 10654 81604 46098
rect 81004 10418 81186 10654
rect 81422 10418 81604 10654
rect 81004 10334 81604 10418
rect 81004 10098 81186 10334
rect 81422 10098 81604 10334
rect 81004 -4106 81604 10098
rect 81004 -4342 81186 -4106
rect 81422 -4342 81604 -4106
rect 81004 -4426 81604 -4342
rect 81004 -4662 81186 -4426
rect 81422 -4662 81604 -4426
rect 81004 -5624 81604 -4662
rect 84604 698254 85204 709922
rect 102604 711418 103204 711440
rect 102604 711182 102786 711418
rect 103022 711182 103204 711418
rect 102604 711098 103204 711182
rect 102604 710862 102786 711098
rect 103022 710862 103204 711098
rect 99004 709538 99604 709560
rect 99004 709302 99186 709538
rect 99422 709302 99604 709538
rect 99004 709218 99604 709302
rect 99004 708982 99186 709218
rect 99422 708982 99604 709218
rect 95404 707658 96004 707680
rect 95404 707422 95586 707658
rect 95822 707422 96004 707658
rect 95404 707338 96004 707422
rect 95404 707102 95586 707338
rect 95822 707102 96004 707338
rect 84604 698018 84786 698254
rect 85022 698018 85204 698254
rect 84604 697934 85204 698018
rect 84604 697698 84786 697934
rect 85022 697698 85204 697934
rect 84604 662254 85204 697698
rect 84604 662018 84786 662254
rect 85022 662018 85204 662254
rect 84604 661934 85204 662018
rect 84604 661698 84786 661934
rect 85022 661698 85204 661934
rect 84604 626254 85204 661698
rect 84604 626018 84786 626254
rect 85022 626018 85204 626254
rect 84604 625934 85204 626018
rect 84604 625698 84786 625934
rect 85022 625698 85204 625934
rect 84604 590254 85204 625698
rect 84604 590018 84786 590254
rect 85022 590018 85204 590254
rect 84604 589934 85204 590018
rect 84604 589698 84786 589934
rect 85022 589698 85204 589934
rect 84604 554254 85204 589698
rect 84604 554018 84786 554254
rect 85022 554018 85204 554254
rect 84604 553934 85204 554018
rect 84604 553698 84786 553934
rect 85022 553698 85204 553934
rect 84604 518254 85204 553698
rect 84604 518018 84786 518254
rect 85022 518018 85204 518254
rect 84604 517934 85204 518018
rect 84604 517698 84786 517934
rect 85022 517698 85204 517934
rect 84604 482254 85204 517698
rect 84604 482018 84786 482254
rect 85022 482018 85204 482254
rect 84604 481934 85204 482018
rect 84604 481698 84786 481934
rect 85022 481698 85204 481934
rect 84604 446254 85204 481698
rect 84604 446018 84786 446254
rect 85022 446018 85204 446254
rect 84604 445934 85204 446018
rect 84604 445698 84786 445934
rect 85022 445698 85204 445934
rect 84604 410254 85204 445698
rect 84604 410018 84786 410254
rect 85022 410018 85204 410254
rect 84604 409934 85204 410018
rect 84604 409698 84786 409934
rect 85022 409698 85204 409934
rect 84604 374254 85204 409698
rect 84604 374018 84786 374254
rect 85022 374018 85204 374254
rect 84604 373934 85204 374018
rect 84604 373698 84786 373934
rect 85022 373698 85204 373934
rect 84604 338254 85204 373698
rect 84604 338018 84786 338254
rect 85022 338018 85204 338254
rect 84604 337934 85204 338018
rect 84604 337698 84786 337934
rect 85022 337698 85204 337934
rect 84604 302254 85204 337698
rect 84604 302018 84786 302254
rect 85022 302018 85204 302254
rect 84604 301934 85204 302018
rect 84604 301698 84786 301934
rect 85022 301698 85204 301934
rect 84604 266254 85204 301698
rect 84604 266018 84786 266254
rect 85022 266018 85204 266254
rect 84604 265934 85204 266018
rect 84604 265698 84786 265934
rect 85022 265698 85204 265934
rect 84604 230254 85204 265698
rect 84604 230018 84786 230254
rect 85022 230018 85204 230254
rect 84604 229934 85204 230018
rect 84604 229698 84786 229934
rect 85022 229698 85204 229934
rect 84604 194254 85204 229698
rect 84604 194018 84786 194254
rect 85022 194018 85204 194254
rect 84604 193934 85204 194018
rect 84604 193698 84786 193934
rect 85022 193698 85204 193934
rect 84604 158254 85204 193698
rect 84604 158018 84786 158254
rect 85022 158018 85204 158254
rect 84604 157934 85204 158018
rect 84604 157698 84786 157934
rect 85022 157698 85204 157934
rect 84604 122254 85204 157698
rect 84604 122018 84786 122254
rect 85022 122018 85204 122254
rect 84604 121934 85204 122018
rect 84604 121698 84786 121934
rect 85022 121698 85204 121934
rect 84604 86254 85204 121698
rect 84604 86018 84786 86254
rect 85022 86018 85204 86254
rect 84604 85934 85204 86018
rect 84604 85698 84786 85934
rect 85022 85698 85204 85934
rect 84604 50254 85204 85698
rect 84604 50018 84786 50254
rect 85022 50018 85204 50254
rect 84604 49934 85204 50018
rect 84604 49698 84786 49934
rect 85022 49698 85204 49934
rect 84604 14254 85204 49698
rect 84604 14018 84786 14254
rect 85022 14018 85204 14254
rect 84604 13934 85204 14018
rect 84604 13698 84786 13934
rect 85022 13698 85204 13934
rect 66604 -7162 66786 -6926
rect 67022 -7162 67204 -6926
rect 66604 -7246 67204 -7162
rect 66604 -7482 66786 -7246
rect 67022 -7482 67204 -7246
rect 66604 -7504 67204 -7482
rect 84604 -5986 85204 13698
rect 91804 705778 92404 705800
rect 91804 705542 91986 705778
rect 92222 705542 92404 705778
rect 91804 705458 92404 705542
rect 91804 705222 91986 705458
rect 92222 705222 92404 705458
rect 91804 669454 92404 705222
rect 91804 669218 91986 669454
rect 92222 669218 92404 669454
rect 91804 669134 92404 669218
rect 91804 668898 91986 669134
rect 92222 668898 92404 669134
rect 91804 633454 92404 668898
rect 91804 633218 91986 633454
rect 92222 633218 92404 633454
rect 91804 633134 92404 633218
rect 91804 632898 91986 633134
rect 92222 632898 92404 633134
rect 91804 597454 92404 632898
rect 91804 597218 91986 597454
rect 92222 597218 92404 597454
rect 91804 597134 92404 597218
rect 91804 596898 91986 597134
rect 92222 596898 92404 597134
rect 91804 561454 92404 596898
rect 91804 561218 91986 561454
rect 92222 561218 92404 561454
rect 91804 561134 92404 561218
rect 91804 560898 91986 561134
rect 92222 560898 92404 561134
rect 91804 525454 92404 560898
rect 91804 525218 91986 525454
rect 92222 525218 92404 525454
rect 91804 525134 92404 525218
rect 91804 524898 91986 525134
rect 92222 524898 92404 525134
rect 91804 489454 92404 524898
rect 91804 489218 91986 489454
rect 92222 489218 92404 489454
rect 91804 489134 92404 489218
rect 91804 488898 91986 489134
rect 92222 488898 92404 489134
rect 91804 453454 92404 488898
rect 91804 453218 91986 453454
rect 92222 453218 92404 453454
rect 91804 453134 92404 453218
rect 91804 452898 91986 453134
rect 92222 452898 92404 453134
rect 91804 417454 92404 452898
rect 91804 417218 91986 417454
rect 92222 417218 92404 417454
rect 91804 417134 92404 417218
rect 91804 416898 91986 417134
rect 92222 416898 92404 417134
rect 91804 381454 92404 416898
rect 91804 381218 91986 381454
rect 92222 381218 92404 381454
rect 91804 381134 92404 381218
rect 91804 380898 91986 381134
rect 92222 380898 92404 381134
rect 91804 345454 92404 380898
rect 91804 345218 91986 345454
rect 92222 345218 92404 345454
rect 91804 345134 92404 345218
rect 91804 344898 91986 345134
rect 92222 344898 92404 345134
rect 91804 309454 92404 344898
rect 91804 309218 91986 309454
rect 92222 309218 92404 309454
rect 91804 309134 92404 309218
rect 91804 308898 91986 309134
rect 92222 308898 92404 309134
rect 91804 273454 92404 308898
rect 91804 273218 91986 273454
rect 92222 273218 92404 273454
rect 91804 273134 92404 273218
rect 91804 272898 91986 273134
rect 92222 272898 92404 273134
rect 91804 237454 92404 272898
rect 91804 237218 91986 237454
rect 92222 237218 92404 237454
rect 91804 237134 92404 237218
rect 91804 236898 91986 237134
rect 92222 236898 92404 237134
rect 91804 201454 92404 236898
rect 91804 201218 91986 201454
rect 92222 201218 92404 201454
rect 91804 201134 92404 201218
rect 91804 200898 91986 201134
rect 92222 200898 92404 201134
rect 91804 165454 92404 200898
rect 91804 165218 91986 165454
rect 92222 165218 92404 165454
rect 91804 165134 92404 165218
rect 91804 164898 91986 165134
rect 92222 164898 92404 165134
rect 91804 129454 92404 164898
rect 91804 129218 91986 129454
rect 92222 129218 92404 129454
rect 91804 129134 92404 129218
rect 91804 128898 91986 129134
rect 92222 128898 92404 129134
rect 91804 93454 92404 128898
rect 91804 93218 91986 93454
rect 92222 93218 92404 93454
rect 91804 93134 92404 93218
rect 91804 92898 91986 93134
rect 92222 92898 92404 93134
rect 91804 57454 92404 92898
rect 91804 57218 91986 57454
rect 92222 57218 92404 57454
rect 91804 57134 92404 57218
rect 91804 56898 91986 57134
rect 92222 56898 92404 57134
rect 91804 21454 92404 56898
rect 91804 21218 91986 21454
rect 92222 21218 92404 21454
rect 91804 21134 92404 21218
rect 91804 20898 91986 21134
rect 92222 20898 92404 21134
rect 91804 -1286 92404 20898
rect 91804 -1522 91986 -1286
rect 92222 -1522 92404 -1286
rect 91804 -1606 92404 -1522
rect 91804 -1842 91986 -1606
rect 92222 -1842 92404 -1606
rect 91804 -1864 92404 -1842
rect 95404 673054 96004 707102
rect 95404 672818 95586 673054
rect 95822 672818 96004 673054
rect 95404 672734 96004 672818
rect 95404 672498 95586 672734
rect 95822 672498 96004 672734
rect 95404 637054 96004 672498
rect 95404 636818 95586 637054
rect 95822 636818 96004 637054
rect 95404 636734 96004 636818
rect 95404 636498 95586 636734
rect 95822 636498 96004 636734
rect 95404 601054 96004 636498
rect 95404 600818 95586 601054
rect 95822 600818 96004 601054
rect 95404 600734 96004 600818
rect 95404 600498 95586 600734
rect 95822 600498 96004 600734
rect 95404 565054 96004 600498
rect 95404 564818 95586 565054
rect 95822 564818 96004 565054
rect 95404 564734 96004 564818
rect 95404 564498 95586 564734
rect 95822 564498 96004 564734
rect 95404 529054 96004 564498
rect 95404 528818 95586 529054
rect 95822 528818 96004 529054
rect 95404 528734 96004 528818
rect 95404 528498 95586 528734
rect 95822 528498 96004 528734
rect 95404 493054 96004 528498
rect 95404 492818 95586 493054
rect 95822 492818 96004 493054
rect 95404 492734 96004 492818
rect 95404 492498 95586 492734
rect 95822 492498 96004 492734
rect 95404 457054 96004 492498
rect 95404 456818 95586 457054
rect 95822 456818 96004 457054
rect 95404 456734 96004 456818
rect 95404 456498 95586 456734
rect 95822 456498 96004 456734
rect 95404 421054 96004 456498
rect 95404 420818 95586 421054
rect 95822 420818 96004 421054
rect 95404 420734 96004 420818
rect 95404 420498 95586 420734
rect 95822 420498 96004 420734
rect 95404 385054 96004 420498
rect 95404 384818 95586 385054
rect 95822 384818 96004 385054
rect 95404 384734 96004 384818
rect 95404 384498 95586 384734
rect 95822 384498 96004 384734
rect 95404 349054 96004 384498
rect 95404 348818 95586 349054
rect 95822 348818 96004 349054
rect 95404 348734 96004 348818
rect 95404 348498 95586 348734
rect 95822 348498 96004 348734
rect 95404 313054 96004 348498
rect 95404 312818 95586 313054
rect 95822 312818 96004 313054
rect 95404 312734 96004 312818
rect 95404 312498 95586 312734
rect 95822 312498 96004 312734
rect 95404 277054 96004 312498
rect 95404 276818 95586 277054
rect 95822 276818 96004 277054
rect 95404 276734 96004 276818
rect 95404 276498 95586 276734
rect 95822 276498 96004 276734
rect 95404 241054 96004 276498
rect 95404 240818 95586 241054
rect 95822 240818 96004 241054
rect 95404 240734 96004 240818
rect 95404 240498 95586 240734
rect 95822 240498 96004 240734
rect 95404 205054 96004 240498
rect 95404 204818 95586 205054
rect 95822 204818 96004 205054
rect 95404 204734 96004 204818
rect 95404 204498 95586 204734
rect 95822 204498 96004 204734
rect 95404 169054 96004 204498
rect 95404 168818 95586 169054
rect 95822 168818 96004 169054
rect 95404 168734 96004 168818
rect 95404 168498 95586 168734
rect 95822 168498 96004 168734
rect 95404 133054 96004 168498
rect 95404 132818 95586 133054
rect 95822 132818 96004 133054
rect 95404 132734 96004 132818
rect 95404 132498 95586 132734
rect 95822 132498 96004 132734
rect 95404 97054 96004 132498
rect 95404 96818 95586 97054
rect 95822 96818 96004 97054
rect 95404 96734 96004 96818
rect 95404 96498 95586 96734
rect 95822 96498 96004 96734
rect 95404 61054 96004 96498
rect 95404 60818 95586 61054
rect 95822 60818 96004 61054
rect 95404 60734 96004 60818
rect 95404 60498 95586 60734
rect 95822 60498 96004 60734
rect 95404 25054 96004 60498
rect 95404 24818 95586 25054
rect 95822 24818 96004 25054
rect 95404 24734 96004 24818
rect 95404 24498 95586 24734
rect 95822 24498 96004 24734
rect 95404 -3166 96004 24498
rect 95404 -3402 95586 -3166
rect 95822 -3402 96004 -3166
rect 95404 -3486 96004 -3402
rect 95404 -3722 95586 -3486
rect 95822 -3722 96004 -3486
rect 95404 -3744 96004 -3722
rect 99004 676654 99604 708982
rect 99004 676418 99186 676654
rect 99422 676418 99604 676654
rect 99004 676334 99604 676418
rect 99004 676098 99186 676334
rect 99422 676098 99604 676334
rect 99004 640654 99604 676098
rect 99004 640418 99186 640654
rect 99422 640418 99604 640654
rect 99004 640334 99604 640418
rect 99004 640098 99186 640334
rect 99422 640098 99604 640334
rect 99004 604654 99604 640098
rect 99004 604418 99186 604654
rect 99422 604418 99604 604654
rect 99004 604334 99604 604418
rect 99004 604098 99186 604334
rect 99422 604098 99604 604334
rect 99004 568654 99604 604098
rect 99004 568418 99186 568654
rect 99422 568418 99604 568654
rect 99004 568334 99604 568418
rect 99004 568098 99186 568334
rect 99422 568098 99604 568334
rect 99004 532654 99604 568098
rect 99004 532418 99186 532654
rect 99422 532418 99604 532654
rect 99004 532334 99604 532418
rect 99004 532098 99186 532334
rect 99422 532098 99604 532334
rect 99004 496654 99604 532098
rect 99004 496418 99186 496654
rect 99422 496418 99604 496654
rect 99004 496334 99604 496418
rect 99004 496098 99186 496334
rect 99422 496098 99604 496334
rect 99004 460654 99604 496098
rect 99004 460418 99186 460654
rect 99422 460418 99604 460654
rect 99004 460334 99604 460418
rect 99004 460098 99186 460334
rect 99422 460098 99604 460334
rect 99004 424654 99604 460098
rect 99004 424418 99186 424654
rect 99422 424418 99604 424654
rect 99004 424334 99604 424418
rect 99004 424098 99186 424334
rect 99422 424098 99604 424334
rect 99004 388654 99604 424098
rect 99004 388418 99186 388654
rect 99422 388418 99604 388654
rect 99004 388334 99604 388418
rect 99004 388098 99186 388334
rect 99422 388098 99604 388334
rect 99004 352654 99604 388098
rect 99004 352418 99186 352654
rect 99422 352418 99604 352654
rect 99004 352334 99604 352418
rect 99004 352098 99186 352334
rect 99422 352098 99604 352334
rect 99004 316654 99604 352098
rect 99004 316418 99186 316654
rect 99422 316418 99604 316654
rect 99004 316334 99604 316418
rect 99004 316098 99186 316334
rect 99422 316098 99604 316334
rect 99004 280654 99604 316098
rect 99004 280418 99186 280654
rect 99422 280418 99604 280654
rect 99004 280334 99604 280418
rect 99004 280098 99186 280334
rect 99422 280098 99604 280334
rect 99004 244654 99604 280098
rect 99004 244418 99186 244654
rect 99422 244418 99604 244654
rect 99004 244334 99604 244418
rect 99004 244098 99186 244334
rect 99422 244098 99604 244334
rect 99004 208654 99604 244098
rect 99004 208418 99186 208654
rect 99422 208418 99604 208654
rect 99004 208334 99604 208418
rect 99004 208098 99186 208334
rect 99422 208098 99604 208334
rect 99004 172654 99604 208098
rect 99004 172418 99186 172654
rect 99422 172418 99604 172654
rect 99004 172334 99604 172418
rect 99004 172098 99186 172334
rect 99422 172098 99604 172334
rect 99004 136654 99604 172098
rect 99004 136418 99186 136654
rect 99422 136418 99604 136654
rect 99004 136334 99604 136418
rect 99004 136098 99186 136334
rect 99422 136098 99604 136334
rect 99004 100654 99604 136098
rect 99004 100418 99186 100654
rect 99422 100418 99604 100654
rect 99004 100334 99604 100418
rect 99004 100098 99186 100334
rect 99422 100098 99604 100334
rect 99004 64654 99604 100098
rect 99004 64418 99186 64654
rect 99422 64418 99604 64654
rect 99004 64334 99604 64418
rect 99004 64098 99186 64334
rect 99422 64098 99604 64334
rect 99004 28654 99604 64098
rect 99004 28418 99186 28654
rect 99422 28418 99604 28654
rect 99004 28334 99604 28418
rect 99004 28098 99186 28334
rect 99422 28098 99604 28334
rect 99004 -5046 99604 28098
rect 99004 -5282 99186 -5046
rect 99422 -5282 99604 -5046
rect 99004 -5366 99604 -5282
rect 99004 -5602 99186 -5366
rect 99422 -5602 99604 -5366
rect 99004 -5624 99604 -5602
rect 102604 680254 103204 710862
rect 120604 710478 121204 711440
rect 120604 710242 120786 710478
rect 121022 710242 121204 710478
rect 120604 710158 121204 710242
rect 120604 709922 120786 710158
rect 121022 709922 121204 710158
rect 117004 708598 117604 709560
rect 117004 708362 117186 708598
rect 117422 708362 117604 708598
rect 117004 708278 117604 708362
rect 117004 708042 117186 708278
rect 117422 708042 117604 708278
rect 113404 706718 114004 707680
rect 113404 706482 113586 706718
rect 113822 706482 114004 706718
rect 113404 706398 114004 706482
rect 113404 706162 113586 706398
rect 113822 706162 114004 706398
rect 102604 680018 102786 680254
rect 103022 680018 103204 680254
rect 102604 679934 103204 680018
rect 102604 679698 102786 679934
rect 103022 679698 103204 679934
rect 102604 644254 103204 679698
rect 102604 644018 102786 644254
rect 103022 644018 103204 644254
rect 102604 643934 103204 644018
rect 102604 643698 102786 643934
rect 103022 643698 103204 643934
rect 102604 608254 103204 643698
rect 102604 608018 102786 608254
rect 103022 608018 103204 608254
rect 102604 607934 103204 608018
rect 102604 607698 102786 607934
rect 103022 607698 103204 607934
rect 102604 572254 103204 607698
rect 109804 704838 110404 705800
rect 109804 704602 109986 704838
rect 110222 704602 110404 704838
rect 109804 704518 110404 704602
rect 109804 704282 109986 704518
rect 110222 704282 110404 704518
rect 109804 687454 110404 704282
rect 109804 687218 109986 687454
rect 110222 687218 110404 687454
rect 109804 687134 110404 687218
rect 109804 686898 109986 687134
rect 110222 686898 110404 687134
rect 109804 651454 110404 686898
rect 109804 651218 109986 651454
rect 110222 651218 110404 651454
rect 109804 651134 110404 651218
rect 109804 650898 109986 651134
rect 110222 650898 110404 651134
rect 109804 615454 110404 650898
rect 109804 615218 109986 615454
rect 110222 615218 110404 615454
rect 109804 615134 110404 615218
rect 109804 614898 109986 615134
rect 110222 614898 110404 615134
rect 109804 598000 110404 614898
rect 113404 691054 114004 706162
rect 113404 690818 113586 691054
rect 113822 690818 114004 691054
rect 113404 690734 114004 690818
rect 113404 690498 113586 690734
rect 113822 690498 114004 690734
rect 113404 655054 114004 690498
rect 113404 654818 113586 655054
rect 113822 654818 114004 655054
rect 113404 654734 114004 654818
rect 113404 654498 113586 654734
rect 113822 654498 114004 654734
rect 113404 619054 114004 654498
rect 113404 618818 113586 619054
rect 113822 618818 114004 619054
rect 113404 618734 114004 618818
rect 113404 618498 113586 618734
rect 113822 618498 114004 618734
rect 113404 598000 114004 618498
rect 117004 694654 117604 708042
rect 117004 694418 117186 694654
rect 117422 694418 117604 694654
rect 117004 694334 117604 694418
rect 117004 694098 117186 694334
rect 117422 694098 117604 694334
rect 117004 658654 117604 694098
rect 117004 658418 117186 658654
rect 117422 658418 117604 658654
rect 117004 658334 117604 658418
rect 117004 658098 117186 658334
rect 117422 658098 117604 658334
rect 117004 622654 117604 658098
rect 117004 622418 117186 622654
rect 117422 622418 117604 622654
rect 117004 622334 117604 622418
rect 117004 622098 117186 622334
rect 117422 622098 117604 622334
rect 117004 598000 117604 622098
rect 120604 698254 121204 709922
rect 138604 711418 139204 711440
rect 138604 711182 138786 711418
rect 139022 711182 139204 711418
rect 138604 711098 139204 711182
rect 138604 710862 138786 711098
rect 139022 710862 139204 711098
rect 135004 709538 135604 709560
rect 135004 709302 135186 709538
rect 135422 709302 135604 709538
rect 135004 709218 135604 709302
rect 135004 708982 135186 709218
rect 135422 708982 135604 709218
rect 131404 707658 132004 707680
rect 131404 707422 131586 707658
rect 131822 707422 132004 707658
rect 131404 707338 132004 707422
rect 131404 707102 131586 707338
rect 131822 707102 132004 707338
rect 120604 698018 120786 698254
rect 121022 698018 121204 698254
rect 120604 697934 121204 698018
rect 120604 697698 120786 697934
rect 121022 697698 121204 697934
rect 120604 662254 121204 697698
rect 120604 662018 120786 662254
rect 121022 662018 121204 662254
rect 120604 661934 121204 662018
rect 120604 661698 120786 661934
rect 121022 661698 121204 661934
rect 120604 626254 121204 661698
rect 120604 626018 120786 626254
rect 121022 626018 121204 626254
rect 120604 625934 121204 626018
rect 120604 625698 120786 625934
rect 121022 625698 121204 625934
rect 120604 598000 121204 625698
rect 127804 705778 128404 705800
rect 127804 705542 127986 705778
rect 128222 705542 128404 705778
rect 127804 705458 128404 705542
rect 127804 705222 127986 705458
rect 128222 705222 128404 705458
rect 127804 669454 128404 705222
rect 127804 669218 127986 669454
rect 128222 669218 128404 669454
rect 127804 669134 128404 669218
rect 127804 668898 127986 669134
rect 128222 668898 128404 669134
rect 127804 633454 128404 668898
rect 127804 633218 127986 633454
rect 128222 633218 128404 633454
rect 127804 633134 128404 633218
rect 127804 632898 127986 633134
rect 128222 632898 128404 633134
rect 127804 598000 128404 632898
rect 131404 673054 132004 707102
rect 131404 672818 131586 673054
rect 131822 672818 132004 673054
rect 131404 672734 132004 672818
rect 131404 672498 131586 672734
rect 131822 672498 132004 672734
rect 131404 637054 132004 672498
rect 131404 636818 131586 637054
rect 131822 636818 132004 637054
rect 131404 636734 132004 636818
rect 131404 636498 131586 636734
rect 131822 636498 132004 636734
rect 131404 601054 132004 636498
rect 131404 600818 131586 601054
rect 131822 600818 132004 601054
rect 131404 600734 132004 600818
rect 131404 600498 131586 600734
rect 131822 600498 132004 600734
rect 131404 598000 132004 600498
rect 135004 676654 135604 708982
rect 135004 676418 135186 676654
rect 135422 676418 135604 676654
rect 135004 676334 135604 676418
rect 135004 676098 135186 676334
rect 135422 676098 135604 676334
rect 135004 640654 135604 676098
rect 135004 640418 135186 640654
rect 135422 640418 135604 640654
rect 135004 640334 135604 640418
rect 135004 640098 135186 640334
rect 135422 640098 135604 640334
rect 135004 604654 135604 640098
rect 135004 604418 135186 604654
rect 135422 604418 135604 604654
rect 135004 604334 135604 604418
rect 135004 604098 135186 604334
rect 135422 604098 135604 604334
rect 135004 598000 135604 604098
rect 138604 680254 139204 710862
rect 156604 710478 157204 711440
rect 156604 710242 156786 710478
rect 157022 710242 157204 710478
rect 156604 710158 157204 710242
rect 156604 709922 156786 710158
rect 157022 709922 157204 710158
rect 153004 708598 153604 709560
rect 153004 708362 153186 708598
rect 153422 708362 153604 708598
rect 153004 708278 153604 708362
rect 153004 708042 153186 708278
rect 153422 708042 153604 708278
rect 149404 706718 150004 707680
rect 149404 706482 149586 706718
rect 149822 706482 150004 706718
rect 149404 706398 150004 706482
rect 149404 706162 149586 706398
rect 149822 706162 150004 706398
rect 138604 680018 138786 680254
rect 139022 680018 139204 680254
rect 138604 679934 139204 680018
rect 138604 679698 138786 679934
rect 139022 679698 139204 679934
rect 138604 644254 139204 679698
rect 138604 644018 138786 644254
rect 139022 644018 139204 644254
rect 138604 643934 139204 644018
rect 138604 643698 138786 643934
rect 139022 643698 139204 643934
rect 138604 608254 139204 643698
rect 138604 608018 138786 608254
rect 139022 608018 139204 608254
rect 138604 607934 139204 608018
rect 138604 607698 138786 607934
rect 139022 607698 139204 607934
rect 138604 598000 139204 607698
rect 145804 704838 146404 705800
rect 145804 704602 145986 704838
rect 146222 704602 146404 704838
rect 145804 704518 146404 704602
rect 145804 704282 145986 704518
rect 146222 704282 146404 704518
rect 145804 687454 146404 704282
rect 145804 687218 145986 687454
rect 146222 687218 146404 687454
rect 145804 687134 146404 687218
rect 145804 686898 145986 687134
rect 146222 686898 146404 687134
rect 145804 651454 146404 686898
rect 145804 651218 145986 651454
rect 146222 651218 146404 651454
rect 145804 651134 146404 651218
rect 145804 650898 145986 651134
rect 146222 650898 146404 651134
rect 145804 615454 146404 650898
rect 145804 615218 145986 615454
rect 146222 615218 146404 615454
rect 145804 615134 146404 615218
rect 145804 614898 145986 615134
rect 146222 614898 146404 615134
rect 145804 598000 146404 614898
rect 149404 691054 150004 706162
rect 149404 690818 149586 691054
rect 149822 690818 150004 691054
rect 149404 690734 150004 690818
rect 149404 690498 149586 690734
rect 149822 690498 150004 690734
rect 149404 655054 150004 690498
rect 149404 654818 149586 655054
rect 149822 654818 150004 655054
rect 149404 654734 150004 654818
rect 149404 654498 149586 654734
rect 149822 654498 150004 654734
rect 149404 619054 150004 654498
rect 149404 618818 149586 619054
rect 149822 618818 150004 619054
rect 149404 618734 150004 618818
rect 149404 618498 149586 618734
rect 149822 618498 150004 618734
rect 149404 598000 150004 618498
rect 153004 694654 153604 708042
rect 153004 694418 153186 694654
rect 153422 694418 153604 694654
rect 153004 694334 153604 694418
rect 153004 694098 153186 694334
rect 153422 694098 153604 694334
rect 153004 658654 153604 694098
rect 153004 658418 153186 658654
rect 153422 658418 153604 658654
rect 153004 658334 153604 658418
rect 153004 658098 153186 658334
rect 153422 658098 153604 658334
rect 153004 622654 153604 658098
rect 153004 622418 153186 622654
rect 153422 622418 153604 622654
rect 153004 622334 153604 622418
rect 153004 622098 153186 622334
rect 153422 622098 153604 622334
rect 153004 598000 153604 622098
rect 156604 698254 157204 709922
rect 174604 711418 175204 711440
rect 174604 711182 174786 711418
rect 175022 711182 175204 711418
rect 174604 711098 175204 711182
rect 174604 710862 174786 711098
rect 175022 710862 175204 711098
rect 171004 709538 171604 709560
rect 171004 709302 171186 709538
rect 171422 709302 171604 709538
rect 171004 709218 171604 709302
rect 171004 708982 171186 709218
rect 171422 708982 171604 709218
rect 167404 707658 168004 707680
rect 167404 707422 167586 707658
rect 167822 707422 168004 707658
rect 167404 707338 168004 707422
rect 167404 707102 167586 707338
rect 167822 707102 168004 707338
rect 156604 698018 156786 698254
rect 157022 698018 157204 698254
rect 156604 697934 157204 698018
rect 156604 697698 156786 697934
rect 157022 697698 157204 697934
rect 156604 662254 157204 697698
rect 156604 662018 156786 662254
rect 157022 662018 157204 662254
rect 156604 661934 157204 662018
rect 156604 661698 156786 661934
rect 157022 661698 157204 661934
rect 156604 626254 157204 661698
rect 156604 626018 156786 626254
rect 157022 626018 157204 626254
rect 156604 625934 157204 626018
rect 156604 625698 156786 625934
rect 157022 625698 157204 625934
rect 156604 598000 157204 625698
rect 163804 705778 164404 705800
rect 163804 705542 163986 705778
rect 164222 705542 164404 705778
rect 163804 705458 164404 705542
rect 163804 705222 163986 705458
rect 164222 705222 164404 705458
rect 163804 669454 164404 705222
rect 163804 669218 163986 669454
rect 164222 669218 164404 669454
rect 163804 669134 164404 669218
rect 163804 668898 163986 669134
rect 164222 668898 164404 669134
rect 163804 633454 164404 668898
rect 163804 633218 163986 633454
rect 164222 633218 164404 633454
rect 163804 633134 164404 633218
rect 163804 632898 163986 633134
rect 164222 632898 164404 633134
rect 163804 598000 164404 632898
rect 167404 673054 168004 707102
rect 167404 672818 167586 673054
rect 167822 672818 168004 673054
rect 167404 672734 168004 672818
rect 167404 672498 167586 672734
rect 167822 672498 168004 672734
rect 167404 637054 168004 672498
rect 167404 636818 167586 637054
rect 167822 636818 168004 637054
rect 167404 636734 168004 636818
rect 167404 636498 167586 636734
rect 167822 636498 168004 636734
rect 167404 601054 168004 636498
rect 167404 600818 167586 601054
rect 167822 600818 168004 601054
rect 167404 600734 168004 600818
rect 167404 600498 167586 600734
rect 167822 600498 168004 600734
rect 167404 598000 168004 600498
rect 171004 676654 171604 708982
rect 171004 676418 171186 676654
rect 171422 676418 171604 676654
rect 171004 676334 171604 676418
rect 171004 676098 171186 676334
rect 171422 676098 171604 676334
rect 171004 640654 171604 676098
rect 171004 640418 171186 640654
rect 171422 640418 171604 640654
rect 171004 640334 171604 640418
rect 171004 640098 171186 640334
rect 171422 640098 171604 640334
rect 171004 604654 171604 640098
rect 171004 604418 171186 604654
rect 171422 604418 171604 604654
rect 171004 604334 171604 604418
rect 171004 604098 171186 604334
rect 171422 604098 171604 604334
rect 171004 598000 171604 604098
rect 174604 680254 175204 710862
rect 192604 710478 193204 711440
rect 192604 710242 192786 710478
rect 193022 710242 193204 710478
rect 192604 710158 193204 710242
rect 192604 709922 192786 710158
rect 193022 709922 193204 710158
rect 189004 708598 189604 709560
rect 189004 708362 189186 708598
rect 189422 708362 189604 708598
rect 189004 708278 189604 708362
rect 189004 708042 189186 708278
rect 189422 708042 189604 708278
rect 185404 706718 186004 707680
rect 185404 706482 185586 706718
rect 185822 706482 186004 706718
rect 185404 706398 186004 706482
rect 185404 706162 185586 706398
rect 185822 706162 186004 706398
rect 174604 680018 174786 680254
rect 175022 680018 175204 680254
rect 174604 679934 175204 680018
rect 174604 679698 174786 679934
rect 175022 679698 175204 679934
rect 174604 644254 175204 679698
rect 174604 644018 174786 644254
rect 175022 644018 175204 644254
rect 174604 643934 175204 644018
rect 174604 643698 174786 643934
rect 175022 643698 175204 643934
rect 174604 608254 175204 643698
rect 174604 608018 174786 608254
rect 175022 608018 175204 608254
rect 174604 607934 175204 608018
rect 174604 607698 174786 607934
rect 175022 607698 175204 607934
rect 174604 598000 175204 607698
rect 181804 704838 182404 705800
rect 181804 704602 181986 704838
rect 182222 704602 182404 704838
rect 181804 704518 182404 704602
rect 181804 704282 181986 704518
rect 182222 704282 182404 704518
rect 181804 687454 182404 704282
rect 181804 687218 181986 687454
rect 182222 687218 182404 687454
rect 181804 687134 182404 687218
rect 181804 686898 181986 687134
rect 182222 686898 182404 687134
rect 181804 651454 182404 686898
rect 181804 651218 181986 651454
rect 182222 651218 182404 651454
rect 181804 651134 182404 651218
rect 181804 650898 181986 651134
rect 182222 650898 182404 651134
rect 181804 615454 182404 650898
rect 181804 615218 181986 615454
rect 182222 615218 182404 615454
rect 181804 615134 182404 615218
rect 181804 614898 181986 615134
rect 182222 614898 182404 615134
rect 181804 598000 182404 614898
rect 185404 691054 186004 706162
rect 185404 690818 185586 691054
rect 185822 690818 186004 691054
rect 185404 690734 186004 690818
rect 185404 690498 185586 690734
rect 185822 690498 186004 690734
rect 185404 655054 186004 690498
rect 185404 654818 185586 655054
rect 185822 654818 186004 655054
rect 185404 654734 186004 654818
rect 185404 654498 185586 654734
rect 185822 654498 186004 654734
rect 185404 619054 186004 654498
rect 185404 618818 185586 619054
rect 185822 618818 186004 619054
rect 185404 618734 186004 618818
rect 185404 618498 185586 618734
rect 185822 618498 186004 618734
rect 185404 598000 186004 618498
rect 189004 694654 189604 708042
rect 189004 694418 189186 694654
rect 189422 694418 189604 694654
rect 189004 694334 189604 694418
rect 189004 694098 189186 694334
rect 189422 694098 189604 694334
rect 189004 658654 189604 694098
rect 189004 658418 189186 658654
rect 189422 658418 189604 658654
rect 189004 658334 189604 658418
rect 189004 658098 189186 658334
rect 189422 658098 189604 658334
rect 189004 622654 189604 658098
rect 189004 622418 189186 622654
rect 189422 622418 189604 622654
rect 189004 622334 189604 622418
rect 189004 622098 189186 622334
rect 189422 622098 189604 622334
rect 189004 598000 189604 622098
rect 192604 698254 193204 709922
rect 210604 711418 211204 711440
rect 210604 711182 210786 711418
rect 211022 711182 211204 711418
rect 210604 711098 211204 711182
rect 210604 710862 210786 711098
rect 211022 710862 211204 711098
rect 207004 709538 207604 709560
rect 207004 709302 207186 709538
rect 207422 709302 207604 709538
rect 207004 709218 207604 709302
rect 207004 708982 207186 709218
rect 207422 708982 207604 709218
rect 203404 707658 204004 707680
rect 203404 707422 203586 707658
rect 203822 707422 204004 707658
rect 203404 707338 204004 707422
rect 203404 707102 203586 707338
rect 203822 707102 204004 707338
rect 192604 698018 192786 698254
rect 193022 698018 193204 698254
rect 192604 697934 193204 698018
rect 192604 697698 192786 697934
rect 193022 697698 193204 697934
rect 192604 662254 193204 697698
rect 192604 662018 192786 662254
rect 193022 662018 193204 662254
rect 192604 661934 193204 662018
rect 192604 661698 192786 661934
rect 193022 661698 193204 661934
rect 192604 626254 193204 661698
rect 192604 626018 192786 626254
rect 193022 626018 193204 626254
rect 192604 625934 193204 626018
rect 192604 625698 192786 625934
rect 193022 625698 193204 625934
rect 192604 598000 193204 625698
rect 199804 705778 200404 705800
rect 199804 705542 199986 705778
rect 200222 705542 200404 705778
rect 199804 705458 200404 705542
rect 199804 705222 199986 705458
rect 200222 705222 200404 705458
rect 199804 669454 200404 705222
rect 199804 669218 199986 669454
rect 200222 669218 200404 669454
rect 199804 669134 200404 669218
rect 199804 668898 199986 669134
rect 200222 668898 200404 669134
rect 199804 633454 200404 668898
rect 199804 633218 199986 633454
rect 200222 633218 200404 633454
rect 199804 633134 200404 633218
rect 199804 632898 199986 633134
rect 200222 632898 200404 633134
rect 199804 598000 200404 632898
rect 203404 673054 204004 707102
rect 203404 672818 203586 673054
rect 203822 672818 204004 673054
rect 203404 672734 204004 672818
rect 203404 672498 203586 672734
rect 203822 672498 204004 672734
rect 203404 637054 204004 672498
rect 203404 636818 203586 637054
rect 203822 636818 204004 637054
rect 203404 636734 204004 636818
rect 203404 636498 203586 636734
rect 203822 636498 204004 636734
rect 203404 601054 204004 636498
rect 203404 600818 203586 601054
rect 203822 600818 204004 601054
rect 203404 600734 204004 600818
rect 203404 600498 203586 600734
rect 203822 600498 204004 600734
rect 203404 598000 204004 600498
rect 207004 676654 207604 708982
rect 207004 676418 207186 676654
rect 207422 676418 207604 676654
rect 207004 676334 207604 676418
rect 207004 676098 207186 676334
rect 207422 676098 207604 676334
rect 207004 640654 207604 676098
rect 207004 640418 207186 640654
rect 207422 640418 207604 640654
rect 207004 640334 207604 640418
rect 207004 640098 207186 640334
rect 207422 640098 207604 640334
rect 207004 604654 207604 640098
rect 207004 604418 207186 604654
rect 207422 604418 207604 604654
rect 207004 604334 207604 604418
rect 207004 604098 207186 604334
rect 207422 604098 207604 604334
rect 207004 598000 207604 604098
rect 210604 680254 211204 710862
rect 228604 710478 229204 711440
rect 228604 710242 228786 710478
rect 229022 710242 229204 710478
rect 228604 710158 229204 710242
rect 228604 709922 228786 710158
rect 229022 709922 229204 710158
rect 225004 708598 225604 709560
rect 225004 708362 225186 708598
rect 225422 708362 225604 708598
rect 225004 708278 225604 708362
rect 225004 708042 225186 708278
rect 225422 708042 225604 708278
rect 221404 706718 222004 707680
rect 221404 706482 221586 706718
rect 221822 706482 222004 706718
rect 221404 706398 222004 706482
rect 221404 706162 221586 706398
rect 221822 706162 222004 706398
rect 210604 680018 210786 680254
rect 211022 680018 211204 680254
rect 210604 679934 211204 680018
rect 210604 679698 210786 679934
rect 211022 679698 211204 679934
rect 210604 644254 211204 679698
rect 210604 644018 210786 644254
rect 211022 644018 211204 644254
rect 210604 643934 211204 644018
rect 210604 643698 210786 643934
rect 211022 643698 211204 643934
rect 210604 608254 211204 643698
rect 210604 608018 210786 608254
rect 211022 608018 211204 608254
rect 210604 607934 211204 608018
rect 210604 607698 210786 607934
rect 211022 607698 211204 607934
rect 210604 598000 211204 607698
rect 217804 704838 218404 705800
rect 217804 704602 217986 704838
rect 218222 704602 218404 704838
rect 217804 704518 218404 704602
rect 217804 704282 217986 704518
rect 218222 704282 218404 704518
rect 217804 687454 218404 704282
rect 217804 687218 217986 687454
rect 218222 687218 218404 687454
rect 217804 687134 218404 687218
rect 217804 686898 217986 687134
rect 218222 686898 218404 687134
rect 217804 651454 218404 686898
rect 217804 651218 217986 651454
rect 218222 651218 218404 651454
rect 217804 651134 218404 651218
rect 217804 650898 217986 651134
rect 218222 650898 218404 651134
rect 217804 615454 218404 650898
rect 217804 615218 217986 615454
rect 218222 615218 218404 615454
rect 217804 615134 218404 615218
rect 217804 614898 217986 615134
rect 218222 614898 218404 615134
rect 217804 598000 218404 614898
rect 221404 691054 222004 706162
rect 221404 690818 221586 691054
rect 221822 690818 222004 691054
rect 221404 690734 222004 690818
rect 221404 690498 221586 690734
rect 221822 690498 222004 690734
rect 221404 655054 222004 690498
rect 221404 654818 221586 655054
rect 221822 654818 222004 655054
rect 221404 654734 222004 654818
rect 221404 654498 221586 654734
rect 221822 654498 222004 654734
rect 221404 619054 222004 654498
rect 221404 618818 221586 619054
rect 221822 618818 222004 619054
rect 221404 618734 222004 618818
rect 221404 618498 221586 618734
rect 221822 618498 222004 618734
rect 221404 598000 222004 618498
rect 225004 694654 225604 708042
rect 225004 694418 225186 694654
rect 225422 694418 225604 694654
rect 225004 694334 225604 694418
rect 225004 694098 225186 694334
rect 225422 694098 225604 694334
rect 225004 658654 225604 694098
rect 225004 658418 225186 658654
rect 225422 658418 225604 658654
rect 225004 658334 225604 658418
rect 225004 658098 225186 658334
rect 225422 658098 225604 658334
rect 225004 622654 225604 658098
rect 225004 622418 225186 622654
rect 225422 622418 225604 622654
rect 225004 622334 225604 622418
rect 225004 622098 225186 622334
rect 225422 622098 225604 622334
rect 225004 598000 225604 622098
rect 228604 698254 229204 709922
rect 246604 711418 247204 711440
rect 246604 711182 246786 711418
rect 247022 711182 247204 711418
rect 246604 711098 247204 711182
rect 246604 710862 246786 711098
rect 247022 710862 247204 711098
rect 243004 709538 243604 709560
rect 243004 709302 243186 709538
rect 243422 709302 243604 709538
rect 243004 709218 243604 709302
rect 243004 708982 243186 709218
rect 243422 708982 243604 709218
rect 239404 707658 240004 707680
rect 239404 707422 239586 707658
rect 239822 707422 240004 707658
rect 239404 707338 240004 707422
rect 239404 707102 239586 707338
rect 239822 707102 240004 707338
rect 228604 698018 228786 698254
rect 229022 698018 229204 698254
rect 228604 697934 229204 698018
rect 228604 697698 228786 697934
rect 229022 697698 229204 697934
rect 228604 662254 229204 697698
rect 228604 662018 228786 662254
rect 229022 662018 229204 662254
rect 228604 661934 229204 662018
rect 228604 661698 228786 661934
rect 229022 661698 229204 661934
rect 228604 626254 229204 661698
rect 228604 626018 228786 626254
rect 229022 626018 229204 626254
rect 228604 625934 229204 626018
rect 228604 625698 228786 625934
rect 229022 625698 229204 625934
rect 228604 598000 229204 625698
rect 235804 705778 236404 705800
rect 235804 705542 235986 705778
rect 236222 705542 236404 705778
rect 235804 705458 236404 705542
rect 235804 705222 235986 705458
rect 236222 705222 236404 705458
rect 235804 669454 236404 705222
rect 235804 669218 235986 669454
rect 236222 669218 236404 669454
rect 235804 669134 236404 669218
rect 235804 668898 235986 669134
rect 236222 668898 236404 669134
rect 235804 633454 236404 668898
rect 235804 633218 235986 633454
rect 236222 633218 236404 633454
rect 235804 633134 236404 633218
rect 235804 632898 235986 633134
rect 236222 632898 236404 633134
rect 235804 598000 236404 632898
rect 239404 673054 240004 707102
rect 239404 672818 239586 673054
rect 239822 672818 240004 673054
rect 239404 672734 240004 672818
rect 239404 672498 239586 672734
rect 239822 672498 240004 672734
rect 239404 637054 240004 672498
rect 239404 636818 239586 637054
rect 239822 636818 240004 637054
rect 239404 636734 240004 636818
rect 239404 636498 239586 636734
rect 239822 636498 240004 636734
rect 239404 601054 240004 636498
rect 239404 600818 239586 601054
rect 239822 600818 240004 601054
rect 239404 600734 240004 600818
rect 239404 600498 239586 600734
rect 239822 600498 240004 600734
rect 239404 598000 240004 600498
rect 243004 676654 243604 708982
rect 243004 676418 243186 676654
rect 243422 676418 243604 676654
rect 243004 676334 243604 676418
rect 243004 676098 243186 676334
rect 243422 676098 243604 676334
rect 243004 640654 243604 676098
rect 243004 640418 243186 640654
rect 243422 640418 243604 640654
rect 243004 640334 243604 640418
rect 243004 640098 243186 640334
rect 243422 640098 243604 640334
rect 243004 604654 243604 640098
rect 243004 604418 243186 604654
rect 243422 604418 243604 604654
rect 243004 604334 243604 604418
rect 243004 604098 243186 604334
rect 243422 604098 243604 604334
rect 243004 598000 243604 604098
rect 246604 680254 247204 710862
rect 264604 710478 265204 711440
rect 264604 710242 264786 710478
rect 265022 710242 265204 710478
rect 264604 710158 265204 710242
rect 264604 709922 264786 710158
rect 265022 709922 265204 710158
rect 261004 708598 261604 709560
rect 261004 708362 261186 708598
rect 261422 708362 261604 708598
rect 261004 708278 261604 708362
rect 261004 708042 261186 708278
rect 261422 708042 261604 708278
rect 257404 706718 258004 707680
rect 257404 706482 257586 706718
rect 257822 706482 258004 706718
rect 257404 706398 258004 706482
rect 257404 706162 257586 706398
rect 257822 706162 258004 706398
rect 246604 680018 246786 680254
rect 247022 680018 247204 680254
rect 246604 679934 247204 680018
rect 246604 679698 246786 679934
rect 247022 679698 247204 679934
rect 246604 644254 247204 679698
rect 246604 644018 246786 644254
rect 247022 644018 247204 644254
rect 246604 643934 247204 644018
rect 246604 643698 246786 643934
rect 247022 643698 247204 643934
rect 246604 608254 247204 643698
rect 246604 608018 246786 608254
rect 247022 608018 247204 608254
rect 246604 607934 247204 608018
rect 246604 607698 246786 607934
rect 247022 607698 247204 607934
rect 246604 598000 247204 607698
rect 253804 704838 254404 705800
rect 253804 704602 253986 704838
rect 254222 704602 254404 704838
rect 253804 704518 254404 704602
rect 253804 704282 253986 704518
rect 254222 704282 254404 704518
rect 253804 687454 254404 704282
rect 253804 687218 253986 687454
rect 254222 687218 254404 687454
rect 253804 687134 254404 687218
rect 253804 686898 253986 687134
rect 254222 686898 254404 687134
rect 253804 651454 254404 686898
rect 253804 651218 253986 651454
rect 254222 651218 254404 651454
rect 253804 651134 254404 651218
rect 253804 650898 253986 651134
rect 254222 650898 254404 651134
rect 253804 615454 254404 650898
rect 253804 615218 253986 615454
rect 254222 615218 254404 615454
rect 253804 615134 254404 615218
rect 253804 614898 253986 615134
rect 254222 614898 254404 615134
rect 253804 598000 254404 614898
rect 257404 691054 258004 706162
rect 257404 690818 257586 691054
rect 257822 690818 258004 691054
rect 257404 690734 258004 690818
rect 257404 690498 257586 690734
rect 257822 690498 258004 690734
rect 257404 655054 258004 690498
rect 257404 654818 257586 655054
rect 257822 654818 258004 655054
rect 257404 654734 258004 654818
rect 257404 654498 257586 654734
rect 257822 654498 258004 654734
rect 257404 619054 258004 654498
rect 257404 618818 257586 619054
rect 257822 618818 258004 619054
rect 257404 618734 258004 618818
rect 257404 618498 257586 618734
rect 257822 618498 258004 618734
rect 257404 598000 258004 618498
rect 261004 694654 261604 708042
rect 261004 694418 261186 694654
rect 261422 694418 261604 694654
rect 261004 694334 261604 694418
rect 261004 694098 261186 694334
rect 261422 694098 261604 694334
rect 261004 658654 261604 694098
rect 261004 658418 261186 658654
rect 261422 658418 261604 658654
rect 261004 658334 261604 658418
rect 261004 658098 261186 658334
rect 261422 658098 261604 658334
rect 261004 622654 261604 658098
rect 261004 622418 261186 622654
rect 261422 622418 261604 622654
rect 261004 622334 261604 622418
rect 261004 622098 261186 622334
rect 261422 622098 261604 622334
rect 261004 598000 261604 622098
rect 264604 698254 265204 709922
rect 282604 711418 283204 711440
rect 282604 711182 282786 711418
rect 283022 711182 283204 711418
rect 282604 711098 283204 711182
rect 282604 710862 282786 711098
rect 283022 710862 283204 711098
rect 279004 709538 279604 709560
rect 279004 709302 279186 709538
rect 279422 709302 279604 709538
rect 279004 709218 279604 709302
rect 279004 708982 279186 709218
rect 279422 708982 279604 709218
rect 275404 707658 276004 707680
rect 275404 707422 275586 707658
rect 275822 707422 276004 707658
rect 275404 707338 276004 707422
rect 275404 707102 275586 707338
rect 275822 707102 276004 707338
rect 264604 698018 264786 698254
rect 265022 698018 265204 698254
rect 264604 697934 265204 698018
rect 264604 697698 264786 697934
rect 265022 697698 265204 697934
rect 264604 662254 265204 697698
rect 264604 662018 264786 662254
rect 265022 662018 265204 662254
rect 264604 661934 265204 662018
rect 264604 661698 264786 661934
rect 265022 661698 265204 661934
rect 264604 626254 265204 661698
rect 264604 626018 264786 626254
rect 265022 626018 265204 626254
rect 264604 625934 265204 626018
rect 264604 625698 264786 625934
rect 265022 625698 265204 625934
rect 264604 598000 265204 625698
rect 271804 705778 272404 705800
rect 271804 705542 271986 705778
rect 272222 705542 272404 705778
rect 271804 705458 272404 705542
rect 271804 705222 271986 705458
rect 272222 705222 272404 705458
rect 271804 669454 272404 705222
rect 271804 669218 271986 669454
rect 272222 669218 272404 669454
rect 271804 669134 272404 669218
rect 271804 668898 271986 669134
rect 272222 668898 272404 669134
rect 271804 633454 272404 668898
rect 271804 633218 271986 633454
rect 272222 633218 272404 633454
rect 271804 633134 272404 633218
rect 271804 632898 271986 633134
rect 272222 632898 272404 633134
rect 271804 598000 272404 632898
rect 275404 673054 276004 707102
rect 275404 672818 275586 673054
rect 275822 672818 276004 673054
rect 275404 672734 276004 672818
rect 275404 672498 275586 672734
rect 275822 672498 276004 672734
rect 275404 637054 276004 672498
rect 275404 636818 275586 637054
rect 275822 636818 276004 637054
rect 275404 636734 276004 636818
rect 275404 636498 275586 636734
rect 275822 636498 276004 636734
rect 275404 601054 276004 636498
rect 275404 600818 275586 601054
rect 275822 600818 276004 601054
rect 275404 600734 276004 600818
rect 275404 600498 275586 600734
rect 275822 600498 276004 600734
rect 275404 598000 276004 600498
rect 279004 676654 279604 708982
rect 279004 676418 279186 676654
rect 279422 676418 279604 676654
rect 279004 676334 279604 676418
rect 279004 676098 279186 676334
rect 279422 676098 279604 676334
rect 279004 640654 279604 676098
rect 279004 640418 279186 640654
rect 279422 640418 279604 640654
rect 279004 640334 279604 640418
rect 279004 640098 279186 640334
rect 279422 640098 279604 640334
rect 279004 604654 279604 640098
rect 279004 604418 279186 604654
rect 279422 604418 279604 604654
rect 279004 604334 279604 604418
rect 279004 604098 279186 604334
rect 279422 604098 279604 604334
rect 279004 598000 279604 604098
rect 282604 680254 283204 710862
rect 300604 710478 301204 711440
rect 300604 710242 300786 710478
rect 301022 710242 301204 710478
rect 300604 710158 301204 710242
rect 300604 709922 300786 710158
rect 301022 709922 301204 710158
rect 297004 708598 297604 709560
rect 297004 708362 297186 708598
rect 297422 708362 297604 708598
rect 297004 708278 297604 708362
rect 297004 708042 297186 708278
rect 297422 708042 297604 708278
rect 293404 706718 294004 707680
rect 293404 706482 293586 706718
rect 293822 706482 294004 706718
rect 293404 706398 294004 706482
rect 293404 706162 293586 706398
rect 293822 706162 294004 706398
rect 282604 680018 282786 680254
rect 283022 680018 283204 680254
rect 282604 679934 283204 680018
rect 282604 679698 282786 679934
rect 283022 679698 283204 679934
rect 282604 644254 283204 679698
rect 282604 644018 282786 644254
rect 283022 644018 283204 644254
rect 282604 643934 283204 644018
rect 282604 643698 282786 643934
rect 283022 643698 283204 643934
rect 282604 608254 283204 643698
rect 282604 608018 282786 608254
rect 283022 608018 283204 608254
rect 282604 607934 283204 608018
rect 282604 607698 282786 607934
rect 283022 607698 283204 607934
rect 282604 598000 283204 607698
rect 289804 704838 290404 705800
rect 289804 704602 289986 704838
rect 290222 704602 290404 704838
rect 289804 704518 290404 704602
rect 289804 704282 289986 704518
rect 290222 704282 290404 704518
rect 289804 687454 290404 704282
rect 289804 687218 289986 687454
rect 290222 687218 290404 687454
rect 289804 687134 290404 687218
rect 289804 686898 289986 687134
rect 290222 686898 290404 687134
rect 289804 651454 290404 686898
rect 289804 651218 289986 651454
rect 290222 651218 290404 651454
rect 289804 651134 290404 651218
rect 289804 650898 289986 651134
rect 290222 650898 290404 651134
rect 289804 615454 290404 650898
rect 289804 615218 289986 615454
rect 290222 615218 290404 615454
rect 289804 615134 290404 615218
rect 289804 614898 289986 615134
rect 290222 614898 290404 615134
rect 289804 598000 290404 614898
rect 293404 691054 294004 706162
rect 293404 690818 293586 691054
rect 293822 690818 294004 691054
rect 293404 690734 294004 690818
rect 293404 690498 293586 690734
rect 293822 690498 294004 690734
rect 293404 655054 294004 690498
rect 293404 654818 293586 655054
rect 293822 654818 294004 655054
rect 293404 654734 294004 654818
rect 293404 654498 293586 654734
rect 293822 654498 294004 654734
rect 293404 619054 294004 654498
rect 293404 618818 293586 619054
rect 293822 618818 294004 619054
rect 293404 618734 294004 618818
rect 293404 618498 293586 618734
rect 293822 618498 294004 618734
rect 293404 598000 294004 618498
rect 297004 694654 297604 708042
rect 297004 694418 297186 694654
rect 297422 694418 297604 694654
rect 297004 694334 297604 694418
rect 297004 694098 297186 694334
rect 297422 694098 297604 694334
rect 297004 658654 297604 694098
rect 297004 658418 297186 658654
rect 297422 658418 297604 658654
rect 297004 658334 297604 658418
rect 297004 658098 297186 658334
rect 297422 658098 297604 658334
rect 297004 622654 297604 658098
rect 297004 622418 297186 622654
rect 297422 622418 297604 622654
rect 297004 622334 297604 622418
rect 297004 622098 297186 622334
rect 297422 622098 297604 622334
rect 297004 598000 297604 622098
rect 300604 698254 301204 709922
rect 318604 711418 319204 711440
rect 318604 711182 318786 711418
rect 319022 711182 319204 711418
rect 318604 711098 319204 711182
rect 318604 710862 318786 711098
rect 319022 710862 319204 711098
rect 315004 709538 315604 709560
rect 315004 709302 315186 709538
rect 315422 709302 315604 709538
rect 315004 709218 315604 709302
rect 315004 708982 315186 709218
rect 315422 708982 315604 709218
rect 311404 707658 312004 707680
rect 311404 707422 311586 707658
rect 311822 707422 312004 707658
rect 311404 707338 312004 707422
rect 311404 707102 311586 707338
rect 311822 707102 312004 707338
rect 300604 698018 300786 698254
rect 301022 698018 301204 698254
rect 300604 697934 301204 698018
rect 300604 697698 300786 697934
rect 301022 697698 301204 697934
rect 300604 662254 301204 697698
rect 300604 662018 300786 662254
rect 301022 662018 301204 662254
rect 300604 661934 301204 662018
rect 300604 661698 300786 661934
rect 301022 661698 301204 661934
rect 300604 626254 301204 661698
rect 300604 626018 300786 626254
rect 301022 626018 301204 626254
rect 300604 625934 301204 626018
rect 300604 625698 300786 625934
rect 301022 625698 301204 625934
rect 300604 598000 301204 625698
rect 307804 705778 308404 705800
rect 307804 705542 307986 705778
rect 308222 705542 308404 705778
rect 307804 705458 308404 705542
rect 307804 705222 307986 705458
rect 308222 705222 308404 705458
rect 307804 669454 308404 705222
rect 307804 669218 307986 669454
rect 308222 669218 308404 669454
rect 307804 669134 308404 669218
rect 307804 668898 307986 669134
rect 308222 668898 308404 669134
rect 307804 633454 308404 668898
rect 307804 633218 307986 633454
rect 308222 633218 308404 633454
rect 307804 633134 308404 633218
rect 307804 632898 307986 633134
rect 308222 632898 308404 633134
rect 307804 598000 308404 632898
rect 311404 673054 312004 707102
rect 311404 672818 311586 673054
rect 311822 672818 312004 673054
rect 311404 672734 312004 672818
rect 311404 672498 311586 672734
rect 311822 672498 312004 672734
rect 311404 637054 312004 672498
rect 311404 636818 311586 637054
rect 311822 636818 312004 637054
rect 311404 636734 312004 636818
rect 311404 636498 311586 636734
rect 311822 636498 312004 636734
rect 311404 601054 312004 636498
rect 311404 600818 311586 601054
rect 311822 600818 312004 601054
rect 311404 600734 312004 600818
rect 311404 600498 311586 600734
rect 311822 600498 312004 600734
rect 311404 598000 312004 600498
rect 315004 676654 315604 708982
rect 315004 676418 315186 676654
rect 315422 676418 315604 676654
rect 315004 676334 315604 676418
rect 315004 676098 315186 676334
rect 315422 676098 315604 676334
rect 315004 640654 315604 676098
rect 315004 640418 315186 640654
rect 315422 640418 315604 640654
rect 315004 640334 315604 640418
rect 315004 640098 315186 640334
rect 315422 640098 315604 640334
rect 315004 604654 315604 640098
rect 315004 604418 315186 604654
rect 315422 604418 315604 604654
rect 315004 604334 315604 604418
rect 315004 604098 315186 604334
rect 315422 604098 315604 604334
rect 315004 598000 315604 604098
rect 318604 680254 319204 710862
rect 336604 710478 337204 711440
rect 336604 710242 336786 710478
rect 337022 710242 337204 710478
rect 336604 710158 337204 710242
rect 336604 709922 336786 710158
rect 337022 709922 337204 710158
rect 333004 708598 333604 709560
rect 333004 708362 333186 708598
rect 333422 708362 333604 708598
rect 333004 708278 333604 708362
rect 333004 708042 333186 708278
rect 333422 708042 333604 708278
rect 329404 706718 330004 707680
rect 329404 706482 329586 706718
rect 329822 706482 330004 706718
rect 329404 706398 330004 706482
rect 329404 706162 329586 706398
rect 329822 706162 330004 706398
rect 318604 680018 318786 680254
rect 319022 680018 319204 680254
rect 318604 679934 319204 680018
rect 318604 679698 318786 679934
rect 319022 679698 319204 679934
rect 318604 644254 319204 679698
rect 318604 644018 318786 644254
rect 319022 644018 319204 644254
rect 318604 643934 319204 644018
rect 318604 643698 318786 643934
rect 319022 643698 319204 643934
rect 318604 608254 319204 643698
rect 318604 608018 318786 608254
rect 319022 608018 319204 608254
rect 318604 607934 319204 608018
rect 318604 607698 318786 607934
rect 319022 607698 319204 607934
rect 318604 598000 319204 607698
rect 325804 704838 326404 705800
rect 325804 704602 325986 704838
rect 326222 704602 326404 704838
rect 325804 704518 326404 704602
rect 325804 704282 325986 704518
rect 326222 704282 326404 704518
rect 325804 687454 326404 704282
rect 325804 687218 325986 687454
rect 326222 687218 326404 687454
rect 325804 687134 326404 687218
rect 325804 686898 325986 687134
rect 326222 686898 326404 687134
rect 325804 651454 326404 686898
rect 325804 651218 325986 651454
rect 326222 651218 326404 651454
rect 325804 651134 326404 651218
rect 325804 650898 325986 651134
rect 326222 650898 326404 651134
rect 325804 615454 326404 650898
rect 325804 615218 325986 615454
rect 326222 615218 326404 615454
rect 325804 615134 326404 615218
rect 325804 614898 325986 615134
rect 326222 614898 326404 615134
rect 325804 598000 326404 614898
rect 329404 691054 330004 706162
rect 329404 690818 329586 691054
rect 329822 690818 330004 691054
rect 329404 690734 330004 690818
rect 329404 690498 329586 690734
rect 329822 690498 330004 690734
rect 329404 655054 330004 690498
rect 329404 654818 329586 655054
rect 329822 654818 330004 655054
rect 329404 654734 330004 654818
rect 329404 654498 329586 654734
rect 329822 654498 330004 654734
rect 329404 619054 330004 654498
rect 329404 618818 329586 619054
rect 329822 618818 330004 619054
rect 329404 618734 330004 618818
rect 329404 618498 329586 618734
rect 329822 618498 330004 618734
rect 329404 598000 330004 618498
rect 333004 694654 333604 708042
rect 333004 694418 333186 694654
rect 333422 694418 333604 694654
rect 333004 694334 333604 694418
rect 333004 694098 333186 694334
rect 333422 694098 333604 694334
rect 333004 658654 333604 694098
rect 333004 658418 333186 658654
rect 333422 658418 333604 658654
rect 333004 658334 333604 658418
rect 333004 658098 333186 658334
rect 333422 658098 333604 658334
rect 333004 622654 333604 658098
rect 333004 622418 333186 622654
rect 333422 622418 333604 622654
rect 333004 622334 333604 622418
rect 333004 622098 333186 622334
rect 333422 622098 333604 622334
rect 333004 598000 333604 622098
rect 336604 698254 337204 709922
rect 354604 711418 355204 711440
rect 354604 711182 354786 711418
rect 355022 711182 355204 711418
rect 354604 711098 355204 711182
rect 354604 710862 354786 711098
rect 355022 710862 355204 711098
rect 351004 709538 351604 709560
rect 351004 709302 351186 709538
rect 351422 709302 351604 709538
rect 351004 709218 351604 709302
rect 351004 708982 351186 709218
rect 351422 708982 351604 709218
rect 347404 707658 348004 707680
rect 347404 707422 347586 707658
rect 347822 707422 348004 707658
rect 347404 707338 348004 707422
rect 347404 707102 347586 707338
rect 347822 707102 348004 707338
rect 336604 698018 336786 698254
rect 337022 698018 337204 698254
rect 336604 697934 337204 698018
rect 336604 697698 336786 697934
rect 337022 697698 337204 697934
rect 336604 662254 337204 697698
rect 336604 662018 336786 662254
rect 337022 662018 337204 662254
rect 336604 661934 337204 662018
rect 336604 661698 336786 661934
rect 337022 661698 337204 661934
rect 336604 626254 337204 661698
rect 336604 626018 336786 626254
rect 337022 626018 337204 626254
rect 336604 625934 337204 626018
rect 336604 625698 336786 625934
rect 337022 625698 337204 625934
rect 336604 598000 337204 625698
rect 343804 705778 344404 705800
rect 343804 705542 343986 705778
rect 344222 705542 344404 705778
rect 343804 705458 344404 705542
rect 343804 705222 343986 705458
rect 344222 705222 344404 705458
rect 343804 669454 344404 705222
rect 343804 669218 343986 669454
rect 344222 669218 344404 669454
rect 343804 669134 344404 669218
rect 343804 668898 343986 669134
rect 344222 668898 344404 669134
rect 343804 633454 344404 668898
rect 343804 633218 343986 633454
rect 344222 633218 344404 633454
rect 343804 633134 344404 633218
rect 343804 632898 343986 633134
rect 344222 632898 344404 633134
rect 343804 598000 344404 632898
rect 347404 673054 348004 707102
rect 347404 672818 347586 673054
rect 347822 672818 348004 673054
rect 347404 672734 348004 672818
rect 347404 672498 347586 672734
rect 347822 672498 348004 672734
rect 347404 637054 348004 672498
rect 347404 636818 347586 637054
rect 347822 636818 348004 637054
rect 347404 636734 348004 636818
rect 347404 636498 347586 636734
rect 347822 636498 348004 636734
rect 347404 601054 348004 636498
rect 347404 600818 347586 601054
rect 347822 600818 348004 601054
rect 347404 600734 348004 600818
rect 347404 600498 347586 600734
rect 347822 600498 348004 600734
rect 347404 598000 348004 600498
rect 351004 676654 351604 708982
rect 351004 676418 351186 676654
rect 351422 676418 351604 676654
rect 351004 676334 351604 676418
rect 351004 676098 351186 676334
rect 351422 676098 351604 676334
rect 351004 640654 351604 676098
rect 351004 640418 351186 640654
rect 351422 640418 351604 640654
rect 351004 640334 351604 640418
rect 351004 640098 351186 640334
rect 351422 640098 351604 640334
rect 351004 604654 351604 640098
rect 351004 604418 351186 604654
rect 351422 604418 351604 604654
rect 351004 604334 351604 604418
rect 351004 604098 351186 604334
rect 351422 604098 351604 604334
rect 351004 598000 351604 604098
rect 354604 680254 355204 710862
rect 372604 710478 373204 711440
rect 372604 710242 372786 710478
rect 373022 710242 373204 710478
rect 372604 710158 373204 710242
rect 372604 709922 372786 710158
rect 373022 709922 373204 710158
rect 369004 708598 369604 709560
rect 369004 708362 369186 708598
rect 369422 708362 369604 708598
rect 369004 708278 369604 708362
rect 369004 708042 369186 708278
rect 369422 708042 369604 708278
rect 365404 706718 366004 707680
rect 365404 706482 365586 706718
rect 365822 706482 366004 706718
rect 365404 706398 366004 706482
rect 365404 706162 365586 706398
rect 365822 706162 366004 706398
rect 354604 680018 354786 680254
rect 355022 680018 355204 680254
rect 354604 679934 355204 680018
rect 354604 679698 354786 679934
rect 355022 679698 355204 679934
rect 354604 644254 355204 679698
rect 354604 644018 354786 644254
rect 355022 644018 355204 644254
rect 354604 643934 355204 644018
rect 354604 643698 354786 643934
rect 355022 643698 355204 643934
rect 354604 608254 355204 643698
rect 354604 608018 354786 608254
rect 355022 608018 355204 608254
rect 354604 607934 355204 608018
rect 354604 607698 354786 607934
rect 355022 607698 355204 607934
rect 354604 598000 355204 607698
rect 361804 704838 362404 705800
rect 361804 704602 361986 704838
rect 362222 704602 362404 704838
rect 361804 704518 362404 704602
rect 361804 704282 361986 704518
rect 362222 704282 362404 704518
rect 361804 687454 362404 704282
rect 361804 687218 361986 687454
rect 362222 687218 362404 687454
rect 361804 687134 362404 687218
rect 361804 686898 361986 687134
rect 362222 686898 362404 687134
rect 361804 651454 362404 686898
rect 361804 651218 361986 651454
rect 362222 651218 362404 651454
rect 361804 651134 362404 651218
rect 361804 650898 361986 651134
rect 362222 650898 362404 651134
rect 361804 615454 362404 650898
rect 361804 615218 361986 615454
rect 362222 615218 362404 615454
rect 361804 615134 362404 615218
rect 361804 614898 361986 615134
rect 362222 614898 362404 615134
rect 361804 598000 362404 614898
rect 365404 691054 366004 706162
rect 365404 690818 365586 691054
rect 365822 690818 366004 691054
rect 365404 690734 366004 690818
rect 365404 690498 365586 690734
rect 365822 690498 366004 690734
rect 365404 655054 366004 690498
rect 365404 654818 365586 655054
rect 365822 654818 366004 655054
rect 365404 654734 366004 654818
rect 365404 654498 365586 654734
rect 365822 654498 366004 654734
rect 365404 619054 366004 654498
rect 365404 618818 365586 619054
rect 365822 618818 366004 619054
rect 365404 618734 366004 618818
rect 365404 618498 365586 618734
rect 365822 618498 366004 618734
rect 365404 598000 366004 618498
rect 369004 694654 369604 708042
rect 369004 694418 369186 694654
rect 369422 694418 369604 694654
rect 369004 694334 369604 694418
rect 369004 694098 369186 694334
rect 369422 694098 369604 694334
rect 369004 658654 369604 694098
rect 369004 658418 369186 658654
rect 369422 658418 369604 658654
rect 369004 658334 369604 658418
rect 369004 658098 369186 658334
rect 369422 658098 369604 658334
rect 369004 622654 369604 658098
rect 369004 622418 369186 622654
rect 369422 622418 369604 622654
rect 369004 622334 369604 622418
rect 369004 622098 369186 622334
rect 369422 622098 369604 622334
rect 369004 598000 369604 622098
rect 372604 698254 373204 709922
rect 390604 711418 391204 711440
rect 390604 711182 390786 711418
rect 391022 711182 391204 711418
rect 390604 711098 391204 711182
rect 390604 710862 390786 711098
rect 391022 710862 391204 711098
rect 387004 709538 387604 709560
rect 387004 709302 387186 709538
rect 387422 709302 387604 709538
rect 387004 709218 387604 709302
rect 387004 708982 387186 709218
rect 387422 708982 387604 709218
rect 383404 707658 384004 707680
rect 383404 707422 383586 707658
rect 383822 707422 384004 707658
rect 383404 707338 384004 707422
rect 383404 707102 383586 707338
rect 383822 707102 384004 707338
rect 372604 698018 372786 698254
rect 373022 698018 373204 698254
rect 372604 697934 373204 698018
rect 372604 697698 372786 697934
rect 373022 697698 373204 697934
rect 372604 662254 373204 697698
rect 372604 662018 372786 662254
rect 373022 662018 373204 662254
rect 372604 661934 373204 662018
rect 372604 661698 372786 661934
rect 373022 661698 373204 661934
rect 372604 626254 373204 661698
rect 372604 626018 372786 626254
rect 373022 626018 373204 626254
rect 372604 625934 373204 626018
rect 372604 625698 372786 625934
rect 373022 625698 373204 625934
rect 372604 598000 373204 625698
rect 379804 705778 380404 705800
rect 379804 705542 379986 705778
rect 380222 705542 380404 705778
rect 379804 705458 380404 705542
rect 379804 705222 379986 705458
rect 380222 705222 380404 705458
rect 379804 669454 380404 705222
rect 379804 669218 379986 669454
rect 380222 669218 380404 669454
rect 379804 669134 380404 669218
rect 379804 668898 379986 669134
rect 380222 668898 380404 669134
rect 379804 633454 380404 668898
rect 379804 633218 379986 633454
rect 380222 633218 380404 633454
rect 379804 633134 380404 633218
rect 379804 632898 379986 633134
rect 380222 632898 380404 633134
rect 379804 598000 380404 632898
rect 383404 673054 384004 707102
rect 383404 672818 383586 673054
rect 383822 672818 384004 673054
rect 383404 672734 384004 672818
rect 383404 672498 383586 672734
rect 383822 672498 384004 672734
rect 383404 637054 384004 672498
rect 383404 636818 383586 637054
rect 383822 636818 384004 637054
rect 383404 636734 384004 636818
rect 383404 636498 383586 636734
rect 383822 636498 384004 636734
rect 383404 601054 384004 636498
rect 383404 600818 383586 601054
rect 383822 600818 384004 601054
rect 383404 600734 384004 600818
rect 383404 600498 383586 600734
rect 383822 600498 384004 600734
rect 383404 598000 384004 600498
rect 387004 676654 387604 708982
rect 387004 676418 387186 676654
rect 387422 676418 387604 676654
rect 387004 676334 387604 676418
rect 387004 676098 387186 676334
rect 387422 676098 387604 676334
rect 387004 640654 387604 676098
rect 387004 640418 387186 640654
rect 387422 640418 387604 640654
rect 387004 640334 387604 640418
rect 387004 640098 387186 640334
rect 387422 640098 387604 640334
rect 387004 604654 387604 640098
rect 387004 604418 387186 604654
rect 387422 604418 387604 604654
rect 387004 604334 387604 604418
rect 387004 604098 387186 604334
rect 387422 604098 387604 604334
rect 387004 598000 387604 604098
rect 390604 680254 391204 710862
rect 408604 710478 409204 711440
rect 408604 710242 408786 710478
rect 409022 710242 409204 710478
rect 408604 710158 409204 710242
rect 408604 709922 408786 710158
rect 409022 709922 409204 710158
rect 405004 708598 405604 709560
rect 405004 708362 405186 708598
rect 405422 708362 405604 708598
rect 405004 708278 405604 708362
rect 405004 708042 405186 708278
rect 405422 708042 405604 708278
rect 401404 706718 402004 707680
rect 401404 706482 401586 706718
rect 401822 706482 402004 706718
rect 401404 706398 402004 706482
rect 401404 706162 401586 706398
rect 401822 706162 402004 706398
rect 390604 680018 390786 680254
rect 391022 680018 391204 680254
rect 390604 679934 391204 680018
rect 390604 679698 390786 679934
rect 391022 679698 391204 679934
rect 390604 644254 391204 679698
rect 390604 644018 390786 644254
rect 391022 644018 391204 644254
rect 390604 643934 391204 644018
rect 390604 643698 390786 643934
rect 391022 643698 391204 643934
rect 390604 608254 391204 643698
rect 390604 608018 390786 608254
rect 391022 608018 391204 608254
rect 390604 607934 391204 608018
rect 390604 607698 390786 607934
rect 391022 607698 391204 607934
rect 390604 598000 391204 607698
rect 397804 704838 398404 705800
rect 397804 704602 397986 704838
rect 398222 704602 398404 704838
rect 397804 704518 398404 704602
rect 397804 704282 397986 704518
rect 398222 704282 398404 704518
rect 397804 687454 398404 704282
rect 397804 687218 397986 687454
rect 398222 687218 398404 687454
rect 397804 687134 398404 687218
rect 397804 686898 397986 687134
rect 398222 686898 398404 687134
rect 397804 651454 398404 686898
rect 397804 651218 397986 651454
rect 398222 651218 398404 651454
rect 397804 651134 398404 651218
rect 397804 650898 397986 651134
rect 398222 650898 398404 651134
rect 397804 615454 398404 650898
rect 397804 615218 397986 615454
rect 398222 615218 398404 615454
rect 397804 615134 398404 615218
rect 397804 614898 397986 615134
rect 398222 614898 398404 615134
rect 397804 598000 398404 614898
rect 401404 691054 402004 706162
rect 401404 690818 401586 691054
rect 401822 690818 402004 691054
rect 401404 690734 402004 690818
rect 401404 690498 401586 690734
rect 401822 690498 402004 690734
rect 401404 655054 402004 690498
rect 401404 654818 401586 655054
rect 401822 654818 402004 655054
rect 401404 654734 402004 654818
rect 401404 654498 401586 654734
rect 401822 654498 402004 654734
rect 401404 619054 402004 654498
rect 401404 618818 401586 619054
rect 401822 618818 402004 619054
rect 401404 618734 402004 618818
rect 401404 618498 401586 618734
rect 401822 618498 402004 618734
rect 401404 598000 402004 618498
rect 405004 694654 405604 708042
rect 405004 694418 405186 694654
rect 405422 694418 405604 694654
rect 405004 694334 405604 694418
rect 405004 694098 405186 694334
rect 405422 694098 405604 694334
rect 405004 658654 405604 694098
rect 405004 658418 405186 658654
rect 405422 658418 405604 658654
rect 405004 658334 405604 658418
rect 405004 658098 405186 658334
rect 405422 658098 405604 658334
rect 405004 622654 405604 658098
rect 405004 622418 405186 622654
rect 405422 622418 405604 622654
rect 405004 622334 405604 622418
rect 405004 622098 405186 622334
rect 405422 622098 405604 622334
rect 405004 598000 405604 622098
rect 408604 698254 409204 709922
rect 426604 711418 427204 711440
rect 426604 711182 426786 711418
rect 427022 711182 427204 711418
rect 426604 711098 427204 711182
rect 426604 710862 426786 711098
rect 427022 710862 427204 711098
rect 423004 709538 423604 709560
rect 423004 709302 423186 709538
rect 423422 709302 423604 709538
rect 423004 709218 423604 709302
rect 423004 708982 423186 709218
rect 423422 708982 423604 709218
rect 419404 707658 420004 707680
rect 419404 707422 419586 707658
rect 419822 707422 420004 707658
rect 419404 707338 420004 707422
rect 419404 707102 419586 707338
rect 419822 707102 420004 707338
rect 408604 698018 408786 698254
rect 409022 698018 409204 698254
rect 408604 697934 409204 698018
rect 408604 697698 408786 697934
rect 409022 697698 409204 697934
rect 408604 662254 409204 697698
rect 408604 662018 408786 662254
rect 409022 662018 409204 662254
rect 408604 661934 409204 662018
rect 408604 661698 408786 661934
rect 409022 661698 409204 661934
rect 408604 626254 409204 661698
rect 408604 626018 408786 626254
rect 409022 626018 409204 626254
rect 408604 625934 409204 626018
rect 408604 625698 408786 625934
rect 409022 625698 409204 625934
rect 408604 598000 409204 625698
rect 415804 705778 416404 705800
rect 415804 705542 415986 705778
rect 416222 705542 416404 705778
rect 415804 705458 416404 705542
rect 415804 705222 415986 705458
rect 416222 705222 416404 705458
rect 415804 669454 416404 705222
rect 415804 669218 415986 669454
rect 416222 669218 416404 669454
rect 415804 669134 416404 669218
rect 415804 668898 415986 669134
rect 416222 668898 416404 669134
rect 415804 633454 416404 668898
rect 415804 633218 415986 633454
rect 416222 633218 416404 633454
rect 415804 633134 416404 633218
rect 415804 632898 415986 633134
rect 416222 632898 416404 633134
rect 415804 598000 416404 632898
rect 419404 673054 420004 707102
rect 419404 672818 419586 673054
rect 419822 672818 420004 673054
rect 419404 672734 420004 672818
rect 419404 672498 419586 672734
rect 419822 672498 420004 672734
rect 419404 637054 420004 672498
rect 419404 636818 419586 637054
rect 419822 636818 420004 637054
rect 419404 636734 420004 636818
rect 419404 636498 419586 636734
rect 419822 636498 420004 636734
rect 419404 601054 420004 636498
rect 419404 600818 419586 601054
rect 419822 600818 420004 601054
rect 419404 600734 420004 600818
rect 419404 600498 419586 600734
rect 419822 600498 420004 600734
rect 419404 598000 420004 600498
rect 423004 676654 423604 708982
rect 423004 676418 423186 676654
rect 423422 676418 423604 676654
rect 423004 676334 423604 676418
rect 423004 676098 423186 676334
rect 423422 676098 423604 676334
rect 423004 640654 423604 676098
rect 423004 640418 423186 640654
rect 423422 640418 423604 640654
rect 423004 640334 423604 640418
rect 423004 640098 423186 640334
rect 423422 640098 423604 640334
rect 423004 604654 423604 640098
rect 423004 604418 423186 604654
rect 423422 604418 423604 604654
rect 423004 604334 423604 604418
rect 423004 604098 423186 604334
rect 423422 604098 423604 604334
rect 423004 598000 423604 604098
rect 426604 680254 427204 710862
rect 444604 710478 445204 711440
rect 444604 710242 444786 710478
rect 445022 710242 445204 710478
rect 444604 710158 445204 710242
rect 444604 709922 444786 710158
rect 445022 709922 445204 710158
rect 441004 708598 441604 709560
rect 441004 708362 441186 708598
rect 441422 708362 441604 708598
rect 441004 708278 441604 708362
rect 441004 708042 441186 708278
rect 441422 708042 441604 708278
rect 437404 706718 438004 707680
rect 437404 706482 437586 706718
rect 437822 706482 438004 706718
rect 437404 706398 438004 706482
rect 437404 706162 437586 706398
rect 437822 706162 438004 706398
rect 426604 680018 426786 680254
rect 427022 680018 427204 680254
rect 426604 679934 427204 680018
rect 426604 679698 426786 679934
rect 427022 679698 427204 679934
rect 426604 644254 427204 679698
rect 426604 644018 426786 644254
rect 427022 644018 427204 644254
rect 426604 643934 427204 644018
rect 426604 643698 426786 643934
rect 427022 643698 427204 643934
rect 426604 608254 427204 643698
rect 426604 608018 426786 608254
rect 427022 608018 427204 608254
rect 426604 607934 427204 608018
rect 426604 607698 426786 607934
rect 427022 607698 427204 607934
rect 426604 598000 427204 607698
rect 433804 704838 434404 705800
rect 433804 704602 433986 704838
rect 434222 704602 434404 704838
rect 433804 704518 434404 704602
rect 433804 704282 433986 704518
rect 434222 704282 434404 704518
rect 433804 687454 434404 704282
rect 433804 687218 433986 687454
rect 434222 687218 434404 687454
rect 433804 687134 434404 687218
rect 433804 686898 433986 687134
rect 434222 686898 434404 687134
rect 433804 651454 434404 686898
rect 433804 651218 433986 651454
rect 434222 651218 434404 651454
rect 433804 651134 434404 651218
rect 433804 650898 433986 651134
rect 434222 650898 434404 651134
rect 433804 615454 434404 650898
rect 433804 615218 433986 615454
rect 434222 615218 434404 615454
rect 433804 615134 434404 615218
rect 433804 614898 433986 615134
rect 434222 614898 434404 615134
rect 433804 598000 434404 614898
rect 437404 691054 438004 706162
rect 437404 690818 437586 691054
rect 437822 690818 438004 691054
rect 437404 690734 438004 690818
rect 437404 690498 437586 690734
rect 437822 690498 438004 690734
rect 437404 655054 438004 690498
rect 437404 654818 437586 655054
rect 437822 654818 438004 655054
rect 437404 654734 438004 654818
rect 437404 654498 437586 654734
rect 437822 654498 438004 654734
rect 437404 619054 438004 654498
rect 437404 618818 437586 619054
rect 437822 618818 438004 619054
rect 437404 618734 438004 618818
rect 437404 618498 437586 618734
rect 437822 618498 438004 618734
rect 437404 598000 438004 618498
rect 441004 694654 441604 708042
rect 441004 694418 441186 694654
rect 441422 694418 441604 694654
rect 441004 694334 441604 694418
rect 441004 694098 441186 694334
rect 441422 694098 441604 694334
rect 441004 658654 441604 694098
rect 441004 658418 441186 658654
rect 441422 658418 441604 658654
rect 441004 658334 441604 658418
rect 441004 658098 441186 658334
rect 441422 658098 441604 658334
rect 441004 622654 441604 658098
rect 441004 622418 441186 622654
rect 441422 622418 441604 622654
rect 441004 622334 441604 622418
rect 441004 622098 441186 622334
rect 441422 622098 441604 622334
rect 441004 598000 441604 622098
rect 444604 698254 445204 709922
rect 462604 711418 463204 711440
rect 462604 711182 462786 711418
rect 463022 711182 463204 711418
rect 462604 711098 463204 711182
rect 462604 710862 462786 711098
rect 463022 710862 463204 711098
rect 459004 709538 459604 709560
rect 459004 709302 459186 709538
rect 459422 709302 459604 709538
rect 459004 709218 459604 709302
rect 459004 708982 459186 709218
rect 459422 708982 459604 709218
rect 455404 707658 456004 707680
rect 455404 707422 455586 707658
rect 455822 707422 456004 707658
rect 455404 707338 456004 707422
rect 455404 707102 455586 707338
rect 455822 707102 456004 707338
rect 444604 698018 444786 698254
rect 445022 698018 445204 698254
rect 444604 697934 445204 698018
rect 444604 697698 444786 697934
rect 445022 697698 445204 697934
rect 444604 662254 445204 697698
rect 444604 662018 444786 662254
rect 445022 662018 445204 662254
rect 444604 661934 445204 662018
rect 444604 661698 444786 661934
rect 445022 661698 445204 661934
rect 444604 626254 445204 661698
rect 444604 626018 444786 626254
rect 445022 626018 445204 626254
rect 444604 625934 445204 626018
rect 444604 625698 444786 625934
rect 445022 625698 445204 625934
rect 444604 598000 445204 625698
rect 451804 705778 452404 705800
rect 451804 705542 451986 705778
rect 452222 705542 452404 705778
rect 451804 705458 452404 705542
rect 451804 705222 451986 705458
rect 452222 705222 452404 705458
rect 451804 669454 452404 705222
rect 451804 669218 451986 669454
rect 452222 669218 452404 669454
rect 451804 669134 452404 669218
rect 451804 668898 451986 669134
rect 452222 668898 452404 669134
rect 451804 633454 452404 668898
rect 451804 633218 451986 633454
rect 452222 633218 452404 633454
rect 451804 633134 452404 633218
rect 451804 632898 451986 633134
rect 452222 632898 452404 633134
rect 451804 597454 452404 632898
rect 451804 597218 451986 597454
rect 452222 597218 452404 597454
rect 451804 597134 452404 597218
rect 451804 596898 451986 597134
rect 452222 596898 452404 597134
rect 102604 572018 102786 572254
rect 103022 572018 103204 572254
rect 102604 571934 103204 572018
rect 102604 571698 102786 571934
rect 103022 571698 103204 571934
rect 102604 536254 103204 571698
rect 102604 536018 102786 536254
rect 103022 536018 103204 536254
rect 102604 535934 103204 536018
rect 102604 535698 102786 535934
rect 103022 535698 103204 535934
rect 102604 500254 103204 535698
rect 102604 500018 102786 500254
rect 103022 500018 103204 500254
rect 102604 499934 103204 500018
rect 102604 499698 102786 499934
rect 103022 499698 103204 499934
rect 102604 464254 103204 499698
rect 102604 464018 102786 464254
rect 103022 464018 103204 464254
rect 102604 463934 103204 464018
rect 102604 463698 102786 463934
rect 103022 463698 103204 463934
rect 102604 428254 103204 463698
rect 102604 428018 102786 428254
rect 103022 428018 103204 428254
rect 102604 427934 103204 428018
rect 102604 427698 102786 427934
rect 103022 427698 103204 427934
rect 102604 392254 103204 427698
rect 102604 392018 102786 392254
rect 103022 392018 103204 392254
rect 102604 391934 103204 392018
rect 102604 391698 102786 391934
rect 103022 391698 103204 391934
rect 102604 356254 103204 391698
rect 102604 356018 102786 356254
rect 103022 356018 103204 356254
rect 102604 355934 103204 356018
rect 102604 355698 102786 355934
rect 103022 355698 103204 355934
rect 102604 320254 103204 355698
rect 102604 320018 102786 320254
rect 103022 320018 103204 320254
rect 102604 319934 103204 320018
rect 102604 319698 102786 319934
rect 103022 319698 103204 319934
rect 102604 284254 103204 319698
rect 102604 284018 102786 284254
rect 103022 284018 103204 284254
rect 102604 283934 103204 284018
rect 102604 283698 102786 283934
rect 103022 283698 103204 283934
rect 102604 248254 103204 283698
rect 102604 248018 102786 248254
rect 103022 248018 103204 248254
rect 102604 247934 103204 248018
rect 102604 247698 102786 247934
rect 103022 247698 103204 247934
rect 102604 212254 103204 247698
rect 123064 583000 133883 588000
rect 123064 582986 132090 583000
rect 123064 582971 130681 582986
rect 123064 582957 129280 582971
rect 123064 582942 127871 582957
rect 123064 582928 126391 582942
rect 123064 582913 124982 582928
rect 123064 582899 123581 582913
rect 123064 582663 123186 582899
rect 123422 582677 123581 582899
rect 123817 582677 123901 582913
rect 124137 582677 124275 582913
rect 124511 582677 124595 582913
rect 124831 582692 124982 582913
rect 125218 582692 125302 582928
rect 125538 582692 125676 582928
rect 125912 582692 125996 582928
rect 126232 582706 126391 582928
rect 126627 582706 126711 582942
rect 126947 582706 127085 582942
rect 127321 582706 127405 582942
rect 127641 582721 127871 582942
rect 128107 582721 128191 582957
rect 128427 582721 128565 582957
rect 128801 582721 128885 582957
rect 129121 582735 129280 582957
rect 129516 582735 129600 582971
rect 129836 582735 129974 582971
rect 130210 582735 130294 582971
rect 130530 582750 130681 582971
rect 130917 582750 131001 582986
rect 131237 582750 131375 582986
rect 131611 582750 131695 582986
rect 131931 582764 132090 582986
rect 132326 582764 132410 583000
rect 132646 582764 132784 583000
rect 133020 582764 133104 583000
rect 133340 582764 133883 583000
rect 131931 582750 133883 582764
rect 130530 582735 133883 582750
rect 129121 582721 133883 582735
rect 127641 582706 133883 582721
rect 126232 582692 133883 582706
rect 124831 582677 133883 582692
rect 123422 582663 133883 582677
rect 123064 546976 133883 582663
rect 123064 546962 132177 546976
rect 123064 546947 130768 546962
rect 123064 546933 129367 546947
rect 123064 546918 127958 546933
rect 123064 546904 126478 546918
rect 123064 546889 125069 546904
rect 123064 546875 123668 546889
rect 123064 546639 123273 546875
rect 123509 546653 123668 546875
rect 123904 546653 123988 546889
rect 124224 546653 124362 546889
rect 124598 546653 124682 546889
rect 124918 546668 125069 546889
rect 125305 546668 125389 546904
rect 125625 546668 125763 546904
rect 125999 546668 126083 546904
rect 126319 546682 126478 546904
rect 126714 546682 126798 546918
rect 127034 546682 127172 546918
rect 127408 546682 127492 546918
rect 127728 546697 127958 546918
rect 128194 546697 128278 546933
rect 128514 546697 128652 546933
rect 128888 546697 128972 546933
rect 129208 546711 129367 546933
rect 129603 546711 129687 546947
rect 129923 546711 130061 546947
rect 130297 546711 130381 546947
rect 130617 546726 130768 546947
rect 131004 546726 131088 546962
rect 131324 546726 131462 546962
rect 131698 546726 131782 546962
rect 132018 546740 132177 546962
rect 132413 546740 132497 546976
rect 132733 546740 132871 546976
rect 133107 546740 133191 546976
rect 133427 546740 133883 546976
rect 132018 546726 133883 546740
rect 130617 546711 133883 546726
rect 129208 546697 133883 546711
rect 127728 546682 133883 546697
rect 126319 546668 133883 546682
rect 124918 546653 133883 546668
rect 123509 546639 133883 546653
rect 123064 510973 133883 546639
rect 123064 510959 132137 510973
rect 123064 510944 130728 510959
rect 123064 510930 129327 510944
rect 123064 510915 127918 510930
rect 123064 510901 126438 510915
rect 123064 510886 125029 510901
rect 123064 510872 123628 510886
rect 123064 510636 123233 510872
rect 123469 510650 123628 510872
rect 123864 510650 123948 510886
rect 124184 510650 124322 510886
rect 124558 510650 124642 510886
rect 124878 510665 125029 510886
rect 125265 510665 125349 510901
rect 125585 510665 125723 510901
rect 125959 510665 126043 510901
rect 126279 510679 126438 510901
rect 126674 510679 126758 510915
rect 126994 510679 127132 510915
rect 127368 510679 127452 510915
rect 127688 510694 127918 510915
rect 128154 510694 128238 510930
rect 128474 510694 128612 510930
rect 128848 510694 128932 510930
rect 129168 510708 129327 510930
rect 129563 510708 129647 510944
rect 129883 510708 130021 510944
rect 130257 510708 130341 510944
rect 130577 510723 130728 510944
rect 130964 510723 131048 510959
rect 131284 510723 131422 510959
rect 131658 510723 131742 510959
rect 131978 510737 132137 510959
rect 132373 510737 132457 510973
rect 132693 510737 132831 510973
rect 133067 510737 133151 510973
rect 133387 510737 133883 510973
rect 131978 510723 133883 510737
rect 130577 510708 133883 510723
rect 129168 510694 133883 510708
rect 127688 510679 133883 510694
rect 126279 510665 133883 510679
rect 124878 510650 133883 510665
rect 123469 510636 133883 510650
rect 123064 473607 133883 510636
rect 123064 473593 132316 473607
rect 123064 473578 130907 473593
rect 123064 473564 129506 473578
rect 123064 473549 128097 473564
rect 123064 473535 126617 473549
rect 123064 473520 125208 473535
rect 123064 473506 123807 473520
rect 123064 473270 123412 473506
rect 123648 473270 123807 473506
rect 123064 473186 123807 473270
rect 123064 472950 123412 473186
rect 123648 472950 123807 473186
rect 123064 472866 123807 472950
rect 123064 472630 123412 472866
rect 123648 472644 123807 472866
rect 124363 472644 124501 473520
rect 125057 472659 125208 473520
rect 125764 472659 125902 473535
rect 126458 472673 126617 473535
rect 127173 472673 127311 473549
rect 127867 472688 128097 473549
rect 128653 472688 128791 473564
rect 129347 472702 129506 473564
rect 130062 472702 130200 473578
rect 130756 472717 130907 473578
rect 131463 472717 131601 473593
rect 132157 472731 132316 473593
rect 132872 472731 133010 473607
rect 133566 472731 133883 473607
rect 132157 472717 133883 472731
rect 130756 472702 133883 472717
rect 129347 472688 133883 472702
rect 127867 472673 133883 472688
rect 126458 472659 133883 472673
rect 125057 472644 133883 472659
rect 123648 472630 133883 472644
rect 123064 465621 133883 472630
rect 123064 465607 132381 465621
rect 123064 465592 130972 465607
rect 123064 465578 129571 465592
rect 123064 465563 128162 465578
rect 123064 465549 126682 465563
rect 123064 465534 125273 465549
rect 123064 465520 123872 465534
rect 123064 465284 123477 465520
rect 123713 465284 123872 465520
rect 123064 465200 123872 465284
rect 123064 464964 123477 465200
rect 123713 464964 123872 465200
rect 123064 464880 123872 464964
rect 123064 464644 123477 464880
rect 123713 464658 123872 464880
rect 124428 464658 124566 465534
rect 125122 464673 125273 465534
rect 125829 464673 125967 465549
rect 126523 464687 126682 465549
rect 127238 464687 127376 465563
rect 127932 464702 128162 465563
rect 128718 464702 128856 465578
rect 129412 464716 129571 465578
rect 130127 464716 130265 465592
rect 130821 464731 130972 465592
rect 131528 464731 131666 465607
rect 132222 464745 132381 465607
rect 132937 464745 133075 465621
rect 133631 464745 133883 465621
rect 132222 464731 133883 464745
rect 130821 464716 133883 464731
rect 129412 464702 133883 464716
rect 127932 464687 133883 464702
rect 126523 464673 133883 464687
rect 125122 464658 133883 464673
rect 123713 464644 133883 464658
rect 123064 457675 133883 464644
rect 123064 457661 132241 457675
rect 123064 457646 130832 457661
rect 123064 457632 129431 457646
rect 123064 457617 128022 457632
rect 123064 457603 126542 457617
rect 123064 457588 125133 457603
rect 123064 457574 123732 457588
rect 123064 457338 123337 457574
rect 123573 457338 123732 457574
rect 123064 457254 123732 457338
rect 123064 457018 123337 457254
rect 123573 457018 123732 457254
rect 123064 456934 123732 457018
rect 123064 456698 123337 456934
rect 123573 456712 123732 456934
rect 124288 456712 124426 457588
rect 124982 456727 125133 457588
rect 125689 456727 125827 457603
rect 126383 456741 126542 457603
rect 127098 456741 127236 457617
rect 127792 456756 128022 457617
rect 128578 456756 128716 457632
rect 129272 456770 129431 457632
rect 129987 456770 130125 457646
rect 130681 456785 130832 457646
rect 131388 456785 131526 457661
rect 132082 456799 132241 457661
rect 132797 456799 132935 457675
rect 133491 456799 133883 457675
rect 132082 456785 133883 456799
rect 130681 456770 133883 456785
rect 129272 456756 133883 456770
rect 127792 456741 133883 456756
rect 126383 456727 133883 456741
rect 124982 456712 133883 456727
rect 123573 456698 133883 456712
rect 123064 449642 133883 456698
rect 123064 449628 132296 449642
rect 123064 449613 130887 449628
rect 123064 449599 129486 449613
rect 123064 449584 128077 449599
rect 123064 449570 126597 449584
rect 123064 449555 125188 449570
rect 123064 449541 123787 449555
rect 123064 449305 123392 449541
rect 123628 449305 123787 449541
rect 123064 449221 123787 449305
rect 123064 448985 123392 449221
rect 123628 448985 123787 449221
rect 123064 448901 123787 448985
rect 123064 448665 123392 448901
rect 123628 448679 123787 448901
rect 124343 448679 124481 449555
rect 125037 448694 125188 449555
rect 125744 448694 125882 449570
rect 126438 448708 126597 449570
rect 127153 448708 127291 449584
rect 127847 448723 128077 449584
rect 128633 448723 128771 449599
rect 129327 448737 129486 449599
rect 130042 448737 130180 449613
rect 130736 448752 130887 449613
rect 131443 448752 131581 449628
rect 132137 448766 132296 449628
rect 132852 448766 132990 449642
rect 133546 448766 133883 449642
rect 132137 448752 133883 448766
rect 130736 448737 133883 448752
rect 129327 448723 133883 448737
rect 127847 448708 133883 448723
rect 126438 448694 133883 448708
rect 125037 448679 133883 448694
rect 123628 448665 133883 448679
rect 123064 441654 133883 448665
rect 123064 441640 132410 441654
rect 123064 441625 131001 441640
rect 123064 441611 129600 441625
rect 123064 441596 128191 441611
rect 123064 441582 126711 441596
rect 123064 441567 125302 441582
rect 123064 441553 123901 441567
rect 123064 441317 123506 441553
rect 123742 441317 123901 441553
rect 123064 441233 123901 441317
rect 123064 440997 123506 441233
rect 123742 440997 123901 441233
rect 123064 440913 123901 440997
rect 123064 440677 123506 440913
rect 123742 440691 123901 440913
rect 124457 440691 124595 441567
rect 125151 440706 125302 441567
rect 125858 440706 125996 441582
rect 126552 440720 126711 441582
rect 127267 440720 127405 441596
rect 127961 440735 128191 441596
rect 128747 440735 128885 441611
rect 129441 440749 129600 441611
rect 130156 440749 130294 441625
rect 130850 440764 131001 441625
rect 131557 440764 131695 441640
rect 132251 440778 132410 441640
rect 132966 440778 133104 441654
rect 133660 440778 133883 441654
rect 132251 440764 133883 440778
rect 130850 440749 133883 440764
rect 129441 440735 133883 440749
rect 127961 440720 133883 440735
rect 126552 440706 133883 440720
rect 125151 440691 133883 440706
rect 123742 440677 133883 440691
rect 123064 433609 133883 440677
rect 123064 433595 132340 433609
rect 123064 433580 130931 433595
rect 123064 433566 129530 433580
rect 123064 433551 128121 433566
rect 123064 433537 126641 433551
rect 123064 433522 125232 433537
rect 123064 433508 123831 433522
rect 123064 433272 123436 433508
rect 123672 433272 123831 433508
rect 123064 433188 123831 433272
rect 123064 432952 123436 433188
rect 123672 432952 123831 433188
rect 123064 432868 123831 432952
rect 123064 432632 123436 432868
rect 123672 432646 123831 432868
rect 124387 432646 124525 433522
rect 125081 432661 125232 433522
rect 125788 432661 125926 433537
rect 126482 432675 126641 433537
rect 127197 432675 127335 433551
rect 127891 432690 128121 433551
rect 128677 432690 128815 433566
rect 129371 432704 129530 433566
rect 130086 432704 130224 433580
rect 130780 432719 130931 433580
rect 131487 432719 131625 433595
rect 132181 432733 132340 433595
rect 132896 432733 133034 433609
rect 133590 432733 133883 433609
rect 132181 432719 133883 432733
rect 130780 432704 133883 432719
rect 129371 432690 133883 432704
rect 127891 432675 133883 432690
rect 126482 432661 133883 432675
rect 125081 432646 133883 432661
rect 123672 432632 133883 432646
rect 123064 425665 133883 432632
rect 123064 425651 132342 425665
rect 123064 425636 130933 425651
rect 123064 425622 129532 425636
rect 123064 425607 128123 425622
rect 123064 425593 126643 425607
rect 123064 425578 125234 425593
rect 123064 425564 123833 425578
rect 123064 425328 123438 425564
rect 123674 425328 123833 425564
rect 123064 425244 123833 425328
rect 123064 425008 123438 425244
rect 123674 425008 123833 425244
rect 123064 424924 123833 425008
rect 123064 424688 123438 424924
rect 123674 424702 123833 424924
rect 124389 424702 124527 425578
rect 125083 424717 125234 425578
rect 125790 424717 125928 425593
rect 126484 424731 126643 425593
rect 127199 424731 127337 425607
rect 127893 424746 128123 425607
rect 128679 424746 128817 425622
rect 129373 424760 129532 425622
rect 130088 424760 130226 425636
rect 130782 424775 130933 425636
rect 131489 424775 131627 425651
rect 132183 424789 132342 425651
rect 132898 424789 133036 425665
rect 133592 424789 133883 425665
rect 132183 424775 133883 424789
rect 130782 424760 133883 424775
rect 129373 424746 133883 424760
rect 127893 424731 133883 424746
rect 126484 424717 133883 424731
rect 125083 424702 133883 424717
rect 123674 424688 133883 424702
rect 123064 417606 133883 424688
rect 123064 417592 132313 417606
rect 123064 417577 130904 417592
rect 123064 417563 129503 417577
rect 123064 417548 128094 417563
rect 123064 417534 126614 417548
rect 123064 417519 125205 417534
rect 123064 417505 123804 417519
rect 123064 417269 123409 417505
rect 123645 417269 123804 417505
rect 123064 417185 123804 417269
rect 123064 416949 123409 417185
rect 123645 416949 123804 417185
rect 123064 416865 123804 416949
rect 123064 416629 123409 416865
rect 123645 416643 123804 416865
rect 124360 416643 124498 417519
rect 125054 416658 125205 417519
rect 125761 416658 125899 417534
rect 126455 416672 126614 417534
rect 127170 416672 127308 417548
rect 127864 416687 128094 417548
rect 128650 416687 128788 417563
rect 129344 416701 129503 417563
rect 130059 416701 130197 417577
rect 130753 416716 130904 417577
rect 131460 416716 131598 417592
rect 132154 416730 132313 417592
rect 132869 416730 133007 417606
rect 133563 416730 133883 417606
rect 132154 416716 133883 416730
rect 130753 416701 133883 416716
rect 129344 416687 133883 416701
rect 127864 416672 133883 416687
rect 126455 416658 133883 416672
rect 125054 416643 133883 416658
rect 123645 416629 133883 416643
rect 123064 409638 133883 416629
rect 123064 409624 132400 409638
rect 123064 409609 130991 409624
rect 123064 409595 129590 409609
rect 123064 409580 128181 409595
rect 123064 409566 126701 409580
rect 123064 409551 125292 409566
rect 123064 409537 123891 409551
rect 123064 409301 123496 409537
rect 123732 409301 123891 409537
rect 123064 409217 123891 409301
rect 123064 408981 123496 409217
rect 123732 408981 123891 409217
rect 123064 408897 123891 408981
rect 123064 408661 123496 408897
rect 123732 408675 123891 408897
rect 124447 408675 124585 409551
rect 125141 408690 125292 409551
rect 125848 408690 125986 409566
rect 126542 408704 126701 409566
rect 127257 408704 127395 409580
rect 127951 408719 128181 409580
rect 128737 408719 128875 409595
rect 129431 408733 129590 409595
rect 130146 408733 130284 409609
rect 130840 408748 130991 409609
rect 131547 408748 131685 409624
rect 132241 408762 132400 409624
rect 132956 408762 133094 409638
rect 133650 408762 133883 409638
rect 132241 408748 133883 408762
rect 130840 408733 133883 408748
rect 129431 408719 133883 408733
rect 127951 408704 133883 408719
rect 126542 408690 133883 408704
rect 125141 408675 133883 408690
rect 123732 408661 133883 408675
rect 123064 401640 133883 408661
rect 123064 401626 132334 401640
rect 123064 401611 130925 401626
rect 123064 401597 129524 401611
rect 123064 401582 128115 401597
rect 123064 401568 126635 401582
rect 123064 401553 125226 401568
rect 123064 401539 123825 401553
rect 123064 401303 123430 401539
rect 123666 401303 123825 401539
rect 123064 401219 123825 401303
rect 123064 400983 123430 401219
rect 123666 400983 123825 401219
rect 123064 400899 123825 400983
rect 123064 400663 123430 400899
rect 123666 400677 123825 400899
rect 124381 400677 124519 401553
rect 125075 400692 125226 401553
rect 125782 400692 125920 401568
rect 126476 400706 126635 401568
rect 127191 400706 127329 401582
rect 127885 400721 128115 401582
rect 128671 400721 128809 401597
rect 129365 400735 129524 401597
rect 130080 400735 130218 401611
rect 130774 400750 130925 401611
rect 131481 400750 131619 401626
rect 132175 400764 132334 401626
rect 132890 400764 133028 401640
rect 133584 400764 133883 401640
rect 132175 400750 133883 400764
rect 130774 400735 133883 400750
rect 129365 400721 133883 400735
rect 127885 400706 133883 400721
rect 126476 400692 133883 400706
rect 125075 400677 133883 400692
rect 123666 400663 133883 400677
rect 123064 393640 133883 400663
rect 123064 393626 132304 393640
rect 123064 393611 130895 393626
rect 123064 393597 129494 393611
rect 123064 393582 128085 393597
rect 123064 393568 126605 393582
rect 123064 393553 125196 393568
rect 123064 393539 123795 393553
rect 123064 393303 123400 393539
rect 123636 393303 123795 393539
rect 123064 393219 123795 393303
rect 123064 392983 123400 393219
rect 123636 392983 123795 393219
rect 123064 392899 123795 392983
rect 123064 392663 123400 392899
rect 123636 392677 123795 392899
rect 124351 392677 124489 393553
rect 125045 392692 125196 393553
rect 125752 392692 125890 393568
rect 126446 392706 126605 393568
rect 127161 392706 127299 393582
rect 127855 392721 128085 393582
rect 128641 392721 128779 393597
rect 129335 392735 129494 393597
rect 130050 392735 130188 393611
rect 130744 392750 130895 393611
rect 131451 392750 131589 393626
rect 132145 392764 132304 393626
rect 132860 392764 132998 393640
rect 133554 392764 133883 393640
rect 132145 392750 133883 392764
rect 130744 392735 133883 392750
rect 129335 392721 133883 392735
rect 127855 392706 133883 392721
rect 126446 392692 133883 392706
rect 125045 392677 133883 392692
rect 123636 392663 133883 392677
rect 123064 385612 133883 392663
rect 123064 385598 132385 385612
rect 123064 385583 130976 385598
rect 123064 385569 129575 385583
rect 123064 385554 128166 385569
rect 123064 385540 126686 385554
rect 123064 385525 125277 385540
rect 123064 385511 123876 385525
rect 123064 385275 123481 385511
rect 123717 385275 123876 385511
rect 123064 385191 123876 385275
rect 123064 384955 123481 385191
rect 123717 384955 123876 385191
rect 123064 384871 123876 384955
rect 123064 384635 123481 384871
rect 123717 384649 123876 384871
rect 124432 384649 124570 385525
rect 125126 384664 125277 385525
rect 125833 384664 125971 385540
rect 126527 384678 126686 385540
rect 127242 384678 127380 385554
rect 127936 384693 128166 385554
rect 128722 384693 128860 385569
rect 129416 384707 129575 385569
rect 130131 384707 130269 385583
rect 130825 384722 130976 385583
rect 131532 384722 131670 385598
rect 132226 384736 132385 385598
rect 132941 384736 133079 385612
rect 133635 384736 133883 385612
rect 132226 384722 133883 384736
rect 130825 384707 133883 384722
rect 129416 384693 133883 384707
rect 127936 384678 133883 384693
rect 126527 384664 133883 384678
rect 125126 384649 133883 384664
rect 123717 384635 133883 384649
rect 123064 377654 133883 384635
rect 123064 377640 132317 377654
rect 123064 377625 130908 377640
rect 123064 377611 129507 377625
rect 123064 377596 128098 377611
rect 123064 377582 126618 377596
rect 123064 377567 125209 377582
rect 123064 377553 123808 377567
rect 123064 377317 123413 377553
rect 123649 377317 123808 377553
rect 123064 377233 123808 377317
rect 123064 376997 123413 377233
rect 123649 376997 123808 377233
rect 123064 376913 123808 376997
rect 123064 376677 123413 376913
rect 123649 376691 123808 376913
rect 124364 376691 124502 377567
rect 125058 376706 125209 377567
rect 125765 376706 125903 377582
rect 126459 376720 126618 377582
rect 127174 376720 127312 377596
rect 127868 376735 128098 377596
rect 128654 376735 128792 377611
rect 129348 376749 129507 377611
rect 130063 376749 130201 377625
rect 130757 376764 130908 377625
rect 131464 376764 131602 377640
rect 132158 376778 132317 377640
rect 132873 376778 133011 377654
rect 133567 376778 133883 377654
rect 132158 376764 133883 376778
rect 130757 376749 133883 376764
rect 129348 376735 133883 376749
rect 127868 376720 133883 376735
rect 126459 376706 133883 376720
rect 125058 376691 133883 376706
rect 123649 376677 133883 376691
rect 123064 369592 133883 376677
rect 123064 369578 132246 369592
rect 123064 369563 130837 369578
rect 123064 369549 129436 369563
rect 123064 369534 128027 369549
rect 123064 369520 126547 369534
rect 123064 369505 125138 369520
rect 123064 369491 123737 369505
rect 123064 369255 123342 369491
rect 123578 369255 123737 369491
rect 123064 369171 123737 369255
rect 123064 368935 123342 369171
rect 123578 368935 123737 369171
rect 123064 368851 123737 368935
rect 123064 368615 123342 368851
rect 123578 368629 123737 368851
rect 124293 368629 124431 369505
rect 124987 368644 125138 369505
rect 125694 368644 125832 369520
rect 126388 368658 126547 369520
rect 127103 368658 127241 369534
rect 127797 368673 128027 369534
rect 128583 368673 128721 369549
rect 129277 368687 129436 369549
rect 129992 368687 130130 369563
rect 130686 368702 130837 369563
rect 131393 368702 131531 369578
rect 132087 368716 132246 369578
rect 132802 368716 132940 369592
rect 133496 368716 133883 369592
rect 132087 368702 133883 368716
rect 130686 368687 133883 368702
rect 129277 368673 133883 368687
rect 127797 368658 133883 368673
rect 126388 368644 133883 368658
rect 124987 368629 133883 368644
rect 123578 368615 133883 368629
rect 123064 361640 133883 368615
rect 123064 361626 132385 361640
rect 123064 361611 130976 361626
rect 123064 361597 129575 361611
rect 123064 361582 128166 361597
rect 123064 361568 126686 361582
rect 123064 361553 125277 361568
rect 123064 361539 123876 361553
rect 123064 361303 123481 361539
rect 123717 361303 123876 361539
rect 123064 361219 123876 361303
rect 123064 360983 123481 361219
rect 123717 360983 123876 361219
rect 123064 360899 123876 360983
rect 123064 360663 123481 360899
rect 123717 360677 123876 360899
rect 124432 360677 124570 361553
rect 125126 360692 125277 361553
rect 125833 360692 125971 361568
rect 126527 360706 126686 361568
rect 127242 360706 127380 361582
rect 127936 360721 128166 361582
rect 128722 360721 128860 361597
rect 129416 360735 129575 361597
rect 130131 360735 130269 361611
rect 130825 360750 130976 361611
rect 131532 360750 131670 361626
rect 132226 360764 132385 361626
rect 132941 360764 133079 361640
rect 133635 360764 133883 361640
rect 132226 360750 133883 360764
rect 130825 360735 133883 360750
rect 129416 360721 133883 360735
rect 127936 360706 133883 360721
rect 126527 360692 133883 360706
rect 125126 360677 133883 360692
rect 123717 360663 133883 360677
rect 123064 353614 133883 360663
rect 123064 353600 132314 353614
rect 123064 353585 130905 353600
rect 123064 353571 129504 353585
rect 123064 353556 128095 353571
rect 123064 353542 126615 353556
rect 123064 353527 125206 353542
rect 123064 353513 123805 353527
rect 123064 353277 123410 353513
rect 123646 353277 123805 353513
rect 123064 353193 123805 353277
rect 123064 352957 123410 353193
rect 123646 352957 123805 353193
rect 123064 352873 123805 352957
rect 123064 352637 123410 352873
rect 123646 352651 123805 352873
rect 124361 352651 124499 353527
rect 125055 352666 125206 353527
rect 125762 352666 125900 353542
rect 126456 352680 126615 353542
rect 127171 352680 127309 353556
rect 127865 352695 128095 353556
rect 128651 352695 128789 353571
rect 129345 352709 129504 353571
rect 130060 352709 130198 353585
rect 130754 352724 130905 353585
rect 131461 352724 131599 353600
rect 132155 352738 132314 353600
rect 132870 352738 133008 353614
rect 133564 352738 133883 353614
rect 132155 352724 133883 352738
rect 130754 352709 133883 352724
rect 129345 352695 133883 352709
rect 127865 352680 133883 352695
rect 126456 352666 133883 352680
rect 125055 352651 133883 352666
rect 123646 352637 133883 352651
rect 123064 345634 133883 352637
rect 123064 345620 132416 345634
rect 123064 345605 131007 345620
rect 123064 345591 129606 345605
rect 123064 345576 128197 345591
rect 123064 345562 126717 345576
rect 123064 345547 125308 345562
rect 123064 345533 123907 345547
rect 123064 345297 123512 345533
rect 123748 345297 123907 345533
rect 123064 345213 123907 345297
rect 123064 344977 123512 345213
rect 123748 344977 123907 345213
rect 123064 344893 123907 344977
rect 123064 344657 123512 344893
rect 123748 344671 123907 344893
rect 124463 344671 124601 345547
rect 125157 344686 125308 345547
rect 125864 344686 126002 345562
rect 126558 344700 126717 345562
rect 127273 344700 127411 345576
rect 127967 344715 128197 345576
rect 128753 344715 128891 345591
rect 129447 344729 129606 345591
rect 130162 344729 130300 345605
rect 130856 344744 131007 345605
rect 131563 344744 131701 345620
rect 132257 344758 132416 345620
rect 132972 344758 133110 345634
rect 133666 344758 133883 345634
rect 132257 344744 133883 344758
rect 130856 344729 133883 344744
rect 129447 344715 133883 344729
rect 127967 344700 133883 344715
rect 126558 344686 133883 344700
rect 125157 344671 133883 344686
rect 123748 344657 133883 344671
rect 123064 330947 133883 344657
rect 123064 330933 132359 330947
rect 123064 330918 130950 330933
rect 123064 330904 129549 330918
rect 123064 330889 128140 330904
rect 123064 330875 126660 330889
rect 123064 330860 125251 330875
rect 123064 330846 123850 330860
rect 123064 330610 123455 330846
rect 123691 330624 123850 330846
rect 124086 330624 124170 330860
rect 124406 330624 124544 330860
rect 124780 330624 124864 330860
rect 125100 330639 125251 330860
rect 125487 330639 125571 330875
rect 125807 330639 125945 330875
rect 126181 330639 126265 330875
rect 126501 330653 126660 330875
rect 126896 330653 126980 330889
rect 127216 330653 127354 330889
rect 127590 330653 127674 330889
rect 127910 330668 128140 330889
rect 128376 330668 128460 330904
rect 128696 330668 128834 330904
rect 129070 330668 129154 330904
rect 129390 330682 129549 330904
rect 129785 330682 129869 330918
rect 130105 330682 130243 330918
rect 130479 330682 130563 330918
rect 130799 330697 130950 330918
rect 131186 330697 131270 330933
rect 131506 330697 131644 330933
rect 131880 330697 131964 330933
rect 132200 330711 132359 330933
rect 132595 330711 132679 330947
rect 132915 330711 133053 330947
rect 133289 330711 133373 330947
rect 133609 330711 133883 330947
rect 132200 330697 133883 330711
rect 130799 330682 133883 330697
rect 129390 330668 133883 330682
rect 127910 330653 133883 330668
rect 126501 330639 133883 330653
rect 125100 330624 133883 330639
rect 123691 330610 133883 330624
rect 123064 294944 133883 330610
rect 123064 294930 132376 294944
rect 123064 294915 130967 294930
rect 123064 294901 129566 294915
rect 123064 294886 128157 294901
rect 123064 294872 126677 294886
rect 123064 294857 125268 294872
rect 123064 294843 123867 294857
rect 123064 294607 123472 294843
rect 123708 294621 123867 294843
rect 124103 294621 124187 294857
rect 124423 294621 124561 294857
rect 124797 294621 124881 294857
rect 125117 294636 125268 294857
rect 125504 294636 125588 294872
rect 125824 294636 125962 294872
rect 126198 294636 126282 294872
rect 126518 294650 126677 294872
rect 126913 294650 126997 294886
rect 127233 294650 127371 294886
rect 127607 294650 127691 294886
rect 127927 294665 128157 294886
rect 128393 294665 128477 294901
rect 128713 294665 128851 294901
rect 129087 294665 129171 294901
rect 129407 294679 129566 294901
rect 129802 294679 129886 294915
rect 130122 294679 130260 294915
rect 130496 294679 130580 294915
rect 130816 294694 130967 294915
rect 131203 294694 131287 294930
rect 131523 294694 131661 294930
rect 131897 294694 131981 294930
rect 132217 294708 132376 294930
rect 132612 294708 132696 294944
rect 132932 294708 133070 294944
rect 133306 294708 133390 294944
rect 133626 294708 133883 294944
rect 132217 294694 133883 294708
rect 130816 294679 133883 294694
rect 129407 294665 133883 294679
rect 127927 294650 133883 294665
rect 126518 294636 133883 294650
rect 125117 294621 133883 294636
rect 123708 294607 133883 294621
rect 123064 258944 133883 294607
rect 123064 258930 132142 258944
rect 123064 258915 130733 258930
rect 123064 258901 129332 258915
rect 123064 258886 127923 258901
rect 123064 258872 126443 258886
rect 123064 258857 125034 258872
rect 123064 258843 123633 258857
rect 123064 258607 123238 258843
rect 123474 258621 123633 258843
rect 123869 258621 123953 258857
rect 124189 258621 124327 258857
rect 124563 258621 124647 258857
rect 124883 258636 125034 258857
rect 125270 258636 125354 258872
rect 125590 258636 125728 258872
rect 125964 258636 126048 258872
rect 126284 258650 126443 258872
rect 126679 258650 126763 258886
rect 126999 258650 127137 258886
rect 127373 258650 127457 258886
rect 127693 258665 127923 258886
rect 128159 258665 128243 258901
rect 128479 258665 128617 258901
rect 128853 258665 128937 258901
rect 129173 258679 129332 258901
rect 129568 258679 129652 258915
rect 129888 258679 130026 258915
rect 130262 258679 130346 258915
rect 130582 258694 130733 258915
rect 130969 258694 131053 258930
rect 131289 258694 131427 258930
rect 131663 258694 131747 258930
rect 131983 258708 132142 258930
rect 132378 258708 132462 258944
rect 132698 258708 132836 258944
rect 133072 258708 133156 258944
rect 133392 258708 133883 258944
rect 131983 258694 133883 258708
rect 130582 258679 133883 258694
rect 129173 258665 133883 258679
rect 127693 258650 133883 258665
rect 126284 258636 133883 258650
rect 124883 258621 133883 258636
rect 123474 258607 133883 258621
rect 123064 236000 133883 258607
rect 140742 579394 151561 588000
rect 140742 579380 149841 579394
rect 140742 579365 148432 579380
rect 140742 579351 147031 579365
rect 140742 579336 145622 579351
rect 140742 579322 144142 579336
rect 140742 579307 142733 579322
rect 140742 579293 141332 579307
rect 140742 579057 140937 579293
rect 141173 579071 141332 579293
rect 141568 579071 141652 579307
rect 141888 579071 142026 579307
rect 142262 579071 142346 579307
rect 142582 579086 142733 579307
rect 142969 579086 143053 579322
rect 143289 579086 143427 579322
rect 143663 579086 143747 579322
rect 143983 579100 144142 579322
rect 144378 579100 144462 579336
rect 144698 579100 144836 579336
rect 145072 579100 145156 579336
rect 145392 579115 145622 579336
rect 145858 579115 145942 579351
rect 146178 579115 146316 579351
rect 146552 579115 146636 579351
rect 146872 579129 147031 579351
rect 147267 579129 147351 579365
rect 147587 579129 147725 579365
rect 147961 579129 148045 579365
rect 148281 579144 148432 579365
rect 148668 579144 148752 579380
rect 148988 579144 149126 579380
rect 149362 579144 149446 579380
rect 149682 579158 149841 579380
rect 150077 579158 150161 579394
rect 150397 579158 150535 579394
rect 150771 579158 150855 579394
rect 151091 579158 151561 579394
rect 149682 579144 151561 579158
rect 148281 579129 151561 579144
rect 146872 579115 151561 579129
rect 145392 579100 151561 579115
rect 143983 579086 151561 579100
rect 142582 579071 151561 579086
rect 141173 579057 151561 579071
rect 140742 543373 151561 579057
rect 140742 543359 149968 543373
rect 140742 543344 148559 543359
rect 140742 543330 147158 543344
rect 140742 543315 145749 543330
rect 140742 543301 144269 543315
rect 140742 543286 142860 543301
rect 140742 543272 141459 543286
rect 140742 543036 141064 543272
rect 141300 543050 141459 543272
rect 141695 543050 141779 543286
rect 142015 543050 142153 543286
rect 142389 543050 142473 543286
rect 142709 543065 142860 543286
rect 143096 543065 143180 543301
rect 143416 543065 143554 543301
rect 143790 543065 143874 543301
rect 144110 543079 144269 543301
rect 144505 543079 144589 543315
rect 144825 543079 144963 543315
rect 145199 543079 145283 543315
rect 145519 543094 145749 543315
rect 145985 543094 146069 543330
rect 146305 543094 146443 543330
rect 146679 543094 146763 543330
rect 146999 543108 147158 543330
rect 147394 543108 147478 543344
rect 147714 543108 147852 543344
rect 148088 543108 148172 543344
rect 148408 543123 148559 543344
rect 148795 543123 148879 543359
rect 149115 543123 149253 543359
rect 149489 543123 149573 543359
rect 149809 543137 149968 543359
rect 150204 543137 150288 543373
rect 150524 543137 150662 543373
rect 150898 543137 150982 543373
rect 151218 543137 151561 543373
rect 149809 543123 151561 543137
rect 148408 543108 151561 543123
rect 146999 543094 151561 543108
rect 145519 543079 151561 543094
rect 144110 543065 151561 543079
rect 142709 543050 151561 543065
rect 141300 543036 151561 543050
rect 140742 507406 151561 543036
rect 140742 507392 150152 507406
rect 140742 507377 148743 507392
rect 140742 507363 147342 507377
rect 140742 507348 145933 507363
rect 140742 507334 144453 507348
rect 140742 507319 143044 507334
rect 140742 507305 141643 507319
rect 140742 507069 141248 507305
rect 141484 507083 141643 507305
rect 141879 507083 141963 507319
rect 142199 507083 142337 507319
rect 142573 507083 142657 507319
rect 142893 507098 143044 507319
rect 143280 507098 143364 507334
rect 143600 507098 143738 507334
rect 143974 507098 144058 507334
rect 144294 507112 144453 507334
rect 144689 507112 144773 507348
rect 145009 507112 145147 507348
rect 145383 507112 145467 507348
rect 145703 507127 145933 507348
rect 146169 507127 146253 507363
rect 146489 507127 146627 507363
rect 146863 507127 146947 507363
rect 147183 507141 147342 507363
rect 147578 507141 147662 507377
rect 147898 507141 148036 507377
rect 148272 507141 148356 507377
rect 148592 507156 148743 507377
rect 148979 507156 149063 507392
rect 149299 507156 149437 507392
rect 149673 507156 149757 507392
rect 149993 507170 150152 507392
rect 150388 507170 150472 507406
rect 150708 507170 150846 507406
rect 151082 507170 151166 507406
rect 151402 507170 151561 507406
rect 149993 507156 151561 507170
rect 148592 507141 151561 507156
rect 147183 507127 151561 507141
rect 145703 507112 151561 507127
rect 144294 507098 151561 507112
rect 142893 507083 151561 507098
rect 141484 507069 151561 507083
rect 140742 471909 151561 507069
rect 140742 471895 149969 471909
rect 140742 471880 148560 471895
rect 140742 471866 147159 471880
rect 140742 471851 145750 471866
rect 140742 471837 144270 471851
rect 140742 471822 142861 471837
rect 140742 471808 141460 471822
rect 140742 471572 141065 471808
rect 141301 471572 141460 471808
rect 140742 471488 141460 471572
rect 140742 471252 141065 471488
rect 141301 471252 141460 471488
rect 140742 471168 141460 471252
rect 140742 470932 141065 471168
rect 141301 470946 141460 471168
rect 142016 470946 142154 471822
rect 142710 470961 142861 471822
rect 143417 470961 143555 471837
rect 144111 470975 144270 471837
rect 144826 470975 144964 471851
rect 145520 470990 145750 471851
rect 146306 470990 146444 471866
rect 147000 471004 147159 471866
rect 147715 471004 147853 471880
rect 148409 471019 148560 471880
rect 149116 471019 149254 471895
rect 149810 471033 149969 471895
rect 150525 471033 150663 471909
rect 151219 471033 151561 471909
rect 149810 471019 151561 471033
rect 148409 471004 151561 471019
rect 147000 470990 151561 471004
rect 145520 470975 151561 470990
rect 144111 470961 151561 470975
rect 142710 470946 151561 470961
rect 141301 470932 151561 470946
rect 140742 463952 151561 470932
rect 140742 463938 149849 463952
rect 140742 463923 148440 463938
rect 140742 463909 147039 463923
rect 140742 463894 145630 463909
rect 140742 463880 144150 463894
rect 140742 463865 142741 463880
rect 140742 463851 141340 463865
rect 140742 463615 140945 463851
rect 141181 463615 141340 463851
rect 140742 463531 141340 463615
rect 140742 463295 140945 463531
rect 141181 463295 141340 463531
rect 140742 463211 141340 463295
rect 140742 462975 140945 463211
rect 141181 462989 141340 463211
rect 141896 462989 142034 463865
rect 142590 463004 142741 463865
rect 143297 463004 143435 463880
rect 143991 463018 144150 463880
rect 144706 463018 144844 463894
rect 145400 463033 145630 463894
rect 146186 463033 146324 463909
rect 146880 463047 147039 463909
rect 147595 463047 147733 463923
rect 148289 463062 148440 463923
rect 148996 463062 149134 463938
rect 149690 463076 149849 463938
rect 150405 463076 150543 463952
rect 151099 463076 151561 463952
rect 149690 463062 151561 463076
rect 148289 463047 151561 463062
rect 146880 463033 151561 463047
rect 145400 463018 151561 463033
rect 143991 463004 151561 463018
rect 142590 462989 151561 463004
rect 141181 462975 151561 462989
rect 140742 455992 151561 462975
rect 140742 455978 149960 455992
rect 140742 455963 148551 455978
rect 140742 455949 147150 455963
rect 140742 455934 145741 455949
rect 140742 455920 144261 455934
rect 140742 455905 142852 455920
rect 140742 455891 141451 455905
rect 140742 455655 141056 455891
rect 141292 455655 141451 455891
rect 140742 455571 141451 455655
rect 140742 455335 141056 455571
rect 141292 455335 141451 455571
rect 140742 455251 141451 455335
rect 140742 455015 141056 455251
rect 141292 455029 141451 455251
rect 142007 455029 142145 455905
rect 142701 455044 142852 455905
rect 143408 455044 143546 455920
rect 144102 455058 144261 455920
rect 144817 455058 144955 455934
rect 145511 455073 145741 455934
rect 146297 455073 146435 455949
rect 146991 455087 147150 455949
rect 147706 455087 147844 455963
rect 148400 455102 148551 455963
rect 149107 455102 149245 455978
rect 149801 455116 149960 455978
rect 150516 455116 150654 455992
rect 151210 455116 151561 455992
rect 149801 455102 151561 455116
rect 148400 455087 151561 455102
rect 146991 455073 151561 455087
rect 145511 455058 151561 455073
rect 144102 455044 151561 455058
rect 142701 455029 151561 455044
rect 141292 455015 151561 455029
rect 140742 447986 151561 455015
rect 140742 447972 150033 447986
rect 140742 447957 148624 447972
rect 140742 447943 147223 447957
rect 140742 447928 145814 447943
rect 140742 447914 144334 447928
rect 140742 447899 142925 447914
rect 140742 447885 141524 447899
rect 140742 447649 141129 447885
rect 141365 447649 141524 447885
rect 140742 447565 141524 447649
rect 140742 447329 141129 447565
rect 141365 447329 141524 447565
rect 140742 447245 141524 447329
rect 140742 447009 141129 447245
rect 141365 447023 141524 447245
rect 142080 447023 142218 447899
rect 142774 447038 142925 447899
rect 143481 447038 143619 447914
rect 144175 447052 144334 447914
rect 144890 447052 145028 447928
rect 145584 447067 145814 447928
rect 146370 447067 146508 447943
rect 147064 447081 147223 447943
rect 147779 447081 147917 447957
rect 148473 447096 148624 447957
rect 149180 447096 149318 447972
rect 149874 447110 150033 447972
rect 150589 447110 150727 447986
rect 151283 447110 151561 447986
rect 149874 447096 151561 447110
rect 148473 447081 151561 447096
rect 147064 447067 151561 447081
rect 145584 447052 151561 447067
rect 144175 447038 151561 447052
rect 142774 447023 151561 447038
rect 141365 447009 151561 447023
rect 140742 440029 151561 447009
rect 140742 440015 150006 440029
rect 140742 440000 148597 440015
rect 140742 439986 147196 440000
rect 140742 439971 145787 439986
rect 140742 439957 144307 439971
rect 140742 439942 142898 439957
rect 140742 439928 141497 439942
rect 140742 439692 141102 439928
rect 141338 439692 141497 439928
rect 140742 439608 141497 439692
rect 140742 439372 141102 439608
rect 141338 439372 141497 439608
rect 140742 439288 141497 439372
rect 140742 439052 141102 439288
rect 141338 439066 141497 439288
rect 142053 439066 142191 439942
rect 142747 439081 142898 439942
rect 143454 439081 143592 439957
rect 144148 439095 144307 439957
rect 144863 439095 145001 439971
rect 145557 439110 145787 439971
rect 146343 439110 146481 439986
rect 147037 439124 147196 439986
rect 147752 439124 147890 440000
rect 148446 439139 148597 440000
rect 149153 439139 149291 440015
rect 149847 439153 150006 440015
rect 150562 439153 150700 440029
rect 151256 439153 151561 440029
rect 149847 439139 151561 439153
rect 148446 439124 151561 439139
rect 147037 439110 151561 439124
rect 145557 439095 151561 439110
rect 144148 439081 151561 439095
rect 142747 439066 151561 439081
rect 141338 439052 151561 439066
rect 140742 431939 151561 439052
rect 140742 431925 149977 431939
rect 140742 431910 148568 431925
rect 140742 431896 147167 431910
rect 140742 431881 145758 431896
rect 140742 431867 144278 431881
rect 140742 431852 142869 431867
rect 140742 431838 141468 431852
rect 140742 431602 141073 431838
rect 141309 431602 141468 431838
rect 140742 431518 141468 431602
rect 140742 431282 141073 431518
rect 141309 431282 141468 431518
rect 140742 431198 141468 431282
rect 140742 430962 141073 431198
rect 141309 430976 141468 431198
rect 142024 430976 142162 431852
rect 142718 430991 142869 431852
rect 143425 430991 143563 431867
rect 144119 431005 144278 431867
rect 144834 431005 144972 431881
rect 145528 431020 145758 431881
rect 146314 431020 146452 431896
rect 147008 431034 147167 431896
rect 147723 431034 147861 431910
rect 148417 431049 148568 431910
rect 149124 431049 149262 431925
rect 149818 431063 149977 431925
rect 150533 431063 150671 431939
rect 151227 431063 151561 431939
rect 149818 431049 151561 431063
rect 148417 431034 151561 431049
rect 147008 431020 151561 431034
rect 145528 431005 151561 431020
rect 144119 430991 151561 431005
rect 142718 430976 151561 430991
rect 141309 430962 151561 430976
rect 140742 423962 151561 430962
rect 140742 423948 150004 423962
rect 140742 423933 148595 423948
rect 140742 423919 147194 423933
rect 140742 423904 145785 423919
rect 140742 423890 144305 423904
rect 140742 423875 142896 423890
rect 140742 423861 141495 423875
rect 140742 423625 141100 423861
rect 141336 423625 141495 423861
rect 140742 423541 141495 423625
rect 140742 423305 141100 423541
rect 141336 423305 141495 423541
rect 140742 423221 141495 423305
rect 140742 422985 141100 423221
rect 141336 422999 141495 423221
rect 142051 422999 142189 423875
rect 142745 423014 142896 423875
rect 143452 423014 143590 423890
rect 144146 423028 144305 423890
rect 144861 423028 144999 423904
rect 145555 423043 145785 423904
rect 146341 423043 146479 423919
rect 147035 423057 147194 423919
rect 147750 423057 147888 423933
rect 148444 423072 148595 423933
rect 149151 423072 149289 423948
rect 149845 423086 150004 423948
rect 150560 423086 150698 423962
rect 151254 423086 151561 423962
rect 149845 423072 151561 423086
rect 148444 423057 151561 423072
rect 147035 423043 151561 423057
rect 145555 423028 151561 423043
rect 144146 423014 151561 423028
rect 142745 422999 151561 423014
rect 141336 422985 151561 422999
rect 140742 416014 151561 422985
rect 140742 416000 149939 416014
rect 140742 415985 148530 416000
rect 140742 415971 147129 415985
rect 140742 415956 145720 415971
rect 140742 415942 144240 415956
rect 140742 415927 142831 415942
rect 140742 415913 141430 415927
rect 140742 415677 141035 415913
rect 141271 415677 141430 415913
rect 140742 415593 141430 415677
rect 140742 415357 141035 415593
rect 141271 415357 141430 415593
rect 140742 415273 141430 415357
rect 140742 415037 141035 415273
rect 141271 415051 141430 415273
rect 141986 415051 142124 415927
rect 142680 415066 142831 415927
rect 143387 415066 143525 415942
rect 144081 415080 144240 415942
rect 144796 415080 144934 415956
rect 145490 415095 145720 415956
rect 146276 415095 146414 415971
rect 146970 415109 147129 415971
rect 147685 415109 147823 415985
rect 148379 415124 148530 415985
rect 149086 415124 149224 416000
rect 149780 415138 149939 416000
rect 150495 415138 150633 416014
rect 151189 415138 151561 416014
rect 149780 415124 151561 415138
rect 148379 415109 151561 415124
rect 146970 415095 151561 415109
rect 145490 415080 151561 415095
rect 144081 415066 151561 415080
rect 142680 415051 151561 415066
rect 141271 415037 151561 415051
rect 140742 407951 151561 415037
rect 140742 407937 149862 407951
rect 140742 407922 148453 407937
rect 140742 407908 147052 407922
rect 140742 407893 145643 407908
rect 140742 407879 144163 407893
rect 140742 407864 142754 407879
rect 140742 407850 141353 407864
rect 140742 407614 140958 407850
rect 141194 407614 141353 407850
rect 140742 407530 141353 407614
rect 140742 407294 140958 407530
rect 141194 407294 141353 407530
rect 140742 407210 141353 407294
rect 140742 406974 140958 407210
rect 141194 406988 141353 407210
rect 141909 406988 142047 407864
rect 142603 407003 142754 407864
rect 143310 407003 143448 407879
rect 144004 407017 144163 407879
rect 144719 407017 144857 407893
rect 145413 407032 145643 407893
rect 146199 407032 146337 407908
rect 146893 407046 147052 407908
rect 147608 407046 147746 407922
rect 148302 407061 148453 407922
rect 149009 407061 149147 407937
rect 149703 407075 149862 407937
rect 150418 407075 150556 407951
rect 151112 407075 151561 407951
rect 149703 407061 151561 407075
rect 148302 407046 151561 407061
rect 146893 407032 151561 407046
rect 145413 407017 151561 407032
rect 144004 407003 151561 407017
rect 142603 406988 151561 407003
rect 141194 406974 151561 406988
rect 140742 399947 151561 406974
rect 140742 399933 149954 399947
rect 140742 399918 148545 399933
rect 140742 399904 147144 399918
rect 140742 399889 145735 399904
rect 140742 399875 144255 399889
rect 140742 399860 142846 399875
rect 140742 399846 141445 399860
rect 140742 399610 141050 399846
rect 141286 399610 141445 399846
rect 140742 399526 141445 399610
rect 140742 399290 141050 399526
rect 141286 399290 141445 399526
rect 140742 399206 141445 399290
rect 140742 398970 141050 399206
rect 141286 398984 141445 399206
rect 142001 398984 142139 399860
rect 142695 398999 142846 399860
rect 143402 398999 143540 399875
rect 144096 399013 144255 399875
rect 144811 399013 144949 399889
rect 145505 399028 145735 399889
rect 146291 399028 146429 399904
rect 146985 399042 147144 399904
rect 147700 399042 147838 399918
rect 148394 399057 148545 399918
rect 149101 399057 149239 399933
rect 149795 399071 149954 399933
rect 150510 399071 150648 399947
rect 151204 399071 151561 399947
rect 149795 399057 151561 399071
rect 148394 399042 151561 399057
rect 146985 399028 151561 399042
rect 145505 399013 151561 399028
rect 144096 398999 151561 399013
rect 142695 398984 151561 398999
rect 141286 398970 151561 398984
rect 140742 391943 151561 398970
rect 140742 391929 149968 391943
rect 140742 391914 148559 391929
rect 140742 391900 147158 391914
rect 140742 391885 145749 391900
rect 140742 391871 144269 391885
rect 140742 391856 142860 391871
rect 140742 391842 141459 391856
rect 140742 391606 141064 391842
rect 141300 391606 141459 391842
rect 140742 391522 141459 391606
rect 140742 391286 141064 391522
rect 141300 391286 141459 391522
rect 140742 391202 141459 391286
rect 140742 390966 141064 391202
rect 141300 390980 141459 391202
rect 142015 390980 142153 391856
rect 142709 390995 142860 391856
rect 143416 390995 143554 391871
rect 144110 391009 144269 391871
rect 144825 391009 144963 391885
rect 145519 391024 145749 391885
rect 146305 391024 146443 391900
rect 146999 391038 147158 391900
rect 147714 391038 147852 391914
rect 148408 391053 148559 391914
rect 149115 391053 149253 391929
rect 149809 391067 149968 391929
rect 150524 391067 150662 391943
rect 151218 391067 151561 391943
rect 149809 391053 151561 391067
rect 148408 391038 151561 391053
rect 146999 391024 151561 391038
rect 145519 391009 151561 391024
rect 144110 390995 151561 391009
rect 142709 390980 151561 390995
rect 141300 390966 151561 390980
rect 140742 383959 151561 390966
rect 140742 383945 149973 383959
rect 140742 383930 148564 383945
rect 140742 383916 147163 383930
rect 140742 383901 145754 383916
rect 140742 383887 144274 383901
rect 140742 383872 142865 383887
rect 140742 383858 141464 383872
rect 140742 383622 141069 383858
rect 141305 383622 141464 383858
rect 140742 383538 141464 383622
rect 140742 383302 141069 383538
rect 141305 383302 141464 383538
rect 140742 383218 141464 383302
rect 140742 382982 141069 383218
rect 141305 382996 141464 383218
rect 142020 382996 142158 383872
rect 142714 383011 142865 383872
rect 143421 383011 143559 383887
rect 144115 383025 144274 383887
rect 144830 383025 144968 383901
rect 145524 383040 145754 383901
rect 146310 383040 146448 383916
rect 147004 383054 147163 383916
rect 147719 383054 147857 383930
rect 148413 383069 148564 383930
rect 149120 383069 149258 383945
rect 149814 383083 149973 383945
rect 150529 383083 150667 383959
rect 151223 383083 151561 383959
rect 149814 383069 151561 383083
rect 148413 383054 151561 383069
rect 147004 383040 151561 383054
rect 145524 383025 151561 383040
rect 144115 383011 151561 383025
rect 142714 382996 151561 383011
rect 141305 382982 151561 382996
rect 140742 375940 151561 382982
rect 140742 375926 149966 375940
rect 140742 375911 148557 375926
rect 140742 375897 147156 375911
rect 140742 375882 145747 375897
rect 140742 375868 144267 375882
rect 140742 375853 142858 375868
rect 140742 375839 141457 375853
rect 140742 375603 141062 375839
rect 141298 375603 141457 375839
rect 140742 375519 141457 375603
rect 140742 375283 141062 375519
rect 141298 375283 141457 375519
rect 140742 375199 141457 375283
rect 140742 374963 141062 375199
rect 141298 374977 141457 375199
rect 142013 374977 142151 375853
rect 142707 374992 142858 375853
rect 143414 374992 143552 375868
rect 144108 375006 144267 375868
rect 144823 375006 144961 375882
rect 145517 375021 145747 375882
rect 146303 375021 146441 375897
rect 146997 375035 147156 375897
rect 147712 375035 147850 375911
rect 148406 375050 148557 375911
rect 149113 375050 149251 375926
rect 149807 375064 149966 375926
rect 150522 375064 150660 375940
rect 151216 375064 151561 375940
rect 149807 375050 151561 375064
rect 148406 375035 151561 375050
rect 146997 375021 151561 375035
rect 145517 375006 151561 375021
rect 144108 374992 151561 375006
rect 142707 374977 151561 374992
rect 141298 374963 151561 374977
rect 140742 368001 151561 374963
rect 140742 367987 149964 368001
rect 140742 367972 148555 367987
rect 140742 367958 147154 367972
rect 140742 367943 145745 367958
rect 140742 367929 144265 367943
rect 140742 367914 142856 367929
rect 140742 367900 141455 367914
rect 140742 367664 141060 367900
rect 141296 367664 141455 367900
rect 140742 367580 141455 367664
rect 140742 367344 141060 367580
rect 141296 367344 141455 367580
rect 140742 367260 141455 367344
rect 140742 367024 141060 367260
rect 141296 367038 141455 367260
rect 142011 367038 142149 367914
rect 142705 367053 142856 367914
rect 143412 367053 143550 367929
rect 144106 367067 144265 367929
rect 144821 367067 144959 367943
rect 145515 367082 145745 367943
rect 146301 367082 146439 367958
rect 146995 367096 147154 367958
rect 147710 367096 147848 367972
rect 148404 367111 148555 367972
rect 149111 367111 149249 367987
rect 149805 367125 149964 367987
rect 150520 367125 150658 368001
rect 151214 367125 151561 368001
rect 149805 367111 151561 367125
rect 148404 367096 151561 367111
rect 146995 367082 151561 367096
rect 145515 367067 151561 367082
rect 144106 367053 151561 367067
rect 142705 367038 151561 367053
rect 141296 367024 151561 367038
rect 140742 359920 151561 367024
rect 140742 359906 149868 359920
rect 140742 359891 148459 359906
rect 140742 359877 147058 359891
rect 140742 359862 145649 359877
rect 140742 359848 144169 359862
rect 140742 359833 142760 359848
rect 140742 359819 141359 359833
rect 140742 359583 140964 359819
rect 141200 359583 141359 359819
rect 140742 359499 141359 359583
rect 140742 359263 140964 359499
rect 141200 359263 141359 359499
rect 140742 359179 141359 359263
rect 140742 358943 140964 359179
rect 141200 358957 141359 359179
rect 141915 358957 142053 359833
rect 142609 358972 142760 359833
rect 143316 358972 143454 359848
rect 144010 358986 144169 359848
rect 144725 358986 144863 359862
rect 145419 359001 145649 359862
rect 146205 359001 146343 359877
rect 146899 359015 147058 359877
rect 147614 359015 147752 359891
rect 148308 359030 148459 359891
rect 149015 359030 149153 359906
rect 149709 359044 149868 359906
rect 150424 359044 150562 359920
rect 151118 359044 151561 359920
rect 149709 359030 151561 359044
rect 148308 359015 151561 359030
rect 146899 359001 151561 359015
rect 145419 358986 151561 359001
rect 144010 358972 151561 358986
rect 142609 358957 151561 358972
rect 141200 358943 151561 358957
rect 140742 351943 151561 358943
rect 140742 351929 149946 351943
rect 140742 351914 148537 351929
rect 140742 351900 147136 351914
rect 140742 351885 145727 351900
rect 140742 351871 144247 351885
rect 140742 351856 142838 351871
rect 140742 351842 141437 351856
rect 140742 351606 141042 351842
rect 141278 351606 141437 351842
rect 140742 351522 141437 351606
rect 140742 351286 141042 351522
rect 141278 351286 141437 351522
rect 140742 351202 141437 351286
rect 140742 350966 141042 351202
rect 141278 350980 141437 351202
rect 141993 350980 142131 351856
rect 142687 350995 142838 351856
rect 143394 350995 143532 351871
rect 144088 351009 144247 351871
rect 144803 351009 144941 351885
rect 145497 351024 145727 351885
rect 146283 351024 146421 351900
rect 146977 351038 147136 351900
rect 147692 351038 147830 351914
rect 148386 351053 148537 351914
rect 149093 351053 149231 351929
rect 149787 351067 149946 351929
rect 150502 351067 150640 351943
rect 151196 351067 151561 351943
rect 149787 351053 151561 351067
rect 148386 351038 151561 351053
rect 146977 351024 151561 351038
rect 145497 351009 151561 351024
rect 144088 350995 151561 351009
rect 142687 350980 151561 350995
rect 141278 350966 151561 350980
rect 140742 343977 151561 350966
rect 407589 564959 418408 574520
rect 407589 564945 416812 564959
rect 407589 564930 415403 564945
rect 407589 564916 414002 564930
rect 407589 564901 412593 564916
rect 407589 564887 411113 564901
rect 407589 564872 409704 564887
rect 407589 564858 408303 564872
rect 407589 564622 407908 564858
rect 408144 564636 408303 564858
rect 408539 564636 408623 564872
rect 408859 564636 408997 564872
rect 409233 564636 409317 564872
rect 409553 564651 409704 564872
rect 409940 564651 410024 564887
rect 410260 564651 410398 564887
rect 410634 564651 410718 564887
rect 410954 564665 411113 564887
rect 411349 564665 411433 564901
rect 411669 564665 411807 564901
rect 412043 564665 412127 564901
rect 412363 564680 412593 564901
rect 412829 564680 412913 564916
rect 413149 564680 413287 564916
rect 413523 564680 413607 564916
rect 413843 564694 414002 564916
rect 414238 564694 414322 564930
rect 414558 564694 414696 564930
rect 414932 564694 415016 564930
rect 415252 564709 415403 564930
rect 415639 564709 415723 564945
rect 415959 564709 416097 564945
rect 416333 564709 416417 564945
rect 416653 564723 416812 564945
rect 417048 564723 417132 564959
rect 417368 564723 417506 564959
rect 417742 564723 417826 564959
rect 418062 564723 418408 564959
rect 416653 564709 418408 564723
rect 415252 564694 418408 564709
rect 413843 564680 418408 564694
rect 412363 564665 418408 564680
rect 410954 564651 418408 564665
rect 409553 564636 418408 564651
rect 408144 564622 418408 564636
rect 407589 528998 418408 564622
rect 407589 528984 416736 528998
rect 407589 528969 415327 528984
rect 407589 528955 413926 528969
rect 407589 528940 412517 528955
rect 407589 528926 411037 528940
rect 407589 528911 409628 528926
rect 407589 528897 408227 528911
rect 407589 528661 407832 528897
rect 408068 528675 408227 528897
rect 408463 528675 408547 528911
rect 408783 528675 408921 528911
rect 409157 528675 409241 528911
rect 409477 528690 409628 528911
rect 409864 528690 409948 528926
rect 410184 528690 410322 528926
rect 410558 528690 410642 528926
rect 410878 528704 411037 528926
rect 411273 528704 411357 528940
rect 411593 528704 411731 528940
rect 411967 528704 412051 528940
rect 412287 528719 412517 528940
rect 412753 528719 412837 528955
rect 413073 528719 413211 528955
rect 413447 528719 413531 528955
rect 413767 528733 413926 528955
rect 414162 528733 414246 528969
rect 414482 528733 414620 528969
rect 414856 528733 414940 528969
rect 415176 528748 415327 528969
rect 415563 528748 415647 528984
rect 415883 528748 416021 528984
rect 416257 528748 416341 528984
rect 416577 528762 416736 528984
rect 416972 528762 417056 528998
rect 417292 528762 417430 528998
rect 417666 528762 417750 528998
rect 417986 528762 418408 528998
rect 416577 528748 418408 528762
rect 415176 528733 418408 528748
rect 413767 528719 418408 528733
rect 412287 528704 418408 528719
rect 410878 528690 418408 528704
rect 409477 528675 418408 528690
rect 408068 528661 418408 528675
rect 407589 492971 418408 528661
rect 407589 492957 416716 492971
rect 407589 492942 415307 492957
rect 407589 492928 413906 492942
rect 407589 492913 412497 492928
rect 407589 492899 411017 492913
rect 407589 492884 409608 492899
rect 407589 492870 408207 492884
rect 407589 492634 407812 492870
rect 408048 492648 408207 492870
rect 408443 492648 408527 492884
rect 408763 492648 408901 492884
rect 409137 492648 409221 492884
rect 409457 492663 409608 492884
rect 409844 492663 409928 492899
rect 410164 492663 410302 492899
rect 410538 492663 410622 492899
rect 410858 492677 411017 492899
rect 411253 492677 411337 492913
rect 411573 492677 411711 492913
rect 411947 492677 412031 492913
rect 412267 492692 412497 492913
rect 412733 492692 412817 492928
rect 413053 492692 413191 492928
rect 413427 492692 413511 492928
rect 413747 492706 413906 492928
rect 414142 492706 414226 492942
rect 414462 492706 414600 492942
rect 414836 492706 414920 492942
rect 415156 492721 415307 492942
rect 415543 492721 415627 492957
rect 415863 492721 416001 492957
rect 416237 492721 416321 492957
rect 416557 492735 416716 492957
rect 416952 492735 417036 492971
rect 417272 492735 417410 492971
rect 417646 492735 417730 492971
rect 417966 492735 418408 492971
rect 416557 492721 418408 492735
rect 415156 492706 418408 492721
rect 413747 492692 418408 492706
rect 412267 492677 418408 492692
rect 410858 492663 418408 492677
rect 409457 492648 418408 492663
rect 408048 492634 418408 492648
rect 407589 469622 418408 492634
rect 407589 469608 416810 469622
rect 407589 469593 415401 469608
rect 407589 469579 414000 469593
rect 407589 469564 412591 469579
rect 407589 469550 411111 469564
rect 407589 469535 409702 469550
rect 407589 469521 408301 469535
rect 407589 469285 407906 469521
rect 408142 469285 408301 469521
rect 407589 469201 408301 469285
rect 407589 468965 407906 469201
rect 408142 468965 408301 469201
rect 407589 468881 408301 468965
rect 407589 468645 407906 468881
rect 408142 468659 408301 468881
rect 408857 468659 408995 469535
rect 409551 468674 409702 469535
rect 410258 468674 410396 469550
rect 410952 468688 411111 469550
rect 411667 468688 411805 469564
rect 412361 468703 412591 469564
rect 413147 468703 413285 469579
rect 413841 468717 414000 469579
rect 414556 468717 414694 469593
rect 415250 468732 415401 469593
rect 415957 468732 416095 469608
rect 416651 468746 416810 469608
rect 417366 468746 417504 469622
rect 418060 468746 418408 469622
rect 416651 468732 418408 468746
rect 415250 468717 418408 468732
rect 413841 468703 418408 468717
rect 412361 468688 418408 468703
rect 410952 468674 418408 468688
rect 409551 468659 418408 468674
rect 408142 468645 418408 468659
rect 407589 461619 418408 468645
rect 407589 461605 416813 461619
rect 407589 461590 415404 461605
rect 407589 461576 414003 461590
rect 407589 461561 412594 461576
rect 407589 461547 411114 461561
rect 407589 461532 409705 461547
rect 407589 461518 408304 461532
rect 407589 461282 407909 461518
rect 408145 461282 408304 461518
rect 407589 461198 408304 461282
rect 407589 460962 407909 461198
rect 408145 460962 408304 461198
rect 407589 460878 408304 460962
rect 407589 460642 407909 460878
rect 408145 460656 408304 460878
rect 408860 460656 408998 461532
rect 409554 460671 409705 461532
rect 410261 460671 410399 461547
rect 410955 460685 411114 461547
rect 411670 460685 411808 461561
rect 412364 460700 412594 461561
rect 413150 460700 413288 461576
rect 413844 460714 414003 461576
rect 414559 460714 414697 461590
rect 415253 460729 415404 461590
rect 415960 460729 416098 461605
rect 416654 460743 416813 461605
rect 417369 460743 417507 461619
rect 418063 460743 418408 461619
rect 416654 460729 418408 460743
rect 415253 460714 418408 460729
rect 413844 460700 418408 460714
rect 412364 460685 418408 460700
rect 410955 460671 418408 460685
rect 409554 460656 418408 460671
rect 408145 460642 418408 460656
rect 407589 453623 418408 460642
rect 407589 453609 416772 453623
rect 407589 453594 415363 453609
rect 407589 453580 413962 453594
rect 407589 453565 412553 453580
rect 407589 453551 411073 453565
rect 407589 453536 409664 453551
rect 407589 453522 408263 453536
rect 407589 453286 407868 453522
rect 408104 453286 408263 453522
rect 407589 453202 408263 453286
rect 407589 452966 407868 453202
rect 408104 452966 408263 453202
rect 407589 452882 408263 452966
rect 407589 452646 407868 452882
rect 408104 452660 408263 452882
rect 408819 452660 408957 453536
rect 409513 452675 409664 453536
rect 410220 452675 410358 453551
rect 410914 452689 411073 453551
rect 411629 452689 411767 453565
rect 412323 452704 412553 453565
rect 413109 452704 413247 453580
rect 413803 452718 413962 453580
rect 414518 452718 414656 453594
rect 415212 452733 415363 453594
rect 415919 452733 416057 453609
rect 416613 452747 416772 453609
rect 417328 452747 417466 453623
rect 418022 452747 418408 453623
rect 416613 452733 418408 452747
rect 415212 452718 418408 452733
rect 413803 452704 418408 452718
rect 412323 452689 418408 452704
rect 410914 452675 418408 452689
rect 409513 452660 418408 452675
rect 408104 452646 418408 452660
rect 407589 445614 418408 452646
rect 407589 445600 416763 445614
rect 407589 445585 415354 445600
rect 407589 445571 413953 445585
rect 407589 445556 412544 445571
rect 407589 445542 411064 445556
rect 407589 445527 409655 445542
rect 407589 445513 408254 445527
rect 407589 445277 407859 445513
rect 408095 445277 408254 445513
rect 407589 445193 408254 445277
rect 407589 444957 407859 445193
rect 408095 444957 408254 445193
rect 407589 444873 408254 444957
rect 407589 444637 407859 444873
rect 408095 444651 408254 444873
rect 408810 444651 408948 445527
rect 409504 444666 409655 445527
rect 410211 444666 410349 445542
rect 410905 444680 411064 445542
rect 411620 444680 411758 445556
rect 412314 444695 412544 445556
rect 413100 444695 413238 445571
rect 413794 444709 413953 445571
rect 414509 444709 414647 445585
rect 415203 444724 415354 445585
rect 415910 444724 416048 445600
rect 416604 444738 416763 445600
rect 417319 444738 417457 445614
rect 418013 444738 418408 445614
rect 416604 444724 418408 444738
rect 415203 444709 418408 444724
rect 413794 444695 418408 444709
rect 412314 444680 418408 444695
rect 410905 444666 418408 444680
rect 409504 444651 418408 444666
rect 408095 444637 418408 444651
rect 407589 437628 418408 444637
rect 407589 437614 416736 437628
rect 407589 437599 415327 437614
rect 407589 437585 413926 437599
rect 407589 437570 412517 437585
rect 407589 437556 411037 437570
rect 407589 437541 409628 437556
rect 407589 437527 408227 437541
rect 407589 437291 407832 437527
rect 408068 437291 408227 437527
rect 407589 437207 408227 437291
rect 407589 436971 407832 437207
rect 408068 436971 408227 437207
rect 407589 436887 408227 436971
rect 407589 436651 407832 436887
rect 408068 436665 408227 436887
rect 408783 436665 408921 437541
rect 409477 436680 409628 437541
rect 410184 436680 410322 437556
rect 410878 436694 411037 437556
rect 411593 436694 411731 437570
rect 412287 436709 412517 437570
rect 413073 436709 413211 437585
rect 413767 436723 413926 437585
rect 414482 436723 414620 437599
rect 415176 436738 415327 437599
rect 415883 436738 416021 437614
rect 416577 436752 416736 437614
rect 417292 436752 417430 437628
rect 417986 436752 418408 437628
rect 416577 436738 418408 436752
rect 415176 436723 418408 436738
rect 413767 436709 418408 436723
rect 412287 436694 418408 436709
rect 410878 436680 418408 436694
rect 409477 436665 418408 436680
rect 408068 436651 418408 436665
rect 407589 429597 418408 436651
rect 407589 429583 416760 429597
rect 407589 429568 415351 429583
rect 407589 429554 413950 429568
rect 407589 429539 412541 429554
rect 407589 429525 411061 429539
rect 407589 429510 409652 429525
rect 407589 429496 408251 429510
rect 407589 429260 407856 429496
rect 408092 429260 408251 429496
rect 407589 429176 408251 429260
rect 407589 428940 407856 429176
rect 408092 428940 408251 429176
rect 407589 428856 408251 428940
rect 407589 428620 407856 428856
rect 408092 428634 408251 428856
rect 408807 428634 408945 429510
rect 409501 428649 409652 429510
rect 410208 428649 410346 429525
rect 410902 428663 411061 429525
rect 411617 428663 411755 429539
rect 412311 428678 412541 429539
rect 413097 428678 413235 429554
rect 413791 428692 413950 429554
rect 414506 428692 414644 429568
rect 415200 428707 415351 429568
rect 415907 428707 416045 429583
rect 416601 428721 416760 429583
rect 417316 428721 417454 429597
rect 418010 428721 418408 429597
rect 416601 428707 418408 428721
rect 415200 428692 418408 428707
rect 413791 428678 418408 428692
rect 412311 428663 418408 428678
rect 410902 428649 418408 428663
rect 409501 428634 418408 428649
rect 408092 428620 418408 428634
rect 407589 421666 418408 428620
rect 407589 421652 416822 421666
rect 407589 421637 415413 421652
rect 407589 421623 414012 421637
rect 407589 421608 412603 421623
rect 407589 421594 411123 421608
rect 407589 421579 409714 421594
rect 407589 421565 408313 421579
rect 407589 421329 407918 421565
rect 408154 421329 408313 421565
rect 407589 421245 408313 421329
rect 407589 421009 407918 421245
rect 408154 421009 408313 421245
rect 407589 420925 408313 421009
rect 407589 420689 407918 420925
rect 408154 420703 408313 420925
rect 408869 420703 409007 421579
rect 409563 420718 409714 421579
rect 410270 420718 410408 421594
rect 410964 420732 411123 421594
rect 411679 420732 411817 421608
rect 412373 420747 412603 421608
rect 413159 420747 413297 421623
rect 413853 420761 414012 421623
rect 414568 420761 414706 421637
rect 415262 420776 415413 421637
rect 415969 420776 416107 421652
rect 416663 420790 416822 421652
rect 417378 420790 417516 421666
rect 418072 420790 418408 421666
rect 416663 420776 418408 420790
rect 415262 420761 418408 420776
rect 413853 420747 418408 420761
rect 412373 420732 418408 420747
rect 410964 420718 418408 420732
rect 409563 420703 418408 420718
rect 408154 420689 418408 420703
rect 407589 413636 418408 420689
rect 407589 413622 416838 413636
rect 407589 413607 415429 413622
rect 407589 413593 414028 413607
rect 407589 413578 412619 413593
rect 407589 413564 411139 413578
rect 407589 413549 409730 413564
rect 407589 413535 408329 413549
rect 407589 413299 407934 413535
rect 408170 413299 408329 413535
rect 407589 413215 408329 413299
rect 407589 412979 407934 413215
rect 408170 412979 408329 413215
rect 407589 412895 408329 412979
rect 407589 412659 407934 412895
rect 408170 412673 408329 412895
rect 408885 412673 409023 413549
rect 409579 412688 409730 413549
rect 410286 412688 410424 413564
rect 410980 412702 411139 413564
rect 411695 412702 411833 413578
rect 412389 412717 412619 413578
rect 413175 412717 413313 413593
rect 413869 412731 414028 413593
rect 414584 412731 414722 413607
rect 415278 412746 415429 413607
rect 415985 412746 416123 413622
rect 416679 412760 416838 413622
rect 417394 412760 417532 413636
rect 418088 412760 418408 413636
rect 416679 412746 418408 412760
rect 415278 412731 418408 412746
rect 413869 412717 418408 412731
rect 412389 412702 418408 412717
rect 410980 412688 418408 412702
rect 409579 412673 418408 412688
rect 408170 412659 418408 412673
rect 407589 405628 418408 412659
rect 407589 405614 416812 405628
rect 407589 405599 415403 405614
rect 407589 405585 414002 405599
rect 407589 405570 412593 405585
rect 407589 405556 411113 405570
rect 407589 405541 409704 405556
rect 407589 405527 408303 405541
rect 407589 405291 407908 405527
rect 408144 405291 408303 405527
rect 407589 405207 408303 405291
rect 407589 404971 407908 405207
rect 408144 404971 408303 405207
rect 407589 404887 408303 404971
rect 407589 404651 407908 404887
rect 408144 404665 408303 404887
rect 408859 404665 408997 405541
rect 409553 404680 409704 405541
rect 410260 404680 410398 405556
rect 410954 404694 411113 405556
rect 411669 404694 411807 405570
rect 412363 404709 412593 405570
rect 413149 404709 413287 405585
rect 413843 404723 414002 405585
rect 414558 404723 414696 405599
rect 415252 404738 415403 405599
rect 415959 404738 416097 405614
rect 416653 404752 416812 405614
rect 417368 404752 417506 405628
rect 418062 404752 418408 405628
rect 416653 404738 418408 404752
rect 415252 404723 418408 404738
rect 413843 404709 418408 404723
rect 412363 404694 418408 404709
rect 410954 404680 418408 404694
rect 409553 404665 418408 404680
rect 408144 404651 418408 404665
rect 407589 397609 418408 404651
rect 407589 397595 416786 397609
rect 407589 397580 415377 397595
rect 407589 397566 413976 397580
rect 407589 397551 412567 397566
rect 407589 397537 411087 397551
rect 407589 397522 409678 397537
rect 407589 397508 408277 397522
rect 407589 397272 407882 397508
rect 408118 397272 408277 397508
rect 407589 397188 408277 397272
rect 407589 396952 407882 397188
rect 408118 396952 408277 397188
rect 407589 396868 408277 396952
rect 407589 396632 407882 396868
rect 408118 396646 408277 396868
rect 408833 396646 408971 397522
rect 409527 396661 409678 397522
rect 410234 396661 410372 397537
rect 410928 396675 411087 397537
rect 411643 396675 411781 397551
rect 412337 396690 412567 397551
rect 413123 396690 413261 397566
rect 413817 396704 413976 397566
rect 414532 396704 414670 397580
rect 415226 396719 415377 397580
rect 415933 396719 416071 397595
rect 416627 396733 416786 397595
rect 417342 396733 417480 397609
rect 418036 396733 418408 397609
rect 416627 396719 418408 396733
rect 415226 396704 418408 396719
rect 413817 396690 418408 396704
rect 412337 396675 418408 396690
rect 410928 396661 418408 396675
rect 409527 396646 418408 396661
rect 408118 396632 418408 396646
rect 407589 389606 418408 396632
rect 407589 389592 416877 389606
rect 407589 389577 415468 389592
rect 407589 389563 414067 389577
rect 407589 389548 412658 389563
rect 407589 389534 411178 389548
rect 407589 389519 409769 389534
rect 407589 389505 408368 389519
rect 407589 389269 407973 389505
rect 408209 389269 408368 389505
rect 407589 389185 408368 389269
rect 407589 388949 407973 389185
rect 408209 388949 408368 389185
rect 407589 388865 408368 388949
rect 407589 388629 407973 388865
rect 408209 388643 408368 388865
rect 408924 388643 409062 389519
rect 409618 388658 409769 389519
rect 410325 388658 410463 389534
rect 411019 388672 411178 389534
rect 411734 388672 411872 389548
rect 412428 388687 412658 389548
rect 413214 388687 413352 389563
rect 413908 388701 414067 389563
rect 414623 388701 414761 389577
rect 415317 388716 415468 389577
rect 416024 388716 416162 389592
rect 416718 388730 416877 389592
rect 417433 388730 417571 389606
rect 418127 388730 418408 389606
rect 416718 388716 418408 388730
rect 415317 388701 418408 388716
rect 413908 388687 418408 388701
rect 412428 388672 418408 388687
rect 411019 388658 418408 388672
rect 409618 388643 418408 388658
rect 408209 388629 418408 388643
rect 407589 381655 418408 388629
rect 407589 381641 416798 381655
rect 407589 381626 415389 381641
rect 407589 381612 413988 381626
rect 407589 381597 412579 381612
rect 407589 381583 411099 381597
rect 407589 381568 409690 381583
rect 407589 381554 408289 381568
rect 407589 381318 407894 381554
rect 408130 381318 408289 381554
rect 407589 381234 408289 381318
rect 407589 380998 407894 381234
rect 408130 380998 408289 381234
rect 407589 380914 408289 380998
rect 407589 380678 407894 380914
rect 408130 380692 408289 380914
rect 408845 380692 408983 381568
rect 409539 380707 409690 381568
rect 410246 380707 410384 381583
rect 410940 380721 411099 381583
rect 411655 380721 411793 381597
rect 412349 380736 412579 381597
rect 413135 380736 413273 381612
rect 413829 380750 413988 381612
rect 414544 380750 414682 381626
rect 415238 380765 415389 381626
rect 415945 380765 416083 381641
rect 416639 380779 416798 381641
rect 417354 380779 417492 381655
rect 418048 380779 418408 381655
rect 416639 380765 418408 380779
rect 415238 380750 418408 380765
rect 413829 380736 418408 380750
rect 412349 380721 418408 380736
rect 410940 380707 418408 380721
rect 409539 380692 418408 380707
rect 408130 380678 418408 380692
rect 407589 373627 418408 380678
rect 407589 373613 416789 373627
rect 407589 373598 415380 373613
rect 407589 373584 413979 373598
rect 407589 373569 412570 373584
rect 407589 373555 411090 373569
rect 407589 373540 409681 373555
rect 407589 373526 408280 373540
rect 407589 373290 407885 373526
rect 408121 373290 408280 373526
rect 407589 373206 408280 373290
rect 407589 372970 407885 373206
rect 408121 372970 408280 373206
rect 407589 372886 408280 372970
rect 407589 372650 407885 372886
rect 408121 372664 408280 372886
rect 408836 372664 408974 373540
rect 409530 372679 409681 373540
rect 410237 372679 410375 373555
rect 410931 372693 411090 373555
rect 411646 372693 411784 373569
rect 412340 372708 412570 373569
rect 413126 372708 413264 373584
rect 413820 372722 413979 373584
rect 414535 372722 414673 373598
rect 415229 372737 415380 373598
rect 415936 372737 416074 373613
rect 416630 372751 416789 373613
rect 417345 372751 417483 373627
rect 418039 372751 418408 373627
rect 416630 372737 418408 372751
rect 415229 372722 418408 372737
rect 413820 372708 418408 372722
rect 412340 372693 418408 372708
rect 410931 372679 418408 372693
rect 409530 372664 418408 372679
rect 408121 372650 418408 372664
rect 407589 365636 418408 372650
rect 407589 365622 416781 365636
rect 407589 365607 415372 365622
rect 407589 365593 413971 365607
rect 407589 365578 412562 365593
rect 407589 365564 411082 365578
rect 407589 365549 409673 365564
rect 407589 365535 408272 365549
rect 407589 365299 407877 365535
rect 408113 365299 408272 365535
rect 407589 365215 408272 365299
rect 407589 364979 407877 365215
rect 408113 364979 408272 365215
rect 407589 364895 408272 364979
rect 407589 364659 407877 364895
rect 408113 364673 408272 364895
rect 408828 364673 408966 365549
rect 409522 364688 409673 365549
rect 410229 364688 410367 365564
rect 410923 364702 411082 365564
rect 411638 364702 411776 365578
rect 412332 364717 412562 365578
rect 413118 364717 413256 365593
rect 413812 364731 413971 365593
rect 414527 364731 414665 365607
rect 415221 364746 415372 365607
rect 415928 364746 416066 365622
rect 416622 364760 416781 365622
rect 417337 364760 417475 365636
rect 418031 364760 418408 365636
rect 416622 364746 418408 364760
rect 415221 364731 418408 364746
rect 413812 364717 418408 364731
rect 412332 364702 418408 364717
rect 410923 364688 418408 364702
rect 409522 364673 418408 364688
rect 408113 364659 418408 364673
rect 407589 357646 418408 364659
rect 407589 357632 416718 357646
rect 407589 357617 415309 357632
rect 407589 357603 413908 357617
rect 407589 357588 412499 357603
rect 407589 357574 411019 357588
rect 407589 357559 409610 357574
rect 407589 357545 408209 357559
rect 407589 357309 407814 357545
rect 408050 357309 408209 357545
rect 407589 357225 408209 357309
rect 407589 356989 407814 357225
rect 408050 356989 408209 357225
rect 407589 356905 408209 356989
rect 407589 356669 407814 356905
rect 408050 356683 408209 356905
rect 408765 356683 408903 357559
rect 409459 356698 409610 357559
rect 410166 356698 410304 357574
rect 410860 356712 411019 357574
rect 411575 356712 411713 357588
rect 412269 356727 412499 357588
rect 413055 356727 413193 357603
rect 413749 356741 413908 357603
rect 414464 356741 414602 357617
rect 415158 356756 415309 357617
rect 415865 356756 416003 357632
rect 416559 356770 416718 357632
rect 417274 356770 417412 357646
rect 417968 356770 418408 357646
rect 416559 356756 418408 356770
rect 415158 356741 418408 356756
rect 413749 356727 418408 356741
rect 412269 356712 418408 356727
rect 410860 356698 418408 356712
rect 409459 356683 418408 356698
rect 408050 356669 418408 356683
rect 407589 349633 418408 356669
rect 407589 349619 416805 349633
rect 407589 349604 415396 349619
rect 407589 349590 413995 349604
rect 407589 349575 412586 349590
rect 407589 349561 411106 349575
rect 407589 349546 409697 349561
rect 407589 349532 408296 349546
rect 407589 349296 407901 349532
rect 408137 349296 408296 349532
rect 407589 349212 408296 349296
rect 407589 348976 407901 349212
rect 408137 348976 408296 349212
rect 407589 348892 408296 348976
rect 407589 348656 407901 348892
rect 408137 348670 408296 348892
rect 408852 348670 408990 349546
rect 409546 348685 409697 349546
rect 410253 348685 410391 349561
rect 410947 348699 411106 349561
rect 411662 348699 411800 349575
rect 412356 348714 412586 349575
rect 413142 348714 413280 349590
rect 413836 348728 413995 349590
rect 414551 348728 414689 349604
rect 415245 348743 415396 349604
rect 415952 348743 416090 349619
rect 416646 348757 416805 349619
rect 417361 348757 417499 349633
rect 418055 348757 418408 349633
rect 416646 348743 418408 348757
rect 415245 348728 418408 348743
rect 413836 348714 418408 348728
rect 412356 348699 418408 348714
rect 410947 348685 418408 348699
rect 409546 348670 418408 348685
rect 408137 348656 418408 348670
rect 389771 344452 389837 344453
rect 389771 344388 389772 344452
rect 389836 344388 389837 344452
rect 389771 344387 389837 344388
rect 140742 343963 150021 343977
rect 140742 343948 148612 343963
rect 140742 343934 147211 343948
rect 140742 343919 145802 343934
rect 140742 343905 144322 343919
rect 140742 343890 142913 343905
rect 140742 343876 141512 343890
rect 140742 343640 141117 343876
rect 141353 343640 141512 343876
rect 140742 343556 141512 343640
rect 140742 343320 141117 343556
rect 141353 343320 141512 343556
rect 140742 343236 141512 343320
rect 140742 343000 141117 343236
rect 141353 343014 141512 343236
rect 142068 343014 142206 343890
rect 142762 343029 142913 343890
rect 143469 343029 143607 343905
rect 144163 343043 144322 343905
rect 144878 343043 145016 343919
rect 145572 343058 145802 343919
rect 146358 343058 146496 343934
rect 147052 343072 147211 343934
rect 147767 343072 147905 343948
rect 148461 343087 148612 343948
rect 149168 343087 149306 343963
rect 149862 343101 150021 343963
rect 150577 343101 150715 343977
rect 151271 343101 151561 343977
rect 149862 343087 151561 343101
rect 148461 343072 151561 343087
rect 147052 343058 151561 343072
rect 145572 343043 151561 343058
rect 144163 343029 151561 343043
rect 142762 343014 151561 343029
rect 141353 343000 151561 343014
rect 140742 327368 151561 343000
rect 140742 327354 150048 327368
rect 140742 327339 148639 327354
rect 140742 327325 147238 327339
rect 140742 327310 145829 327325
rect 140742 327296 144349 327310
rect 140742 327281 142940 327296
rect 140742 327267 141539 327281
rect 140742 327031 141144 327267
rect 141380 327045 141539 327267
rect 141775 327045 141859 327281
rect 142095 327045 142233 327281
rect 142469 327045 142553 327281
rect 142789 327060 142940 327281
rect 143176 327060 143260 327296
rect 143496 327060 143634 327296
rect 143870 327060 143954 327296
rect 144190 327074 144349 327296
rect 144585 327074 144669 327310
rect 144905 327074 145043 327310
rect 145279 327074 145363 327310
rect 145599 327089 145829 327310
rect 146065 327089 146149 327325
rect 146385 327089 146523 327325
rect 146759 327089 146843 327325
rect 147079 327103 147238 327325
rect 147474 327103 147558 327339
rect 147794 327103 147932 327339
rect 148168 327103 148252 327339
rect 148488 327118 148639 327339
rect 148875 327118 148959 327354
rect 149195 327118 149333 327354
rect 149569 327118 149653 327354
rect 149889 327132 150048 327354
rect 150284 327132 150368 327368
rect 150604 327132 150742 327368
rect 150978 327132 151062 327368
rect 151298 327132 151561 327368
rect 149889 327118 151561 327132
rect 148488 327103 151561 327118
rect 147079 327089 151561 327103
rect 145599 327074 151561 327089
rect 144190 327060 151561 327074
rect 142789 327045 151561 327060
rect 141380 327031 151561 327045
rect 140742 291335 151561 327031
rect 140742 291321 149921 291335
rect 140742 291306 148512 291321
rect 140742 291292 147111 291306
rect 140742 291277 145702 291292
rect 140742 291263 144222 291277
rect 140742 291248 142813 291263
rect 140742 291234 141412 291248
rect 140742 290998 141017 291234
rect 141253 291012 141412 291234
rect 141648 291012 141732 291248
rect 141968 291012 142106 291248
rect 142342 291012 142426 291248
rect 142662 291027 142813 291248
rect 143049 291027 143133 291263
rect 143369 291027 143507 291263
rect 143743 291027 143827 291263
rect 144063 291041 144222 291263
rect 144458 291041 144542 291277
rect 144778 291041 144916 291277
rect 145152 291041 145236 291277
rect 145472 291056 145702 291277
rect 145938 291056 146022 291292
rect 146258 291056 146396 291292
rect 146632 291056 146716 291292
rect 146952 291070 147111 291292
rect 147347 291070 147431 291306
rect 147667 291070 147805 291306
rect 148041 291070 148125 291306
rect 148361 291085 148512 291306
rect 148748 291085 148832 291321
rect 149068 291085 149206 291321
rect 149442 291085 149526 291321
rect 149762 291099 149921 291321
rect 150157 291099 150241 291335
rect 150477 291099 150615 291335
rect 150851 291099 150935 291335
rect 151171 291099 151561 291335
rect 149762 291085 151561 291099
rect 148361 291070 151561 291085
rect 146952 291056 151561 291070
rect 145472 291041 151561 291056
rect 144063 291027 151561 291041
rect 142662 291012 151561 291027
rect 141253 290998 151561 291012
rect 140742 255325 151561 290998
rect 140742 255311 149949 255325
rect 140742 255296 148540 255311
rect 140742 255282 147139 255296
rect 140742 255267 145730 255282
rect 140742 255253 144250 255267
rect 140742 255238 142841 255253
rect 140742 255224 141440 255238
rect 140742 254988 141045 255224
rect 141281 255002 141440 255224
rect 141676 255002 141760 255238
rect 141996 255002 142134 255238
rect 142370 255002 142454 255238
rect 142690 255017 142841 255238
rect 143077 255017 143161 255253
rect 143397 255017 143535 255253
rect 143771 255017 143855 255253
rect 144091 255031 144250 255253
rect 144486 255031 144570 255267
rect 144806 255031 144944 255267
rect 145180 255031 145264 255267
rect 145500 255046 145730 255267
rect 145966 255046 146050 255282
rect 146286 255046 146424 255282
rect 146660 255046 146744 255282
rect 146980 255060 147139 255282
rect 147375 255060 147459 255296
rect 147695 255060 147833 255296
rect 148069 255060 148153 255296
rect 148389 255075 148540 255296
rect 148776 255075 148860 255311
rect 149096 255075 149234 255311
rect 149470 255075 149554 255311
rect 149790 255089 149949 255311
rect 150185 255089 150269 255325
rect 150505 255089 150643 255325
rect 150879 255089 150963 255325
rect 151199 255089 151561 255325
rect 149790 255075 151561 255089
rect 148389 255060 151561 255075
rect 146980 255046 151561 255060
rect 145500 255031 151561 255046
rect 144091 255017 151561 255031
rect 142690 255002 151561 255017
rect 141281 254988 151561 255002
rect 140742 236000 151561 254988
rect 102604 212018 102786 212254
rect 103022 212018 103204 212254
rect 102604 211934 103204 212018
rect 102604 211698 102786 211934
rect 103022 211698 103204 211934
rect 102604 176254 103204 211698
rect 102604 176018 102786 176254
rect 103022 176018 103204 176254
rect 102604 175934 103204 176018
rect 102604 175698 102786 175934
rect 103022 175698 103204 175934
rect 102604 140254 103204 175698
rect 102604 140018 102786 140254
rect 103022 140018 103204 140254
rect 102604 139934 103204 140018
rect 102604 139698 102786 139934
rect 103022 139698 103204 139934
rect 102604 104254 103204 139698
rect 102604 104018 102786 104254
rect 103022 104018 103204 104254
rect 102604 103934 103204 104018
rect 102604 103698 102786 103934
rect 103022 103698 103204 103934
rect 102604 68254 103204 103698
rect 102604 68018 102786 68254
rect 103022 68018 103204 68254
rect 102604 67934 103204 68018
rect 102604 67698 102786 67934
rect 103022 67698 103204 67934
rect 102604 32254 103204 67698
rect 102604 32018 102786 32254
rect 103022 32018 103204 32254
rect 102604 31934 103204 32018
rect 102604 31698 102786 31934
rect 103022 31698 103204 31934
rect 84604 -6222 84786 -5986
rect 85022 -6222 85204 -5986
rect 84604 -6306 85204 -6222
rect 84604 -6542 84786 -6306
rect 85022 -6542 85204 -6306
rect 84604 -7504 85204 -6542
rect 102604 -6926 103204 31698
rect 109804 183454 110404 218000
rect 109804 183218 109986 183454
rect 110222 183218 110404 183454
rect 109804 183134 110404 183218
rect 109804 182898 109986 183134
rect 110222 182898 110404 183134
rect 109804 147454 110404 182898
rect 109804 147218 109986 147454
rect 110222 147218 110404 147454
rect 109804 147134 110404 147218
rect 109804 146898 109986 147134
rect 110222 146898 110404 147134
rect 109804 111454 110404 146898
rect 109804 111218 109986 111454
rect 110222 111218 110404 111454
rect 109804 111134 110404 111218
rect 109804 110898 109986 111134
rect 110222 110898 110404 111134
rect 109804 75454 110404 110898
rect 109804 75218 109986 75454
rect 110222 75218 110404 75454
rect 109804 75134 110404 75218
rect 109804 74898 109986 75134
rect 110222 74898 110404 75134
rect 109804 39454 110404 74898
rect 109804 39218 109986 39454
rect 110222 39218 110404 39454
rect 109804 39134 110404 39218
rect 109804 38898 109986 39134
rect 110222 38898 110404 39134
rect 109804 3454 110404 38898
rect 109804 3218 109986 3454
rect 110222 3218 110404 3454
rect 109804 3134 110404 3218
rect 109804 2898 109986 3134
rect 110222 2898 110404 3134
rect 109804 -346 110404 2898
rect 109804 -582 109986 -346
rect 110222 -582 110404 -346
rect 109804 -666 110404 -582
rect 109804 -902 109986 -666
rect 110222 -902 110404 -666
rect 109804 -1864 110404 -902
rect 113404 187054 114004 218000
rect 113404 186818 113586 187054
rect 113822 186818 114004 187054
rect 113404 186734 114004 186818
rect 113404 186498 113586 186734
rect 113822 186498 114004 186734
rect 113404 151054 114004 186498
rect 113404 150818 113586 151054
rect 113822 150818 114004 151054
rect 113404 150734 114004 150818
rect 113404 150498 113586 150734
rect 113822 150498 114004 150734
rect 113404 115054 114004 150498
rect 113404 114818 113586 115054
rect 113822 114818 114004 115054
rect 113404 114734 114004 114818
rect 113404 114498 113586 114734
rect 113822 114498 114004 114734
rect 113404 79054 114004 114498
rect 113404 78818 113586 79054
rect 113822 78818 114004 79054
rect 113404 78734 114004 78818
rect 113404 78498 113586 78734
rect 113822 78498 114004 78734
rect 113404 43054 114004 78498
rect 113404 42818 113586 43054
rect 113822 42818 114004 43054
rect 113404 42734 114004 42818
rect 113404 42498 113586 42734
rect 113822 42498 114004 42734
rect 113404 7054 114004 42498
rect 113404 6818 113586 7054
rect 113822 6818 114004 7054
rect 113404 6734 114004 6818
rect 113404 6498 113586 6734
rect 113822 6498 114004 6734
rect 113404 -2226 114004 6498
rect 113404 -2462 113586 -2226
rect 113822 -2462 114004 -2226
rect 113404 -2546 114004 -2462
rect 113404 -2782 113586 -2546
rect 113822 -2782 114004 -2546
rect 113404 -3744 114004 -2782
rect 117004 190654 117604 218000
rect 117004 190418 117186 190654
rect 117422 190418 117604 190654
rect 117004 190334 117604 190418
rect 117004 190098 117186 190334
rect 117422 190098 117604 190334
rect 117004 154654 117604 190098
rect 117004 154418 117186 154654
rect 117422 154418 117604 154654
rect 117004 154334 117604 154418
rect 117004 154098 117186 154334
rect 117422 154098 117604 154334
rect 117004 118654 117604 154098
rect 117004 118418 117186 118654
rect 117422 118418 117604 118654
rect 117004 118334 117604 118418
rect 117004 118098 117186 118334
rect 117422 118098 117604 118334
rect 117004 82654 117604 118098
rect 117004 82418 117186 82654
rect 117422 82418 117604 82654
rect 117004 82334 117604 82418
rect 117004 82098 117186 82334
rect 117422 82098 117604 82334
rect 117004 46654 117604 82098
rect 117004 46418 117186 46654
rect 117422 46418 117604 46654
rect 117004 46334 117604 46418
rect 117004 46098 117186 46334
rect 117422 46098 117604 46334
rect 117004 10654 117604 46098
rect 117004 10418 117186 10654
rect 117422 10418 117604 10654
rect 117004 10334 117604 10418
rect 117004 10098 117186 10334
rect 117422 10098 117604 10334
rect 117004 -4106 117604 10098
rect 117004 -4342 117186 -4106
rect 117422 -4342 117604 -4106
rect 117004 -4426 117604 -4342
rect 117004 -4662 117186 -4426
rect 117422 -4662 117604 -4426
rect 117004 -5624 117604 -4662
rect 120604 194254 121204 218000
rect 120604 194018 120786 194254
rect 121022 194018 121204 194254
rect 120604 193934 121204 194018
rect 120604 193698 120786 193934
rect 121022 193698 121204 193934
rect 120604 158254 121204 193698
rect 120604 158018 120786 158254
rect 121022 158018 121204 158254
rect 120604 157934 121204 158018
rect 120604 157698 120786 157934
rect 121022 157698 121204 157934
rect 120604 122254 121204 157698
rect 120604 122018 120786 122254
rect 121022 122018 121204 122254
rect 120604 121934 121204 122018
rect 120604 121698 120786 121934
rect 121022 121698 121204 121934
rect 120604 86254 121204 121698
rect 120604 86018 120786 86254
rect 121022 86018 121204 86254
rect 120604 85934 121204 86018
rect 120604 85698 120786 85934
rect 121022 85698 121204 85934
rect 120604 50254 121204 85698
rect 120604 50018 120786 50254
rect 121022 50018 121204 50254
rect 120604 49934 121204 50018
rect 120604 49698 120786 49934
rect 121022 49698 121204 49934
rect 120604 14254 121204 49698
rect 120604 14018 120786 14254
rect 121022 14018 121204 14254
rect 120604 13934 121204 14018
rect 120604 13698 120786 13934
rect 121022 13698 121204 13934
rect 102604 -7162 102786 -6926
rect 103022 -7162 103204 -6926
rect 102604 -7246 103204 -7162
rect 102604 -7482 102786 -7246
rect 103022 -7482 103204 -7246
rect 102604 -7504 103204 -7482
rect 120604 -5986 121204 13698
rect 127804 201454 128404 218000
rect 127804 201218 127986 201454
rect 128222 201218 128404 201454
rect 127804 201134 128404 201218
rect 127804 200898 127986 201134
rect 128222 200898 128404 201134
rect 127804 165454 128404 200898
rect 127804 165218 127986 165454
rect 128222 165218 128404 165454
rect 127804 165134 128404 165218
rect 127804 164898 127986 165134
rect 128222 164898 128404 165134
rect 127804 129454 128404 164898
rect 127804 129218 127986 129454
rect 128222 129218 128404 129454
rect 127804 129134 128404 129218
rect 127804 128898 127986 129134
rect 128222 128898 128404 129134
rect 127804 93454 128404 128898
rect 127804 93218 127986 93454
rect 128222 93218 128404 93454
rect 127804 93134 128404 93218
rect 127804 92898 127986 93134
rect 128222 92898 128404 93134
rect 127804 57454 128404 92898
rect 127804 57218 127986 57454
rect 128222 57218 128404 57454
rect 127804 57134 128404 57218
rect 127804 56898 127986 57134
rect 128222 56898 128404 57134
rect 127804 21454 128404 56898
rect 127804 21218 127986 21454
rect 128222 21218 128404 21454
rect 127804 21134 128404 21218
rect 127804 20898 127986 21134
rect 128222 20898 128404 21134
rect 127804 -1286 128404 20898
rect 127804 -1522 127986 -1286
rect 128222 -1522 128404 -1286
rect 127804 -1606 128404 -1522
rect 127804 -1842 127986 -1606
rect 128222 -1842 128404 -1606
rect 127804 -1864 128404 -1842
rect 131404 205054 132004 218000
rect 131404 204818 131586 205054
rect 131822 204818 132004 205054
rect 131404 204734 132004 204818
rect 131404 204498 131586 204734
rect 131822 204498 132004 204734
rect 131404 169054 132004 204498
rect 131404 168818 131586 169054
rect 131822 168818 132004 169054
rect 131404 168734 132004 168818
rect 131404 168498 131586 168734
rect 131822 168498 132004 168734
rect 131404 133054 132004 168498
rect 131404 132818 131586 133054
rect 131822 132818 132004 133054
rect 131404 132734 132004 132818
rect 131404 132498 131586 132734
rect 131822 132498 132004 132734
rect 131404 97054 132004 132498
rect 131404 96818 131586 97054
rect 131822 96818 132004 97054
rect 131404 96734 132004 96818
rect 131404 96498 131586 96734
rect 131822 96498 132004 96734
rect 131404 61054 132004 96498
rect 131404 60818 131586 61054
rect 131822 60818 132004 61054
rect 131404 60734 132004 60818
rect 131404 60498 131586 60734
rect 131822 60498 132004 60734
rect 131404 25054 132004 60498
rect 131404 24818 131586 25054
rect 131822 24818 132004 25054
rect 131404 24734 132004 24818
rect 131404 24498 131586 24734
rect 131822 24498 132004 24734
rect 131404 -3166 132004 24498
rect 131404 -3402 131586 -3166
rect 131822 -3402 132004 -3166
rect 131404 -3486 132004 -3402
rect 131404 -3722 131586 -3486
rect 131822 -3722 132004 -3486
rect 131404 -3744 132004 -3722
rect 135004 208654 135604 218000
rect 135004 208418 135186 208654
rect 135422 208418 135604 208654
rect 135004 208334 135604 208418
rect 135004 208098 135186 208334
rect 135422 208098 135604 208334
rect 135004 172654 135604 208098
rect 135004 172418 135186 172654
rect 135422 172418 135604 172654
rect 135004 172334 135604 172418
rect 135004 172098 135186 172334
rect 135422 172098 135604 172334
rect 135004 136654 135604 172098
rect 135004 136418 135186 136654
rect 135422 136418 135604 136654
rect 135004 136334 135604 136418
rect 135004 136098 135186 136334
rect 135422 136098 135604 136334
rect 135004 100654 135604 136098
rect 135004 100418 135186 100654
rect 135422 100418 135604 100654
rect 135004 100334 135604 100418
rect 135004 100098 135186 100334
rect 135422 100098 135604 100334
rect 135004 64654 135604 100098
rect 135004 64418 135186 64654
rect 135422 64418 135604 64654
rect 135004 64334 135604 64418
rect 135004 64098 135186 64334
rect 135422 64098 135604 64334
rect 135004 28654 135604 64098
rect 135004 28418 135186 28654
rect 135422 28418 135604 28654
rect 135004 28334 135604 28418
rect 135004 28098 135186 28334
rect 135422 28098 135604 28334
rect 135004 -5046 135604 28098
rect 135004 -5282 135186 -5046
rect 135422 -5282 135604 -5046
rect 135004 -5366 135604 -5282
rect 135004 -5602 135186 -5366
rect 135422 -5602 135604 -5366
rect 135004 -5624 135604 -5602
rect 138604 212254 139204 218000
rect 138604 212018 138786 212254
rect 139022 212018 139204 212254
rect 138604 211934 139204 212018
rect 138604 211698 138786 211934
rect 139022 211698 139204 211934
rect 138604 176254 139204 211698
rect 138604 176018 138786 176254
rect 139022 176018 139204 176254
rect 138604 175934 139204 176018
rect 138604 175698 138786 175934
rect 139022 175698 139204 175934
rect 138604 140254 139204 175698
rect 138604 140018 138786 140254
rect 139022 140018 139204 140254
rect 138604 139934 139204 140018
rect 138604 139698 138786 139934
rect 139022 139698 139204 139934
rect 138604 104254 139204 139698
rect 138604 104018 138786 104254
rect 139022 104018 139204 104254
rect 138604 103934 139204 104018
rect 138604 103698 138786 103934
rect 139022 103698 139204 103934
rect 138604 68254 139204 103698
rect 138604 68018 138786 68254
rect 139022 68018 139204 68254
rect 138604 67934 139204 68018
rect 138604 67698 138786 67934
rect 139022 67698 139204 67934
rect 138604 32254 139204 67698
rect 138604 32018 138786 32254
rect 139022 32018 139204 32254
rect 138604 31934 139204 32018
rect 138604 31698 138786 31934
rect 139022 31698 139204 31934
rect 120604 -6222 120786 -5986
rect 121022 -6222 121204 -5986
rect 120604 -6306 121204 -6222
rect 120604 -6542 120786 -6306
rect 121022 -6542 121204 -6306
rect 120604 -7504 121204 -6542
rect 138604 -6926 139204 31698
rect 145804 183454 146404 218000
rect 145804 183218 145986 183454
rect 146222 183218 146404 183454
rect 145804 183134 146404 183218
rect 145804 182898 145986 183134
rect 146222 182898 146404 183134
rect 145804 147454 146404 182898
rect 145804 147218 145986 147454
rect 146222 147218 146404 147454
rect 145804 147134 146404 147218
rect 145804 146898 145986 147134
rect 146222 146898 146404 147134
rect 145804 111454 146404 146898
rect 145804 111218 145986 111454
rect 146222 111218 146404 111454
rect 145804 111134 146404 111218
rect 145804 110898 145986 111134
rect 146222 110898 146404 111134
rect 145804 75454 146404 110898
rect 145804 75218 145986 75454
rect 146222 75218 146404 75454
rect 145804 75134 146404 75218
rect 145804 74898 145986 75134
rect 146222 74898 146404 75134
rect 145804 39454 146404 74898
rect 145804 39218 145986 39454
rect 146222 39218 146404 39454
rect 145804 39134 146404 39218
rect 145804 38898 145986 39134
rect 146222 38898 146404 39134
rect 145804 3454 146404 38898
rect 145804 3218 145986 3454
rect 146222 3218 146404 3454
rect 145804 3134 146404 3218
rect 145804 2898 145986 3134
rect 146222 2898 146404 3134
rect 145804 -346 146404 2898
rect 145804 -582 145986 -346
rect 146222 -582 146404 -346
rect 145804 -666 146404 -582
rect 145804 -902 145986 -666
rect 146222 -902 146404 -666
rect 145804 -1864 146404 -902
rect 149404 187054 150004 218000
rect 149404 186818 149586 187054
rect 149822 186818 150004 187054
rect 149404 186734 150004 186818
rect 149404 186498 149586 186734
rect 149822 186498 150004 186734
rect 149404 151054 150004 186498
rect 149404 150818 149586 151054
rect 149822 150818 150004 151054
rect 149404 150734 150004 150818
rect 149404 150498 149586 150734
rect 149822 150498 150004 150734
rect 149404 115054 150004 150498
rect 149404 114818 149586 115054
rect 149822 114818 150004 115054
rect 149404 114734 150004 114818
rect 149404 114498 149586 114734
rect 149822 114498 150004 114734
rect 149404 79054 150004 114498
rect 149404 78818 149586 79054
rect 149822 78818 150004 79054
rect 149404 78734 150004 78818
rect 149404 78498 149586 78734
rect 149822 78498 150004 78734
rect 149404 43054 150004 78498
rect 149404 42818 149586 43054
rect 149822 42818 150004 43054
rect 149404 42734 150004 42818
rect 149404 42498 149586 42734
rect 149822 42498 150004 42734
rect 149404 7054 150004 42498
rect 149404 6818 149586 7054
rect 149822 6818 150004 7054
rect 149404 6734 150004 6818
rect 149404 6498 149586 6734
rect 149822 6498 150004 6734
rect 149404 -2226 150004 6498
rect 149404 -2462 149586 -2226
rect 149822 -2462 150004 -2226
rect 149404 -2546 150004 -2462
rect 149404 -2782 149586 -2546
rect 149822 -2782 150004 -2546
rect 149404 -3744 150004 -2782
rect 153004 190654 153604 218000
rect 153004 190418 153186 190654
rect 153422 190418 153604 190654
rect 153004 190334 153604 190418
rect 153004 190098 153186 190334
rect 153422 190098 153604 190334
rect 153004 154654 153604 190098
rect 153004 154418 153186 154654
rect 153422 154418 153604 154654
rect 153004 154334 153604 154418
rect 153004 154098 153186 154334
rect 153422 154098 153604 154334
rect 153004 118654 153604 154098
rect 153004 118418 153186 118654
rect 153422 118418 153604 118654
rect 153004 118334 153604 118418
rect 153004 118098 153186 118334
rect 153422 118098 153604 118334
rect 153004 82654 153604 118098
rect 153004 82418 153186 82654
rect 153422 82418 153604 82654
rect 153004 82334 153604 82418
rect 153004 82098 153186 82334
rect 153422 82098 153604 82334
rect 153004 46654 153604 82098
rect 153004 46418 153186 46654
rect 153422 46418 153604 46654
rect 153004 46334 153604 46418
rect 153004 46098 153186 46334
rect 153422 46098 153604 46334
rect 153004 10654 153604 46098
rect 153004 10418 153186 10654
rect 153422 10418 153604 10654
rect 153004 10334 153604 10418
rect 153004 10098 153186 10334
rect 153422 10098 153604 10334
rect 153004 -4106 153604 10098
rect 153004 -4342 153186 -4106
rect 153422 -4342 153604 -4106
rect 153004 -4426 153604 -4342
rect 153004 -4662 153186 -4426
rect 153422 -4662 153604 -4426
rect 153004 -5624 153604 -4662
rect 156604 194254 157204 218000
rect 156604 194018 156786 194254
rect 157022 194018 157204 194254
rect 156604 193934 157204 194018
rect 156604 193698 156786 193934
rect 157022 193698 157204 193934
rect 156604 158254 157204 193698
rect 156604 158018 156786 158254
rect 157022 158018 157204 158254
rect 156604 157934 157204 158018
rect 156604 157698 156786 157934
rect 157022 157698 157204 157934
rect 156604 122254 157204 157698
rect 156604 122018 156786 122254
rect 157022 122018 157204 122254
rect 156604 121934 157204 122018
rect 156604 121698 156786 121934
rect 157022 121698 157204 121934
rect 156604 86254 157204 121698
rect 156604 86018 156786 86254
rect 157022 86018 157204 86254
rect 156604 85934 157204 86018
rect 156604 85698 156786 85934
rect 157022 85698 157204 85934
rect 156604 50254 157204 85698
rect 156604 50018 156786 50254
rect 157022 50018 157204 50254
rect 156604 49934 157204 50018
rect 156604 49698 156786 49934
rect 157022 49698 157204 49934
rect 156604 14254 157204 49698
rect 156604 14018 156786 14254
rect 157022 14018 157204 14254
rect 156604 13934 157204 14018
rect 156604 13698 156786 13934
rect 157022 13698 157204 13934
rect 138604 -7162 138786 -6926
rect 139022 -7162 139204 -6926
rect 138604 -7246 139204 -7162
rect 138604 -7482 138786 -7246
rect 139022 -7482 139204 -7246
rect 138604 -7504 139204 -7482
rect 156604 -5986 157204 13698
rect 163804 201454 164404 218000
rect 163804 201218 163986 201454
rect 164222 201218 164404 201454
rect 163804 201134 164404 201218
rect 163804 200898 163986 201134
rect 164222 200898 164404 201134
rect 163804 165454 164404 200898
rect 163804 165218 163986 165454
rect 164222 165218 164404 165454
rect 163804 165134 164404 165218
rect 163804 164898 163986 165134
rect 164222 164898 164404 165134
rect 163804 129454 164404 164898
rect 163804 129218 163986 129454
rect 164222 129218 164404 129454
rect 163804 129134 164404 129218
rect 163804 128898 163986 129134
rect 164222 128898 164404 129134
rect 163804 93454 164404 128898
rect 163804 93218 163986 93454
rect 164222 93218 164404 93454
rect 163804 93134 164404 93218
rect 163804 92898 163986 93134
rect 164222 92898 164404 93134
rect 163804 57454 164404 92898
rect 163804 57218 163986 57454
rect 164222 57218 164404 57454
rect 163804 57134 164404 57218
rect 163804 56898 163986 57134
rect 164222 56898 164404 57134
rect 163804 21454 164404 56898
rect 163804 21218 163986 21454
rect 164222 21218 164404 21454
rect 163804 21134 164404 21218
rect 163804 20898 163986 21134
rect 164222 20898 164404 21134
rect 163804 -1286 164404 20898
rect 163804 -1522 163986 -1286
rect 164222 -1522 164404 -1286
rect 163804 -1606 164404 -1522
rect 163804 -1842 163986 -1606
rect 164222 -1842 164404 -1606
rect 163804 -1864 164404 -1842
rect 167404 205054 168004 218000
rect 167404 204818 167586 205054
rect 167822 204818 168004 205054
rect 167404 204734 168004 204818
rect 167404 204498 167586 204734
rect 167822 204498 168004 204734
rect 167404 169054 168004 204498
rect 167404 168818 167586 169054
rect 167822 168818 168004 169054
rect 167404 168734 168004 168818
rect 167404 168498 167586 168734
rect 167822 168498 168004 168734
rect 167404 133054 168004 168498
rect 167404 132818 167586 133054
rect 167822 132818 168004 133054
rect 167404 132734 168004 132818
rect 167404 132498 167586 132734
rect 167822 132498 168004 132734
rect 167404 97054 168004 132498
rect 167404 96818 167586 97054
rect 167822 96818 168004 97054
rect 167404 96734 168004 96818
rect 167404 96498 167586 96734
rect 167822 96498 168004 96734
rect 167404 61054 168004 96498
rect 167404 60818 167586 61054
rect 167822 60818 168004 61054
rect 167404 60734 168004 60818
rect 167404 60498 167586 60734
rect 167822 60498 168004 60734
rect 167404 25054 168004 60498
rect 167404 24818 167586 25054
rect 167822 24818 168004 25054
rect 167404 24734 168004 24818
rect 167404 24498 167586 24734
rect 167822 24498 168004 24734
rect 167404 -3166 168004 24498
rect 167404 -3402 167586 -3166
rect 167822 -3402 168004 -3166
rect 167404 -3486 168004 -3402
rect 167404 -3722 167586 -3486
rect 167822 -3722 168004 -3486
rect 167404 -3744 168004 -3722
rect 171004 208654 171604 218000
rect 171004 208418 171186 208654
rect 171422 208418 171604 208654
rect 171004 208334 171604 208418
rect 171004 208098 171186 208334
rect 171422 208098 171604 208334
rect 171004 172654 171604 208098
rect 171004 172418 171186 172654
rect 171422 172418 171604 172654
rect 171004 172334 171604 172418
rect 171004 172098 171186 172334
rect 171422 172098 171604 172334
rect 171004 136654 171604 172098
rect 171004 136418 171186 136654
rect 171422 136418 171604 136654
rect 171004 136334 171604 136418
rect 171004 136098 171186 136334
rect 171422 136098 171604 136334
rect 171004 100654 171604 136098
rect 171004 100418 171186 100654
rect 171422 100418 171604 100654
rect 171004 100334 171604 100418
rect 171004 100098 171186 100334
rect 171422 100098 171604 100334
rect 171004 64654 171604 100098
rect 171004 64418 171186 64654
rect 171422 64418 171604 64654
rect 171004 64334 171604 64418
rect 171004 64098 171186 64334
rect 171422 64098 171604 64334
rect 171004 28654 171604 64098
rect 171004 28418 171186 28654
rect 171422 28418 171604 28654
rect 171004 28334 171604 28418
rect 171004 28098 171186 28334
rect 171422 28098 171604 28334
rect 171004 -5046 171604 28098
rect 171004 -5282 171186 -5046
rect 171422 -5282 171604 -5046
rect 171004 -5366 171604 -5282
rect 171004 -5602 171186 -5366
rect 171422 -5602 171604 -5366
rect 171004 -5624 171604 -5602
rect 174604 212254 175204 218000
rect 174604 212018 174786 212254
rect 175022 212018 175204 212254
rect 174604 211934 175204 212018
rect 174604 211698 174786 211934
rect 175022 211698 175204 211934
rect 174604 176254 175204 211698
rect 174604 176018 174786 176254
rect 175022 176018 175204 176254
rect 174604 175934 175204 176018
rect 174604 175698 174786 175934
rect 175022 175698 175204 175934
rect 174604 140254 175204 175698
rect 174604 140018 174786 140254
rect 175022 140018 175204 140254
rect 174604 139934 175204 140018
rect 174604 139698 174786 139934
rect 175022 139698 175204 139934
rect 174604 104254 175204 139698
rect 174604 104018 174786 104254
rect 175022 104018 175204 104254
rect 174604 103934 175204 104018
rect 174604 103698 174786 103934
rect 175022 103698 175204 103934
rect 174604 68254 175204 103698
rect 174604 68018 174786 68254
rect 175022 68018 175204 68254
rect 174604 67934 175204 68018
rect 174604 67698 174786 67934
rect 175022 67698 175204 67934
rect 174604 32254 175204 67698
rect 174604 32018 174786 32254
rect 175022 32018 175204 32254
rect 174604 31934 175204 32018
rect 174604 31698 174786 31934
rect 175022 31698 175204 31934
rect 156604 -6222 156786 -5986
rect 157022 -6222 157204 -5986
rect 156604 -6306 157204 -6222
rect 156604 -6542 156786 -6306
rect 157022 -6542 157204 -6306
rect 156604 -7504 157204 -6542
rect 174604 -6926 175204 31698
rect 181804 183454 182404 218000
rect 181804 183218 181986 183454
rect 182222 183218 182404 183454
rect 181804 183134 182404 183218
rect 181804 182898 181986 183134
rect 182222 182898 182404 183134
rect 181804 147454 182404 182898
rect 181804 147218 181986 147454
rect 182222 147218 182404 147454
rect 181804 147134 182404 147218
rect 181804 146898 181986 147134
rect 182222 146898 182404 147134
rect 181804 111454 182404 146898
rect 181804 111218 181986 111454
rect 182222 111218 182404 111454
rect 181804 111134 182404 111218
rect 181804 110898 181986 111134
rect 182222 110898 182404 111134
rect 181804 75454 182404 110898
rect 181804 75218 181986 75454
rect 182222 75218 182404 75454
rect 181804 75134 182404 75218
rect 181804 74898 181986 75134
rect 182222 74898 182404 75134
rect 181804 39454 182404 74898
rect 181804 39218 181986 39454
rect 182222 39218 182404 39454
rect 181804 39134 182404 39218
rect 181804 38898 181986 39134
rect 182222 38898 182404 39134
rect 181804 3454 182404 38898
rect 181804 3218 181986 3454
rect 182222 3218 182404 3454
rect 181804 3134 182404 3218
rect 181804 2898 181986 3134
rect 182222 2898 182404 3134
rect 181804 -346 182404 2898
rect 181804 -582 181986 -346
rect 182222 -582 182404 -346
rect 181804 -666 182404 -582
rect 181804 -902 181986 -666
rect 182222 -902 182404 -666
rect 181804 -1864 182404 -902
rect 185404 187054 186004 218000
rect 185404 186818 185586 187054
rect 185822 186818 186004 187054
rect 185404 186734 186004 186818
rect 185404 186498 185586 186734
rect 185822 186498 186004 186734
rect 185404 151054 186004 186498
rect 185404 150818 185586 151054
rect 185822 150818 186004 151054
rect 185404 150734 186004 150818
rect 185404 150498 185586 150734
rect 185822 150498 186004 150734
rect 185404 115054 186004 150498
rect 185404 114818 185586 115054
rect 185822 114818 186004 115054
rect 185404 114734 186004 114818
rect 185404 114498 185586 114734
rect 185822 114498 186004 114734
rect 185404 79054 186004 114498
rect 185404 78818 185586 79054
rect 185822 78818 186004 79054
rect 185404 78734 186004 78818
rect 185404 78498 185586 78734
rect 185822 78498 186004 78734
rect 185404 43054 186004 78498
rect 185404 42818 185586 43054
rect 185822 42818 186004 43054
rect 185404 42734 186004 42818
rect 185404 42498 185586 42734
rect 185822 42498 186004 42734
rect 185404 7054 186004 42498
rect 185404 6818 185586 7054
rect 185822 6818 186004 7054
rect 185404 6734 186004 6818
rect 185404 6498 185586 6734
rect 185822 6498 186004 6734
rect 185404 -2226 186004 6498
rect 185404 -2462 185586 -2226
rect 185822 -2462 186004 -2226
rect 185404 -2546 186004 -2462
rect 185404 -2782 185586 -2546
rect 185822 -2782 186004 -2546
rect 185404 -3744 186004 -2782
rect 189004 190654 189604 218000
rect 189004 190418 189186 190654
rect 189422 190418 189604 190654
rect 189004 190334 189604 190418
rect 189004 190098 189186 190334
rect 189422 190098 189604 190334
rect 189004 154654 189604 190098
rect 189004 154418 189186 154654
rect 189422 154418 189604 154654
rect 189004 154334 189604 154418
rect 189004 154098 189186 154334
rect 189422 154098 189604 154334
rect 189004 118654 189604 154098
rect 189004 118418 189186 118654
rect 189422 118418 189604 118654
rect 189004 118334 189604 118418
rect 189004 118098 189186 118334
rect 189422 118098 189604 118334
rect 189004 82654 189604 118098
rect 189004 82418 189186 82654
rect 189422 82418 189604 82654
rect 189004 82334 189604 82418
rect 189004 82098 189186 82334
rect 189422 82098 189604 82334
rect 189004 46654 189604 82098
rect 189004 46418 189186 46654
rect 189422 46418 189604 46654
rect 189004 46334 189604 46418
rect 189004 46098 189186 46334
rect 189422 46098 189604 46334
rect 189004 10654 189604 46098
rect 189004 10418 189186 10654
rect 189422 10418 189604 10654
rect 189004 10334 189604 10418
rect 189004 10098 189186 10334
rect 189422 10098 189604 10334
rect 189004 -4106 189604 10098
rect 189004 -4342 189186 -4106
rect 189422 -4342 189604 -4106
rect 189004 -4426 189604 -4342
rect 189004 -4662 189186 -4426
rect 189422 -4662 189604 -4426
rect 189004 -5624 189604 -4662
rect 192604 194254 193204 218000
rect 192604 194018 192786 194254
rect 193022 194018 193204 194254
rect 192604 193934 193204 194018
rect 192604 193698 192786 193934
rect 193022 193698 193204 193934
rect 192604 158254 193204 193698
rect 192604 158018 192786 158254
rect 193022 158018 193204 158254
rect 192604 157934 193204 158018
rect 192604 157698 192786 157934
rect 193022 157698 193204 157934
rect 192604 122254 193204 157698
rect 192604 122018 192786 122254
rect 193022 122018 193204 122254
rect 192604 121934 193204 122018
rect 192604 121698 192786 121934
rect 193022 121698 193204 121934
rect 192604 86254 193204 121698
rect 192604 86018 192786 86254
rect 193022 86018 193204 86254
rect 192604 85934 193204 86018
rect 192604 85698 192786 85934
rect 193022 85698 193204 85934
rect 192604 50254 193204 85698
rect 192604 50018 192786 50254
rect 193022 50018 193204 50254
rect 192604 49934 193204 50018
rect 192604 49698 192786 49934
rect 193022 49698 193204 49934
rect 192604 14254 193204 49698
rect 192604 14018 192786 14254
rect 193022 14018 193204 14254
rect 192604 13934 193204 14018
rect 192604 13698 192786 13934
rect 193022 13698 193204 13934
rect 174604 -7162 174786 -6926
rect 175022 -7162 175204 -6926
rect 174604 -7246 175204 -7162
rect 174604 -7482 174786 -7246
rect 175022 -7482 175204 -7246
rect 174604 -7504 175204 -7482
rect 192604 -5986 193204 13698
rect 199804 201454 200404 218000
rect 199804 201218 199986 201454
rect 200222 201218 200404 201454
rect 199804 201134 200404 201218
rect 199804 200898 199986 201134
rect 200222 200898 200404 201134
rect 199804 165454 200404 200898
rect 199804 165218 199986 165454
rect 200222 165218 200404 165454
rect 199804 165134 200404 165218
rect 199804 164898 199986 165134
rect 200222 164898 200404 165134
rect 199804 129454 200404 164898
rect 199804 129218 199986 129454
rect 200222 129218 200404 129454
rect 199804 129134 200404 129218
rect 199804 128898 199986 129134
rect 200222 128898 200404 129134
rect 199804 93454 200404 128898
rect 199804 93218 199986 93454
rect 200222 93218 200404 93454
rect 199804 93134 200404 93218
rect 199804 92898 199986 93134
rect 200222 92898 200404 93134
rect 199804 57454 200404 92898
rect 199804 57218 199986 57454
rect 200222 57218 200404 57454
rect 199804 57134 200404 57218
rect 199804 56898 199986 57134
rect 200222 56898 200404 57134
rect 199804 21454 200404 56898
rect 199804 21218 199986 21454
rect 200222 21218 200404 21454
rect 199804 21134 200404 21218
rect 199804 20898 199986 21134
rect 200222 20898 200404 21134
rect 199804 -1286 200404 20898
rect 199804 -1522 199986 -1286
rect 200222 -1522 200404 -1286
rect 199804 -1606 200404 -1522
rect 199804 -1842 199986 -1606
rect 200222 -1842 200404 -1606
rect 199804 -1864 200404 -1842
rect 203404 205054 204004 218000
rect 203404 204818 203586 205054
rect 203822 204818 204004 205054
rect 203404 204734 204004 204818
rect 203404 204498 203586 204734
rect 203822 204498 204004 204734
rect 203404 169054 204004 204498
rect 203404 168818 203586 169054
rect 203822 168818 204004 169054
rect 203404 168734 204004 168818
rect 203404 168498 203586 168734
rect 203822 168498 204004 168734
rect 203404 133054 204004 168498
rect 203404 132818 203586 133054
rect 203822 132818 204004 133054
rect 203404 132734 204004 132818
rect 203404 132498 203586 132734
rect 203822 132498 204004 132734
rect 203404 97054 204004 132498
rect 203404 96818 203586 97054
rect 203822 96818 204004 97054
rect 203404 96734 204004 96818
rect 203404 96498 203586 96734
rect 203822 96498 204004 96734
rect 203404 61054 204004 96498
rect 203404 60818 203586 61054
rect 203822 60818 204004 61054
rect 203404 60734 204004 60818
rect 203404 60498 203586 60734
rect 203822 60498 204004 60734
rect 203404 25054 204004 60498
rect 203404 24818 203586 25054
rect 203822 24818 204004 25054
rect 203404 24734 204004 24818
rect 203404 24498 203586 24734
rect 203822 24498 204004 24734
rect 203404 -3166 204004 24498
rect 203404 -3402 203586 -3166
rect 203822 -3402 204004 -3166
rect 203404 -3486 204004 -3402
rect 203404 -3722 203586 -3486
rect 203822 -3722 204004 -3486
rect 203404 -3744 204004 -3722
rect 207004 208654 207604 218000
rect 207004 208418 207186 208654
rect 207422 208418 207604 208654
rect 207004 208334 207604 208418
rect 207004 208098 207186 208334
rect 207422 208098 207604 208334
rect 207004 172654 207604 208098
rect 207004 172418 207186 172654
rect 207422 172418 207604 172654
rect 207004 172334 207604 172418
rect 207004 172098 207186 172334
rect 207422 172098 207604 172334
rect 207004 136654 207604 172098
rect 207004 136418 207186 136654
rect 207422 136418 207604 136654
rect 207004 136334 207604 136418
rect 207004 136098 207186 136334
rect 207422 136098 207604 136334
rect 207004 100654 207604 136098
rect 207004 100418 207186 100654
rect 207422 100418 207604 100654
rect 207004 100334 207604 100418
rect 207004 100098 207186 100334
rect 207422 100098 207604 100334
rect 207004 64654 207604 100098
rect 207004 64418 207186 64654
rect 207422 64418 207604 64654
rect 207004 64334 207604 64418
rect 207004 64098 207186 64334
rect 207422 64098 207604 64334
rect 207004 28654 207604 64098
rect 207004 28418 207186 28654
rect 207422 28418 207604 28654
rect 207004 28334 207604 28418
rect 207004 28098 207186 28334
rect 207422 28098 207604 28334
rect 207004 -5046 207604 28098
rect 207004 -5282 207186 -5046
rect 207422 -5282 207604 -5046
rect 207004 -5366 207604 -5282
rect 207004 -5602 207186 -5366
rect 207422 -5602 207604 -5366
rect 207004 -5624 207604 -5602
rect 210604 212254 211204 218000
rect 210604 212018 210786 212254
rect 211022 212018 211204 212254
rect 210604 211934 211204 212018
rect 210604 211698 210786 211934
rect 211022 211698 211204 211934
rect 210604 176254 211204 211698
rect 210604 176018 210786 176254
rect 211022 176018 211204 176254
rect 210604 175934 211204 176018
rect 210604 175698 210786 175934
rect 211022 175698 211204 175934
rect 210604 140254 211204 175698
rect 210604 140018 210786 140254
rect 211022 140018 211204 140254
rect 210604 139934 211204 140018
rect 210604 139698 210786 139934
rect 211022 139698 211204 139934
rect 210604 104254 211204 139698
rect 210604 104018 210786 104254
rect 211022 104018 211204 104254
rect 210604 103934 211204 104018
rect 210604 103698 210786 103934
rect 211022 103698 211204 103934
rect 210604 68254 211204 103698
rect 210604 68018 210786 68254
rect 211022 68018 211204 68254
rect 210604 67934 211204 68018
rect 210604 67698 210786 67934
rect 211022 67698 211204 67934
rect 210604 32254 211204 67698
rect 210604 32018 210786 32254
rect 211022 32018 211204 32254
rect 210604 31934 211204 32018
rect 210604 31698 210786 31934
rect 211022 31698 211204 31934
rect 192604 -6222 192786 -5986
rect 193022 -6222 193204 -5986
rect 192604 -6306 193204 -6222
rect 192604 -6542 192786 -6306
rect 193022 -6542 193204 -6306
rect 192604 -7504 193204 -6542
rect 210604 -6926 211204 31698
rect 217804 183454 218404 218000
rect 217804 183218 217986 183454
rect 218222 183218 218404 183454
rect 217804 183134 218404 183218
rect 217804 182898 217986 183134
rect 218222 182898 218404 183134
rect 217804 147454 218404 182898
rect 217804 147218 217986 147454
rect 218222 147218 218404 147454
rect 217804 147134 218404 147218
rect 217804 146898 217986 147134
rect 218222 146898 218404 147134
rect 217804 111454 218404 146898
rect 217804 111218 217986 111454
rect 218222 111218 218404 111454
rect 217804 111134 218404 111218
rect 217804 110898 217986 111134
rect 218222 110898 218404 111134
rect 217804 75454 218404 110898
rect 217804 75218 217986 75454
rect 218222 75218 218404 75454
rect 217804 75134 218404 75218
rect 217804 74898 217986 75134
rect 218222 74898 218404 75134
rect 217804 39454 218404 74898
rect 217804 39218 217986 39454
rect 218222 39218 218404 39454
rect 217804 39134 218404 39218
rect 217804 38898 217986 39134
rect 218222 38898 218404 39134
rect 217804 3454 218404 38898
rect 217804 3218 217986 3454
rect 218222 3218 218404 3454
rect 217804 3134 218404 3218
rect 217804 2898 217986 3134
rect 218222 2898 218404 3134
rect 217804 -346 218404 2898
rect 217804 -582 217986 -346
rect 218222 -582 218404 -346
rect 217804 -666 218404 -582
rect 217804 -902 217986 -666
rect 218222 -902 218404 -666
rect 217804 -1864 218404 -902
rect 221404 187054 222004 218000
rect 221404 186818 221586 187054
rect 221822 186818 222004 187054
rect 221404 186734 222004 186818
rect 221404 186498 221586 186734
rect 221822 186498 222004 186734
rect 221404 151054 222004 186498
rect 221404 150818 221586 151054
rect 221822 150818 222004 151054
rect 221404 150734 222004 150818
rect 221404 150498 221586 150734
rect 221822 150498 222004 150734
rect 221404 115054 222004 150498
rect 221404 114818 221586 115054
rect 221822 114818 222004 115054
rect 221404 114734 222004 114818
rect 221404 114498 221586 114734
rect 221822 114498 222004 114734
rect 221404 79054 222004 114498
rect 221404 78818 221586 79054
rect 221822 78818 222004 79054
rect 221404 78734 222004 78818
rect 221404 78498 221586 78734
rect 221822 78498 222004 78734
rect 221404 43054 222004 78498
rect 221404 42818 221586 43054
rect 221822 42818 222004 43054
rect 221404 42734 222004 42818
rect 221404 42498 221586 42734
rect 221822 42498 222004 42734
rect 221404 7054 222004 42498
rect 221404 6818 221586 7054
rect 221822 6818 222004 7054
rect 221404 6734 222004 6818
rect 221404 6498 221586 6734
rect 221822 6498 222004 6734
rect 221404 -2226 222004 6498
rect 221404 -2462 221586 -2226
rect 221822 -2462 222004 -2226
rect 221404 -2546 222004 -2462
rect 221404 -2782 221586 -2546
rect 221822 -2782 222004 -2546
rect 221404 -3744 222004 -2782
rect 225004 190654 225604 218000
rect 225004 190418 225186 190654
rect 225422 190418 225604 190654
rect 225004 190334 225604 190418
rect 225004 190098 225186 190334
rect 225422 190098 225604 190334
rect 225004 154654 225604 190098
rect 225004 154418 225186 154654
rect 225422 154418 225604 154654
rect 225004 154334 225604 154418
rect 225004 154098 225186 154334
rect 225422 154098 225604 154334
rect 225004 118654 225604 154098
rect 225004 118418 225186 118654
rect 225422 118418 225604 118654
rect 225004 118334 225604 118418
rect 225004 118098 225186 118334
rect 225422 118098 225604 118334
rect 225004 82654 225604 118098
rect 225004 82418 225186 82654
rect 225422 82418 225604 82654
rect 225004 82334 225604 82418
rect 225004 82098 225186 82334
rect 225422 82098 225604 82334
rect 225004 46654 225604 82098
rect 225004 46418 225186 46654
rect 225422 46418 225604 46654
rect 225004 46334 225604 46418
rect 225004 46098 225186 46334
rect 225422 46098 225604 46334
rect 225004 10654 225604 46098
rect 225004 10418 225186 10654
rect 225422 10418 225604 10654
rect 225004 10334 225604 10418
rect 225004 10098 225186 10334
rect 225422 10098 225604 10334
rect 225004 -4106 225604 10098
rect 225004 -4342 225186 -4106
rect 225422 -4342 225604 -4106
rect 225004 -4426 225604 -4342
rect 225004 -4662 225186 -4426
rect 225422 -4662 225604 -4426
rect 225004 -5624 225604 -4662
rect 228604 194254 229204 218000
rect 228604 194018 228786 194254
rect 229022 194018 229204 194254
rect 228604 193934 229204 194018
rect 228604 193698 228786 193934
rect 229022 193698 229204 193934
rect 228604 158254 229204 193698
rect 228604 158018 228786 158254
rect 229022 158018 229204 158254
rect 228604 157934 229204 158018
rect 228604 157698 228786 157934
rect 229022 157698 229204 157934
rect 228604 122254 229204 157698
rect 228604 122018 228786 122254
rect 229022 122018 229204 122254
rect 228604 121934 229204 122018
rect 228604 121698 228786 121934
rect 229022 121698 229204 121934
rect 228604 86254 229204 121698
rect 228604 86018 228786 86254
rect 229022 86018 229204 86254
rect 228604 85934 229204 86018
rect 228604 85698 228786 85934
rect 229022 85698 229204 85934
rect 228604 50254 229204 85698
rect 228604 50018 228786 50254
rect 229022 50018 229204 50254
rect 228604 49934 229204 50018
rect 228604 49698 228786 49934
rect 229022 49698 229204 49934
rect 228604 14254 229204 49698
rect 228604 14018 228786 14254
rect 229022 14018 229204 14254
rect 228604 13934 229204 14018
rect 228604 13698 228786 13934
rect 229022 13698 229204 13934
rect 210604 -7162 210786 -6926
rect 211022 -7162 211204 -6926
rect 210604 -7246 211204 -7162
rect 210604 -7482 210786 -7246
rect 211022 -7482 211204 -7246
rect 210604 -7504 211204 -7482
rect 228604 -5986 229204 13698
rect 235804 201454 236404 218000
rect 235804 201218 235986 201454
rect 236222 201218 236404 201454
rect 235804 201134 236404 201218
rect 235804 200898 235986 201134
rect 236222 200898 236404 201134
rect 235804 165454 236404 200898
rect 235804 165218 235986 165454
rect 236222 165218 236404 165454
rect 235804 165134 236404 165218
rect 235804 164898 235986 165134
rect 236222 164898 236404 165134
rect 235804 129454 236404 164898
rect 235804 129218 235986 129454
rect 236222 129218 236404 129454
rect 235804 129134 236404 129218
rect 235804 128898 235986 129134
rect 236222 128898 236404 129134
rect 235804 93454 236404 128898
rect 235804 93218 235986 93454
rect 236222 93218 236404 93454
rect 235804 93134 236404 93218
rect 235804 92898 235986 93134
rect 236222 92898 236404 93134
rect 235804 57454 236404 92898
rect 235804 57218 235986 57454
rect 236222 57218 236404 57454
rect 235804 57134 236404 57218
rect 235804 56898 235986 57134
rect 236222 56898 236404 57134
rect 235804 21454 236404 56898
rect 235804 21218 235986 21454
rect 236222 21218 236404 21454
rect 235804 21134 236404 21218
rect 235804 20898 235986 21134
rect 236222 20898 236404 21134
rect 235804 -1286 236404 20898
rect 235804 -1522 235986 -1286
rect 236222 -1522 236404 -1286
rect 235804 -1606 236404 -1522
rect 235804 -1842 235986 -1606
rect 236222 -1842 236404 -1606
rect 235804 -1864 236404 -1842
rect 239404 205054 240004 218000
rect 239404 204818 239586 205054
rect 239822 204818 240004 205054
rect 239404 204734 240004 204818
rect 239404 204498 239586 204734
rect 239822 204498 240004 204734
rect 239404 169054 240004 204498
rect 239404 168818 239586 169054
rect 239822 168818 240004 169054
rect 239404 168734 240004 168818
rect 239404 168498 239586 168734
rect 239822 168498 240004 168734
rect 239404 133054 240004 168498
rect 239404 132818 239586 133054
rect 239822 132818 240004 133054
rect 239404 132734 240004 132818
rect 239404 132498 239586 132734
rect 239822 132498 240004 132734
rect 239404 97054 240004 132498
rect 239404 96818 239586 97054
rect 239822 96818 240004 97054
rect 239404 96734 240004 96818
rect 239404 96498 239586 96734
rect 239822 96498 240004 96734
rect 239404 61054 240004 96498
rect 239404 60818 239586 61054
rect 239822 60818 240004 61054
rect 239404 60734 240004 60818
rect 239404 60498 239586 60734
rect 239822 60498 240004 60734
rect 239404 25054 240004 60498
rect 239404 24818 239586 25054
rect 239822 24818 240004 25054
rect 239404 24734 240004 24818
rect 239404 24498 239586 24734
rect 239822 24498 240004 24734
rect 239404 -3166 240004 24498
rect 239404 -3402 239586 -3166
rect 239822 -3402 240004 -3166
rect 239404 -3486 240004 -3402
rect 239404 -3722 239586 -3486
rect 239822 -3722 240004 -3486
rect 239404 -3744 240004 -3722
rect 243004 208654 243604 218000
rect 243004 208418 243186 208654
rect 243422 208418 243604 208654
rect 243004 208334 243604 208418
rect 243004 208098 243186 208334
rect 243422 208098 243604 208334
rect 243004 172654 243604 208098
rect 243004 172418 243186 172654
rect 243422 172418 243604 172654
rect 243004 172334 243604 172418
rect 243004 172098 243186 172334
rect 243422 172098 243604 172334
rect 243004 136654 243604 172098
rect 243004 136418 243186 136654
rect 243422 136418 243604 136654
rect 243004 136334 243604 136418
rect 243004 136098 243186 136334
rect 243422 136098 243604 136334
rect 243004 100654 243604 136098
rect 243004 100418 243186 100654
rect 243422 100418 243604 100654
rect 243004 100334 243604 100418
rect 243004 100098 243186 100334
rect 243422 100098 243604 100334
rect 243004 64654 243604 100098
rect 243004 64418 243186 64654
rect 243422 64418 243604 64654
rect 243004 64334 243604 64418
rect 243004 64098 243186 64334
rect 243422 64098 243604 64334
rect 243004 28654 243604 64098
rect 243004 28418 243186 28654
rect 243422 28418 243604 28654
rect 243004 28334 243604 28418
rect 243004 28098 243186 28334
rect 243422 28098 243604 28334
rect 243004 -5046 243604 28098
rect 243004 -5282 243186 -5046
rect 243422 -5282 243604 -5046
rect 243004 -5366 243604 -5282
rect 243004 -5602 243186 -5366
rect 243422 -5602 243604 -5366
rect 243004 -5624 243604 -5602
rect 246604 212254 247204 218000
rect 246604 212018 246786 212254
rect 247022 212018 247204 212254
rect 246604 211934 247204 212018
rect 246604 211698 246786 211934
rect 247022 211698 247204 211934
rect 246604 176254 247204 211698
rect 246604 176018 246786 176254
rect 247022 176018 247204 176254
rect 246604 175934 247204 176018
rect 246604 175698 246786 175934
rect 247022 175698 247204 175934
rect 246604 140254 247204 175698
rect 246604 140018 246786 140254
rect 247022 140018 247204 140254
rect 246604 139934 247204 140018
rect 246604 139698 246786 139934
rect 247022 139698 247204 139934
rect 246604 104254 247204 139698
rect 246604 104018 246786 104254
rect 247022 104018 247204 104254
rect 246604 103934 247204 104018
rect 246604 103698 246786 103934
rect 247022 103698 247204 103934
rect 246604 68254 247204 103698
rect 246604 68018 246786 68254
rect 247022 68018 247204 68254
rect 246604 67934 247204 68018
rect 246604 67698 246786 67934
rect 247022 67698 247204 67934
rect 246604 32254 247204 67698
rect 246604 32018 246786 32254
rect 247022 32018 247204 32254
rect 246604 31934 247204 32018
rect 246604 31698 246786 31934
rect 247022 31698 247204 31934
rect 228604 -6222 228786 -5986
rect 229022 -6222 229204 -5986
rect 228604 -6306 229204 -6222
rect 228604 -6542 228786 -6306
rect 229022 -6542 229204 -6306
rect 228604 -7504 229204 -6542
rect 246604 -6926 247204 31698
rect 253804 183454 254404 218000
rect 253804 183218 253986 183454
rect 254222 183218 254404 183454
rect 253804 183134 254404 183218
rect 253804 182898 253986 183134
rect 254222 182898 254404 183134
rect 253804 147454 254404 182898
rect 253804 147218 253986 147454
rect 254222 147218 254404 147454
rect 253804 147134 254404 147218
rect 253804 146898 253986 147134
rect 254222 146898 254404 147134
rect 253804 111454 254404 146898
rect 253804 111218 253986 111454
rect 254222 111218 254404 111454
rect 253804 111134 254404 111218
rect 253804 110898 253986 111134
rect 254222 110898 254404 111134
rect 253804 75454 254404 110898
rect 253804 75218 253986 75454
rect 254222 75218 254404 75454
rect 253804 75134 254404 75218
rect 253804 74898 253986 75134
rect 254222 74898 254404 75134
rect 253804 39454 254404 74898
rect 253804 39218 253986 39454
rect 254222 39218 254404 39454
rect 253804 39134 254404 39218
rect 253804 38898 253986 39134
rect 254222 38898 254404 39134
rect 253804 3454 254404 38898
rect 253804 3218 253986 3454
rect 254222 3218 254404 3454
rect 253804 3134 254404 3218
rect 253804 2898 253986 3134
rect 254222 2898 254404 3134
rect 253804 -346 254404 2898
rect 253804 -582 253986 -346
rect 254222 -582 254404 -346
rect 253804 -666 254404 -582
rect 253804 -902 253986 -666
rect 254222 -902 254404 -666
rect 253804 -1864 254404 -902
rect 257404 187054 258004 218000
rect 257404 186818 257586 187054
rect 257822 186818 258004 187054
rect 257404 186734 258004 186818
rect 257404 186498 257586 186734
rect 257822 186498 258004 186734
rect 257404 151054 258004 186498
rect 257404 150818 257586 151054
rect 257822 150818 258004 151054
rect 257404 150734 258004 150818
rect 257404 150498 257586 150734
rect 257822 150498 258004 150734
rect 257404 115054 258004 150498
rect 257404 114818 257586 115054
rect 257822 114818 258004 115054
rect 257404 114734 258004 114818
rect 257404 114498 257586 114734
rect 257822 114498 258004 114734
rect 257404 79054 258004 114498
rect 257404 78818 257586 79054
rect 257822 78818 258004 79054
rect 257404 78734 258004 78818
rect 257404 78498 257586 78734
rect 257822 78498 258004 78734
rect 257404 43054 258004 78498
rect 257404 42818 257586 43054
rect 257822 42818 258004 43054
rect 257404 42734 258004 42818
rect 257404 42498 257586 42734
rect 257822 42498 258004 42734
rect 257404 7054 258004 42498
rect 257404 6818 257586 7054
rect 257822 6818 258004 7054
rect 257404 6734 258004 6818
rect 257404 6498 257586 6734
rect 257822 6498 258004 6734
rect 257404 -2226 258004 6498
rect 257404 -2462 257586 -2226
rect 257822 -2462 258004 -2226
rect 257404 -2546 258004 -2462
rect 257404 -2782 257586 -2546
rect 257822 -2782 258004 -2546
rect 257404 -3744 258004 -2782
rect 261004 190654 261604 218000
rect 261004 190418 261186 190654
rect 261422 190418 261604 190654
rect 261004 190334 261604 190418
rect 261004 190098 261186 190334
rect 261422 190098 261604 190334
rect 261004 154654 261604 190098
rect 261004 154418 261186 154654
rect 261422 154418 261604 154654
rect 261004 154334 261604 154418
rect 261004 154098 261186 154334
rect 261422 154098 261604 154334
rect 261004 118654 261604 154098
rect 261004 118418 261186 118654
rect 261422 118418 261604 118654
rect 261004 118334 261604 118418
rect 261004 118098 261186 118334
rect 261422 118098 261604 118334
rect 261004 82654 261604 118098
rect 261004 82418 261186 82654
rect 261422 82418 261604 82654
rect 261004 82334 261604 82418
rect 261004 82098 261186 82334
rect 261422 82098 261604 82334
rect 261004 46654 261604 82098
rect 261004 46418 261186 46654
rect 261422 46418 261604 46654
rect 261004 46334 261604 46418
rect 261004 46098 261186 46334
rect 261422 46098 261604 46334
rect 261004 10654 261604 46098
rect 261004 10418 261186 10654
rect 261422 10418 261604 10654
rect 261004 10334 261604 10418
rect 261004 10098 261186 10334
rect 261422 10098 261604 10334
rect 261004 -4106 261604 10098
rect 261004 -4342 261186 -4106
rect 261422 -4342 261604 -4106
rect 261004 -4426 261604 -4342
rect 261004 -4662 261186 -4426
rect 261422 -4662 261604 -4426
rect 261004 -5624 261604 -4662
rect 264604 194254 265204 218000
rect 264604 194018 264786 194254
rect 265022 194018 265204 194254
rect 264604 193934 265204 194018
rect 264604 193698 264786 193934
rect 265022 193698 265204 193934
rect 264604 158254 265204 193698
rect 264604 158018 264786 158254
rect 265022 158018 265204 158254
rect 264604 157934 265204 158018
rect 264604 157698 264786 157934
rect 265022 157698 265204 157934
rect 264604 122254 265204 157698
rect 264604 122018 264786 122254
rect 265022 122018 265204 122254
rect 264604 121934 265204 122018
rect 264604 121698 264786 121934
rect 265022 121698 265204 121934
rect 264604 86254 265204 121698
rect 264604 86018 264786 86254
rect 265022 86018 265204 86254
rect 264604 85934 265204 86018
rect 264604 85698 264786 85934
rect 265022 85698 265204 85934
rect 264604 50254 265204 85698
rect 264604 50018 264786 50254
rect 265022 50018 265204 50254
rect 264604 49934 265204 50018
rect 264604 49698 264786 49934
rect 265022 49698 265204 49934
rect 264604 14254 265204 49698
rect 264604 14018 264786 14254
rect 265022 14018 265204 14254
rect 264604 13934 265204 14018
rect 264604 13698 264786 13934
rect 265022 13698 265204 13934
rect 246604 -7162 246786 -6926
rect 247022 -7162 247204 -6926
rect 246604 -7246 247204 -7162
rect 246604 -7482 246786 -7246
rect 247022 -7482 247204 -7246
rect 246604 -7504 247204 -7482
rect 264604 -5986 265204 13698
rect 271804 201454 272404 218000
rect 271804 201218 271986 201454
rect 272222 201218 272404 201454
rect 271804 201134 272404 201218
rect 271804 200898 271986 201134
rect 272222 200898 272404 201134
rect 271804 165454 272404 200898
rect 271804 165218 271986 165454
rect 272222 165218 272404 165454
rect 271804 165134 272404 165218
rect 271804 164898 271986 165134
rect 272222 164898 272404 165134
rect 271804 129454 272404 164898
rect 271804 129218 271986 129454
rect 272222 129218 272404 129454
rect 271804 129134 272404 129218
rect 271804 128898 271986 129134
rect 272222 128898 272404 129134
rect 271804 93454 272404 128898
rect 271804 93218 271986 93454
rect 272222 93218 272404 93454
rect 271804 93134 272404 93218
rect 271804 92898 271986 93134
rect 272222 92898 272404 93134
rect 271804 57454 272404 92898
rect 271804 57218 271986 57454
rect 272222 57218 272404 57454
rect 271804 57134 272404 57218
rect 271804 56898 271986 57134
rect 272222 56898 272404 57134
rect 271804 21454 272404 56898
rect 271804 21218 271986 21454
rect 272222 21218 272404 21454
rect 271804 21134 272404 21218
rect 271804 20898 271986 21134
rect 272222 20898 272404 21134
rect 271804 -1286 272404 20898
rect 271804 -1522 271986 -1286
rect 272222 -1522 272404 -1286
rect 271804 -1606 272404 -1522
rect 271804 -1842 271986 -1606
rect 272222 -1842 272404 -1606
rect 271804 -1864 272404 -1842
rect 275404 205054 276004 218000
rect 275404 204818 275586 205054
rect 275822 204818 276004 205054
rect 275404 204734 276004 204818
rect 275404 204498 275586 204734
rect 275822 204498 276004 204734
rect 275404 169054 276004 204498
rect 275404 168818 275586 169054
rect 275822 168818 276004 169054
rect 275404 168734 276004 168818
rect 275404 168498 275586 168734
rect 275822 168498 276004 168734
rect 275404 133054 276004 168498
rect 275404 132818 275586 133054
rect 275822 132818 276004 133054
rect 275404 132734 276004 132818
rect 275404 132498 275586 132734
rect 275822 132498 276004 132734
rect 275404 97054 276004 132498
rect 275404 96818 275586 97054
rect 275822 96818 276004 97054
rect 275404 96734 276004 96818
rect 275404 96498 275586 96734
rect 275822 96498 276004 96734
rect 275404 61054 276004 96498
rect 275404 60818 275586 61054
rect 275822 60818 276004 61054
rect 275404 60734 276004 60818
rect 275404 60498 275586 60734
rect 275822 60498 276004 60734
rect 275404 25054 276004 60498
rect 275404 24818 275586 25054
rect 275822 24818 276004 25054
rect 275404 24734 276004 24818
rect 275404 24498 275586 24734
rect 275822 24498 276004 24734
rect 275404 -3166 276004 24498
rect 275404 -3402 275586 -3166
rect 275822 -3402 276004 -3166
rect 275404 -3486 276004 -3402
rect 275404 -3722 275586 -3486
rect 275822 -3722 276004 -3486
rect 275404 -3744 276004 -3722
rect 279004 208654 279604 218000
rect 279004 208418 279186 208654
rect 279422 208418 279604 208654
rect 279004 208334 279604 208418
rect 279004 208098 279186 208334
rect 279422 208098 279604 208334
rect 279004 172654 279604 208098
rect 279004 172418 279186 172654
rect 279422 172418 279604 172654
rect 279004 172334 279604 172418
rect 279004 172098 279186 172334
rect 279422 172098 279604 172334
rect 279004 136654 279604 172098
rect 279004 136418 279186 136654
rect 279422 136418 279604 136654
rect 279004 136334 279604 136418
rect 279004 136098 279186 136334
rect 279422 136098 279604 136334
rect 279004 100654 279604 136098
rect 279004 100418 279186 100654
rect 279422 100418 279604 100654
rect 279004 100334 279604 100418
rect 279004 100098 279186 100334
rect 279422 100098 279604 100334
rect 279004 64654 279604 100098
rect 279004 64418 279186 64654
rect 279422 64418 279604 64654
rect 279004 64334 279604 64418
rect 279004 64098 279186 64334
rect 279422 64098 279604 64334
rect 279004 28654 279604 64098
rect 279004 28418 279186 28654
rect 279422 28418 279604 28654
rect 279004 28334 279604 28418
rect 279004 28098 279186 28334
rect 279422 28098 279604 28334
rect 279004 -5046 279604 28098
rect 279004 -5282 279186 -5046
rect 279422 -5282 279604 -5046
rect 279004 -5366 279604 -5282
rect 279004 -5602 279186 -5366
rect 279422 -5602 279604 -5366
rect 279004 -5624 279604 -5602
rect 282604 212254 283204 218000
rect 282604 212018 282786 212254
rect 283022 212018 283204 212254
rect 282604 211934 283204 212018
rect 282604 211698 282786 211934
rect 283022 211698 283204 211934
rect 282604 176254 283204 211698
rect 282604 176018 282786 176254
rect 283022 176018 283204 176254
rect 282604 175934 283204 176018
rect 282604 175698 282786 175934
rect 283022 175698 283204 175934
rect 282604 140254 283204 175698
rect 282604 140018 282786 140254
rect 283022 140018 283204 140254
rect 282604 139934 283204 140018
rect 282604 139698 282786 139934
rect 283022 139698 283204 139934
rect 282604 104254 283204 139698
rect 282604 104018 282786 104254
rect 283022 104018 283204 104254
rect 282604 103934 283204 104018
rect 282604 103698 282786 103934
rect 283022 103698 283204 103934
rect 282604 68254 283204 103698
rect 282604 68018 282786 68254
rect 283022 68018 283204 68254
rect 282604 67934 283204 68018
rect 282604 67698 282786 67934
rect 283022 67698 283204 67934
rect 282604 32254 283204 67698
rect 282604 32018 282786 32254
rect 283022 32018 283204 32254
rect 282604 31934 283204 32018
rect 282604 31698 282786 31934
rect 283022 31698 283204 31934
rect 264604 -6222 264786 -5986
rect 265022 -6222 265204 -5986
rect 264604 -6306 265204 -6222
rect 264604 -6542 264786 -6306
rect 265022 -6542 265204 -6306
rect 264604 -7504 265204 -6542
rect 282604 -6926 283204 31698
rect 289804 183454 290404 218000
rect 289804 183218 289986 183454
rect 290222 183218 290404 183454
rect 289804 183134 290404 183218
rect 289804 182898 289986 183134
rect 290222 182898 290404 183134
rect 289804 147454 290404 182898
rect 289804 147218 289986 147454
rect 290222 147218 290404 147454
rect 289804 147134 290404 147218
rect 289804 146898 289986 147134
rect 290222 146898 290404 147134
rect 289804 111454 290404 146898
rect 289804 111218 289986 111454
rect 290222 111218 290404 111454
rect 289804 111134 290404 111218
rect 289804 110898 289986 111134
rect 290222 110898 290404 111134
rect 289804 75454 290404 110898
rect 289804 75218 289986 75454
rect 290222 75218 290404 75454
rect 289804 75134 290404 75218
rect 289804 74898 289986 75134
rect 290222 74898 290404 75134
rect 289804 39454 290404 74898
rect 289804 39218 289986 39454
rect 290222 39218 290404 39454
rect 289804 39134 290404 39218
rect 289804 38898 289986 39134
rect 290222 38898 290404 39134
rect 289804 3454 290404 38898
rect 289804 3218 289986 3454
rect 290222 3218 290404 3454
rect 289804 3134 290404 3218
rect 289804 2898 289986 3134
rect 290222 2898 290404 3134
rect 289804 -346 290404 2898
rect 289804 -582 289986 -346
rect 290222 -582 290404 -346
rect 289804 -666 290404 -582
rect 289804 -902 289986 -666
rect 290222 -902 290404 -666
rect 289804 -1864 290404 -902
rect 293404 187054 294004 218000
rect 293404 186818 293586 187054
rect 293822 186818 294004 187054
rect 293404 186734 294004 186818
rect 293404 186498 293586 186734
rect 293822 186498 294004 186734
rect 293404 151054 294004 186498
rect 293404 150818 293586 151054
rect 293822 150818 294004 151054
rect 293404 150734 294004 150818
rect 293404 150498 293586 150734
rect 293822 150498 294004 150734
rect 293404 115054 294004 150498
rect 293404 114818 293586 115054
rect 293822 114818 294004 115054
rect 293404 114734 294004 114818
rect 293404 114498 293586 114734
rect 293822 114498 294004 114734
rect 293404 79054 294004 114498
rect 293404 78818 293586 79054
rect 293822 78818 294004 79054
rect 293404 78734 294004 78818
rect 293404 78498 293586 78734
rect 293822 78498 294004 78734
rect 293404 43054 294004 78498
rect 293404 42818 293586 43054
rect 293822 42818 294004 43054
rect 293404 42734 294004 42818
rect 293404 42498 293586 42734
rect 293822 42498 294004 42734
rect 293404 7054 294004 42498
rect 293404 6818 293586 7054
rect 293822 6818 294004 7054
rect 293404 6734 294004 6818
rect 293404 6498 293586 6734
rect 293822 6498 294004 6734
rect 293404 -2226 294004 6498
rect 293404 -2462 293586 -2226
rect 293822 -2462 294004 -2226
rect 293404 -2546 294004 -2462
rect 293404 -2782 293586 -2546
rect 293822 -2782 294004 -2546
rect 293404 -3744 294004 -2782
rect 297004 190654 297604 218000
rect 297004 190418 297186 190654
rect 297422 190418 297604 190654
rect 297004 190334 297604 190418
rect 297004 190098 297186 190334
rect 297422 190098 297604 190334
rect 297004 154654 297604 190098
rect 297004 154418 297186 154654
rect 297422 154418 297604 154654
rect 297004 154334 297604 154418
rect 297004 154098 297186 154334
rect 297422 154098 297604 154334
rect 297004 118654 297604 154098
rect 297004 118418 297186 118654
rect 297422 118418 297604 118654
rect 297004 118334 297604 118418
rect 297004 118098 297186 118334
rect 297422 118098 297604 118334
rect 297004 82654 297604 118098
rect 297004 82418 297186 82654
rect 297422 82418 297604 82654
rect 297004 82334 297604 82418
rect 297004 82098 297186 82334
rect 297422 82098 297604 82334
rect 297004 46654 297604 82098
rect 297004 46418 297186 46654
rect 297422 46418 297604 46654
rect 297004 46334 297604 46418
rect 297004 46098 297186 46334
rect 297422 46098 297604 46334
rect 297004 10654 297604 46098
rect 297004 10418 297186 10654
rect 297422 10418 297604 10654
rect 297004 10334 297604 10418
rect 297004 10098 297186 10334
rect 297422 10098 297604 10334
rect 297004 -4106 297604 10098
rect 297004 -4342 297186 -4106
rect 297422 -4342 297604 -4106
rect 297004 -4426 297604 -4342
rect 297004 -4662 297186 -4426
rect 297422 -4662 297604 -4426
rect 297004 -5624 297604 -4662
rect 300604 194254 301204 218000
rect 300604 194018 300786 194254
rect 301022 194018 301204 194254
rect 300604 193934 301204 194018
rect 300604 193698 300786 193934
rect 301022 193698 301204 193934
rect 300604 158254 301204 193698
rect 300604 158018 300786 158254
rect 301022 158018 301204 158254
rect 300604 157934 301204 158018
rect 300604 157698 300786 157934
rect 301022 157698 301204 157934
rect 300604 122254 301204 157698
rect 300604 122018 300786 122254
rect 301022 122018 301204 122254
rect 300604 121934 301204 122018
rect 300604 121698 300786 121934
rect 301022 121698 301204 121934
rect 300604 86254 301204 121698
rect 300604 86018 300786 86254
rect 301022 86018 301204 86254
rect 300604 85934 301204 86018
rect 300604 85698 300786 85934
rect 301022 85698 301204 85934
rect 300604 50254 301204 85698
rect 300604 50018 300786 50254
rect 301022 50018 301204 50254
rect 300604 49934 301204 50018
rect 300604 49698 300786 49934
rect 301022 49698 301204 49934
rect 300604 14254 301204 49698
rect 300604 14018 300786 14254
rect 301022 14018 301204 14254
rect 300604 13934 301204 14018
rect 300604 13698 300786 13934
rect 301022 13698 301204 13934
rect 282604 -7162 282786 -6926
rect 283022 -7162 283204 -6926
rect 282604 -7246 283204 -7162
rect 282604 -7482 282786 -7246
rect 283022 -7482 283204 -7246
rect 282604 -7504 283204 -7482
rect 300604 -5986 301204 13698
rect 307804 201454 308404 218000
rect 307804 201218 307986 201454
rect 308222 201218 308404 201454
rect 307804 201134 308404 201218
rect 307804 200898 307986 201134
rect 308222 200898 308404 201134
rect 307804 165454 308404 200898
rect 307804 165218 307986 165454
rect 308222 165218 308404 165454
rect 307804 165134 308404 165218
rect 307804 164898 307986 165134
rect 308222 164898 308404 165134
rect 307804 129454 308404 164898
rect 307804 129218 307986 129454
rect 308222 129218 308404 129454
rect 307804 129134 308404 129218
rect 307804 128898 307986 129134
rect 308222 128898 308404 129134
rect 307804 93454 308404 128898
rect 307804 93218 307986 93454
rect 308222 93218 308404 93454
rect 307804 93134 308404 93218
rect 307804 92898 307986 93134
rect 308222 92898 308404 93134
rect 307804 57454 308404 92898
rect 307804 57218 307986 57454
rect 308222 57218 308404 57454
rect 307804 57134 308404 57218
rect 307804 56898 307986 57134
rect 308222 56898 308404 57134
rect 307804 21454 308404 56898
rect 307804 21218 307986 21454
rect 308222 21218 308404 21454
rect 307804 21134 308404 21218
rect 307804 20898 307986 21134
rect 308222 20898 308404 21134
rect 307804 -1286 308404 20898
rect 307804 -1522 307986 -1286
rect 308222 -1522 308404 -1286
rect 307804 -1606 308404 -1522
rect 307804 -1842 307986 -1606
rect 308222 -1842 308404 -1606
rect 307804 -1864 308404 -1842
rect 311404 205054 312004 218000
rect 311404 204818 311586 205054
rect 311822 204818 312004 205054
rect 311404 204734 312004 204818
rect 311404 204498 311586 204734
rect 311822 204498 312004 204734
rect 311404 169054 312004 204498
rect 311404 168818 311586 169054
rect 311822 168818 312004 169054
rect 311404 168734 312004 168818
rect 311404 168498 311586 168734
rect 311822 168498 312004 168734
rect 311404 133054 312004 168498
rect 311404 132818 311586 133054
rect 311822 132818 312004 133054
rect 311404 132734 312004 132818
rect 311404 132498 311586 132734
rect 311822 132498 312004 132734
rect 311404 97054 312004 132498
rect 311404 96818 311586 97054
rect 311822 96818 312004 97054
rect 311404 96734 312004 96818
rect 311404 96498 311586 96734
rect 311822 96498 312004 96734
rect 311404 61054 312004 96498
rect 311404 60818 311586 61054
rect 311822 60818 312004 61054
rect 311404 60734 312004 60818
rect 311404 60498 311586 60734
rect 311822 60498 312004 60734
rect 311404 25054 312004 60498
rect 311404 24818 311586 25054
rect 311822 24818 312004 25054
rect 311404 24734 312004 24818
rect 311404 24498 311586 24734
rect 311822 24498 312004 24734
rect 311404 -3166 312004 24498
rect 311404 -3402 311586 -3166
rect 311822 -3402 312004 -3166
rect 311404 -3486 312004 -3402
rect 311404 -3722 311586 -3486
rect 311822 -3722 312004 -3486
rect 311404 -3744 312004 -3722
rect 315004 208654 315604 218000
rect 315004 208418 315186 208654
rect 315422 208418 315604 208654
rect 315004 208334 315604 208418
rect 315004 208098 315186 208334
rect 315422 208098 315604 208334
rect 315004 172654 315604 208098
rect 315004 172418 315186 172654
rect 315422 172418 315604 172654
rect 315004 172334 315604 172418
rect 315004 172098 315186 172334
rect 315422 172098 315604 172334
rect 315004 136654 315604 172098
rect 315004 136418 315186 136654
rect 315422 136418 315604 136654
rect 315004 136334 315604 136418
rect 315004 136098 315186 136334
rect 315422 136098 315604 136334
rect 315004 100654 315604 136098
rect 315004 100418 315186 100654
rect 315422 100418 315604 100654
rect 315004 100334 315604 100418
rect 315004 100098 315186 100334
rect 315422 100098 315604 100334
rect 315004 64654 315604 100098
rect 315004 64418 315186 64654
rect 315422 64418 315604 64654
rect 315004 64334 315604 64418
rect 315004 64098 315186 64334
rect 315422 64098 315604 64334
rect 315004 28654 315604 64098
rect 315004 28418 315186 28654
rect 315422 28418 315604 28654
rect 315004 28334 315604 28418
rect 315004 28098 315186 28334
rect 315422 28098 315604 28334
rect 315004 -5046 315604 28098
rect 315004 -5282 315186 -5046
rect 315422 -5282 315604 -5046
rect 315004 -5366 315604 -5282
rect 315004 -5602 315186 -5366
rect 315422 -5602 315604 -5366
rect 315004 -5624 315604 -5602
rect 318604 212254 319204 218000
rect 318604 212018 318786 212254
rect 319022 212018 319204 212254
rect 318604 211934 319204 212018
rect 318604 211698 318786 211934
rect 319022 211698 319204 211934
rect 318604 176254 319204 211698
rect 318604 176018 318786 176254
rect 319022 176018 319204 176254
rect 318604 175934 319204 176018
rect 318604 175698 318786 175934
rect 319022 175698 319204 175934
rect 318604 140254 319204 175698
rect 318604 140018 318786 140254
rect 319022 140018 319204 140254
rect 318604 139934 319204 140018
rect 318604 139698 318786 139934
rect 319022 139698 319204 139934
rect 318604 104254 319204 139698
rect 318604 104018 318786 104254
rect 319022 104018 319204 104254
rect 318604 103934 319204 104018
rect 318604 103698 318786 103934
rect 319022 103698 319204 103934
rect 318604 68254 319204 103698
rect 318604 68018 318786 68254
rect 319022 68018 319204 68254
rect 318604 67934 319204 68018
rect 318604 67698 318786 67934
rect 319022 67698 319204 67934
rect 318604 32254 319204 67698
rect 318604 32018 318786 32254
rect 319022 32018 319204 32254
rect 318604 31934 319204 32018
rect 318604 31698 318786 31934
rect 319022 31698 319204 31934
rect 300604 -6222 300786 -5986
rect 301022 -6222 301204 -5986
rect 300604 -6306 301204 -6222
rect 300604 -6542 300786 -6306
rect 301022 -6542 301204 -6306
rect 300604 -7504 301204 -6542
rect 318604 -6926 319204 31698
rect 325804 183454 326404 218000
rect 325804 183218 325986 183454
rect 326222 183218 326404 183454
rect 325804 183134 326404 183218
rect 325804 182898 325986 183134
rect 326222 182898 326404 183134
rect 325804 147454 326404 182898
rect 325804 147218 325986 147454
rect 326222 147218 326404 147454
rect 325804 147134 326404 147218
rect 325804 146898 325986 147134
rect 326222 146898 326404 147134
rect 325804 111454 326404 146898
rect 325804 111218 325986 111454
rect 326222 111218 326404 111454
rect 325804 111134 326404 111218
rect 325804 110898 325986 111134
rect 326222 110898 326404 111134
rect 325804 75454 326404 110898
rect 325804 75218 325986 75454
rect 326222 75218 326404 75454
rect 325804 75134 326404 75218
rect 325804 74898 325986 75134
rect 326222 74898 326404 75134
rect 325804 39454 326404 74898
rect 325804 39218 325986 39454
rect 326222 39218 326404 39454
rect 325804 39134 326404 39218
rect 325804 38898 325986 39134
rect 326222 38898 326404 39134
rect 325804 3454 326404 38898
rect 325804 3218 325986 3454
rect 326222 3218 326404 3454
rect 325804 3134 326404 3218
rect 325804 2898 325986 3134
rect 326222 2898 326404 3134
rect 325804 -346 326404 2898
rect 325804 -582 325986 -346
rect 326222 -582 326404 -346
rect 325804 -666 326404 -582
rect 325804 -902 325986 -666
rect 326222 -902 326404 -666
rect 325804 -1864 326404 -902
rect 329404 187054 330004 218000
rect 329404 186818 329586 187054
rect 329822 186818 330004 187054
rect 329404 186734 330004 186818
rect 329404 186498 329586 186734
rect 329822 186498 330004 186734
rect 329404 151054 330004 186498
rect 329404 150818 329586 151054
rect 329822 150818 330004 151054
rect 329404 150734 330004 150818
rect 329404 150498 329586 150734
rect 329822 150498 330004 150734
rect 329404 115054 330004 150498
rect 329404 114818 329586 115054
rect 329822 114818 330004 115054
rect 329404 114734 330004 114818
rect 329404 114498 329586 114734
rect 329822 114498 330004 114734
rect 329404 79054 330004 114498
rect 329404 78818 329586 79054
rect 329822 78818 330004 79054
rect 329404 78734 330004 78818
rect 329404 78498 329586 78734
rect 329822 78498 330004 78734
rect 329404 43054 330004 78498
rect 329404 42818 329586 43054
rect 329822 42818 330004 43054
rect 329404 42734 330004 42818
rect 329404 42498 329586 42734
rect 329822 42498 330004 42734
rect 329404 7054 330004 42498
rect 329404 6818 329586 7054
rect 329822 6818 330004 7054
rect 329404 6734 330004 6818
rect 329404 6498 329586 6734
rect 329822 6498 330004 6734
rect 329404 -2226 330004 6498
rect 329404 -2462 329586 -2226
rect 329822 -2462 330004 -2226
rect 329404 -2546 330004 -2462
rect 329404 -2782 329586 -2546
rect 329822 -2782 330004 -2546
rect 329404 -3744 330004 -2782
rect 333004 190654 333604 218000
rect 333004 190418 333186 190654
rect 333422 190418 333604 190654
rect 333004 190334 333604 190418
rect 333004 190098 333186 190334
rect 333422 190098 333604 190334
rect 333004 154654 333604 190098
rect 333004 154418 333186 154654
rect 333422 154418 333604 154654
rect 333004 154334 333604 154418
rect 333004 154098 333186 154334
rect 333422 154098 333604 154334
rect 333004 118654 333604 154098
rect 333004 118418 333186 118654
rect 333422 118418 333604 118654
rect 333004 118334 333604 118418
rect 333004 118098 333186 118334
rect 333422 118098 333604 118334
rect 333004 82654 333604 118098
rect 333004 82418 333186 82654
rect 333422 82418 333604 82654
rect 333004 82334 333604 82418
rect 333004 82098 333186 82334
rect 333422 82098 333604 82334
rect 333004 46654 333604 82098
rect 333004 46418 333186 46654
rect 333422 46418 333604 46654
rect 333004 46334 333604 46418
rect 333004 46098 333186 46334
rect 333422 46098 333604 46334
rect 333004 10654 333604 46098
rect 333004 10418 333186 10654
rect 333422 10418 333604 10654
rect 333004 10334 333604 10418
rect 333004 10098 333186 10334
rect 333422 10098 333604 10334
rect 333004 -4106 333604 10098
rect 333004 -4342 333186 -4106
rect 333422 -4342 333604 -4106
rect 333004 -4426 333604 -4342
rect 333004 -4662 333186 -4426
rect 333422 -4662 333604 -4426
rect 333004 -5624 333604 -4662
rect 336604 194254 337204 218000
rect 336604 194018 336786 194254
rect 337022 194018 337204 194254
rect 336604 193934 337204 194018
rect 336604 193698 336786 193934
rect 337022 193698 337204 193934
rect 336604 158254 337204 193698
rect 336604 158018 336786 158254
rect 337022 158018 337204 158254
rect 336604 157934 337204 158018
rect 336604 157698 336786 157934
rect 337022 157698 337204 157934
rect 336604 122254 337204 157698
rect 336604 122018 336786 122254
rect 337022 122018 337204 122254
rect 336604 121934 337204 122018
rect 336604 121698 336786 121934
rect 337022 121698 337204 121934
rect 336604 86254 337204 121698
rect 336604 86018 336786 86254
rect 337022 86018 337204 86254
rect 336604 85934 337204 86018
rect 336604 85698 336786 85934
rect 337022 85698 337204 85934
rect 336604 50254 337204 85698
rect 336604 50018 336786 50254
rect 337022 50018 337204 50254
rect 336604 49934 337204 50018
rect 336604 49698 336786 49934
rect 337022 49698 337204 49934
rect 336604 14254 337204 49698
rect 336604 14018 336786 14254
rect 337022 14018 337204 14254
rect 336604 13934 337204 14018
rect 336604 13698 336786 13934
rect 337022 13698 337204 13934
rect 318604 -7162 318786 -6926
rect 319022 -7162 319204 -6926
rect 318604 -7246 319204 -7162
rect 318604 -7482 318786 -7246
rect 319022 -7482 319204 -7246
rect 318604 -7504 319204 -7482
rect 336604 -5986 337204 13698
rect 343804 201454 344404 218000
rect 343804 201218 343986 201454
rect 344222 201218 344404 201454
rect 343804 201134 344404 201218
rect 343804 200898 343986 201134
rect 344222 200898 344404 201134
rect 343804 165454 344404 200898
rect 343804 165218 343986 165454
rect 344222 165218 344404 165454
rect 343804 165134 344404 165218
rect 343804 164898 343986 165134
rect 344222 164898 344404 165134
rect 343804 129454 344404 164898
rect 343804 129218 343986 129454
rect 344222 129218 344404 129454
rect 343804 129134 344404 129218
rect 343804 128898 343986 129134
rect 344222 128898 344404 129134
rect 343804 93454 344404 128898
rect 343804 93218 343986 93454
rect 344222 93218 344404 93454
rect 343804 93134 344404 93218
rect 343804 92898 343986 93134
rect 344222 92898 344404 93134
rect 343804 57454 344404 92898
rect 343804 57218 343986 57454
rect 344222 57218 344404 57454
rect 343804 57134 344404 57218
rect 343804 56898 343986 57134
rect 344222 56898 344404 57134
rect 343804 21454 344404 56898
rect 343804 21218 343986 21454
rect 344222 21218 344404 21454
rect 343804 21134 344404 21218
rect 343804 20898 343986 21134
rect 344222 20898 344404 21134
rect 343804 -1286 344404 20898
rect 343804 -1522 343986 -1286
rect 344222 -1522 344404 -1286
rect 343804 -1606 344404 -1522
rect 343804 -1842 343986 -1606
rect 344222 -1842 344404 -1606
rect 343804 -1864 344404 -1842
rect 347404 205054 348004 218000
rect 347404 204818 347586 205054
rect 347822 204818 348004 205054
rect 347404 204734 348004 204818
rect 347404 204498 347586 204734
rect 347822 204498 348004 204734
rect 347404 169054 348004 204498
rect 347404 168818 347586 169054
rect 347822 168818 348004 169054
rect 347404 168734 348004 168818
rect 347404 168498 347586 168734
rect 347822 168498 348004 168734
rect 347404 133054 348004 168498
rect 347404 132818 347586 133054
rect 347822 132818 348004 133054
rect 347404 132734 348004 132818
rect 347404 132498 347586 132734
rect 347822 132498 348004 132734
rect 347404 97054 348004 132498
rect 347404 96818 347586 97054
rect 347822 96818 348004 97054
rect 347404 96734 348004 96818
rect 347404 96498 347586 96734
rect 347822 96498 348004 96734
rect 347404 61054 348004 96498
rect 347404 60818 347586 61054
rect 347822 60818 348004 61054
rect 347404 60734 348004 60818
rect 347404 60498 347586 60734
rect 347822 60498 348004 60734
rect 347404 25054 348004 60498
rect 347404 24818 347586 25054
rect 347822 24818 348004 25054
rect 347404 24734 348004 24818
rect 347404 24498 347586 24734
rect 347822 24498 348004 24734
rect 347404 -3166 348004 24498
rect 347404 -3402 347586 -3166
rect 347822 -3402 348004 -3166
rect 347404 -3486 348004 -3402
rect 347404 -3722 347586 -3486
rect 347822 -3722 348004 -3486
rect 347404 -3744 348004 -3722
rect 351004 208654 351604 218000
rect 351004 208418 351186 208654
rect 351422 208418 351604 208654
rect 351004 208334 351604 208418
rect 351004 208098 351186 208334
rect 351422 208098 351604 208334
rect 351004 172654 351604 208098
rect 351004 172418 351186 172654
rect 351422 172418 351604 172654
rect 351004 172334 351604 172418
rect 351004 172098 351186 172334
rect 351422 172098 351604 172334
rect 351004 136654 351604 172098
rect 351004 136418 351186 136654
rect 351422 136418 351604 136654
rect 351004 136334 351604 136418
rect 351004 136098 351186 136334
rect 351422 136098 351604 136334
rect 351004 100654 351604 136098
rect 351004 100418 351186 100654
rect 351422 100418 351604 100654
rect 351004 100334 351604 100418
rect 351004 100098 351186 100334
rect 351422 100098 351604 100334
rect 351004 64654 351604 100098
rect 351004 64418 351186 64654
rect 351422 64418 351604 64654
rect 351004 64334 351604 64418
rect 351004 64098 351186 64334
rect 351422 64098 351604 64334
rect 351004 28654 351604 64098
rect 351004 28418 351186 28654
rect 351422 28418 351604 28654
rect 351004 28334 351604 28418
rect 351004 28098 351186 28334
rect 351422 28098 351604 28334
rect 351004 -5046 351604 28098
rect 351004 -5282 351186 -5046
rect 351422 -5282 351604 -5046
rect 351004 -5366 351604 -5282
rect 351004 -5602 351186 -5366
rect 351422 -5602 351604 -5366
rect 351004 -5624 351604 -5602
rect 354604 212254 355204 218000
rect 354604 212018 354786 212254
rect 355022 212018 355204 212254
rect 354604 211934 355204 212018
rect 354604 211698 354786 211934
rect 355022 211698 355204 211934
rect 354604 176254 355204 211698
rect 354604 176018 354786 176254
rect 355022 176018 355204 176254
rect 354604 175934 355204 176018
rect 354604 175698 354786 175934
rect 355022 175698 355204 175934
rect 354604 140254 355204 175698
rect 354604 140018 354786 140254
rect 355022 140018 355204 140254
rect 354604 139934 355204 140018
rect 354604 139698 354786 139934
rect 355022 139698 355204 139934
rect 354604 104254 355204 139698
rect 354604 104018 354786 104254
rect 355022 104018 355204 104254
rect 354604 103934 355204 104018
rect 354604 103698 354786 103934
rect 355022 103698 355204 103934
rect 354604 68254 355204 103698
rect 354604 68018 354786 68254
rect 355022 68018 355204 68254
rect 354604 67934 355204 68018
rect 354604 67698 354786 67934
rect 355022 67698 355204 67934
rect 354604 32254 355204 67698
rect 354604 32018 354786 32254
rect 355022 32018 355204 32254
rect 354604 31934 355204 32018
rect 354604 31698 354786 31934
rect 355022 31698 355204 31934
rect 336604 -6222 336786 -5986
rect 337022 -6222 337204 -5986
rect 336604 -6306 337204 -6222
rect 336604 -6542 336786 -6306
rect 337022 -6542 337204 -6306
rect 336604 -7504 337204 -6542
rect 354604 -6926 355204 31698
rect 361804 183454 362404 218000
rect 361804 183218 361986 183454
rect 362222 183218 362404 183454
rect 361804 183134 362404 183218
rect 361804 182898 361986 183134
rect 362222 182898 362404 183134
rect 361804 147454 362404 182898
rect 361804 147218 361986 147454
rect 362222 147218 362404 147454
rect 361804 147134 362404 147218
rect 361804 146898 361986 147134
rect 362222 146898 362404 147134
rect 361804 111454 362404 146898
rect 361804 111218 361986 111454
rect 362222 111218 362404 111454
rect 361804 111134 362404 111218
rect 361804 110898 361986 111134
rect 362222 110898 362404 111134
rect 361804 75454 362404 110898
rect 361804 75218 361986 75454
rect 362222 75218 362404 75454
rect 361804 75134 362404 75218
rect 361804 74898 361986 75134
rect 362222 74898 362404 75134
rect 361804 39454 362404 74898
rect 361804 39218 361986 39454
rect 362222 39218 362404 39454
rect 361804 39134 362404 39218
rect 361804 38898 361986 39134
rect 362222 38898 362404 39134
rect 361804 3454 362404 38898
rect 361804 3218 361986 3454
rect 362222 3218 362404 3454
rect 361804 3134 362404 3218
rect 361804 2898 361986 3134
rect 362222 2898 362404 3134
rect 361804 -346 362404 2898
rect 361804 -582 361986 -346
rect 362222 -582 362404 -346
rect 361804 -666 362404 -582
rect 361804 -902 361986 -666
rect 362222 -902 362404 -666
rect 361804 -1864 362404 -902
rect 365404 187054 366004 218000
rect 365404 186818 365586 187054
rect 365822 186818 366004 187054
rect 365404 186734 366004 186818
rect 365404 186498 365586 186734
rect 365822 186498 366004 186734
rect 365404 151054 366004 186498
rect 365404 150818 365586 151054
rect 365822 150818 366004 151054
rect 365404 150734 366004 150818
rect 365404 150498 365586 150734
rect 365822 150498 366004 150734
rect 365404 115054 366004 150498
rect 365404 114818 365586 115054
rect 365822 114818 366004 115054
rect 365404 114734 366004 114818
rect 365404 114498 365586 114734
rect 365822 114498 366004 114734
rect 365404 79054 366004 114498
rect 365404 78818 365586 79054
rect 365822 78818 366004 79054
rect 365404 78734 366004 78818
rect 365404 78498 365586 78734
rect 365822 78498 366004 78734
rect 365404 43054 366004 78498
rect 365404 42818 365586 43054
rect 365822 42818 366004 43054
rect 365404 42734 366004 42818
rect 365404 42498 365586 42734
rect 365822 42498 366004 42734
rect 365404 7054 366004 42498
rect 365404 6818 365586 7054
rect 365822 6818 366004 7054
rect 365404 6734 366004 6818
rect 365404 6498 365586 6734
rect 365822 6498 366004 6734
rect 365404 -2226 366004 6498
rect 365404 -2462 365586 -2226
rect 365822 -2462 366004 -2226
rect 365404 -2546 366004 -2462
rect 365404 -2782 365586 -2546
rect 365822 -2782 366004 -2546
rect 365404 -3744 366004 -2782
rect 369004 190654 369604 218000
rect 369004 190418 369186 190654
rect 369422 190418 369604 190654
rect 369004 190334 369604 190418
rect 369004 190098 369186 190334
rect 369422 190098 369604 190334
rect 369004 154654 369604 190098
rect 369004 154418 369186 154654
rect 369422 154418 369604 154654
rect 369004 154334 369604 154418
rect 369004 154098 369186 154334
rect 369422 154098 369604 154334
rect 369004 118654 369604 154098
rect 369004 118418 369186 118654
rect 369422 118418 369604 118654
rect 369004 118334 369604 118418
rect 369004 118098 369186 118334
rect 369422 118098 369604 118334
rect 369004 82654 369604 118098
rect 369004 82418 369186 82654
rect 369422 82418 369604 82654
rect 369004 82334 369604 82418
rect 369004 82098 369186 82334
rect 369422 82098 369604 82334
rect 369004 46654 369604 82098
rect 369004 46418 369186 46654
rect 369422 46418 369604 46654
rect 369004 46334 369604 46418
rect 369004 46098 369186 46334
rect 369422 46098 369604 46334
rect 369004 10654 369604 46098
rect 369004 10418 369186 10654
rect 369422 10418 369604 10654
rect 369004 10334 369604 10418
rect 369004 10098 369186 10334
rect 369422 10098 369604 10334
rect 369004 -4106 369604 10098
rect 369004 -4342 369186 -4106
rect 369422 -4342 369604 -4106
rect 369004 -4426 369604 -4342
rect 369004 -4662 369186 -4426
rect 369422 -4662 369604 -4426
rect 369004 -5624 369604 -4662
rect 372604 194254 373204 218000
rect 372604 194018 372786 194254
rect 373022 194018 373204 194254
rect 372604 193934 373204 194018
rect 372604 193698 372786 193934
rect 373022 193698 373204 193934
rect 372604 158254 373204 193698
rect 372604 158018 372786 158254
rect 373022 158018 373204 158254
rect 372604 157934 373204 158018
rect 372604 157698 372786 157934
rect 373022 157698 373204 157934
rect 372604 122254 373204 157698
rect 372604 122018 372786 122254
rect 373022 122018 373204 122254
rect 372604 121934 373204 122018
rect 372604 121698 372786 121934
rect 373022 121698 373204 121934
rect 372604 86254 373204 121698
rect 372604 86018 372786 86254
rect 373022 86018 373204 86254
rect 372604 85934 373204 86018
rect 372604 85698 372786 85934
rect 373022 85698 373204 85934
rect 372604 50254 373204 85698
rect 372604 50018 372786 50254
rect 373022 50018 373204 50254
rect 372604 49934 373204 50018
rect 372604 49698 372786 49934
rect 373022 49698 373204 49934
rect 372604 14254 373204 49698
rect 372604 14018 372786 14254
rect 373022 14018 373204 14254
rect 372604 13934 373204 14018
rect 372604 13698 372786 13934
rect 373022 13698 373204 13934
rect 354604 -7162 354786 -6926
rect 355022 -7162 355204 -6926
rect 354604 -7246 355204 -7162
rect 354604 -7482 354786 -7246
rect 355022 -7482 355204 -7246
rect 354604 -7504 355204 -7482
rect 372604 -5986 373204 13698
rect 379804 201454 380404 218000
rect 379804 201218 379986 201454
rect 380222 201218 380404 201454
rect 379804 201134 380404 201218
rect 379804 200898 379986 201134
rect 380222 200898 380404 201134
rect 379804 165454 380404 200898
rect 379804 165218 379986 165454
rect 380222 165218 380404 165454
rect 379804 165134 380404 165218
rect 379804 164898 379986 165134
rect 380222 164898 380404 165134
rect 379804 129454 380404 164898
rect 379804 129218 379986 129454
rect 380222 129218 380404 129454
rect 379804 129134 380404 129218
rect 379804 128898 379986 129134
rect 380222 128898 380404 129134
rect 379804 93454 380404 128898
rect 379804 93218 379986 93454
rect 380222 93218 380404 93454
rect 379804 93134 380404 93218
rect 379804 92898 379986 93134
rect 380222 92898 380404 93134
rect 379804 57454 380404 92898
rect 379804 57218 379986 57454
rect 380222 57218 380404 57454
rect 379804 57134 380404 57218
rect 379804 56898 379986 57134
rect 380222 56898 380404 57134
rect 379804 21454 380404 56898
rect 379804 21218 379986 21454
rect 380222 21218 380404 21454
rect 379804 21134 380404 21218
rect 379804 20898 379986 21134
rect 380222 20898 380404 21134
rect 379804 -1286 380404 20898
rect 379804 -1522 379986 -1286
rect 380222 -1522 380404 -1286
rect 379804 -1606 380404 -1522
rect 379804 -1842 379986 -1606
rect 380222 -1842 380404 -1606
rect 379804 -1864 380404 -1842
rect 383404 205054 384004 218000
rect 383404 204818 383586 205054
rect 383822 204818 384004 205054
rect 383404 204734 384004 204818
rect 383404 204498 383586 204734
rect 383822 204498 384004 204734
rect 383404 169054 384004 204498
rect 383404 168818 383586 169054
rect 383822 168818 384004 169054
rect 383404 168734 384004 168818
rect 383404 168498 383586 168734
rect 383822 168498 384004 168734
rect 383404 133054 384004 168498
rect 383404 132818 383586 133054
rect 383822 132818 384004 133054
rect 383404 132734 384004 132818
rect 383404 132498 383586 132734
rect 383822 132498 384004 132734
rect 383404 97054 384004 132498
rect 383404 96818 383586 97054
rect 383822 96818 384004 97054
rect 383404 96734 384004 96818
rect 383404 96498 383586 96734
rect 383822 96498 384004 96734
rect 383404 61054 384004 96498
rect 383404 60818 383586 61054
rect 383822 60818 384004 61054
rect 383404 60734 384004 60818
rect 383404 60498 383586 60734
rect 383822 60498 384004 60734
rect 383404 25054 384004 60498
rect 383404 24818 383586 25054
rect 383822 24818 384004 25054
rect 383404 24734 384004 24818
rect 383404 24498 383586 24734
rect 383822 24498 384004 24734
rect 383404 -3166 384004 24498
rect 383404 -3402 383586 -3166
rect 383822 -3402 384004 -3166
rect 383404 -3486 384004 -3402
rect 383404 -3722 383586 -3486
rect 383822 -3722 384004 -3486
rect 383404 -3744 384004 -3722
rect 387004 208654 387604 218000
rect 387004 208418 387186 208654
rect 387422 208418 387604 208654
rect 387004 208334 387604 208418
rect 387004 208098 387186 208334
rect 387422 208098 387604 208334
rect 387004 172654 387604 208098
rect 387004 172418 387186 172654
rect 387422 172418 387604 172654
rect 387004 172334 387604 172418
rect 387004 172098 387186 172334
rect 387422 172098 387604 172334
rect 387004 136654 387604 172098
rect 387004 136418 387186 136654
rect 387422 136418 387604 136654
rect 387004 136334 387604 136418
rect 387004 136098 387186 136334
rect 387422 136098 387604 136334
rect 387004 100654 387604 136098
rect 387004 100418 387186 100654
rect 387422 100418 387604 100654
rect 387004 100334 387604 100418
rect 387004 100098 387186 100334
rect 387422 100098 387604 100334
rect 387004 64654 387604 100098
rect 387004 64418 387186 64654
rect 387422 64418 387604 64654
rect 387004 64334 387604 64418
rect 387004 64098 387186 64334
rect 387422 64098 387604 64334
rect 387004 28654 387604 64098
rect 389774 31789 389834 344387
rect 407589 312960 418408 348656
rect 407589 312946 416821 312960
rect 407589 312931 415412 312946
rect 407589 312917 414011 312931
rect 407589 312902 412602 312917
rect 407589 312888 411122 312902
rect 407589 312873 409713 312888
rect 407589 312859 408312 312873
rect 407589 312623 407917 312859
rect 408153 312637 408312 312859
rect 408548 312637 408632 312873
rect 408868 312637 409006 312873
rect 409242 312637 409326 312873
rect 409562 312652 409713 312873
rect 409949 312652 410033 312888
rect 410269 312652 410407 312888
rect 410643 312652 410727 312888
rect 410963 312666 411122 312888
rect 411358 312666 411442 312902
rect 411678 312666 411816 312902
rect 412052 312666 412136 312902
rect 412372 312681 412602 312902
rect 412838 312681 412922 312917
rect 413158 312681 413296 312917
rect 413532 312681 413616 312917
rect 413852 312695 414011 312917
rect 414247 312695 414331 312931
rect 414567 312695 414705 312931
rect 414941 312695 415025 312931
rect 415261 312710 415412 312931
rect 415648 312710 415732 312946
rect 415968 312710 416106 312946
rect 416342 312710 416426 312946
rect 416662 312724 416821 312946
rect 417057 312724 417141 312960
rect 417377 312724 417515 312960
rect 417751 312724 417835 312960
rect 418071 312724 418408 312960
rect 416662 312710 418408 312724
rect 415261 312695 418408 312710
rect 413852 312681 418408 312695
rect 412372 312666 418408 312681
rect 410963 312652 418408 312666
rect 409562 312637 418408 312652
rect 408153 312623 418408 312637
rect 407589 276941 418408 312623
rect 407589 276927 416796 276941
rect 407589 276912 415387 276927
rect 407589 276898 413986 276912
rect 407589 276883 412577 276898
rect 407589 276869 411097 276883
rect 407589 276854 409688 276869
rect 407589 276840 408287 276854
rect 407589 276604 407892 276840
rect 408128 276618 408287 276840
rect 408523 276618 408607 276854
rect 408843 276618 408981 276854
rect 409217 276618 409301 276854
rect 409537 276633 409688 276854
rect 409924 276633 410008 276869
rect 410244 276633 410382 276869
rect 410618 276633 410702 276869
rect 410938 276647 411097 276869
rect 411333 276647 411417 276883
rect 411653 276647 411791 276883
rect 412027 276647 412111 276883
rect 412347 276662 412577 276883
rect 412813 276662 412897 276898
rect 413133 276662 413271 276898
rect 413507 276662 413591 276898
rect 413827 276676 413986 276898
rect 414222 276676 414306 276912
rect 414542 276676 414680 276912
rect 414916 276676 415000 276912
rect 415236 276691 415387 276912
rect 415623 276691 415707 276927
rect 415943 276691 416081 276927
rect 416317 276691 416401 276927
rect 416637 276705 416796 276927
rect 417032 276705 417116 276941
rect 417352 276705 417490 276941
rect 417726 276705 417810 276941
rect 418046 276705 418408 276941
rect 416637 276691 418408 276705
rect 415236 276676 418408 276691
rect 413827 276662 418408 276676
rect 412347 276647 418408 276662
rect 410938 276633 418408 276647
rect 409537 276618 418408 276633
rect 408128 276604 418408 276618
rect 407589 240943 418408 276604
rect 407589 240929 416782 240943
rect 407589 240914 415373 240929
rect 407589 240900 413972 240914
rect 407589 240885 412563 240900
rect 407589 240871 411083 240885
rect 407589 240856 409674 240871
rect 407589 240842 408273 240856
rect 407589 240606 407878 240842
rect 408114 240620 408273 240842
rect 408509 240620 408593 240856
rect 408829 240620 408967 240856
rect 409203 240620 409287 240856
rect 409523 240635 409674 240856
rect 409910 240635 409994 240871
rect 410230 240635 410368 240871
rect 410604 240635 410688 240871
rect 410924 240649 411083 240871
rect 411319 240649 411403 240885
rect 411639 240649 411777 240885
rect 412013 240649 412097 240885
rect 412333 240664 412563 240885
rect 412799 240664 412883 240900
rect 413119 240664 413257 240900
rect 413493 240664 413577 240900
rect 413813 240678 413972 240900
rect 414208 240678 414292 240914
rect 414528 240678 414666 240914
rect 414902 240678 414986 240914
rect 415222 240693 415373 240914
rect 415609 240693 415693 240929
rect 415929 240693 416067 240929
rect 416303 240693 416387 240929
rect 416623 240707 416782 240929
rect 417018 240707 417102 240943
rect 417338 240707 417476 240943
rect 417712 240707 417796 240943
rect 418032 240707 418408 240943
rect 416623 240693 418408 240707
rect 415222 240678 418408 240693
rect 413813 240664 418408 240678
rect 412333 240649 418408 240664
rect 410924 240635 418408 240649
rect 409523 240620 418408 240635
rect 408114 240606 418408 240620
rect 407589 234520 418408 240606
rect 425267 561359 436086 574520
rect 425267 561345 434457 561359
rect 425267 561330 433048 561345
rect 425267 561316 431647 561330
rect 425267 561301 430238 561316
rect 425267 561287 428758 561301
rect 425267 561272 427349 561287
rect 425267 561258 425948 561272
rect 425267 561022 425553 561258
rect 425789 561036 425948 561258
rect 426184 561036 426268 561272
rect 426504 561036 426642 561272
rect 426878 561036 426962 561272
rect 427198 561051 427349 561272
rect 427585 561051 427669 561287
rect 427905 561051 428043 561287
rect 428279 561051 428363 561287
rect 428599 561065 428758 561287
rect 428994 561065 429078 561301
rect 429314 561065 429452 561301
rect 429688 561065 429772 561301
rect 430008 561080 430238 561301
rect 430474 561080 430558 561316
rect 430794 561080 430932 561316
rect 431168 561080 431252 561316
rect 431488 561094 431647 561316
rect 431883 561094 431967 561330
rect 432203 561094 432341 561330
rect 432577 561094 432661 561330
rect 432897 561109 433048 561330
rect 433284 561109 433368 561345
rect 433604 561109 433742 561345
rect 433978 561109 434062 561345
rect 434298 561123 434457 561345
rect 434693 561123 434777 561359
rect 435013 561123 435151 561359
rect 435387 561123 435471 561359
rect 435707 561123 436086 561359
rect 434298 561109 436086 561123
rect 432897 561094 436086 561109
rect 431488 561080 436086 561094
rect 430008 561065 436086 561080
rect 428599 561051 436086 561065
rect 427198 561036 436086 561051
rect 425789 561022 436086 561036
rect 425267 525366 436086 561022
rect 425267 525352 434596 525366
rect 425267 525337 433187 525352
rect 425267 525323 431786 525337
rect 425267 525308 430377 525323
rect 425267 525294 428897 525308
rect 425267 525279 427488 525294
rect 425267 525265 426087 525279
rect 425267 525029 425692 525265
rect 425928 525043 426087 525265
rect 426323 525043 426407 525279
rect 426643 525043 426781 525279
rect 427017 525043 427101 525279
rect 427337 525058 427488 525279
rect 427724 525058 427808 525294
rect 428044 525058 428182 525294
rect 428418 525058 428502 525294
rect 428738 525072 428897 525294
rect 429133 525072 429217 525308
rect 429453 525072 429591 525308
rect 429827 525072 429911 525308
rect 430147 525087 430377 525308
rect 430613 525087 430697 525323
rect 430933 525087 431071 525323
rect 431307 525087 431391 525323
rect 431627 525101 431786 525323
rect 432022 525101 432106 525337
rect 432342 525101 432480 525337
rect 432716 525101 432800 525337
rect 433036 525116 433187 525337
rect 433423 525116 433507 525352
rect 433743 525116 433881 525352
rect 434117 525116 434201 525352
rect 434437 525130 434596 525352
rect 434832 525130 434916 525366
rect 435152 525130 435290 525366
rect 435526 525130 435610 525366
rect 435846 525130 436086 525366
rect 434437 525116 436086 525130
rect 433036 525101 436086 525116
rect 431627 525087 436086 525101
rect 430147 525072 436086 525087
rect 428738 525058 436086 525072
rect 427337 525043 436086 525058
rect 425928 525029 436086 525043
rect 425267 489373 436086 525029
rect 425267 489359 434595 489373
rect 425267 489344 433186 489359
rect 425267 489330 431785 489344
rect 425267 489315 430376 489330
rect 425267 489301 428896 489315
rect 425267 489286 427487 489301
rect 425267 489272 426086 489286
rect 425267 489036 425691 489272
rect 425927 489050 426086 489272
rect 426322 489050 426406 489286
rect 426642 489050 426780 489286
rect 427016 489050 427100 489286
rect 427336 489065 427487 489286
rect 427723 489065 427807 489301
rect 428043 489065 428181 489301
rect 428417 489065 428501 489301
rect 428737 489079 428896 489301
rect 429132 489079 429216 489315
rect 429452 489079 429590 489315
rect 429826 489079 429910 489315
rect 430146 489094 430376 489315
rect 430612 489094 430696 489330
rect 430932 489094 431070 489330
rect 431306 489094 431390 489330
rect 431626 489108 431785 489330
rect 432021 489108 432105 489344
rect 432341 489108 432479 489344
rect 432715 489108 432799 489344
rect 433035 489123 433186 489344
rect 433422 489123 433506 489359
rect 433742 489123 433880 489359
rect 434116 489123 434200 489359
rect 434436 489137 434595 489359
rect 434831 489137 434915 489373
rect 435151 489137 435289 489373
rect 435525 489137 435609 489373
rect 435845 489137 436086 489373
rect 434436 489123 436086 489137
rect 433035 489108 436086 489123
rect 431626 489094 436086 489108
rect 430146 489079 436086 489094
rect 428737 489065 436086 489079
rect 427336 489050 436086 489065
rect 425927 489036 436086 489050
rect 425267 467943 436086 489036
rect 425267 467929 434602 467943
rect 425267 467914 433193 467929
rect 425267 467900 431792 467914
rect 425267 467885 430383 467900
rect 425267 467871 428903 467885
rect 425267 467856 427494 467871
rect 425267 467842 426093 467856
rect 425267 467606 425698 467842
rect 425934 467606 426093 467842
rect 425267 467522 426093 467606
rect 425267 467286 425698 467522
rect 425934 467286 426093 467522
rect 425267 467202 426093 467286
rect 425267 466966 425698 467202
rect 425934 466980 426093 467202
rect 426649 466980 426787 467856
rect 427343 466995 427494 467856
rect 428050 466995 428188 467871
rect 428744 467009 428903 467871
rect 429459 467009 429597 467885
rect 430153 467024 430383 467885
rect 430939 467024 431077 467900
rect 431633 467038 431792 467900
rect 432348 467038 432486 467914
rect 433042 467053 433193 467914
rect 433749 467053 433887 467929
rect 434443 467067 434602 467929
rect 435158 467067 435296 467943
rect 435852 467067 436086 467943
rect 434443 467053 436086 467067
rect 433042 467038 436086 467053
rect 431633 467024 436086 467038
rect 430153 467009 436086 467024
rect 428744 466995 436086 467009
rect 427343 466980 436086 466995
rect 425934 466966 436086 466980
rect 425267 451956 436086 466966
rect 425267 451942 434479 451956
rect 425267 451927 433070 451942
rect 425267 451913 431669 451927
rect 425267 451898 430260 451913
rect 425267 451884 428780 451898
rect 425267 451869 427371 451884
rect 425267 451855 425970 451869
rect 425267 451619 425575 451855
rect 425811 451619 425970 451855
rect 425267 451535 425970 451619
rect 425267 451299 425575 451535
rect 425811 451299 425970 451535
rect 425267 451215 425970 451299
rect 425267 450979 425575 451215
rect 425811 450993 425970 451215
rect 426526 450993 426664 451869
rect 427220 451008 427371 451869
rect 427927 451008 428065 451884
rect 428621 451022 428780 451884
rect 429336 451022 429474 451898
rect 430030 451037 430260 451898
rect 430816 451037 430954 451913
rect 431510 451051 431669 451913
rect 432225 451051 432363 451927
rect 432919 451066 433070 451927
rect 433626 451066 433764 451942
rect 434320 451080 434479 451942
rect 435035 451080 435173 451956
rect 435729 451080 436086 451956
rect 434320 451066 436086 451080
rect 432919 451051 436086 451066
rect 431510 451037 436086 451051
rect 430030 451022 436086 451037
rect 428621 451008 436086 451022
rect 427220 450993 436086 451008
rect 425811 450979 436086 450993
rect 425267 443960 436086 450979
rect 425267 443946 434604 443960
rect 425267 443931 433195 443946
rect 425267 443917 431794 443931
rect 425267 443902 430385 443917
rect 425267 443888 428905 443902
rect 425267 443873 427496 443888
rect 425267 443859 426095 443873
rect 425267 443623 425700 443859
rect 425936 443623 426095 443859
rect 425267 443539 426095 443623
rect 425267 443303 425700 443539
rect 425936 443303 426095 443539
rect 425267 443219 426095 443303
rect 425267 442983 425700 443219
rect 425936 442997 426095 443219
rect 426651 442997 426789 443873
rect 427345 443012 427496 443873
rect 428052 443012 428190 443888
rect 428746 443026 428905 443888
rect 429461 443026 429599 443902
rect 430155 443041 430385 443902
rect 430941 443041 431079 443917
rect 431635 443055 431794 443917
rect 432350 443055 432488 443931
rect 433044 443070 433195 443931
rect 433751 443070 433889 443946
rect 434445 443084 434604 443946
rect 435160 443084 435298 443960
rect 435854 443084 436086 443960
rect 434445 443070 436086 443084
rect 433044 443055 436086 443070
rect 431635 443041 436086 443055
rect 430155 443026 436086 443041
rect 428746 443012 436086 443026
rect 427345 442997 436086 443012
rect 425936 442983 436086 442997
rect 425267 435927 436086 442983
rect 425267 435913 434518 435927
rect 425267 435898 433109 435913
rect 425267 435884 431708 435898
rect 425267 435869 430299 435884
rect 425267 435855 428819 435869
rect 425267 435840 427410 435855
rect 425267 435826 426009 435840
rect 425267 435590 425614 435826
rect 425850 435590 426009 435826
rect 425267 435506 426009 435590
rect 425267 435270 425614 435506
rect 425850 435270 426009 435506
rect 425267 435186 426009 435270
rect 425267 434950 425614 435186
rect 425850 434964 426009 435186
rect 426565 434964 426703 435840
rect 427259 434979 427410 435840
rect 427966 434979 428104 435855
rect 428660 434993 428819 435855
rect 429375 434993 429513 435869
rect 430069 435008 430299 435869
rect 430855 435008 430993 435884
rect 431549 435022 431708 435884
rect 432264 435022 432402 435898
rect 432958 435037 433109 435898
rect 433665 435037 433803 435913
rect 434359 435051 434518 435913
rect 435074 435051 435212 435927
rect 435768 435051 436086 435927
rect 434359 435037 436086 435051
rect 432958 435022 436086 435037
rect 431549 435008 436086 435022
rect 430069 434993 436086 435008
rect 428660 434979 436086 434993
rect 427259 434964 436086 434979
rect 425850 434950 436086 434964
rect 425267 427890 436086 434950
rect 425267 427876 434521 427890
rect 425267 427861 433112 427876
rect 425267 427847 431711 427861
rect 425267 427832 430302 427847
rect 425267 427818 428822 427832
rect 425267 427803 427413 427818
rect 425267 427789 426012 427803
rect 425267 427553 425617 427789
rect 425853 427553 426012 427789
rect 425267 427469 426012 427553
rect 425267 427233 425617 427469
rect 425853 427233 426012 427469
rect 425267 427149 426012 427233
rect 425267 426913 425617 427149
rect 425853 426927 426012 427149
rect 426568 426927 426706 427803
rect 427262 426942 427413 427803
rect 427969 426942 428107 427818
rect 428663 426956 428822 427818
rect 429378 426956 429516 427832
rect 430072 426971 430302 427832
rect 430858 426971 430996 427847
rect 431552 426985 431711 427847
rect 432267 426985 432405 427861
rect 432961 427000 433112 427861
rect 433668 427000 433806 427876
rect 434362 427014 434521 427876
rect 435077 427014 435215 427890
rect 435771 427014 436086 427890
rect 434362 427000 436086 427014
rect 432961 426985 436086 427000
rect 431552 426971 436086 426985
rect 430072 426956 436086 426971
rect 428663 426942 436086 426956
rect 427262 426927 436086 426942
rect 425853 426913 436086 426927
rect 425267 419955 436086 426913
rect 425267 419941 434535 419955
rect 425267 419926 433126 419941
rect 425267 419912 431725 419926
rect 425267 419897 430316 419912
rect 425267 419883 428836 419897
rect 425267 419868 427427 419883
rect 425267 419854 426026 419868
rect 425267 419618 425631 419854
rect 425867 419618 426026 419854
rect 425267 419534 426026 419618
rect 425267 419298 425631 419534
rect 425867 419298 426026 419534
rect 425267 419214 426026 419298
rect 425267 418978 425631 419214
rect 425867 418992 426026 419214
rect 426582 418992 426720 419868
rect 427276 419007 427427 419868
rect 427983 419007 428121 419883
rect 428677 419021 428836 419883
rect 429392 419021 429530 419897
rect 430086 419036 430316 419897
rect 430872 419036 431010 419912
rect 431566 419050 431725 419912
rect 432281 419050 432419 419926
rect 432975 419065 433126 419926
rect 433682 419065 433820 419941
rect 434376 419079 434535 419941
rect 435091 419079 435229 419955
rect 435785 419079 436086 419955
rect 434376 419065 436086 419079
rect 432975 419050 436086 419065
rect 431566 419036 436086 419050
rect 430086 419021 436086 419036
rect 428677 419007 436086 419021
rect 427276 418992 436086 419007
rect 425867 418978 436086 418992
rect 425267 411966 436086 418978
rect 425267 411952 434435 411966
rect 425267 411937 433026 411952
rect 425267 411923 431625 411937
rect 425267 411908 430216 411923
rect 425267 411894 428736 411908
rect 425267 411879 427327 411894
rect 425267 411865 425926 411879
rect 425267 411629 425531 411865
rect 425767 411629 425926 411865
rect 425267 411545 425926 411629
rect 425267 411309 425531 411545
rect 425767 411309 425926 411545
rect 425267 411225 425926 411309
rect 425267 410989 425531 411225
rect 425767 411003 425926 411225
rect 426482 411003 426620 411879
rect 427176 411018 427327 411879
rect 427883 411018 428021 411894
rect 428577 411032 428736 411894
rect 429292 411032 429430 411908
rect 429986 411047 430216 411908
rect 430772 411047 430910 411923
rect 431466 411061 431625 411923
rect 432181 411061 432319 411937
rect 432875 411076 433026 411937
rect 433582 411076 433720 411952
rect 434276 411090 434435 411952
rect 434991 411090 435129 411966
rect 435685 411090 436086 411966
rect 434276 411076 436086 411090
rect 432875 411061 436086 411076
rect 431466 411047 436086 411061
rect 429986 411032 436086 411047
rect 428577 411018 436086 411032
rect 427176 411003 436086 411018
rect 425767 410989 436086 411003
rect 425267 403941 436086 410989
rect 425267 403927 434580 403941
rect 425267 403912 433171 403927
rect 425267 403898 431770 403912
rect 425267 403883 430361 403898
rect 425267 403869 428881 403883
rect 425267 403854 427472 403869
rect 425267 403840 426071 403854
rect 425267 403604 425676 403840
rect 425912 403604 426071 403840
rect 425267 403520 426071 403604
rect 425267 403284 425676 403520
rect 425912 403284 426071 403520
rect 425267 403200 426071 403284
rect 425267 402964 425676 403200
rect 425912 402978 426071 403200
rect 426627 402978 426765 403854
rect 427321 402993 427472 403854
rect 428028 402993 428166 403869
rect 428722 403007 428881 403869
rect 429437 403007 429575 403883
rect 430131 403022 430361 403883
rect 430917 403022 431055 403898
rect 431611 403036 431770 403898
rect 432326 403036 432464 403912
rect 433020 403051 433171 403912
rect 433727 403051 433865 403927
rect 434421 403065 434580 403927
rect 435136 403065 435274 403941
rect 435830 403065 436086 403941
rect 434421 403051 436086 403065
rect 433020 403036 436086 403051
rect 431611 403022 436086 403036
rect 430131 403007 436086 403022
rect 428722 402993 436086 403007
rect 427321 402978 436086 402993
rect 425912 402964 436086 402978
rect 425267 395913 436086 402964
rect 425267 395899 434560 395913
rect 425267 395884 433151 395899
rect 425267 395870 431750 395884
rect 425267 395855 430341 395870
rect 425267 395841 428861 395855
rect 425267 395826 427452 395841
rect 425267 395812 426051 395826
rect 425267 395576 425656 395812
rect 425892 395576 426051 395812
rect 425267 395492 426051 395576
rect 425267 395256 425656 395492
rect 425892 395256 426051 395492
rect 425267 395172 426051 395256
rect 425267 394936 425656 395172
rect 425892 394950 426051 395172
rect 426607 394950 426745 395826
rect 427301 394965 427452 395826
rect 428008 394965 428146 395841
rect 428702 394979 428861 395841
rect 429417 394979 429555 395855
rect 430111 394994 430341 395855
rect 430897 394994 431035 395870
rect 431591 395008 431750 395870
rect 432306 395008 432444 395884
rect 433000 395023 433151 395884
rect 433707 395023 433845 395899
rect 434401 395037 434560 395899
rect 435116 395037 435254 395913
rect 435810 395037 436086 395913
rect 434401 395023 436086 395037
rect 433000 395008 436086 395023
rect 431591 394994 436086 395008
rect 430111 394979 436086 394994
rect 428702 394965 436086 394979
rect 427301 394950 436086 394965
rect 425892 394936 436086 394950
rect 425267 387922 436086 394936
rect 425267 387908 434579 387922
rect 425267 387893 433170 387908
rect 425267 387879 431769 387893
rect 425267 387864 430360 387879
rect 425267 387850 428880 387864
rect 425267 387835 427471 387850
rect 425267 387821 426070 387835
rect 425267 387585 425675 387821
rect 425911 387585 426070 387821
rect 425267 387501 426070 387585
rect 425267 387265 425675 387501
rect 425911 387265 426070 387501
rect 425267 387181 426070 387265
rect 425267 386945 425675 387181
rect 425911 386959 426070 387181
rect 426626 386959 426764 387835
rect 427320 386974 427471 387835
rect 428027 386974 428165 387850
rect 428721 386988 428880 387850
rect 429436 386988 429574 387864
rect 430130 387003 430360 387864
rect 430916 387003 431054 387879
rect 431610 387017 431769 387879
rect 432325 387017 432463 387893
rect 433019 387032 433170 387893
rect 433726 387032 433864 387908
rect 434420 387046 434579 387908
rect 435135 387046 435273 387922
rect 435829 387046 436086 387922
rect 434420 387032 436086 387046
rect 433019 387017 436086 387032
rect 431610 387003 436086 387017
rect 430130 386988 436086 387003
rect 428721 386974 436086 386988
rect 427320 386959 436086 386974
rect 425911 386945 436086 386959
rect 425267 379945 436086 386945
rect 425267 379931 434543 379945
rect 425267 379916 433134 379931
rect 425267 379902 431733 379916
rect 425267 379887 430324 379902
rect 425267 379873 428844 379887
rect 425267 379858 427435 379873
rect 425267 379844 426034 379858
rect 425267 379608 425639 379844
rect 425875 379608 426034 379844
rect 425267 379524 426034 379608
rect 425267 379288 425639 379524
rect 425875 379288 426034 379524
rect 425267 379204 426034 379288
rect 425267 378968 425639 379204
rect 425875 378982 426034 379204
rect 426590 378982 426728 379858
rect 427284 378997 427435 379858
rect 427991 378997 428129 379873
rect 428685 379011 428844 379873
rect 429400 379011 429538 379887
rect 430094 379026 430324 379887
rect 430880 379026 431018 379902
rect 431574 379040 431733 379902
rect 432289 379040 432427 379916
rect 432983 379055 433134 379916
rect 433690 379055 433828 379931
rect 434384 379069 434543 379931
rect 435099 379069 435237 379945
rect 435793 379069 436086 379945
rect 434384 379055 436086 379069
rect 432983 379040 436086 379055
rect 431574 379026 436086 379040
rect 430094 379011 436086 379026
rect 428685 378997 436086 379011
rect 427284 378982 436086 378997
rect 425875 378968 436086 378982
rect 425267 371957 436086 378968
rect 425267 371943 434531 371957
rect 425267 371928 433122 371943
rect 425267 371914 431721 371928
rect 425267 371899 430312 371914
rect 425267 371885 428832 371899
rect 425267 371870 427423 371885
rect 425267 371856 426022 371870
rect 425267 371620 425627 371856
rect 425863 371620 426022 371856
rect 425267 371536 426022 371620
rect 425267 371300 425627 371536
rect 425863 371300 426022 371536
rect 425267 371216 426022 371300
rect 425267 370980 425627 371216
rect 425863 370994 426022 371216
rect 426578 370994 426716 371870
rect 427272 371009 427423 371870
rect 427979 371009 428117 371885
rect 428673 371023 428832 371885
rect 429388 371023 429526 371899
rect 430082 371038 430312 371899
rect 430868 371038 431006 371914
rect 431562 371052 431721 371914
rect 432277 371052 432415 371928
rect 432971 371067 433122 371928
rect 433678 371067 433816 371943
rect 434372 371081 434531 371943
rect 435087 371081 435225 371957
rect 435781 371081 436086 371957
rect 434372 371067 436086 371081
rect 432971 371052 436086 371067
rect 431562 371038 436086 371052
rect 430082 371023 436086 371038
rect 428673 371009 436086 371023
rect 427272 370994 436086 371009
rect 425863 370980 436086 370994
rect 425267 363967 436086 370980
rect 425267 363953 434519 363967
rect 425267 363938 433110 363953
rect 425267 363924 431709 363938
rect 425267 363909 430300 363924
rect 425267 363895 428820 363909
rect 425267 363880 427411 363895
rect 425267 363866 426010 363880
rect 425267 363630 425615 363866
rect 425851 363630 426010 363866
rect 425267 363546 426010 363630
rect 425267 363310 425615 363546
rect 425851 363310 426010 363546
rect 425267 363226 426010 363310
rect 425267 362990 425615 363226
rect 425851 363004 426010 363226
rect 426566 363004 426704 363880
rect 427260 363019 427411 363880
rect 427967 363019 428105 363895
rect 428661 363033 428820 363895
rect 429376 363033 429514 363909
rect 430070 363048 430300 363909
rect 430856 363048 430994 363924
rect 431550 363062 431709 363924
rect 432265 363062 432403 363938
rect 432959 363077 433110 363938
rect 433666 363077 433804 363953
rect 434360 363091 434519 363953
rect 435075 363091 435213 363967
rect 435769 363091 436086 363967
rect 434360 363077 436086 363091
rect 432959 363062 436086 363077
rect 431550 363048 436086 363062
rect 430070 363033 436086 363048
rect 428661 363019 436086 363033
rect 427260 363004 436086 363019
rect 425851 362990 436086 363004
rect 425267 355958 436086 362990
rect 425267 355944 434568 355958
rect 425267 355929 433159 355944
rect 425267 355915 431758 355929
rect 425267 355900 430349 355915
rect 425267 355886 428869 355900
rect 425267 355871 427460 355886
rect 425267 355857 426059 355871
rect 425267 355621 425664 355857
rect 425900 355621 426059 355857
rect 425267 355537 426059 355621
rect 425267 355301 425664 355537
rect 425900 355301 426059 355537
rect 425267 355217 426059 355301
rect 425267 354981 425664 355217
rect 425900 354995 426059 355217
rect 426615 354995 426753 355871
rect 427309 355010 427460 355871
rect 428016 355010 428154 355886
rect 428710 355024 428869 355886
rect 429425 355024 429563 355900
rect 430119 355039 430349 355900
rect 430905 355039 431043 355915
rect 431599 355053 431758 355915
rect 432314 355053 432452 355929
rect 433008 355068 433159 355929
rect 433715 355068 433853 355944
rect 434409 355082 434568 355944
rect 435124 355082 435262 355958
rect 435818 355082 436086 355958
rect 434409 355068 436086 355082
rect 433008 355053 436086 355068
rect 431599 355039 436086 355053
rect 430119 355024 436086 355039
rect 428710 355010 436086 355024
rect 427309 354995 436086 355010
rect 425900 354981 436086 354995
rect 425267 347996 436086 354981
rect 425267 347982 434595 347996
rect 425267 347967 433186 347982
rect 425267 347953 431785 347967
rect 425267 347938 430376 347953
rect 425267 347924 428896 347938
rect 425267 347909 427487 347924
rect 425267 347895 426086 347909
rect 425267 347659 425691 347895
rect 425927 347659 426086 347895
rect 425267 347575 426086 347659
rect 425267 347339 425691 347575
rect 425927 347339 426086 347575
rect 425267 347255 426086 347339
rect 425267 347019 425691 347255
rect 425927 347033 426086 347255
rect 426642 347033 426780 347909
rect 427336 347048 427487 347909
rect 428043 347048 428181 347924
rect 428737 347062 428896 347924
rect 429452 347062 429590 347938
rect 430146 347077 430376 347938
rect 430932 347077 431070 347953
rect 431626 347091 431785 347953
rect 432341 347091 432479 347967
rect 433035 347106 433186 347967
rect 433742 347106 433880 347982
rect 434436 347120 434595 347982
rect 435151 347120 435289 347996
rect 435845 347120 436086 347996
rect 434436 347106 436086 347120
rect 433035 347091 436086 347106
rect 431626 347077 436086 347091
rect 430146 347062 436086 347077
rect 428737 347048 436086 347062
rect 427336 347033 436086 347048
rect 425927 347019 436086 347033
rect 425267 309371 436086 347019
rect 425267 309357 434539 309371
rect 425267 309342 433130 309357
rect 425267 309328 431729 309342
rect 425267 309313 430320 309328
rect 425267 309299 428840 309313
rect 425267 309284 427431 309299
rect 425267 309270 426030 309284
rect 425267 309034 425635 309270
rect 425871 309048 426030 309270
rect 426266 309048 426350 309284
rect 426586 309048 426724 309284
rect 426960 309048 427044 309284
rect 427280 309063 427431 309284
rect 427667 309063 427751 309299
rect 427987 309063 428125 309299
rect 428361 309063 428445 309299
rect 428681 309077 428840 309299
rect 429076 309077 429160 309313
rect 429396 309077 429534 309313
rect 429770 309077 429854 309313
rect 430090 309092 430320 309313
rect 430556 309092 430640 309328
rect 430876 309092 431014 309328
rect 431250 309092 431334 309328
rect 431570 309106 431729 309328
rect 431965 309106 432049 309342
rect 432285 309106 432423 309342
rect 432659 309106 432743 309342
rect 432979 309121 433130 309342
rect 433366 309121 433450 309357
rect 433686 309121 433824 309357
rect 434060 309121 434144 309357
rect 434380 309135 434539 309357
rect 434775 309135 434859 309371
rect 435095 309135 435233 309371
rect 435469 309135 435553 309371
rect 435789 309135 436086 309371
rect 434380 309121 436086 309135
rect 432979 309106 436086 309121
rect 431570 309092 436086 309106
rect 430090 309077 436086 309092
rect 428681 309063 436086 309077
rect 427280 309048 436086 309063
rect 425871 309034 436086 309048
rect 425267 273350 436086 309034
rect 425267 273336 434590 273350
rect 425267 273321 433181 273336
rect 425267 273307 431780 273321
rect 425267 273292 430371 273307
rect 425267 273278 428891 273292
rect 425267 273263 427482 273278
rect 425267 273249 426081 273263
rect 425267 273013 425686 273249
rect 425922 273027 426081 273249
rect 426317 273027 426401 273263
rect 426637 273027 426775 273263
rect 427011 273027 427095 273263
rect 427331 273042 427482 273263
rect 427718 273042 427802 273278
rect 428038 273042 428176 273278
rect 428412 273042 428496 273278
rect 428732 273056 428891 273278
rect 429127 273056 429211 273292
rect 429447 273056 429585 273292
rect 429821 273056 429905 273292
rect 430141 273071 430371 273292
rect 430607 273071 430691 273307
rect 430927 273071 431065 273307
rect 431301 273071 431385 273307
rect 431621 273085 431780 273307
rect 432016 273085 432100 273321
rect 432336 273085 432474 273321
rect 432710 273085 432794 273321
rect 433030 273100 433181 273321
rect 433417 273100 433501 273336
rect 433737 273100 433875 273336
rect 434111 273100 434195 273336
rect 434431 273114 434590 273336
rect 434826 273114 434910 273350
rect 435146 273114 435284 273350
rect 435520 273114 435604 273350
rect 435840 273114 436086 273350
rect 434431 273100 436086 273114
rect 433030 273085 436086 273100
rect 431621 273071 436086 273085
rect 430141 273056 436086 273071
rect 428732 273042 436086 273056
rect 427331 273027 436086 273042
rect 425922 273013 436086 273027
rect 425267 237395 436086 273013
rect 425267 237381 434622 237395
rect 425267 237366 433213 237381
rect 425267 237352 431812 237366
rect 425267 237337 430403 237352
rect 425267 237323 428923 237337
rect 425267 237308 427514 237323
rect 425267 237294 426113 237308
rect 425267 237058 425718 237294
rect 425954 237072 426113 237294
rect 426349 237072 426433 237308
rect 426669 237072 426807 237308
rect 427043 237072 427127 237308
rect 427363 237087 427514 237308
rect 427750 237087 427834 237323
rect 428070 237087 428208 237323
rect 428444 237087 428528 237323
rect 428764 237101 428923 237323
rect 429159 237101 429243 237337
rect 429479 237101 429617 237337
rect 429853 237101 429937 237337
rect 430173 237116 430403 237337
rect 430639 237116 430723 237352
rect 430959 237116 431097 237352
rect 431333 237116 431417 237352
rect 431653 237130 431812 237352
rect 432048 237130 432132 237366
rect 432368 237130 432506 237366
rect 432742 237130 432826 237366
rect 433062 237145 433213 237366
rect 433449 237145 433533 237381
rect 433769 237145 433907 237381
rect 434143 237145 434227 237381
rect 434463 237159 434622 237381
rect 434858 237159 434942 237395
rect 435178 237159 435316 237395
rect 435552 237159 435636 237395
rect 435872 237159 436086 237395
rect 434463 237145 436086 237159
rect 433062 237130 436086 237145
rect 431653 237116 436086 237130
rect 430173 237101 436086 237116
rect 428764 237087 436086 237101
rect 427363 237072 436086 237087
rect 425954 237058 436086 237072
rect 425267 234520 436086 237058
rect 451804 561454 452404 596898
rect 451804 561218 451986 561454
rect 452222 561218 452404 561454
rect 451804 561134 452404 561218
rect 451804 560898 451986 561134
rect 452222 560898 452404 561134
rect 451804 525454 452404 560898
rect 451804 525218 451986 525454
rect 452222 525218 452404 525454
rect 451804 525134 452404 525218
rect 451804 524898 451986 525134
rect 452222 524898 452404 525134
rect 451804 489454 452404 524898
rect 451804 489218 451986 489454
rect 452222 489218 452404 489454
rect 451804 489134 452404 489218
rect 451804 488898 451986 489134
rect 452222 488898 452404 489134
rect 451804 453454 452404 488898
rect 451804 453218 451986 453454
rect 452222 453218 452404 453454
rect 451804 453134 452404 453218
rect 451804 452898 451986 453134
rect 452222 452898 452404 453134
rect 451804 417454 452404 452898
rect 451804 417218 451986 417454
rect 452222 417218 452404 417454
rect 451804 417134 452404 417218
rect 451804 416898 451986 417134
rect 452222 416898 452404 417134
rect 451804 381454 452404 416898
rect 451804 381218 451986 381454
rect 452222 381218 452404 381454
rect 451804 381134 452404 381218
rect 451804 380898 451986 381134
rect 452222 380898 452404 381134
rect 451804 345454 452404 380898
rect 451804 345218 451986 345454
rect 452222 345218 452404 345454
rect 451804 345134 452404 345218
rect 451804 344898 451986 345134
rect 452222 344898 452404 345134
rect 451804 309454 452404 344898
rect 451804 309218 451986 309454
rect 452222 309218 452404 309454
rect 451804 309134 452404 309218
rect 451804 308898 451986 309134
rect 452222 308898 452404 309134
rect 451804 273454 452404 308898
rect 451804 273218 451986 273454
rect 452222 273218 452404 273454
rect 451804 273134 452404 273218
rect 451804 272898 451986 273134
rect 452222 272898 452404 273134
rect 451804 237454 452404 272898
rect 451804 237218 451986 237454
rect 452222 237218 452404 237454
rect 451804 237134 452404 237218
rect 451804 236898 451986 237134
rect 452222 236898 452404 237134
rect 390604 212254 391204 218000
rect 390604 212018 390786 212254
rect 391022 212018 391204 212254
rect 390604 211934 391204 212018
rect 390604 211698 390786 211934
rect 391022 211698 391204 211934
rect 390604 176254 391204 211698
rect 390604 176018 390786 176254
rect 391022 176018 391204 176254
rect 390604 175934 391204 176018
rect 390604 175698 390786 175934
rect 391022 175698 391204 175934
rect 390604 140254 391204 175698
rect 390604 140018 390786 140254
rect 391022 140018 391204 140254
rect 390604 139934 391204 140018
rect 390604 139698 390786 139934
rect 391022 139698 391204 139934
rect 390604 104254 391204 139698
rect 390604 104018 390786 104254
rect 391022 104018 391204 104254
rect 390604 103934 391204 104018
rect 390604 103698 390786 103934
rect 391022 103698 391204 103934
rect 390604 68254 391204 103698
rect 390604 68018 390786 68254
rect 391022 68018 391204 68254
rect 390604 67934 391204 68018
rect 390604 67698 390786 67934
rect 391022 67698 391204 67934
rect 390604 32254 391204 67698
rect 390604 32018 390786 32254
rect 391022 32018 391204 32254
rect 390604 31934 391204 32018
rect 389771 31788 389837 31789
rect 389771 31724 389772 31788
rect 389836 31724 389837 31788
rect 389771 31723 389837 31724
rect 387004 28418 387186 28654
rect 387422 28418 387604 28654
rect 387004 28334 387604 28418
rect 387004 28098 387186 28334
rect 387422 28098 387604 28334
rect 387004 -5046 387604 28098
rect 387004 -5282 387186 -5046
rect 387422 -5282 387604 -5046
rect 387004 -5366 387604 -5282
rect 387004 -5602 387186 -5366
rect 387422 -5602 387604 -5366
rect 387004 -5624 387604 -5602
rect 390604 31698 390786 31934
rect 391022 31698 391204 31934
rect 372604 -6222 372786 -5986
rect 373022 -6222 373204 -5986
rect 372604 -6306 373204 -6222
rect 372604 -6542 372786 -6306
rect 373022 -6542 373204 -6306
rect 372604 -7504 373204 -6542
rect 390604 -6926 391204 31698
rect 397804 183454 398404 218000
rect 397804 183218 397986 183454
rect 398222 183218 398404 183454
rect 397804 183134 398404 183218
rect 397804 182898 397986 183134
rect 398222 182898 398404 183134
rect 397804 147454 398404 182898
rect 397804 147218 397986 147454
rect 398222 147218 398404 147454
rect 397804 147134 398404 147218
rect 397804 146898 397986 147134
rect 398222 146898 398404 147134
rect 397804 111454 398404 146898
rect 397804 111218 397986 111454
rect 398222 111218 398404 111454
rect 397804 111134 398404 111218
rect 397804 110898 397986 111134
rect 398222 110898 398404 111134
rect 397804 75454 398404 110898
rect 397804 75218 397986 75454
rect 398222 75218 398404 75454
rect 397804 75134 398404 75218
rect 397804 74898 397986 75134
rect 398222 74898 398404 75134
rect 397804 39454 398404 74898
rect 397804 39218 397986 39454
rect 398222 39218 398404 39454
rect 397804 39134 398404 39218
rect 397804 38898 397986 39134
rect 398222 38898 398404 39134
rect 397804 3454 398404 38898
rect 397804 3218 397986 3454
rect 398222 3218 398404 3454
rect 397804 3134 398404 3218
rect 397804 2898 397986 3134
rect 398222 2898 398404 3134
rect 397804 -346 398404 2898
rect 397804 -582 397986 -346
rect 398222 -582 398404 -346
rect 397804 -666 398404 -582
rect 397804 -902 397986 -666
rect 398222 -902 398404 -666
rect 397804 -1864 398404 -902
rect 401404 187054 402004 218000
rect 401404 186818 401586 187054
rect 401822 186818 402004 187054
rect 401404 186734 402004 186818
rect 401404 186498 401586 186734
rect 401822 186498 402004 186734
rect 401404 151054 402004 186498
rect 401404 150818 401586 151054
rect 401822 150818 402004 151054
rect 401404 150734 402004 150818
rect 401404 150498 401586 150734
rect 401822 150498 402004 150734
rect 401404 115054 402004 150498
rect 401404 114818 401586 115054
rect 401822 114818 402004 115054
rect 401404 114734 402004 114818
rect 401404 114498 401586 114734
rect 401822 114498 402004 114734
rect 401404 79054 402004 114498
rect 401404 78818 401586 79054
rect 401822 78818 402004 79054
rect 401404 78734 402004 78818
rect 401404 78498 401586 78734
rect 401822 78498 402004 78734
rect 401404 43054 402004 78498
rect 401404 42818 401586 43054
rect 401822 42818 402004 43054
rect 401404 42734 402004 42818
rect 401404 42498 401586 42734
rect 401822 42498 402004 42734
rect 401404 7054 402004 42498
rect 401404 6818 401586 7054
rect 401822 6818 402004 7054
rect 401404 6734 402004 6818
rect 401404 6498 401586 6734
rect 401822 6498 402004 6734
rect 401404 -2226 402004 6498
rect 401404 -2462 401586 -2226
rect 401822 -2462 402004 -2226
rect 401404 -2546 402004 -2462
rect 401404 -2782 401586 -2546
rect 401822 -2782 402004 -2546
rect 401404 -3744 402004 -2782
rect 405004 190654 405604 218000
rect 405004 190418 405186 190654
rect 405422 190418 405604 190654
rect 405004 190334 405604 190418
rect 405004 190098 405186 190334
rect 405422 190098 405604 190334
rect 405004 154654 405604 190098
rect 405004 154418 405186 154654
rect 405422 154418 405604 154654
rect 405004 154334 405604 154418
rect 405004 154098 405186 154334
rect 405422 154098 405604 154334
rect 405004 118654 405604 154098
rect 405004 118418 405186 118654
rect 405422 118418 405604 118654
rect 405004 118334 405604 118418
rect 405004 118098 405186 118334
rect 405422 118098 405604 118334
rect 405004 82654 405604 118098
rect 405004 82418 405186 82654
rect 405422 82418 405604 82654
rect 405004 82334 405604 82418
rect 405004 82098 405186 82334
rect 405422 82098 405604 82334
rect 405004 46654 405604 82098
rect 405004 46418 405186 46654
rect 405422 46418 405604 46654
rect 405004 46334 405604 46418
rect 405004 46098 405186 46334
rect 405422 46098 405604 46334
rect 405004 10654 405604 46098
rect 405004 10418 405186 10654
rect 405422 10418 405604 10654
rect 405004 10334 405604 10418
rect 405004 10098 405186 10334
rect 405422 10098 405604 10334
rect 405004 -4106 405604 10098
rect 405004 -4342 405186 -4106
rect 405422 -4342 405604 -4106
rect 405004 -4426 405604 -4342
rect 405004 -4662 405186 -4426
rect 405422 -4662 405604 -4426
rect 405004 -5624 405604 -4662
rect 408604 194254 409204 218000
rect 408604 194018 408786 194254
rect 409022 194018 409204 194254
rect 408604 193934 409204 194018
rect 408604 193698 408786 193934
rect 409022 193698 409204 193934
rect 408604 158254 409204 193698
rect 408604 158018 408786 158254
rect 409022 158018 409204 158254
rect 408604 157934 409204 158018
rect 408604 157698 408786 157934
rect 409022 157698 409204 157934
rect 408604 122254 409204 157698
rect 408604 122018 408786 122254
rect 409022 122018 409204 122254
rect 408604 121934 409204 122018
rect 408604 121698 408786 121934
rect 409022 121698 409204 121934
rect 408604 86254 409204 121698
rect 408604 86018 408786 86254
rect 409022 86018 409204 86254
rect 408604 85934 409204 86018
rect 408604 85698 408786 85934
rect 409022 85698 409204 85934
rect 408604 50254 409204 85698
rect 408604 50018 408786 50254
rect 409022 50018 409204 50254
rect 408604 49934 409204 50018
rect 408604 49698 408786 49934
rect 409022 49698 409204 49934
rect 408604 14254 409204 49698
rect 408604 14018 408786 14254
rect 409022 14018 409204 14254
rect 408604 13934 409204 14018
rect 408604 13698 408786 13934
rect 409022 13698 409204 13934
rect 390604 -7162 390786 -6926
rect 391022 -7162 391204 -6926
rect 390604 -7246 391204 -7162
rect 390604 -7482 390786 -7246
rect 391022 -7482 391204 -7246
rect 390604 -7504 391204 -7482
rect 408604 -5986 409204 13698
rect 415804 201454 416404 218000
rect 415804 201218 415986 201454
rect 416222 201218 416404 201454
rect 415804 201134 416404 201218
rect 415804 200898 415986 201134
rect 416222 200898 416404 201134
rect 415804 165454 416404 200898
rect 415804 165218 415986 165454
rect 416222 165218 416404 165454
rect 415804 165134 416404 165218
rect 415804 164898 415986 165134
rect 416222 164898 416404 165134
rect 415804 129454 416404 164898
rect 415804 129218 415986 129454
rect 416222 129218 416404 129454
rect 415804 129134 416404 129218
rect 415804 128898 415986 129134
rect 416222 128898 416404 129134
rect 415804 93454 416404 128898
rect 415804 93218 415986 93454
rect 416222 93218 416404 93454
rect 415804 93134 416404 93218
rect 415804 92898 415986 93134
rect 416222 92898 416404 93134
rect 415804 57454 416404 92898
rect 415804 57218 415986 57454
rect 416222 57218 416404 57454
rect 415804 57134 416404 57218
rect 415804 56898 415986 57134
rect 416222 56898 416404 57134
rect 415804 21454 416404 56898
rect 415804 21218 415986 21454
rect 416222 21218 416404 21454
rect 415804 21134 416404 21218
rect 415804 20898 415986 21134
rect 416222 20898 416404 21134
rect 415804 -1286 416404 20898
rect 415804 -1522 415986 -1286
rect 416222 -1522 416404 -1286
rect 415804 -1606 416404 -1522
rect 415804 -1842 415986 -1606
rect 416222 -1842 416404 -1606
rect 415804 -1864 416404 -1842
rect 419404 205054 420004 218000
rect 419404 204818 419586 205054
rect 419822 204818 420004 205054
rect 419404 204734 420004 204818
rect 419404 204498 419586 204734
rect 419822 204498 420004 204734
rect 419404 169054 420004 204498
rect 419404 168818 419586 169054
rect 419822 168818 420004 169054
rect 419404 168734 420004 168818
rect 419404 168498 419586 168734
rect 419822 168498 420004 168734
rect 419404 133054 420004 168498
rect 419404 132818 419586 133054
rect 419822 132818 420004 133054
rect 419404 132734 420004 132818
rect 419404 132498 419586 132734
rect 419822 132498 420004 132734
rect 419404 97054 420004 132498
rect 419404 96818 419586 97054
rect 419822 96818 420004 97054
rect 419404 96734 420004 96818
rect 419404 96498 419586 96734
rect 419822 96498 420004 96734
rect 419404 61054 420004 96498
rect 419404 60818 419586 61054
rect 419822 60818 420004 61054
rect 419404 60734 420004 60818
rect 419404 60498 419586 60734
rect 419822 60498 420004 60734
rect 419404 25054 420004 60498
rect 419404 24818 419586 25054
rect 419822 24818 420004 25054
rect 419404 24734 420004 24818
rect 419404 24498 419586 24734
rect 419822 24498 420004 24734
rect 419404 -3166 420004 24498
rect 419404 -3402 419586 -3166
rect 419822 -3402 420004 -3166
rect 419404 -3486 420004 -3402
rect 419404 -3722 419586 -3486
rect 419822 -3722 420004 -3486
rect 419404 -3744 420004 -3722
rect 423004 208654 423604 218000
rect 423004 208418 423186 208654
rect 423422 208418 423604 208654
rect 423004 208334 423604 208418
rect 423004 208098 423186 208334
rect 423422 208098 423604 208334
rect 423004 172654 423604 208098
rect 423004 172418 423186 172654
rect 423422 172418 423604 172654
rect 423004 172334 423604 172418
rect 423004 172098 423186 172334
rect 423422 172098 423604 172334
rect 423004 136654 423604 172098
rect 423004 136418 423186 136654
rect 423422 136418 423604 136654
rect 423004 136334 423604 136418
rect 423004 136098 423186 136334
rect 423422 136098 423604 136334
rect 423004 100654 423604 136098
rect 423004 100418 423186 100654
rect 423422 100418 423604 100654
rect 423004 100334 423604 100418
rect 423004 100098 423186 100334
rect 423422 100098 423604 100334
rect 423004 64654 423604 100098
rect 423004 64418 423186 64654
rect 423422 64418 423604 64654
rect 423004 64334 423604 64418
rect 423004 64098 423186 64334
rect 423422 64098 423604 64334
rect 423004 28654 423604 64098
rect 423004 28418 423186 28654
rect 423422 28418 423604 28654
rect 423004 28334 423604 28418
rect 423004 28098 423186 28334
rect 423422 28098 423604 28334
rect 423004 -5046 423604 28098
rect 423004 -5282 423186 -5046
rect 423422 -5282 423604 -5046
rect 423004 -5366 423604 -5282
rect 423004 -5602 423186 -5366
rect 423422 -5602 423604 -5366
rect 423004 -5624 423604 -5602
rect 426604 212254 427204 218000
rect 426604 212018 426786 212254
rect 427022 212018 427204 212254
rect 426604 211934 427204 212018
rect 426604 211698 426786 211934
rect 427022 211698 427204 211934
rect 426604 176254 427204 211698
rect 426604 176018 426786 176254
rect 427022 176018 427204 176254
rect 426604 175934 427204 176018
rect 426604 175698 426786 175934
rect 427022 175698 427204 175934
rect 426604 140254 427204 175698
rect 426604 140018 426786 140254
rect 427022 140018 427204 140254
rect 426604 139934 427204 140018
rect 426604 139698 426786 139934
rect 427022 139698 427204 139934
rect 426604 104254 427204 139698
rect 426604 104018 426786 104254
rect 427022 104018 427204 104254
rect 426604 103934 427204 104018
rect 426604 103698 426786 103934
rect 427022 103698 427204 103934
rect 426604 68254 427204 103698
rect 426604 68018 426786 68254
rect 427022 68018 427204 68254
rect 426604 67934 427204 68018
rect 426604 67698 426786 67934
rect 427022 67698 427204 67934
rect 426604 32254 427204 67698
rect 426604 32018 426786 32254
rect 427022 32018 427204 32254
rect 426604 31934 427204 32018
rect 426604 31698 426786 31934
rect 427022 31698 427204 31934
rect 408604 -6222 408786 -5986
rect 409022 -6222 409204 -5986
rect 408604 -6306 409204 -6222
rect 408604 -6542 408786 -6306
rect 409022 -6542 409204 -6306
rect 408604 -7504 409204 -6542
rect 426604 -6926 427204 31698
rect 433804 183454 434404 218000
rect 433804 183218 433986 183454
rect 434222 183218 434404 183454
rect 433804 183134 434404 183218
rect 433804 182898 433986 183134
rect 434222 182898 434404 183134
rect 433804 147454 434404 182898
rect 433804 147218 433986 147454
rect 434222 147218 434404 147454
rect 433804 147134 434404 147218
rect 433804 146898 433986 147134
rect 434222 146898 434404 147134
rect 433804 111454 434404 146898
rect 433804 111218 433986 111454
rect 434222 111218 434404 111454
rect 433804 111134 434404 111218
rect 433804 110898 433986 111134
rect 434222 110898 434404 111134
rect 433804 75454 434404 110898
rect 433804 75218 433986 75454
rect 434222 75218 434404 75454
rect 433804 75134 434404 75218
rect 433804 74898 433986 75134
rect 434222 74898 434404 75134
rect 433804 39454 434404 74898
rect 433804 39218 433986 39454
rect 434222 39218 434404 39454
rect 433804 39134 434404 39218
rect 433804 38898 433986 39134
rect 434222 38898 434404 39134
rect 433804 3454 434404 38898
rect 433804 3218 433986 3454
rect 434222 3218 434404 3454
rect 433804 3134 434404 3218
rect 433804 2898 433986 3134
rect 434222 2898 434404 3134
rect 433804 -346 434404 2898
rect 433804 -582 433986 -346
rect 434222 -582 434404 -346
rect 433804 -666 434404 -582
rect 433804 -902 433986 -666
rect 434222 -902 434404 -666
rect 433804 -1864 434404 -902
rect 437404 187054 438004 218000
rect 437404 186818 437586 187054
rect 437822 186818 438004 187054
rect 437404 186734 438004 186818
rect 437404 186498 437586 186734
rect 437822 186498 438004 186734
rect 437404 151054 438004 186498
rect 437404 150818 437586 151054
rect 437822 150818 438004 151054
rect 437404 150734 438004 150818
rect 437404 150498 437586 150734
rect 437822 150498 438004 150734
rect 437404 115054 438004 150498
rect 437404 114818 437586 115054
rect 437822 114818 438004 115054
rect 437404 114734 438004 114818
rect 437404 114498 437586 114734
rect 437822 114498 438004 114734
rect 437404 79054 438004 114498
rect 437404 78818 437586 79054
rect 437822 78818 438004 79054
rect 437404 78734 438004 78818
rect 437404 78498 437586 78734
rect 437822 78498 438004 78734
rect 437404 43054 438004 78498
rect 437404 42818 437586 43054
rect 437822 42818 438004 43054
rect 437404 42734 438004 42818
rect 437404 42498 437586 42734
rect 437822 42498 438004 42734
rect 437404 7054 438004 42498
rect 437404 6818 437586 7054
rect 437822 6818 438004 7054
rect 437404 6734 438004 6818
rect 437404 6498 437586 6734
rect 437822 6498 438004 6734
rect 437404 -2226 438004 6498
rect 437404 -2462 437586 -2226
rect 437822 -2462 438004 -2226
rect 437404 -2546 438004 -2462
rect 437404 -2782 437586 -2546
rect 437822 -2782 438004 -2546
rect 437404 -3744 438004 -2782
rect 441004 190654 441604 218000
rect 441004 190418 441186 190654
rect 441422 190418 441604 190654
rect 441004 190334 441604 190418
rect 441004 190098 441186 190334
rect 441422 190098 441604 190334
rect 441004 154654 441604 190098
rect 441004 154418 441186 154654
rect 441422 154418 441604 154654
rect 441004 154334 441604 154418
rect 441004 154098 441186 154334
rect 441422 154098 441604 154334
rect 441004 118654 441604 154098
rect 441004 118418 441186 118654
rect 441422 118418 441604 118654
rect 441004 118334 441604 118418
rect 441004 118098 441186 118334
rect 441422 118098 441604 118334
rect 441004 82654 441604 118098
rect 441004 82418 441186 82654
rect 441422 82418 441604 82654
rect 441004 82334 441604 82418
rect 441004 82098 441186 82334
rect 441422 82098 441604 82334
rect 441004 46654 441604 82098
rect 441004 46418 441186 46654
rect 441422 46418 441604 46654
rect 441004 46334 441604 46418
rect 441004 46098 441186 46334
rect 441422 46098 441604 46334
rect 441004 10654 441604 46098
rect 441004 10418 441186 10654
rect 441422 10418 441604 10654
rect 441004 10334 441604 10418
rect 441004 10098 441186 10334
rect 441422 10098 441604 10334
rect 441004 -4106 441604 10098
rect 441004 -4342 441186 -4106
rect 441422 -4342 441604 -4106
rect 441004 -4426 441604 -4342
rect 441004 -4662 441186 -4426
rect 441422 -4662 441604 -4426
rect 441004 -5624 441604 -4662
rect 444604 194254 445204 218000
rect 444604 194018 444786 194254
rect 445022 194018 445204 194254
rect 444604 193934 445204 194018
rect 444604 193698 444786 193934
rect 445022 193698 445204 193934
rect 444604 158254 445204 193698
rect 444604 158018 444786 158254
rect 445022 158018 445204 158254
rect 444604 157934 445204 158018
rect 444604 157698 444786 157934
rect 445022 157698 445204 157934
rect 444604 122254 445204 157698
rect 444604 122018 444786 122254
rect 445022 122018 445204 122254
rect 444604 121934 445204 122018
rect 444604 121698 444786 121934
rect 445022 121698 445204 121934
rect 444604 86254 445204 121698
rect 444604 86018 444786 86254
rect 445022 86018 445204 86254
rect 444604 85934 445204 86018
rect 444604 85698 444786 85934
rect 445022 85698 445204 85934
rect 444604 50254 445204 85698
rect 444604 50018 444786 50254
rect 445022 50018 445204 50254
rect 444604 49934 445204 50018
rect 444604 49698 444786 49934
rect 445022 49698 445204 49934
rect 444604 14254 445204 49698
rect 444604 14018 444786 14254
rect 445022 14018 445204 14254
rect 444604 13934 445204 14018
rect 444604 13698 444786 13934
rect 445022 13698 445204 13934
rect 426604 -7162 426786 -6926
rect 427022 -7162 427204 -6926
rect 426604 -7246 427204 -7162
rect 426604 -7482 426786 -7246
rect 427022 -7482 427204 -7246
rect 426604 -7504 427204 -7482
rect 444604 -5986 445204 13698
rect 451804 201454 452404 236898
rect 451804 201218 451986 201454
rect 452222 201218 452404 201454
rect 451804 201134 452404 201218
rect 451804 200898 451986 201134
rect 452222 200898 452404 201134
rect 451804 165454 452404 200898
rect 451804 165218 451986 165454
rect 452222 165218 452404 165454
rect 451804 165134 452404 165218
rect 451804 164898 451986 165134
rect 452222 164898 452404 165134
rect 451804 129454 452404 164898
rect 451804 129218 451986 129454
rect 452222 129218 452404 129454
rect 451804 129134 452404 129218
rect 451804 128898 451986 129134
rect 452222 128898 452404 129134
rect 451804 93454 452404 128898
rect 451804 93218 451986 93454
rect 452222 93218 452404 93454
rect 451804 93134 452404 93218
rect 451804 92898 451986 93134
rect 452222 92898 452404 93134
rect 451804 57454 452404 92898
rect 451804 57218 451986 57454
rect 452222 57218 452404 57454
rect 451804 57134 452404 57218
rect 451804 56898 451986 57134
rect 452222 56898 452404 57134
rect 451804 21454 452404 56898
rect 451804 21218 451986 21454
rect 452222 21218 452404 21454
rect 451804 21134 452404 21218
rect 451804 20898 451986 21134
rect 452222 20898 452404 21134
rect 451804 -1286 452404 20898
rect 451804 -1522 451986 -1286
rect 452222 -1522 452404 -1286
rect 451804 -1606 452404 -1522
rect 451804 -1842 451986 -1606
rect 452222 -1842 452404 -1606
rect 451804 -1864 452404 -1842
rect 455404 673054 456004 707102
rect 455404 672818 455586 673054
rect 455822 672818 456004 673054
rect 455404 672734 456004 672818
rect 455404 672498 455586 672734
rect 455822 672498 456004 672734
rect 455404 637054 456004 672498
rect 455404 636818 455586 637054
rect 455822 636818 456004 637054
rect 455404 636734 456004 636818
rect 455404 636498 455586 636734
rect 455822 636498 456004 636734
rect 455404 601054 456004 636498
rect 455404 600818 455586 601054
rect 455822 600818 456004 601054
rect 455404 600734 456004 600818
rect 455404 600498 455586 600734
rect 455822 600498 456004 600734
rect 455404 565054 456004 600498
rect 455404 564818 455586 565054
rect 455822 564818 456004 565054
rect 455404 564734 456004 564818
rect 455404 564498 455586 564734
rect 455822 564498 456004 564734
rect 455404 529054 456004 564498
rect 455404 528818 455586 529054
rect 455822 528818 456004 529054
rect 455404 528734 456004 528818
rect 455404 528498 455586 528734
rect 455822 528498 456004 528734
rect 455404 493054 456004 528498
rect 455404 492818 455586 493054
rect 455822 492818 456004 493054
rect 455404 492734 456004 492818
rect 455404 492498 455586 492734
rect 455822 492498 456004 492734
rect 455404 457054 456004 492498
rect 455404 456818 455586 457054
rect 455822 456818 456004 457054
rect 455404 456734 456004 456818
rect 455404 456498 455586 456734
rect 455822 456498 456004 456734
rect 455404 421054 456004 456498
rect 455404 420818 455586 421054
rect 455822 420818 456004 421054
rect 455404 420734 456004 420818
rect 455404 420498 455586 420734
rect 455822 420498 456004 420734
rect 455404 385054 456004 420498
rect 455404 384818 455586 385054
rect 455822 384818 456004 385054
rect 455404 384734 456004 384818
rect 455404 384498 455586 384734
rect 455822 384498 456004 384734
rect 455404 349054 456004 384498
rect 455404 348818 455586 349054
rect 455822 348818 456004 349054
rect 455404 348734 456004 348818
rect 455404 348498 455586 348734
rect 455822 348498 456004 348734
rect 455404 313054 456004 348498
rect 455404 312818 455586 313054
rect 455822 312818 456004 313054
rect 455404 312734 456004 312818
rect 455404 312498 455586 312734
rect 455822 312498 456004 312734
rect 455404 277054 456004 312498
rect 455404 276818 455586 277054
rect 455822 276818 456004 277054
rect 455404 276734 456004 276818
rect 455404 276498 455586 276734
rect 455822 276498 456004 276734
rect 455404 241054 456004 276498
rect 455404 240818 455586 241054
rect 455822 240818 456004 241054
rect 455404 240734 456004 240818
rect 455404 240498 455586 240734
rect 455822 240498 456004 240734
rect 455404 205054 456004 240498
rect 455404 204818 455586 205054
rect 455822 204818 456004 205054
rect 455404 204734 456004 204818
rect 455404 204498 455586 204734
rect 455822 204498 456004 204734
rect 455404 169054 456004 204498
rect 455404 168818 455586 169054
rect 455822 168818 456004 169054
rect 455404 168734 456004 168818
rect 455404 168498 455586 168734
rect 455822 168498 456004 168734
rect 455404 133054 456004 168498
rect 455404 132818 455586 133054
rect 455822 132818 456004 133054
rect 455404 132734 456004 132818
rect 455404 132498 455586 132734
rect 455822 132498 456004 132734
rect 455404 97054 456004 132498
rect 455404 96818 455586 97054
rect 455822 96818 456004 97054
rect 455404 96734 456004 96818
rect 455404 96498 455586 96734
rect 455822 96498 456004 96734
rect 455404 61054 456004 96498
rect 455404 60818 455586 61054
rect 455822 60818 456004 61054
rect 455404 60734 456004 60818
rect 455404 60498 455586 60734
rect 455822 60498 456004 60734
rect 455404 25054 456004 60498
rect 455404 24818 455586 25054
rect 455822 24818 456004 25054
rect 455404 24734 456004 24818
rect 455404 24498 455586 24734
rect 455822 24498 456004 24734
rect 455404 -3166 456004 24498
rect 455404 -3402 455586 -3166
rect 455822 -3402 456004 -3166
rect 455404 -3486 456004 -3402
rect 455404 -3722 455586 -3486
rect 455822 -3722 456004 -3486
rect 455404 -3744 456004 -3722
rect 459004 676654 459604 708982
rect 459004 676418 459186 676654
rect 459422 676418 459604 676654
rect 459004 676334 459604 676418
rect 459004 676098 459186 676334
rect 459422 676098 459604 676334
rect 459004 640654 459604 676098
rect 459004 640418 459186 640654
rect 459422 640418 459604 640654
rect 459004 640334 459604 640418
rect 459004 640098 459186 640334
rect 459422 640098 459604 640334
rect 459004 604654 459604 640098
rect 459004 604418 459186 604654
rect 459422 604418 459604 604654
rect 459004 604334 459604 604418
rect 459004 604098 459186 604334
rect 459422 604098 459604 604334
rect 459004 568654 459604 604098
rect 459004 568418 459186 568654
rect 459422 568418 459604 568654
rect 459004 568334 459604 568418
rect 459004 568098 459186 568334
rect 459422 568098 459604 568334
rect 459004 532654 459604 568098
rect 459004 532418 459186 532654
rect 459422 532418 459604 532654
rect 459004 532334 459604 532418
rect 459004 532098 459186 532334
rect 459422 532098 459604 532334
rect 459004 496654 459604 532098
rect 459004 496418 459186 496654
rect 459422 496418 459604 496654
rect 459004 496334 459604 496418
rect 459004 496098 459186 496334
rect 459422 496098 459604 496334
rect 459004 460654 459604 496098
rect 459004 460418 459186 460654
rect 459422 460418 459604 460654
rect 459004 460334 459604 460418
rect 459004 460098 459186 460334
rect 459422 460098 459604 460334
rect 459004 424654 459604 460098
rect 459004 424418 459186 424654
rect 459422 424418 459604 424654
rect 459004 424334 459604 424418
rect 459004 424098 459186 424334
rect 459422 424098 459604 424334
rect 459004 388654 459604 424098
rect 459004 388418 459186 388654
rect 459422 388418 459604 388654
rect 459004 388334 459604 388418
rect 459004 388098 459186 388334
rect 459422 388098 459604 388334
rect 459004 352654 459604 388098
rect 459004 352418 459186 352654
rect 459422 352418 459604 352654
rect 459004 352334 459604 352418
rect 459004 352098 459186 352334
rect 459422 352098 459604 352334
rect 459004 316654 459604 352098
rect 459004 316418 459186 316654
rect 459422 316418 459604 316654
rect 459004 316334 459604 316418
rect 459004 316098 459186 316334
rect 459422 316098 459604 316334
rect 459004 280654 459604 316098
rect 459004 280418 459186 280654
rect 459422 280418 459604 280654
rect 459004 280334 459604 280418
rect 459004 280098 459186 280334
rect 459422 280098 459604 280334
rect 459004 244654 459604 280098
rect 459004 244418 459186 244654
rect 459422 244418 459604 244654
rect 459004 244334 459604 244418
rect 459004 244098 459186 244334
rect 459422 244098 459604 244334
rect 459004 208654 459604 244098
rect 459004 208418 459186 208654
rect 459422 208418 459604 208654
rect 459004 208334 459604 208418
rect 459004 208098 459186 208334
rect 459422 208098 459604 208334
rect 459004 172654 459604 208098
rect 459004 172418 459186 172654
rect 459422 172418 459604 172654
rect 459004 172334 459604 172418
rect 459004 172098 459186 172334
rect 459422 172098 459604 172334
rect 459004 136654 459604 172098
rect 459004 136418 459186 136654
rect 459422 136418 459604 136654
rect 459004 136334 459604 136418
rect 459004 136098 459186 136334
rect 459422 136098 459604 136334
rect 459004 100654 459604 136098
rect 459004 100418 459186 100654
rect 459422 100418 459604 100654
rect 459004 100334 459604 100418
rect 459004 100098 459186 100334
rect 459422 100098 459604 100334
rect 459004 64654 459604 100098
rect 459004 64418 459186 64654
rect 459422 64418 459604 64654
rect 459004 64334 459604 64418
rect 459004 64098 459186 64334
rect 459422 64098 459604 64334
rect 459004 28654 459604 64098
rect 459004 28418 459186 28654
rect 459422 28418 459604 28654
rect 459004 28334 459604 28418
rect 459004 28098 459186 28334
rect 459422 28098 459604 28334
rect 459004 -5046 459604 28098
rect 459004 -5282 459186 -5046
rect 459422 -5282 459604 -5046
rect 459004 -5366 459604 -5282
rect 459004 -5602 459186 -5366
rect 459422 -5602 459604 -5366
rect 459004 -5624 459604 -5602
rect 462604 680254 463204 710862
rect 480604 710478 481204 711440
rect 480604 710242 480786 710478
rect 481022 710242 481204 710478
rect 480604 710158 481204 710242
rect 480604 709922 480786 710158
rect 481022 709922 481204 710158
rect 477004 708598 477604 709560
rect 477004 708362 477186 708598
rect 477422 708362 477604 708598
rect 477004 708278 477604 708362
rect 477004 708042 477186 708278
rect 477422 708042 477604 708278
rect 473404 706718 474004 707680
rect 473404 706482 473586 706718
rect 473822 706482 474004 706718
rect 473404 706398 474004 706482
rect 473404 706162 473586 706398
rect 473822 706162 474004 706398
rect 462604 680018 462786 680254
rect 463022 680018 463204 680254
rect 462604 679934 463204 680018
rect 462604 679698 462786 679934
rect 463022 679698 463204 679934
rect 462604 644254 463204 679698
rect 462604 644018 462786 644254
rect 463022 644018 463204 644254
rect 462604 643934 463204 644018
rect 462604 643698 462786 643934
rect 463022 643698 463204 643934
rect 462604 608254 463204 643698
rect 462604 608018 462786 608254
rect 463022 608018 463204 608254
rect 462604 607934 463204 608018
rect 462604 607698 462786 607934
rect 463022 607698 463204 607934
rect 462604 572254 463204 607698
rect 462604 572018 462786 572254
rect 463022 572018 463204 572254
rect 462604 571934 463204 572018
rect 462604 571698 462786 571934
rect 463022 571698 463204 571934
rect 462604 536254 463204 571698
rect 462604 536018 462786 536254
rect 463022 536018 463204 536254
rect 462604 535934 463204 536018
rect 462604 535698 462786 535934
rect 463022 535698 463204 535934
rect 462604 500254 463204 535698
rect 462604 500018 462786 500254
rect 463022 500018 463204 500254
rect 462604 499934 463204 500018
rect 462604 499698 462786 499934
rect 463022 499698 463204 499934
rect 462604 464254 463204 499698
rect 462604 464018 462786 464254
rect 463022 464018 463204 464254
rect 462604 463934 463204 464018
rect 462604 463698 462786 463934
rect 463022 463698 463204 463934
rect 462604 428254 463204 463698
rect 462604 428018 462786 428254
rect 463022 428018 463204 428254
rect 462604 427934 463204 428018
rect 462604 427698 462786 427934
rect 463022 427698 463204 427934
rect 462604 392254 463204 427698
rect 462604 392018 462786 392254
rect 463022 392018 463204 392254
rect 462604 391934 463204 392018
rect 462604 391698 462786 391934
rect 463022 391698 463204 391934
rect 462604 356254 463204 391698
rect 462604 356018 462786 356254
rect 463022 356018 463204 356254
rect 462604 355934 463204 356018
rect 462604 355698 462786 355934
rect 463022 355698 463204 355934
rect 462604 320254 463204 355698
rect 462604 320018 462786 320254
rect 463022 320018 463204 320254
rect 462604 319934 463204 320018
rect 462604 319698 462786 319934
rect 463022 319698 463204 319934
rect 462604 284254 463204 319698
rect 462604 284018 462786 284254
rect 463022 284018 463204 284254
rect 462604 283934 463204 284018
rect 462604 283698 462786 283934
rect 463022 283698 463204 283934
rect 462604 248254 463204 283698
rect 462604 248018 462786 248254
rect 463022 248018 463204 248254
rect 462604 247934 463204 248018
rect 462604 247698 462786 247934
rect 463022 247698 463204 247934
rect 462604 212254 463204 247698
rect 462604 212018 462786 212254
rect 463022 212018 463204 212254
rect 462604 211934 463204 212018
rect 462604 211698 462786 211934
rect 463022 211698 463204 211934
rect 462604 176254 463204 211698
rect 462604 176018 462786 176254
rect 463022 176018 463204 176254
rect 462604 175934 463204 176018
rect 462604 175698 462786 175934
rect 463022 175698 463204 175934
rect 462604 140254 463204 175698
rect 462604 140018 462786 140254
rect 463022 140018 463204 140254
rect 462604 139934 463204 140018
rect 462604 139698 462786 139934
rect 463022 139698 463204 139934
rect 462604 104254 463204 139698
rect 462604 104018 462786 104254
rect 463022 104018 463204 104254
rect 462604 103934 463204 104018
rect 462604 103698 462786 103934
rect 463022 103698 463204 103934
rect 462604 68254 463204 103698
rect 462604 68018 462786 68254
rect 463022 68018 463204 68254
rect 462604 67934 463204 68018
rect 462604 67698 462786 67934
rect 463022 67698 463204 67934
rect 462604 32254 463204 67698
rect 462604 32018 462786 32254
rect 463022 32018 463204 32254
rect 462604 31934 463204 32018
rect 462604 31698 462786 31934
rect 463022 31698 463204 31934
rect 444604 -6222 444786 -5986
rect 445022 -6222 445204 -5986
rect 444604 -6306 445204 -6222
rect 444604 -6542 444786 -6306
rect 445022 -6542 445204 -6306
rect 444604 -7504 445204 -6542
rect 462604 -6926 463204 31698
rect 469804 704838 470404 705800
rect 469804 704602 469986 704838
rect 470222 704602 470404 704838
rect 469804 704518 470404 704602
rect 469804 704282 469986 704518
rect 470222 704282 470404 704518
rect 469804 687454 470404 704282
rect 469804 687218 469986 687454
rect 470222 687218 470404 687454
rect 469804 687134 470404 687218
rect 469804 686898 469986 687134
rect 470222 686898 470404 687134
rect 469804 651454 470404 686898
rect 469804 651218 469986 651454
rect 470222 651218 470404 651454
rect 469804 651134 470404 651218
rect 469804 650898 469986 651134
rect 470222 650898 470404 651134
rect 469804 615454 470404 650898
rect 469804 615218 469986 615454
rect 470222 615218 470404 615454
rect 469804 615134 470404 615218
rect 469804 614898 469986 615134
rect 470222 614898 470404 615134
rect 469804 579454 470404 614898
rect 469804 579218 469986 579454
rect 470222 579218 470404 579454
rect 469804 579134 470404 579218
rect 469804 578898 469986 579134
rect 470222 578898 470404 579134
rect 469804 543454 470404 578898
rect 469804 543218 469986 543454
rect 470222 543218 470404 543454
rect 469804 543134 470404 543218
rect 469804 542898 469986 543134
rect 470222 542898 470404 543134
rect 469804 507454 470404 542898
rect 469804 507218 469986 507454
rect 470222 507218 470404 507454
rect 469804 507134 470404 507218
rect 469804 506898 469986 507134
rect 470222 506898 470404 507134
rect 469804 471454 470404 506898
rect 469804 471218 469986 471454
rect 470222 471218 470404 471454
rect 469804 471134 470404 471218
rect 469804 470898 469986 471134
rect 470222 470898 470404 471134
rect 469804 435454 470404 470898
rect 469804 435218 469986 435454
rect 470222 435218 470404 435454
rect 469804 435134 470404 435218
rect 469804 434898 469986 435134
rect 470222 434898 470404 435134
rect 469804 399454 470404 434898
rect 469804 399218 469986 399454
rect 470222 399218 470404 399454
rect 469804 399134 470404 399218
rect 469804 398898 469986 399134
rect 470222 398898 470404 399134
rect 469804 363454 470404 398898
rect 469804 363218 469986 363454
rect 470222 363218 470404 363454
rect 469804 363134 470404 363218
rect 469804 362898 469986 363134
rect 470222 362898 470404 363134
rect 469804 327454 470404 362898
rect 469804 327218 469986 327454
rect 470222 327218 470404 327454
rect 469804 327134 470404 327218
rect 469804 326898 469986 327134
rect 470222 326898 470404 327134
rect 469804 291454 470404 326898
rect 469804 291218 469986 291454
rect 470222 291218 470404 291454
rect 469804 291134 470404 291218
rect 469804 290898 469986 291134
rect 470222 290898 470404 291134
rect 469804 255454 470404 290898
rect 469804 255218 469986 255454
rect 470222 255218 470404 255454
rect 469804 255134 470404 255218
rect 469804 254898 469986 255134
rect 470222 254898 470404 255134
rect 469804 219454 470404 254898
rect 469804 219218 469986 219454
rect 470222 219218 470404 219454
rect 469804 219134 470404 219218
rect 469804 218898 469986 219134
rect 470222 218898 470404 219134
rect 469804 183454 470404 218898
rect 469804 183218 469986 183454
rect 470222 183218 470404 183454
rect 469804 183134 470404 183218
rect 469804 182898 469986 183134
rect 470222 182898 470404 183134
rect 469804 147454 470404 182898
rect 469804 147218 469986 147454
rect 470222 147218 470404 147454
rect 469804 147134 470404 147218
rect 469804 146898 469986 147134
rect 470222 146898 470404 147134
rect 469804 111454 470404 146898
rect 469804 111218 469986 111454
rect 470222 111218 470404 111454
rect 469804 111134 470404 111218
rect 469804 110898 469986 111134
rect 470222 110898 470404 111134
rect 469804 75454 470404 110898
rect 469804 75218 469986 75454
rect 470222 75218 470404 75454
rect 469804 75134 470404 75218
rect 469804 74898 469986 75134
rect 470222 74898 470404 75134
rect 469804 39454 470404 74898
rect 469804 39218 469986 39454
rect 470222 39218 470404 39454
rect 469804 39134 470404 39218
rect 469804 38898 469986 39134
rect 470222 38898 470404 39134
rect 469804 3454 470404 38898
rect 469804 3218 469986 3454
rect 470222 3218 470404 3454
rect 469804 3134 470404 3218
rect 469804 2898 469986 3134
rect 470222 2898 470404 3134
rect 469804 -346 470404 2898
rect 469804 -582 469986 -346
rect 470222 -582 470404 -346
rect 469804 -666 470404 -582
rect 469804 -902 469986 -666
rect 470222 -902 470404 -666
rect 469804 -1864 470404 -902
rect 473404 691054 474004 706162
rect 473404 690818 473586 691054
rect 473822 690818 474004 691054
rect 473404 690734 474004 690818
rect 473404 690498 473586 690734
rect 473822 690498 474004 690734
rect 473404 655054 474004 690498
rect 473404 654818 473586 655054
rect 473822 654818 474004 655054
rect 473404 654734 474004 654818
rect 473404 654498 473586 654734
rect 473822 654498 474004 654734
rect 473404 619054 474004 654498
rect 473404 618818 473586 619054
rect 473822 618818 474004 619054
rect 473404 618734 474004 618818
rect 473404 618498 473586 618734
rect 473822 618498 474004 618734
rect 473404 583054 474004 618498
rect 473404 582818 473586 583054
rect 473822 582818 474004 583054
rect 473404 582734 474004 582818
rect 473404 582498 473586 582734
rect 473822 582498 474004 582734
rect 473404 547054 474004 582498
rect 473404 546818 473586 547054
rect 473822 546818 474004 547054
rect 473404 546734 474004 546818
rect 473404 546498 473586 546734
rect 473822 546498 474004 546734
rect 473404 511054 474004 546498
rect 473404 510818 473586 511054
rect 473822 510818 474004 511054
rect 473404 510734 474004 510818
rect 473404 510498 473586 510734
rect 473822 510498 474004 510734
rect 473404 475054 474004 510498
rect 473404 474818 473586 475054
rect 473822 474818 474004 475054
rect 473404 474734 474004 474818
rect 473404 474498 473586 474734
rect 473822 474498 474004 474734
rect 473404 439054 474004 474498
rect 473404 438818 473586 439054
rect 473822 438818 474004 439054
rect 473404 438734 474004 438818
rect 473404 438498 473586 438734
rect 473822 438498 474004 438734
rect 473404 403054 474004 438498
rect 473404 402818 473586 403054
rect 473822 402818 474004 403054
rect 473404 402734 474004 402818
rect 473404 402498 473586 402734
rect 473822 402498 474004 402734
rect 473404 367054 474004 402498
rect 473404 366818 473586 367054
rect 473822 366818 474004 367054
rect 473404 366734 474004 366818
rect 473404 366498 473586 366734
rect 473822 366498 474004 366734
rect 473404 331054 474004 366498
rect 473404 330818 473586 331054
rect 473822 330818 474004 331054
rect 473404 330734 474004 330818
rect 473404 330498 473586 330734
rect 473822 330498 474004 330734
rect 473404 295054 474004 330498
rect 473404 294818 473586 295054
rect 473822 294818 474004 295054
rect 473404 294734 474004 294818
rect 473404 294498 473586 294734
rect 473822 294498 474004 294734
rect 473404 259054 474004 294498
rect 473404 258818 473586 259054
rect 473822 258818 474004 259054
rect 473404 258734 474004 258818
rect 473404 258498 473586 258734
rect 473822 258498 474004 258734
rect 473404 223054 474004 258498
rect 473404 222818 473586 223054
rect 473822 222818 474004 223054
rect 473404 222734 474004 222818
rect 473404 222498 473586 222734
rect 473822 222498 474004 222734
rect 473404 187054 474004 222498
rect 473404 186818 473586 187054
rect 473822 186818 474004 187054
rect 473404 186734 474004 186818
rect 473404 186498 473586 186734
rect 473822 186498 474004 186734
rect 473404 151054 474004 186498
rect 473404 150818 473586 151054
rect 473822 150818 474004 151054
rect 473404 150734 474004 150818
rect 473404 150498 473586 150734
rect 473822 150498 474004 150734
rect 473404 115054 474004 150498
rect 473404 114818 473586 115054
rect 473822 114818 474004 115054
rect 473404 114734 474004 114818
rect 473404 114498 473586 114734
rect 473822 114498 474004 114734
rect 473404 79054 474004 114498
rect 473404 78818 473586 79054
rect 473822 78818 474004 79054
rect 473404 78734 474004 78818
rect 473404 78498 473586 78734
rect 473822 78498 474004 78734
rect 473404 43054 474004 78498
rect 473404 42818 473586 43054
rect 473822 42818 474004 43054
rect 473404 42734 474004 42818
rect 473404 42498 473586 42734
rect 473822 42498 474004 42734
rect 473404 7054 474004 42498
rect 473404 6818 473586 7054
rect 473822 6818 474004 7054
rect 473404 6734 474004 6818
rect 473404 6498 473586 6734
rect 473822 6498 474004 6734
rect 473404 -2226 474004 6498
rect 473404 -2462 473586 -2226
rect 473822 -2462 474004 -2226
rect 473404 -2546 474004 -2462
rect 473404 -2782 473586 -2546
rect 473822 -2782 474004 -2546
rect 473404 -3744 474004 -2782
rect 477004 694654 477604 708042
rect 477004 694418 477186 694654
rect 477422 694418 477604 694654
rect 477004 694334 477604 694418
rect 477004 694098 477186 694334
rect 477422 694098 477604 694334
rect 477004 658654 477604 694098
rect 477004 658418 477186 658654
rect 477422 658418 477604 658654
rect 477004 658334 477604 658418
rect 477004 658098 477186 658334
rect 477422 658098 477604 658334
rect 477004 622654 477604 658098
rect 477004 622418 477186 622654
rect 477422 622418 477604 622654
rect 477004 622334 477604 622418
rect 477004 622098 477186 622334
rect 477422 622098 477604 622334
rect 477004 586654 477604 622098
rect 477004 586418 477186 586654
rect 477422 586418 477604 586654
rect 477004 586334 477604 586418
rect 477004 586098 477186 586334
rect 477422 586098 477604 586334
rect 477004 550654 477604 586098
rect 477004 550418 477186 550654
rect 477422 550418 477604 550654
rect 477004 550334 477604 550418
rect 477004 550098 477186 550334
rect 477422 550098 477604 550334
rect 477004 514654 477604 550098
rect 477004 514418 477186 514654
rect 477422 514418 477604 514654
rect 477004 514334 477604 514418
rect 477004 514098 477186 514334
rect 477422 514098 477604 514334
rect 477004 478654 477604 514098
rect 477004 478418 477186 478654
rect 477422 478418 477604 478654
rect 477004 478334 477604 478418
rect 477004 478098 477186 478334
rect 477422 478098 477604 478334
rect 477004 442654 477604 478098
rect 477004 442418 477186 442654
rect 477422 442418 477604 442654
rect 477004 442334 477604 442418
rect 477004 442098 477186 442334
rect 477422 442098 477604 442334
rect 477004 406654 477604 442098
rect 477004 406418 477186 406654
rect 477422 406418 477604 406654
rect 477004 406334 477604 406418
rect 477004 406098 477186 406334
rect 477422 406098 477604 406334
rect 477004 370654 477604 406098
rect 477004 370418 477186 370654
rect 477422 370418 477604 370654
rect 477004 370334 477604 370418
rect 477004 370098 477186 370334
rect 477422 370098 477604 370334
rect 477004 334654 477604 370098
rect 477004 334418 477186 334654
rect 477422 334418 477604 334654
rect 477004 334334 477604 334418
rect 477004 334098 477186 334334
rect 477422 334098 477604 334334
rect 477004 298654 477604 334098
rect 477004 298418 477186 298654
rect 477422 298418 477604 298654
rect 477004 298334 477604 298418
rect 477004 298098 477186 298334
rect 477422 298098 477604 298334
rect 477004 262654 477604 298098
rect 477004 262418 477186 262654
rect 477422 262418 477604 262654
rect 477004 262334 477604 262418
rect 477004 262098 477186 262334
rect 477422 262098 477604 262334
rect 477004 226654 477604 262098
rect 477004 226418 477186 226654
rect 477422 226418 477604 226654
rect 477004 226334 477604 226418
rect 477004 226098 477186 226334
rect 477422 226098 477604 226334
rect 477004 190654 477604 226098
rect 477004 190418 477186 190654
rect 477422 190418 477604 190654
rect 477004 190334 477604 190418
rect 477004 190098 477186 190334
rect 477422 190098 477604 190334
rect 477004 154654 477604 190098
rect 477004 154418 477186 154654
rect 477422 154418 477604 154654
rect 477004 154334 477604 154418
rect 477004 154098 477186 154334
rect 477422 154098 477604 154334
rect 477004 118654 477604 154098
rect 477004 118418 477186 118654
rect 477422 118418 477604 118654
rect 477004 118334 477604 118418
rect 477004 118098 477186 118334
rect 477422 118098 477604 118334
rect 477004 82654 477604 118098
rect 477004 82418 477186 82654
rect 477422 82418 477604 82654
rect 477004 82334 477604 82418
rect 477004 82098 477186 82334
rect 477422 82098 477604 82334
rect 477004 46654 477604 82098
rect 477004 46418 477186 46654
rect 477422 46418 477604 46654
rect 477004 46334 477604 46418
rect 477004 46098 477186 46334
rect 477422 46098 477604 46334
rect 477004 10654 477604 46098
rect 477004 10418 477186 10654
rect 477422 10418 477604 10654
rect 477004 10334 477604 10418
rect 477004 10098 477186 10334
rect 477422 10098 477604 10334
rect 477004 -4106 477604 10098
rect 477004 -4342 477186 -4106
rect 477422 -4342 477604 -4106
rect 477004 -4426 477604 -4342
rect 477004 -4662 477186 -4426
rect 477422 -4662 477604 -4426
rect 477004 -5624 477604 -4662
rect 480604 698254 481204 709922
rect 498604 711418 499204 711440
rect 498604 711182 498786 711418
rect 499022 711182 499204 711418
rect 498604 711098 499204 711182
rect 498604 710862 498786 711098
rect 499022 710862 499204 711098
rect 495004 709538 495604 709560
rect 495004 709302 495186 709538
rect 495422 709302 495604 709538
rect 495004 709218 495604 709302
rect 495004 708982 495186 709218
rect 495422 708982 495604 709218
rect 491404 707658 492004 707680
rect 491404 707422 491586 707658
rect 491822 707422 492004 707658
rect 491404 707338 492004 707422
rect 491404 707102 491586 707338
rect 491822 707102 492004 707338
rect 480604 698018 480786 698254
rect 481022 698018 481204 698254
rect 480604 697934 481204 698018
rect 480604 697698 480786 697934
rect 481022 697698 481204 697934
rect 480604 662254 481204 697698
rect 480604 662018 480786 662254
rect 481022 662018 481204 662254
rect 480604 661934 481204 662018
rect 480604 661698 480786 661934
rect 481022 661698 481204 661934
rect 480604 626254 481204 661698
rect 480604 626018 480786 626254
rect 481022 626018 481204 626254
rect 480604 625934 481204 626018
rect 480604 625698 480786 625934
rect 481022 625698 481204 625934
rect 480604 590254 481204 625698
rect 480604 590018 480786 590254
rect 481022 590018 481204 590254
rect 480604 589934 481204 590018
rect 480604 589698 480786 589934
rect 481022 589698 481204 589934
rect 480604 554254 481204 589698
rect 480604 554018 480786 554254
rect 481022 554018 481204 554254
rect 480604 553934 481204 554018
rect 480604 553698 480786 553934
rect 481022 553698 481204 553934
rect 480604 518254 481204 553698
rect 480604 518018 480786 518254
rect 481022 518018 481204 518254
rect 480604 517934 481204 518018
rect 480604 517698 480786 517934
rect 481022 517698 481204 517934
rect 480604 482254 481204 517698
rect 480604 482018 480786 482254
rect 481022 482018 481204 482254
rect 480604 481934 481204 482018
rect 480604 481698 480786 481934
rect 481022 481698 481204 481934
rect 480604 446254 481204 481698
rect 480604 446018 480786 446254
rect 481022 446018 481204 446254
rect 480604 445934 481204 446018
rect 480604 445698 480786 445934
rect 481022 445698 481204 445934
rect 480604 410254 481204 445698
rect 480604 410018 480786 410254
rect 481022 410018 481204 410254
rect 480604 409934 481204 410018
rect 480604 409698 480786 409934
rect 481022 409698 481204 409934
rect 480604 374254 481204 409698
rect 480604 374018 480786 374254
rect 481022 374018 481204 374254
rect 480604 373934 481204 374018
rect 480604 373698 480786 373934
rect 481022 373698 481204 373934
rect 480604 338254 481204 373698
rect 480604 338018 480786 338254
rect 481022 338018 481204 338254
rect 480604 337934 481204 338018
rect 480604 337698 480786 337934
rect 481022 337698 481204 337934
rect 480604 302254 481204 337698
rect 480604 302018 480786 302254
rect 481022 302018 481204 302254
rect 480604 301934 481204 302018
rect 480604 301698 480786 301934
rect 481022 301698 481204 301934
rect 480604 266254 481204 301698
rect 480604 266018 480786 266254
rect 481022 266018 481204 266254
rect 480604 265934 481204 266018
rect 480604 265698 480786 265934
rect 481022 265698 481204 265934
rect 480604 230254 481204 265698
rect 480604 230018 480786 230254
rect 481022 230018 481204 230254
rect 480604 229934 481204 230018
rect 480604 229698 480786 229934
rect 481022 229698 481204 229934
rect 480604 194254 481204 229698
rect 480604 194018 480786 194254
rect 481022 194018 481204 194254
rect 480604 193934 481204 194018
rect 480604 193698 480786 193934
rect 481022 193698 481204 193934
rect 480604 158254 481204 193698
rect 480604 158018 480786 158254
rect 481022 158018 481204 158254
rect 480604 157934 481204 158018
rect 480604 157698 480786 157934
rect 481022 157698 481204 157934
rect 480604 122254 481204 157698
rect 480604 122018 480786 122254
rect 481022 122018 481204 122254
rect 480604 121934 481204 122018
rect 480604 121698 480786 121934
rect 481022 121698 481204 121934
rect 480604 86254 481204 121698
rect 480604 86018 480786 86254
rect 481022 86018 481204 86254
rect 480604 85934 481204 86018
rect 480604 85698 480786 85934
rect 481022 85698 481204 85934
rect 480604 50254 481204 85698
rect 480604 50018 480786 50254
rect 481022 50018 481204 50254
rect 480604 49934 481204 50018
rect 480604 49698 480786 49934
rect 481022 49698 481204 49934
rect 480604 14254 481204 49698
rect 480604 14018 480786 14254
rect 481022 14018 481204 14254
rect 480604 13934 481204 14018
rect 480604 13698 480786 13934
rect 481022 13698 481204 13934
rect 462604 -7162 462786 -6926
rect 463022 -7162 463204 -6926
rect 462604 -7246 463204 -7162
rect 462604 -7482 462786 -7246
rect 463022 -7482 463204 -7246
rect 462604 -7504 463204 -7482
rect 480604 -5986 481204 13698
rect 487804 705778 488404 705800
rect 487804 705542 487986 705778
rect 488222 705542 488404 705778
rect 487804 705458 488404 705542
rect 487804 705222 487986 705458
rect 488222 705222 488404 705458
rect 487804 669454 488404 705222
rect 487804 669218 487986 669454
rect 488222 669218 488404 669454
rect 487804 669134 488404 669218
rect 487804 668898 487986 669134
rect 488222 668898 488404 669134
rect 487804 633454 488404 668898
rect 487804 633218 487986 633454
rect 488222 633218 488404 633454
rect 487804 633134 488404 633218
rect 487804 632898 487986 633134
rect 488222 632898 488404 633134
rect 487804 597454 488404 632898
rect 487804 597218 487986 597454
rect 488222 597218 488404 597454
rect 487804 597134 488404 597218
rect 487804 596898 487986 597134
rect 488222 596898 488404 597134
rect 487804 561454 488404 596898
rect 487804 561218 487986 561454
rect 488222 561218 488404 561454
rect 487804 561134 488404 561218
rect 487804 560898 487986 561134
rect 488222 560898 488404 561134
rect 487804 525454 488404 560898
rect 487804 525218 487986 525454
rect 488222 525218 488404 525454
rect 487804 525134 488404 525218
rect 487804 524898 487986 525134
rect 488222 524898 488404 525134
rect 487804 489454 488404 524898
rect 487804 489218 487986 489454
rect 488222 489218 488404 489454
rect 487804 489134 488404 489218
rect 487804 488898 487986 489134
rect 488222 488898 488404 489134
rect 487804 453454 488404 488898
rect 487804 453218 487986 453454
rect 488222 453218 488404 453454
rect 487804 453134 488404 453218
rect 487804 452898 487986 453134
rect 488222 452898 488404 453134
rect 487804 417454 488404 452898
rect 487804 417218 487986 417454
rect 488222 417218 488404 417454
rect 487804 417134 488404 417218
rect 487804 416898 487986 417134
rect 488222 416898 488404 417134
rect 487804 381454 488404 416898
rect 487804 381218 487986 381454
rect 488222 381218 488404 381454
rect 487804 381134 488404 381218
rect 487804 380898 487986 381134
rect 488222 380898 488404 381134
rect 487804 345454 488404 380898
rect 487804 345218 487986 345454
rect 488222 345218 488404 345454
rect 487804 345134 488404 345218
rect 487804 344898 487986 345134
rect 488222 344898 488404 345134
rect 487804 309454 488404 344898
rect 487804 309218 487986 309454
rect 488222 309218 488404 309454
rect 487804 309134 488404 309218
rect 487804 308898 487986 309134
rect 488222 308898 488404 309134
rect 487804 273454 488404 308898
rect 487804 273218 487986 273454
rect 488222 273218 488404 273454
rect 487804 273134 488404 273218
rect 487804 272898 487986 273134
rect 488222 272898 488404 273134
rect 487804 237454 488404 272898
rect 487804 237218 487986 237454
rect 488222 237218 488404 237454
rect 487804 237134 488404 237218
rect 487804 236898 487986 237134
rect 488222 236898 488404 237134
rect 487804 201454 488404 236898
rect 487804 201218 487986 201454
rect 488222 201218 488404 201454
rect 487804 201134 488404 201218
rect 487804 200898 487986 201134
rect 488222 200898 488404 201134
rect 487804 165454 488404 200898
rect 487804 165218 487986 165454
rect 488222 165218 488404 165454
rect 487804 165134 488404 165218
rect 487804 164898 487986 165134
rect 488222 164898 488404 165134
rect 487804 129454 488404 164898
rect 487804 129218 487986 129454
rect 488222 129218 488404 129454
rect 487804 129134 488404 129218
rect 487804 128898 487986 129134
rect 488222 128898 488404 129134
rect 487804 93454 488404 128898
rect 487804 93218 487986 93454
rect 488222 93218 488404 93454
rect 487804 93134 488404 93218
rect 487804 92898 487986 93134
rect 488222 92898 488404 93134
rect 487804 57454 488404 92898
rect 487804 57218 487986 57454
rect 488222 57218 488404 57454
rect 487804 57134 488404 57218
rect 487804 56898 487986 57134
rect 488222 56898 488404 57134
rect 487804 21454 488404 56898
rect 487804 21218 487986 21454
rect 488222 21218 488404 21454
rect 487804 21134 488404 21218
rect 487804 20898 487986 21134
rect 488222 20898 488404 21134
rect 487804 -1286 488404 20898
rect 487804 -1522 487986 -1286
rect 488222 -1522 488404 -1286
rect 487804 -1606 488404 -1522
rect 487804 -1842 487986 -1606
rect 488222 -1842 488404 -1606
rect 487804 -1864 488404 -1842
rect 491404 673054 492004 707102
rect 491404 672818 491586 673054
rect 491822 672818 492004 673054
rect 491404 672734 492004 672818
rect 491404 672498 491586 672734
rect 491822 672498 492004 672734
rect 491404 637054 492004 672498
rect 491404 636818 491586 637054
rect 491822 636818 492004 637054
rect 491404 636734 492004 636818
rect 491404 636498 491586 636734
rect 491822 636498 492004 636734
rect 491404 601054 492004 636498
rect 491404 600818 491586 601054
rect 491822 600818 492004 601054
rect 491404 600734 492004 600818
rect 491404 600498 491586 600734
rect 491822 600498 492004 600734
rect 491404 565054 492004 600498
rect 491404 564818 491586 565054
rect 491822 564818 492004 565054
rect 491404 564734 492004 564818
rect 491404 564498 491586 564734
rect 491822 564498 492004 564734
rect 491404 529054 492004 564498
rect 491404 528818 491586 529054
rect 491822 528818 492004 529054
rect 491404 528734 492004 528818
rect 491404 528498 491586 528734
rect 491822 528498 492004 528734
rect 491404 493054 492004 528498
rect 491404 492818 491586 493054
rect 491822 492818 492004 493054
rect 491404 492734 492004 492818
rect 491404 492498 491586 492734
rect 491822 492498 492004 492734
rect 491404 457054 492004 492498
rect 491404 456818 491586 457054
rect 491822 456818 492004 457054
rect 491404 456734 492004 456818
rect 491404 456498 491586 456734
rect 491822 456498 492004 456734
rect 491404 421054 492004 456498
rect 491404 420818 491586 421054
rect 491822 420818 492004 421054
rect 491404 420734 492004 420818
rect 491404 420498 491586 420734
rect 491822 420498 492004 420734
rect 491404 385054 492004 420498
rect 491404 384818 491586 385054
rect 491822 384818 492004 385054
rect 491404 384734 492004 384818
rect 491404 384498 491586 384734
rect 491822 384498 492004 384734
rect 491404 349054 492004 384498
rect 491404 348818 491586 349054
rect 491822 348818 492004 349054
rect 491404 348734 492004 348818
rect 491404 348498 491586 348734
rect 491822 348498 492004 348734
rect 491404 313054 492004 348498
rect 491404 312818 491586 313054
rect 491822 312818 492004 313054
rect 491404 312734 492004 312818
rect 491404 312498 491586 312734
rect 491822 312498 492004 312734
rect 491404 277054 492004 312498
rect 491404 276818 491586 277054
rect 491822 276818 492004 277054
rect 491404 276734 492004 276818
rect 491404 276498 491586 276734
rect 491822 276498 492004 276734
rect 491404 241054 492004 276498
rect 491404 240818 491586 241054
rect 491822 240818 492004 241054
rect 491404 240734 492004 240818
rect 491404 240498 491586 240734
rect 491822 240498 492004 240734
rect 491404 205054 492004 240498
rect 491404 204818 491586 205054
rect 491822 204818 492004 205054
rect 491404 204734 492004 204818
rect 491404 204498 491586 204734
rect 491822 204498 492004 204734
rect 491404 169054 492004 204498
rect 491404 168818 491586 169054
rect 491822 168818 492004 169054
rect 491404 168734 492004 168818
rect 491404 168498 491586 168734
rect 491822 168498 492004 168734
rect 491404 133054 492004 168498
rect 491404 132818 491586 133054
rect 491822 132818 492004 133054
rect 491404 132734 492004 132818
rect 491404 132498 491586 132734
rect 491822 132498 492004 132734
rect 491404 97054 492004 132498
rect 491404 96818 491586 97054
rect 491822 96818 492004 97054
rect 491404 96734 492004 96818
rect 491404 96498 491586 96734
rect 491822 96498 492004 96734
rect 491404 61054 492004 96498
rect 491404 60818 491586 61054
rect 491822 60818 492004 61054
rect 491404 60734 492004 60818
rect 491404 60498 491586 60734
rect 491822 60498 492004 60734
rect 491404 25054 492004 60498
rect 491404 24818 491586 25054
rect 491822 24818 492004 25054
rect 491404 24734 492004 24818
rect 491404 24498 491586 24734
rect 491822 24498 492004 24734
rect 491404 -3166 492004 24498
rect 491404 -3402 491586 -3166
rect 491822 -3402 492004 -3166
rect 491404 -3486 492004 -3402
rect 491404 -3722 491586 -3486
rect 491822 -3722 492004 -3486
rect 491404 -3744 492004 -3722
rect 495004 676654 495604 708982
rect 495004 676418 495186 676654
rect 495422 676418 495604 676654
rect 495004 676334 495604 676418
rect 495004 676098 495186 676334
rect 495422 676098 495604 676334
rect 495004 640654 495604 676098
rect 495004 640418 495186 640654
rect 495422 640418 495604 640654
rect 495004 640334 495604 640418
rect 495004 640098 495186 640334
rect 495422 640098 495604 640334
rect 495004 604654 495604 640098
rect 495004 604418 495186 604654
rect 495422 604418 495604 604654
rect 495004 604334 495604 604418
rect 495004 604098 495186 604334
rect 495422 604098 495604 604334
rect 495004 568654 495604 604098
rect 495004 568418 495186 568654
rect 495422 568418 495604 568654
rect 495004 568334 495604 568418
rect 495004 568098 495186 568334
rect 495422 568098 495604 568334
rect 495004 532654 495604 568098
rect 495004 532418 495186 532654
rect 495422 532418 495604 532654
rect 495004 532334 495604 532418
rect 495004 532098 495186 532334
rect 495422 532098 495604 532334
rect 495004 496654 495604 532098
rect 495004 496418 495186 496654
rect 495422 496418 495604 496654
rect 495004 496334 495604 496418
rect 495004 496098 495186 496334
rect 495422 496098 495604 496334
rect 495004 460654 495604 496098
rect 495004 460418 495186 460654
rect 495422 460418 495604 460654
rect 495004 460334 495604 460418
rect 495004 460098 495186 460334
rect 495422 460098 495604 460334
rect 495004 424654 495604 460098
rect 495004 424418 495186 424654
rect 495422 424418 495604 424654
rect 495004 424334 495604 424418
rect 495004 424098 495186 424334
rect 495422 424098 495604 424334
rect 495004 388654 495604 424098
rect 495004 388418 495186 388654
rect 495422 388418 495604 388654
rect 495004 388334 495604 388418
rect 495004 388098 495186 388334
rect 495422 388098 495604 388334
rect 495004 352654 495604 388098
rect 495004 352418 495186 352654
rect 495422 352418 495604 352654
rect 495004 352334 495604 352418
rect 495004 352098 495186 352334
rect 495422 352098 495604 352334
rect 495004 316654 495604 352098
rect 495004 316418 495186 316654
rect 495422 316418 495604 316654
rect 495004 316334 495604 316418
rect 495004 316098 495186 316334
rect 495422 316098 495604 316334
rect 495004 280654 495604 316098
rect 495004 280418 495186 280654
rect 495422 280418 495604 280654
rect 495004 280334 495604 280418
rect 495004 280098 495186 280334
rect 495422 280098 495604 280334
rect 495004 244654 495604 280098
rect 495004 244418 495186 244654
rect 495422 244418 495604 244654
rect 495004 244334 495604 244418
rect 495004 244098 495186 244334
rect 495422 244098 495604 244334
rect 495004 208654 495604 244098
rect 495004 208418 495186 208654
rect 495422 208418 495604 208654
rect 495004 208334 495604 208418
rect 495004 208098 495186 208334
rect 495422 208098 495604 208334
rect 495004 172654 495604 208098
rect 495004 172418 495186 172654
rect 495422 172418 495604 172654
rect 495004 172334 495604 172418
rect 495004 172098 495186 172334
rect 495422 172098 495604 172334
rect 495004 136654 495604 172098
rect 495004 136418 495186 136654
rect 495422 136418 495604 136654
rect 495004 136334 495604 136418
rect 495004 136098 495186 136334
rect 495422 136098 495604 136334
rect 495004 100654 495604 136098
rect 495004 100418 495186 100654
rect 495422 100418 495604 100654
rect 495004 100334 495604 100418
rect 495004 100098 495186 100334
rect 495422 100098 495604 100334
rect 495004 64654 495604 100098
rect 495004 64418 495186 64654
rect 495422 64418 495604 64654
rect 495004 64334 495604 64418
rect 495004 64098 495186 64334
rect 495422 64098 495604 64334
rect 495004 28654 495604 64098
rect 495004 28418 495186 28654
rect 495422 28418 495604 28654
rect 495004 28334 495604 28418
rect 495004 28098 495186 28334
rect 495422 28098 495604 28334
rect 495004 -5046 495604 28098
rect 495004 -5282 495186 -5046
rect 495422 -5282 495604 -5046
rect 495004 -5366 495604 -5282
rect 495004 -5602 495186 -5366
rect 495422 -5602 495604 -5366
rect 495004 -5624 495604 -5602
rect 498604 680254 499204 710862
rect 516604 710478 517204 711440
rect 516604 710242 516786 710478
rect 517022 710242 517204 710478
rect 516604 710158 517204 710242
rect 516604 709922 516786 710158
rect 517022 709922 517204 710158
rect 513004 708598 513604 709560
rect 513004 708362 513186 708598
rect 513422 708362 513604 708598
rect 513004 708278 513604 708362
rect 513004 708042 513186 708278
rect 513422 708042 513604 708278
rect 509404 706718 510004 707680
rect 509404 706482 509586 706718
rect 509822 706482 510004 706718
rect 509404 706398 510004 706482
rect 509404 706162 509586 706398
rect 509822 706162 510004 706398
rect 498604 680018 498786 680254
rect 499022 680018 499204 680254
rect 498604 679934 499204 680018
rect 498604 679698 498786 679934
rect 499022 679698 499204 679934
rect 498604 644254 499204 679698
rect 498604 644018 498786 644254
rect 499022 644018 499204 644254
rect 498604 643934 499204 644018
rect 498604 643698 498786 643934
rect 499022 643698 499204 643934
rect 498604 608254 499204 643698
rect 498604 608018 498786 608254
rect 499022 608018 499204 608254
rect 498604 607934 499204 608018
rect 498604 607698 498786 607934
rect 499022 607698 499204 607934
rect 498604 572254 499204 607698
rect 498604 572018 498786 572254
rect 499022 572018 499204 572254
rect 498604 571934 499204 572018
rect 498604 571698 498786 571934
rect 499022 571698 499204 571934
rect 498604 536254 499204 571698
rect 498604 536018 498786 536254
rect 499022 536018 499204 536254
rect 498604 535934 499204 536018
rect 498604 535698 498786 535934
rect 499022 535698 499204 535934
rect 498604 500254 499204 535698
rect 498604 500018 498786 500254
rect 499022 500018 499204 500254
rect 498604 499934 499204 500018
rect 498604 499698 498786 499934
rect 499022 499698 499204 499934
rect 498604 464254 499204 499698
rect 498604 464018 498786 464254
rect 499022 464018 499204 464254
rect 498604 463934 499204 464018
rect 498604 463698 498786 463934
rect 499022 463698 499204 463934
rect 498604 428254 499204 463698
rect 498604 428018 498786 428254
rect 499022 428018 499204 428254
rect 498604 427934 499204 428018
rect 498604 427698 498786 427934
rect 499022 427698 499204 427934
rect 498604 392254 499204 427698
rect 498604 392018 498786 392254
rect 499022 392018 499204 392254
rect 498604 391934 499204 392018
rect 498604 391698 498786 391934
rect 499022 391698 499204 391934
rect 498604 356254 499204 391698
rect 498604 356018 498786 356254
rect 499022 356018 499204 356254
rect 498604 355934 499204 356018
rect 498604 355698 498786 355934
rect 499022 355698 499204 355934
rect 498604 320254 499204 355698
rect 498604 320018 498786 320254
rect 499022 320018 499204 320254
rect 498604 319934 499204 320018
rect 498604 319698 498786 319934
rect 499022 319698 499204 319934
rect 498604 284254 499204 319698
rect 498604 284018 498786 284254
rect 499022 284018 499204 284254
rect 498604 283934 499204 284018
rect 498604 283698 498786 283934
rect 499022 283698 499204 283934
rect 498604 248254 499204 283698
rect 498604 248018 498786 248254
rect 499022 248018 499204 248254
rect 498604 247934 499204 248018
rect 498604 247698 498786 247934
rect 499022 247698 499204 247934
rect 498604 212254 499204 247698
rect 498604 212018 498786 212254
rect 499022 212018 499204 212254
rect 498604 211934 499204 212018
rect 498604 211698 498786 211934
rect 499022 211698 499204 211934
rect 498604 176254 499204 211698
rect 498604 176018 498786 176254
rect 499022 176018 499204 176254
rect 498604 175934 499204 176018
rect 498604 175698 498786 175934
rect 499022 175698 499204 175934
rect 498604 140254 499204 175698
rect 498604 140018 498786 140254
rect 499022 140018 499204 140254
rect 498604 139934 499204 140018
rect 498604 139698 498786 139934
rect 499022 139698 499204 139934
rect 498604 104254 499204 139698
rect 498604 104018 498786 104254
rect 499022 104018 499204 104254
rect 498604 103934 499204 104018
rect 498604 103698 498786 103934
rect 499022 103698 499204 103934
rect 498604 68254 499204 103698
rect 498604 68018 498786 68254
rect 499022 68018 499204 68254
rect 498604 67934 499204 68018
rect 498604 67698 498786 67934
rect 499022 67698 499204 67934
rect 498604 32254 499204 67698
rect 498604 32018 498786 32254
rect 499022 32018 499204 32254
rect 498604 31934 499204 32018
rect 498604 31698 498786 31934
rect 499022 31698 499204 31934
rect 480604 -6222 480786 -5986
rect 481022 -6222 481204 -5986
rect 480604 -6306 481204 -6222
rect 480604 -6542 480786 -6306
rect 481022 -6542 481204 -6306
rect 480604 -7504 481204 -6542
rect 498604 -6926 499204 31698
rect 505804 704838 506404 705800
rect 505804 704602 505986 704838
rect 506222 704602 506404 704838
rect 505804 704518 506404 704602
rect 505804 704282 505986 704518
rect 506222 704282 506404 704518
rect 505804 687454 506404 704282
rect 505804 687218 505986 687454
rect 506222 687218 506404 687454
rect 505804 687134 506404 687218
rect 505804 686898 505986 687134
rect 506222 686898 506404 687134
rect 505804 651454 506404 686898
rect 505804 651218 505986 651454
rect 506222 651218 506404 651454
rect 505804 651134 506404 651218
rect 505804 650898 505986 651134
rect 506222 650898 506404 651134
rect 505804 615454 506404 650898
rect 505804 615218 505986 615454
rect 506222 615218 506404 615454
rect 505804 615134 506404 615218
rect 505804 614898 505986 615134
rect 506222 614898 506404 615134
rect 505804 579454 506404 614898
rect 505804 579218 505986 579454
rect 506222 579218 506404 579454
rect 505804 579134 506404 579218
rect 505804 578898 505986 579134
rect 506222 578898 506404 579134
rect 505804 543454 506404 578898
rect 505804 543218 505986 543454
rect 506222 543218 506404 543454
rect 505804 543134 506404 543218
rect 505804 542898 505986 543134
rect 506222 542898 506404 543134
rect 505804 507454 506404 542898
rect 505804 507218 505986 507454
rect 506222 507218 506404 507454
rect 505804 507134 506404 507218
rect 505804 506898 505986 507134
rect 506222 506898 506404 507134
rect 505804 471454 506404 506898
rect 505804 471218 505986 471454
rect 506222 471218 506404 471454
rect 505804 471134 506404 471218
rect 505804 470898 505986 471134
rect 506222 470898 506404 471134
rect 505804 435454 506404 470898
rect 505804 435218 505986 435454
rect 506222 435218 506404 435454
rect 505804 435134 506404 435218
rect 505804 434898 505986 435134
rect 506222 434898 506404 435134
rect 505804 399454 506404 434898
rect 505804 399218 505986 399454
rect 506222 399218 506404 399454
rect 505804 399134 506404 399218
rect 505804 398898 505986 399134
rect 506222 398898 506404 399134
rect 505804 363454 506404 398898
rect 505804 363218 505986 363454
rect 506222 363218 506404 363454
rect 505804 363134 506404 363218
rect 505804 362898 505986 363134
rect 506222 362898 506404 363134
rect 505804 327454 506404 362898
rect 505804 327218 505986 327454
rect 506222 327218 506404 327454
rect 505804 327134 506404 327218
rect 505804 326898 505986 327134
rect 506222 326898 506404 327134
rect 505804 291454 506404 326898
rect 505804 291218 505986 291454
rect 506222 291218 506404 291454
rect 505804 291134 506404 291218
rect 505804 290898 505986 291134
rect 506222 290898 506404 291134
rect 505804 255454 506404 290898
rect 505804 255218 505986 255454
rect 506222 255218 506404 255454
rect 505804 255134 506404 255218
rect 505804 254898 505986 255134
rect 506222 254898 506404 255134
rect 505804 219454 506404 254898
rect 505804 219218 505986 219454
rect 506222 219218 506404 219454
rect 505804 219134 506404 219218
rect 505804 218898 505986 219134
rect 506222 218898 506404 219134
rect 505804 183454 506404 218898
rect 505804 183218 505986 183454
rect 506222 183218 506404 183454
rect 505804 183134 506404 183218
rect 505804 182898 505986 183134
rect 506222 182898 506404 183134
rect 505804 147454 506404 182898
rect 505804 147218 505986 147454
rect 506222 147218 506404 147454
rect 505804 147134 506404 147218
rect 505804 146898 505986 147134
rect 506222 146898 506404 147134
rect 505804 111454 506404 146898
rect 505804 111218 505986 111454
rect 506222 111218 506404 111454
rect 505804 111134 506404 111218
rect 505804 110898 505986 111134
rect 506222 110898 506404 111134
rect 505804 75454 506404 110898
rect 505804 75218 505986 75454
rect 506222 75218 506404 75454
rect 505804 75134 506404 75218
rect 505804 74898 505986 75134
rect 506222 74898 506404 75134
rect 505804 39454 506404 74898
rect 505804 39218 505986 39454
rect 506222 39218 506404 39454
rect 505804 39134 506404 39218
rect 505804 38898 505986 39134
rect 506222 38898 506404 39134
rect 505804 3454 506404 38898
rect 505804 3218 505986 3454
rect 506222 3218 506404 3454
rect 505804 3134 506404 3218
rect 505804 2898 505986 3134
rect 506222 2898 506404 3134
rect 505804 -346 506404 2898
rect 505804 -582 505986 -346
rect 506222 -582 506404 -346
rect 505804 -666 506404 -582
rect 505804 -902 505986 -666
rect 506222 -902 506404 -666
rect 505804 -1864 506404 -902
rect 509404 691054 510004 706162
rect 509404 690818 509586 691054
rect 509822 690818 510004 691054
rect 509404 690734 510004 690818
rect 509404 690498 509586 690734
rect 509822 690498 510004 690734
rect 509404 655054 510004 690498
rect 509404 654818 509586 655054
rect 509822 654818 510004 655054
rect 509404 654734 510004 654818
rect 509404 654498 509586 654734
rect 509822 654498 510004 654734
rect 509404 619054 510004 654498
rect 509404 618818 509586 619054
rect 509822 618818 510004 619054
rect 509404 618734 510004 618818
rect 509404 618498 509586 618734
rect 509822 618498 510004 618734
rect 509404 583054 510004 618498
rect 509404 582818 509586 583054
rect 509822 582818 510004 583054
rect 509404 582734 510004 582818
rect 509404 582498 509586 582734
rect 509822 582498 510004 582734
rect 509404 547054 510004 582498
rect 509404 546818 509586 547054
rect 509822 546818 510004 547054
rect 509404 546734 510004 546818
rect 509404 546498 509586 546734
rect 509822 546498 510004 546734
rect 509404 511054 510004 546498
rect 509404 510818 509586 511054
rect 509822 510818 510004 511054
rect 509404 510734 510004 510818
rect 509404 510498 509586 510734
rect 509822 510498 510004 510734
rect 509404 475054 510004 510498
rect 509404 474818 509586 475054
rect 509822 474818 510004 475054
rect 509404 474734 510004 474818
rect 509404 474498 509586 474734
rect 509822 474498 510004 474734
rect 509404 439054 510004 474498
rect 509404 438818 509586 439054
rect 509822 438818 510004 439054
rect 509404 438734 510004 438818
rect 509404 438498 509586 438734
rect 509822 438498 510004 438734
rect 509404 403054 510004 438498
rect 509404 402818 509586 403054
rect 509822 402818 510004 403054
rect 509404 402734 510004 402818
rect 509404 402498 509586 402734
rect 509822 402498 510004 402734
rect 509404 367054 510004 402498
rect 509404 366818 509586 367054
rect 509822 366818 510004 367054
rect 509404 366734 510004 366818
rect 509404 366498 509586 366734
rect 509822 366498 510004 366734
rect 509404 331054 510004 366498
rect 509404 330818 509586 331054
rect 509822 330818 510004 331054
rect 509404 330734 510004 330818
rect 509404 330498 509586 330734
rect 509822 330498 510004 330734
rect 509404 295054 510004 330498
rect 509404 294818 509586 295054
rect 509822 294818 510004 295054
rect 509404 294734 510004 294818
rect 509404 294498 509586 294734
rect 509822 294498 510004 294734
rect 509404 259054 510004 294498
rect 509404 258818 509586 259054
rect 509822 258818 510004 259054
rect 509404 258734 510004 258818
rect 509404 258498 509586 258734
rect 509822 258498 510004 258734
rect 509404 223054 510004 258498
rect 509404 222818 509586 223054
rect 509822 222818 510004 223054
rect 509404 222734 510004 222818
rect 509404 222498 509586 222734
rect 509822 222498 510004 222734
rect 509404 187054 510004 222498
rect 509404 186818 509586 187054
rect 509822 186818 510004 187054
rect 509404 186734 510004 186818
rect 509404 186498 509586 186734
rect 509822 186498 510004 186734
rect 509404 151054 510004 186498
rect 509404 150818 509586 151054
rect 509822 150818 510004 151054
rect 509404 150734 510004 150818
rect 509404 150498 509586 150734
rect 509822 150498 510004 150734
rect 509404 115054 510004 150498
rect 509404 114818 509586 115054
rect 509822 114818 510004 115054
rect 509404 114734 510004 114818
rect 509404 114498 509586 114734
rect 509822 114498 510004 114734
rect 509404 79054 510004 114498
rect 509404 78818 509586 79054
rect 509822 78818 510004 79054
rect 509404 78734 510004 78818
rect 509404 78498 509586 78734
rect 509822 78498 510004 78734
rect 509404 43054 510004 78498
rect 509404 42818 509586 43054
rect 509822 42818 510004 43054
rect 509404 42734 510004 42818
rect 509404 42498 509586 42734
rect 509822 42498 510004 42734
rect 509404 7054 510004 42498
rect 509404 6818 509586 7054
rect 509822 6818 510004 7054
rect 509404 6734 510004 6818
rect 509404 6498 509586 6734
rect 509822 6498 510004 6734
rect 509404 -2226 510004 6498
rect 509404 -2462 509586 -2226
rect 509822 -2462 510004 -2226
rect 509404 -2546 510004 -2462
rect 509404 -2782 509586 -2546
rect 509822 -2782 510004 -2546
rect 509404 -3744 510004 -2782
rect 513004 694654 513604 708042
rect 513004 694418 513186 694654
rect 513422 694418 513604 694654
rect 513004 694334 513604 694418
rect 513004 694098 513186 694334
rect 513422 694098 513604 694334
rect 513004 658654 513604 694098
rect 513004 658418 513186 658654
rect 513422 658418 513604 658654
rect 513004 658334 513604 658418
rect 513004 658098 513186 658334
rect 513422 658098 513604 658334
rect 513004 622654 513604 658098
rect 513004 622418 513186 622654
rect 513422 622418 513604 622654
rect 513004 622334 513604 622418
rect 513004 622098 513186 622334
rect 513422 622098 513604 622334
rect 513004 586654 513604 622098
rect 513004 586418 513186 586654
rect 513422 586418 513604 586654
rect 513004 586334 513604 586418
rect 513004 586098 513186 586334
rect 513422 586098 513604 586334
rect 513004 550654 513604 586098
rect 513004 550418 513186 550654
rect 513422 550418 513604 550654
rect 513004 550334 513604 550418
rect 513004 550098 513186 550334
rect 513422 550098 513604 550334
rect 513004 514654 513604 550098
rect 513004 514418 513186 514654
rect 513422 514418 513604 514654
rect 513004 514334 513604 514418
rect 513004 514098 513186 514334
rect 513422 514098 513604 514334
rect 513004 478654 513604 514098
rect 513004 478418 513186 478654
rect 513422 478418 513604 478654
rect 513004 478334 513604 478418
rect 513004 478098 513186 478334
rect 513422 478098 513604 478334
rect 513004 442654 513604 478098
rect 513004 442418 513186 442654
rect 513422 442418 513604 442654
rect 513004 442334 513604 442418
rect 513004 442098 513186 442334
rect 513422 442098 513604 442334
rect 513004 406654 513604 442098
rect 513004 406418 513186 406654
rect 513422 406418 513604 406654
rect 513004 406334 513604 406418
rect 513004 406098 513186 406334
rect 513422 406098 513604 406334
rect 513004 370654 513604 406098
rect 513004 370418 513186 370654
rect 513422 370418 513604 370654
rect 513004 370334 513604 370418
rect 513004 370098 513186 370334
rect 513422 370098 513604 370334
rect 513004 334654 513604 370098
rect 513004 334418 513186 334654
rect 513422 334418 513604 334654
rect 513004 334334 513604 334418
rect 513004 334098 513186 334334
rect 513422 334098 513604 334334
rect 513004 298654 513604 334098
rect 513004 298418 513186 298654
rect 513422 298418 513604 298654
rect 513004 298334 513604 298418
rect 513004 298098 513186 298334
rect 513422 298098 513604 298334
rect 513004 262654 513604 298098
rect 513004 262418 513186 262654
rect 513422 262418 513604 262654
rect 513004 262334 513604 262418
rect 513004 262098 513186 262334
rect 513422 262098 513604 262334
rect 513004 226654 513604 262098
rect 513004 226418 513186 226654
rect 513422 226418 513604 226654
rect 513004 226334 513604 226418
rect 513004 226098 513186 226334
rect 513422 226098 513604 226334
rect 513004 190654 513604 226098
rect 513004 190418 513186 190654
rect 513422 190418 513604 190654
rect 513004 190334 513604 190418
rect 513004 190098 513186 190334
rect 513422 190098 513604 190334
rect 513004 154654 513604 190098
rect 513004 154418 513186 154654
rect 513422 154418 513604 154654
rect 513004 154334 513604 154418
rect 513004 154098 513186 154334
rect 513422 154098 513604 154334
rect 513004 118654 513604 154098
rect 513004 118418 513186 118654
rect 513422 118418 513604 118654
rect 513004 118334 513604 118418
rect 513004 118098 513186 118334
rect 513422 118098 513604 118334
rect 513004 82654 513604 118098
rect 513004 82418 513186 82654
rect 513422 82418 513604 82654
rect 513004 82334 513604 82418
rect 513004 82098 513186 82334
rect 513422 82098 513604 82334
rect 513004 46654 513604 82098
rect 513004 46418 513186 46654
rect 513422 46418 513604 46654
rect 513004 46334 513604 46418
rect 513004 46098 513186 46334
rect 513422 46098 513604 46334
rect 513004 10654 513604 46098
rect 513004 10418 513186 10654
rect 513422 10418 513604 10654
rect 513004 10334 513604 10418
rect 513004 10098 513186 10334
rect 513422 10098 513604 10334
rect 513004 -4106 513604 10098
rect 513004 -4342 513186 -4106
rect 513422 -4342 513604 -4106
rect 513004 -4426 513604 -4342
rect 513004 -4662 513186 -4426
rect 513422 -4662 513604 -4426
rect 513004 -5624 513604 -4662
rect 516604 698254 517204 709922
rect 534604 711418 535204 711440
rect 534604 711182 534786 711418
rect 535022 711182 535204 711418
rect 534604 711098 535204 711182
rect 534604 710862 534786 711098
rect 535022 710862 535204 711098
rect 531004 709538 531604 709560
rect 531004 709302 531186 709538
rect 531422 709302 531604 709538
rect 531004 709218 531604 709302
rect 531004 708982 531186 709218
rect 531422 708982 531604 709218
rect 527404 707658 528004 707680
rect 527404 707422 527586 707658
rect 527822 707422 528004 707658
rect 527404 707338 528004 707422
rect 527404 707102 527586 707338
rect 527822 707102 528004 707338
rect 516604 698018 516786 698254
rect 517022 698018 517204 698254
rect 516604 697934 517204 698018
rect 516604 697698 516786 697934
rect 517022 697698 517204 697934
rect 516604 662254 517204 697698
rect 516604 662018 516786 662254
rect 517022 662018 517204 662254
rect 516604 661934 517204 662018
rect 516604 661698 516786 661934
rect 517022 661698 517204 661934
rect 516604 626254 517204 661698
rect 516604 626018 516786 626254
rect 517022 626018 517204 626254
rect 516604 625934 517204 626018
rect 516604 625698 516786 625934
rect 517022 625698 517204 625934
rect 516604 590254 517204 625698
rect 516604 590018 516786 590254
rect 517022 590018 517204 590254
rect 516604 589934 517204 590018
rect 516604 589698 516786 589934
rect 517022 589698 517204 589934
rect 516604 554254 517204 589698
rect 516604 554018 516786 554254
rect 517022 554018 517204 554254
rect 516604 553934 517204 554018
rect 516604 553698 516786 553934
rect 517022 553698 517204 553934
rect 516604 518254 517204 553698
rect 516604 518018 516786 518254
rect 517022 518018 517204 518254
rect 516604 517934 517204 518018
rect 516604 517698 516786 517934
rect 517022 517698 517204 517934
rect 516604 482254 517204 517698
rect 516604 482018 516786 482254
rect 517022 482018 517204 482254
rect 516604 481934 517204 482018
rect 516604 481698 516786 481934
rect 517022 481698 517204 481934
rect 516604 446254 517204 481698
rect 516604 446018 516786 446254
rect 517022 446018 517204 446254
rect 516604 445934 517204 446018
rect 516604 445698 516786 445934
rect 517022 445698 517204 445934
rect 516604 410254 517204 445698
rect 516604 410018 516786 410254
rect 517022 410018 517204 410254
rect 516604 409934 517204 410018
rect 516604 409698 516786 409934
rect 517022 409698 517204 409934
rect 516604 374254 517204 409698
rect 516604 374018 516786 374254
rect 517022 374018 517204 374254
rect 516604 373934 517204 374018
rect 516604 373698 516786 373934
rect 517022 373698 517204 373934
rect 516604 338254 517204 373698
rect 516604 338018 516786 338254
rect 517022 338018 517204 338254
rect 516604 337934 517204 338018
rect 516604 337698 516786 337934
rect 517022 337698 517204 337934
rect 516604 302254 517204 337698
rect 516604 302018 516786 302254
rect 517022 302018 517204 302254
rect 516604 301934 517204 302018
rect 516604 301698 516786 301934
rect 517022 301698 517204 301934
rect 516604 266254 517204 301698
rect 516604 266018 516786 266254
rect 517022 266018 517204 266254
rect 516604 265934 517204 266018
rect 516604 265698 516786 265934
rect 517022 265698 517204 265934
rect 516604 230254 517204 265698
rect 516604 230018 516786 230254
rect 517022 230018 517204 230254
rect 516604 229934 517204 230018
rect 516604 229698 516786 229934
rect 517022 229698 517204 229934
rect 516604 194254 517204 229698
rect 516604 194018 516786 194254
rect 517022 194018 517204 194254
rect 516604 193934 517204 194018
rect 516604 193698 516786 193934
rect 517022 193698 517204 193934
rect 516604 158254 517204 193698
rect 516604 158018 516786 158254
rect 517022 158018 517204 158254
rect 516604 157934 517204 158018
rect 516604 157698 516786 157934
rect 517022 157698 517204 157934
rect 516604 122254 517204 157698
rect 516604 122018 516786 122254
rect 517022 122018 517204 122254
rect 516604 121934 517204 122018
rect 516604 121698 516786 121934
rect 517022 121698 517204 121934
rect 516604 86254 517204 121698
rect 516604 86018 516786 86254
rect 517022 86018 517204 86254
rect 516604 85934 517204 86018
rect 516604 85698 516786 85934
rect 517022 85698 517204 85934
rect 516604 50254 517204 85698
rect 516604 50018 516786 50254
rect 517022 50018 517204 50254
rect 516604 49934 517204 50018
rect 516604 49698 516786 49934
rect 517022 49698 517204 49934
rect 516604 14254 517204 49698
rect 516604 14018 516786 14254
rect 517022 14018 517204 14254
rect 516604 13934 517204 14018
rect 516604 13698 516786 13934
rect 517022 13698 517204 13934
rect 498604 -7162 498786 -6926
rect 499022 -7162 499204 -6926
rect 498604 -7246 499204 -7162
rect 498604 -7482 498786 -7246
rect 499022 -7482 499204 -7246
rect 498604 -7504 499204 -7482
rect 516604 -5986 517204 13698
rect 523804 705778 524404 705800
rect 523804 705542 523986 705778
rect 524222 705542 524404 705778
rect 523804 705458 524404 705542
rect 523804 705222 523986 705458
rect 524222 705222 524404 705458
rect 523804 669454 524404 705222
rect 523804 669218 523986 669454
rect 524222 669218 524404 669454
rect 523804 669134 524404 669218
rect 523804 668898 523986 669134
rect 524222 668898 524404 669134
rect 523804 633454 524404 668898
rect 523804 633218 523986 633454
rect 524222 633218 524404 633454
rect 523804 633134 524404 633218
rect 523804 632898 523986 633134
rect 524222 632898 524404 633134
rect 523804 597454 524404 632898
rect 523804 597218 523986 597454
rect 524222 597218 524404 597454
rect 523804 597134 524404 597218
rect 523804 596898 523986 597134
rect 524222 596898 524404 597134
rect 523804 561454 524404 596898
rect 523804 561218 523986 561454
rect 524222 561218 524404 561454
rect 523804 561134 524404 561218
rect 523804 560898 523986 561134
rect 524222 560898 524404 561134
rect 523804 525454 524404 560898
rect 523804 525218 523986 525454
rect 524222 525218 524404 525454
rect 523804 525134 524404 525218
rect 523804 524898 523986 525134
rect 524222 524898 524404 525134
rect 523804 489454 524404 524898
rect 523804 489218 523986 489454
rect 524222 489218 524404 489454
rect 523804 489134 524404 489218
rect 523804 488898 523986 489134
rect 524222 488898 524404 489134
rect 523804 453454 524404 488898
rect 523804 453218 523986 453454
rect 524222 453218 524404 453454
rect 523804 453134 524404 453218
rect 523804 452898 523986 453134
rect 524222 452898 524404 453134
rect 523804 417454 524404 452898
rect 523804 417218 523986 417454
rect 524222 417218 524404 417454
rect 523804 417134 524404 417218
rect 523804 416898 523986 417134
rect 524222 416898 524404 417134
rect 523804 381454 524404 416898
rect 523804 381218 523986 381454
rect 524222 381218 524404 381454
rect 523804 381134 524404 381218
rect 523804 380898 523986 381134
rect 524222 380898 524404 381134
rect 523804 345454 524404 380898
rect 523804 345218 523986 345454
rect 524222 345218 524404 345454
rect 523804 345134 524404 345218
rect 523804 344898 523986 345134
rect 524222 344898 524404 345134
rect 523804 309454 524404 344898
rect 523804 309218 523986 309454
rect 524222 309218 524404 309454
rect 523804 309134 524404 309218
rect 523804 308898 523986 309134
rect 524222 308898 524404 309134
rect 523804 273454 524404 308898
rect 523804 273218 523986 273454
rect 524222 273218 524404 273454
rect 523804 273134 524404 273218
rect 523804 272898 523986 273134
rect 524222 272898 524404 273134
rect 523804 237454 524404 272898
rect 523804 237218 523986 237454
rect 524222 237218 524404 237454
rect 523804 237134 524404 237218
rect 523804 236898 523986 237134
rect 524222 236898 524404 237134
rect 523804 201454 524404 236898
rect 523804 201218 523986 201454
rect 524222 201218 524404 201454
rect 523804 201134 524404 201218
rect 523804 200898 523986 201134
rect 524222 200898 524404 201134
rect 523804 165454 524404 200898
rect 523804 165218 523986 165454
rect 524222 165218 524404 165454
rect 523804 165134 524404 165218
rect 523804 164898 523986 165134
rect 524222 164898 524404 165134
rect 523804 129454 524404 164898
rect 523804 129218 523986 129454
rect 524222 129218 524404 129454
rect 523804 129134 524404 129218
rect 523804 128898 523986 129134
rect 524222 128898 524404 129134
rect 523804 93454 524404 128898
rect 523804 93218 523986 93454
rect 524222 93218 524404 93454
rect 523804 93134 524404 93218
rect 523804 92898 523986 93134
rect 524222 92898 524404 93134
rect 523804 57454 524404 92898
rect 523804 57218 523986 57454
rect 524222 57218 524404 57454
rect 523804 57134 524404 57218
rect 523804 56898 523986 57134
rect 524222 56898 524404 57134
rect 523804 21454 524404 56898
rect 523804 21218 523986 21454
rect 524222 21218 524404 21454
rect 523804 21134 524404 21218
rect 523804 20898 523986 21134
rect 524222 20898 524404 21134
rect 523804 -1286 524404 20898
rect 523804 -1522 523986 -1286
rect 524222 -1522 524404 -1286
rect 523804 -1606 524404 -1522
rect 523804 -1842 523986 -1606
rect 524222 -1842 524404 -1606
rect 523804 -1864 524404 -1842
rect 527404 673054 528004 707102
rect 527404 672818 527586 673054
rect 527822 672818 528004 673054
rect 527404 672734 528004 672818
rect 527404 672498 527586 672734
rect 527822 672498 528004 672734
rect 527404 637054 528004 672498
rect 527404 636818 527586 637054
rect 527822 636818 528004 637054
rect 527404 636734 528004 636818
rect 527404 636498 527586 636734
rect 527822 636498 528004 636734
rect 527404 601054 528004 636498
rect 527404 600818 527586 601054
rect 527822 600818 528004 601054
rect 527404 600734 528004 600818
rect 527404 600498 527586 600734
rect 527822 600498 528004 600734
rect 527404 565054 528004 600498
rect 527404 564818 527586 565054
rect 527822 564818 528004 565054
rect 527404 564734 528004 564818
rect 527404 564498 527586 564734
rect 527822 564498 528004 564734
rect 527404 529054 528004 564498
rect 527404 528818 527586 529054
rect 527822 528818 528004 529054
rect 527404 528734 528004 528818
rect 527404 528498 527586 528734
rect 527822 528498 528004 528734
rect 527404 493054 528004 528498
rect 527404 492818 527586 493054
rect 527822 492818 528004 493054
rect 527404 492734 528004 492818
rect 527404 492498 527586 492734
rect 527822 492498 528004 492734
rect 527404 457054 528004 492498
rect 527404 456818 527586 457054
rect 527822 456818 528004 457054
rect 527404 456734 528004 456818
rect 527404 456498 527586 456734
rect 527822 456498 528004 456734
rect 527404 421054 528004 456498
rect 527404 420818 527586 421054
rect 527822 420818 528004 421054
rect 527404 420734 528004 420818
rect 527404 420498 527586 420734
rect 527822 420498 528004 420734
rect 527404 385054 528004 420498
rect 527404 384818 527586 385054
rect 527822 384818 528004 385054
rect 527404 384734 528004 384818
rect 527404 384498 527586 384734
rect 527822 384498 528004 384734
rect 527404 349054 528004 384498
rect 527404 348818 527586 349054
rect 527822 348818 528004 349054
rect 527404 348734 528004 348818
rect 527404 348498 527586 348734
rect 527822 348498 528004 348734
rect 527404 313054 528004 348498
rect 527404 312818 527586 313054
rect 527822 312818 528004 313054
rect 527404 312734 528004 312818
rect 527404 312498 527586 312734
rect 527822 312498 528004 312734
rect 527404 277054 528004 312498
rect 527404 276818 527586 277054
rect 527822 276818 528004 277054
rect 527404 276734 528004 276818
rect 527404 276498 527586 276734
rect 527822 276498 528004 276734
rect 527404 241054 528004 276498
rect 527404 240818 527586 241054
rect 527822 240818 528004 241054
rect 527404 240734 528004 240818
rect 527404 240498 527586 240734
rect 527822 240498 528004 240734
rect 527404 205054 528004 240498
rect 527404 204818 527586 205054
rect 527822 204818 528004 205054
rect 527404 204734 528004 204818
rect 527404 204498 527586 204734
rect 527822 204498 528004 204734
rect 527404 169054 528004 204498
rect 527404 168818 527586 169054
rect 527822 168818 528004 169054
rect 527404 168734 528004 168818
rect 527404 168498 527586 168734
rect 527822 168498 528004 168734
rect 527404 133054 528004 168498
rect 527404 132818 527586 133054
rect 527822 132818 528004 133054
rect 527404 132734 528004 132818
rect 527404 132498 527586 132734
rect 527822 132498 528004 132734
rect 527404 97054 528004 132498
rect 527404 96818 527586 97054
rect 527822 96818 528004 97054
rect 527404 96734 528004 96818
rect 527404 96498 527586 96734
rect 527822 96498 528004 96734
rect 527404 61054 528004 96498
rect 527404 60818 527586 61054
rect 527822 60818 528004 61054
rect 527404 60734 528004 60818
rect 527404 60498 527586 60734
rect 527822 60498 528004 60734
rect 527404 25054 528004 60498
rect 527404 24818 527586 25054
rect 527822 24818 528004 25054
rect 527404 24734 528004 24818
rect 527404 24498 527586 24734
rect 527822 24498 528004 24734
rect 527404 -3166 528004 24498
rect 527404 -3402 527586 -3166
rect 527822 -3402 528004 -3166
rect 527404 -3486 528004 -3402
rect 527404 -3722 527586 -3486
rect 527822 -3722 528004 -3486
rect 527404 -3744 528004 -3722
rect 531004 676654 531604 708982
rect 531004 676418 531186 676654
rect 531422 676418 531604 676654
rect 531004 676334 531604 676418
rect 531004 676098 531186 676334
rect 531422 676098 531604 676334
rect 531004 640654 531604 676098
rect 531004 640418 531186 640654
rect 531422 640418 531604 640654
rect 531004 640334 531604 640418
rect 531004 640098 531186 640334
rect 531422 640098 531604 640334
rect 531004 604654 531604 640098
rect 531004 604418 531186 604654
rect 531422 604418 531604 604654
rect 531004 604334 531604 604418
rect 531004 604098 531186 604334
rect 531422 604098 531604 604334
rect 531004 568654 531604 604098
rect 531004 568418 531186 568654
rect 531422 568418 531604 568654
rect 531004 568334 531604 568418
rect 531004 568098 531186 568334
rect 531422 568098 531604 568334
rect 531004 532654 531604 568098
rect 531004 532418 531186 532654
rect 531422 532418 531604 532654
rect 531004 532334 531604 532418
rect 531004 532098 531186 532334
rect 531422 532098 531604 532334
rect 531004 496654 531604 532098
rect 531004 496418 531186 496654
rect 531422 496418 531604 496654
rect 531004 496334 531604 496418
rect 531004 496098 531186 496334
rect 531422 496098 531604 496334
rect 531004 460654 531604 496098
rect 531004 460418 531186 460654
rect 531422 460418 531604 460654
rect 531004 460334 531604 460418
rect 531004 460098 531186 460334
rect 531422 460098 531604 460334
rect 531004 424654 531604 460098
rect 531004 424418 531186 424654
rect 531422 424418 531604 424654
rect 531004 424334 531604 424418
rect 531004 424098 531186 424334
rect 531422 424098 531604 424334
rect 531004 388654 531604 424098
rect 531004 388418 531186 388654
rect 531422 388418 531604 388654
rect 531004 388334 531604 388418
rect 531004 388098 531186 388334
rect 531422 388098 531604 388334
rect 531004 352654 531604 388098
rect 531004 352418 531186 352654
rect 531422 352418 531604 352654
rect 531004 352334 531604 352418
rect 531004 352098 531186 352334
rect 531422 352098 531604 352334
rect 531004 316654 531604 352098
rect 531004 316418 531186 316654
rect 531422 316418 531604 316654
rect 531004 316334 531604 316418
rect 531004 316098 531186 316334
rect 531422 316098 531604 316334
rect 531004 280654 531604 316098
rect 531004 280418 531186 280654
rect 531422 280418 531604 280654
rect 531004 280334 531604 280418
rect 531004 280098 531186 280334
rect 531422 280098 531604 280334
rect 531004 244654 531604 280098
rect 531004 244418 531186 244654
rect 531422 244418 531604 244654
rect 531004 244334 531604 244418
rect 531004 244098 531186 244334
rect 531422 244098 531604 244334
rect 531004 208654 531604 244098
rect 531004 208418 531186 208654
rect 531422 208418 531604 208654
rect 531004 208334 531604 208418
rect 531004 208098 531186 208334
rect 531422 208098 531604 208334
rect 531004 172654 531604 208098
rect 531004 172418 531186 172654
rect 531422 172418 531604 172654
rect 531004 172334 531604 172418
rect 531004 172098 531186 172334
rect 531422 172098 531604 172334
rect 531004 136654 531604 172098
rect 531004 136418 531186 136654
rect 531422 136418 531604 136654
rect 531004 136334 531604 136418
rect 531004 136098 531186 136334
rect 531422 136098 531604 136334
rect 531004 100654 531604 136098
rect 531004 100418 531186 100654
rect 531422 100418 531604 100654
rect 531004 100334 531604 100418
rect 531004 100098 531186 100334
rect 531422 100098 531604 100334
rect 531004 64654 531604 100098
rect 531004 64418 531186 64654
rect 531422 64418 531604 64654
rect 531004 64334 531604 64418
rect 531004 64098 531186 64334
rect 531422 64098 531604 64334
rect 531004 28654 531604 64098
rect 531004 28418 531186 28654
rect 531422 28418 531604 28654
rect 531004 28334 531604 28418
rect 531004 28098 531186 28334
rect 531422 28098 531604 28334
rect 531004 -5046 531604 28098
rect 531004 -5282 531186 -5046
rect 531422 -5282 531604 -5046
rect 531004 -5366 531604 -5282
rect 531004 -5602 531186 -5366
rect 531422 -5602 531604 -5366
rect 531004 -5624 531604 -5602
rect 534604 680254 535204 710862
rect 552604 710478 553204 711440
rect 552604 710242 552786 710478
rect 553022 710242 553204 710478
rect 552604 710158 553204 710242
rect 552604 709922 552786 710158
rect 553022 709922 553204 710158
rect 549004 708598 549604 709560
rect 549004 708362 549186 708598
rect 549422 708362 549604 708598
rect 549004 708278 549604 708362
rect 549004 708042 549186 708278
rect 549422 708042 549604 708278
rect 545404 706718 546004 707680
rect 545404 706482 545586 706718
rect 545822 706482 546004 706718
rect 545404 706398 546004 706482
rect 545404 706162 545586 706398
rect 545822 706162 546004 706398
rect 534604 680018 534786 680254
rect 535022 680018 535204 680254
rect 534604 679934 535204 680018
rect 534604 679698 534786 679934
rect 535022 679698 535204 679934
rect 534604 644254 535204 679698
rect 534604 644018 534786 644254
rect 535022 644018 535204 644254
rect 534604 643934 535204 644018
rect 534604 643698 534786 643934
rect 535022 643698 535204 643934
rect 534604 608254 535204 643698
rect 534604 608018 534786 608254
rect 535022 608018 535204 608254
rect 534604 607934 535204 608018
rect 534604 607698 534786 607934
rect 535022 607698 535204 607934
rect 534604 572254 535204 607698
rect 534604 572018 534786 572254
rect 535022 572018 535204 572254
rect 534604 571934 535204 572018
rect 534604 571698 534786 571934
rect 535022 571698 535204 571934
rect 534604 536254 535204 571698
rect 534604 536018 534786 536254
rect 535022 536018 535204 536254
rect 534604 535934 535204 536018
rect 534604 535698 534786 535934
rect 535022 535698 535204 535934
rect 534604 500254 535204 535698
rect 534604 500018 534786 500254
rect 535022 500018 535204 500254
rect 534604 499934 535204 500018
rect 534604 499698 534786 499934
rect 535022 499698 535204 499934
rect 534604 464254 535204 499698
rect 534604 464018 534786 464254
rect 535022 464018 535204 464254
rect 534604 463934 535204 464018
rect 534604 463698 534786 463934
rect 535022 463698 535204 463934
rect 534604 428254 535204 463698
rect 534604 428018 534786 428254
rect 535022 428018 535204 428254
rect 534604 427934 535204 428018
rect 534604 427698 534786 427934
rect 535022 427698 535204 427934
rect 534604 392254 535204 427698
rect 534604 392018 534786 392254
rect 535022 392018 535204 392254
rect 534604 391934 535204 392018
rect 534604 391698 534786 391934
rect 535022 391698 535204 391934
rect 534604 356254 535204 391698
rect 534604 356018 534786 356254
rect 535022 356018 535204 356254
rect 534604 355934 535204 356018
rect 534604 355698 534786 355934
rect 535022 355698 535204 355934
rect 534604 320254 535204 355698
rect 534604 320018 534786 320254
rect 535022 320018 535204 320254
rect 534604 319934 535204 320018
rect 534604 319698 534786 319934
rect 535022 319698 535204 319934
rect 534604 284254 535204 319698
rect 534604 284018 534786 284254
rect 535022 284018 535204 284254
rect 534604 283934 535204 284018
rect 534604 283698 534786 283934
rect 535022 283698 535204 283934
rect 534604 248254 535204 283698
rect 534604 248018 534786 248254
rect 535022 248018 535204 248254
rect 534604 247934 535204 248018
rect 534604 247698 534786 247934
rect 535022 247698 535204 247934
rect 534604 212254 535204 247698
rect 534604 212018 534786 212254
rect 535022 212018 535204 212254
rect 534604 211934 535204 212018
rect 534604 211698 534786 211934
rect 535022 211698 535204 211934
rect 534604 176254 535204 211698
rect 534604 176018 534786 176254
rect 535022 176018 535204 176254
rect 534604 175934 535204 176018
rect 534604 175698 534786 175934
rect 535022 175698 535204 175934
rect 534604 140254 535204 175698
rect 534604 140018 534786 140254
rect 535022 140018 535204 140254
rect 534604 139934 535204 140018
rect 534604 139698 534786 139934
rect 535022 139698 535204 139934
rect 534604 104254 535204 139698
rect 534604 104018 534786 104254
rect 535022 104018 535204 104254
rect 534604 103934 535204 104018
rect 534604 103698 534786 103934
rect 535022 103698 535204 103934
rect 534604 68254 535204 103698
rect 534604 68018 534786 68254
rect 535022 68018 535204 68254
rect 534604 67934 535204 68018
rect 534604 67698 534786 67934
rect 535022 67698 535204 67934
rect 534604 32254 535204 67698
rect 534604 32018 534786 32254
rect 535022 32018 535204 32254
rect 534604 31934 535204 32018
rect 534604 31698 534786 31934
rect 535022 31698 535204 31934
rect 516604 -6222 516786 -5986
rect 517022 -6222 517204 -5986
rect 516604 -6306 517204 -6222
rect 516604 -6542 516786 -6306
rect 517022 -6542 517204 -6306
rect 516604 -7504 517204 -6542
rect 534604 -6926 535204 31698
rect 541804 704838 542404 705800
rect 541804 704602 541986 704838
rect 542222 704602 542404 704838
rect 541804 704518 542404 704602
rect 541804 704282 541986 704518
rect 542222 704282 542404 704518
rect 541804 687454 542404 704282
rect 541804 687218 541986 687454
rect 542222 687218 542404 687454
rect 541804 687134 542404 687218
rect 541804 686898 541986 687134
rect 542222 686898 542404 687134
rect 541804 651454 542404 686898
rect 541804 651218 541986 651454
rect 542222 651218 542404 651454
rect 541804 651134 542404 651218
rect 541804 650898 541986 651134
rect 542222 650898 542404 651134
rect 541804 615454 542404 650898
rect 541804 615218 541986 615454
rect 542222 615218 542404 615454
rect 541804 615134 542404 615218
rect 541804 614898 541986 615134
rect 542222 614898 542404 615134
rect 541804 579454 542404 614898
rect 541804 579218 541986 579454
rect 542222 579218 542404 579454
rect 541804 579134 542404 579218
rect 541804 578898 541986 579134
rect 542222 578898 542404 579134
rect 541804 543454 542404 578898
rect 541804 543218 541986 543454
rect 542222 543218 542404 543454
rect 541804 543134 542404 543218
rect 541804 542898 541986 543134
rect 542222 542898 542404 543134
rect 541804 507454 542404 542898
rect 541804 507218 541986 507454
rect 542222 507218 542404 507454
rect 541804 507134 542404 507218
rect 541804 506898 541986 507134
rect 542222 506898 542404 507134
rect 541804 471454 542404 506898
rect 541804 471218 541986 471454
rect 542222 471218 542404 471454
rect 541804 471134 542404 471218
rect 541804 470898 541986 471134
rect 542222 470898 542404 471134
rect 541804 435454 542404 470898
rect 541804 435218 541986 435454
rect 542222 435218 542404 435454
rect 541804 435134 542404 435218
rect 541804 434898 541986 435134
rect 542222 434898 542404 435134
rect 541804 399454 542404 434898
rect 541804 399218 541986 399454
rect 542222 399218 542404 399454
rect 541804 399134 542404 399218
rect 541804 398898 541986 399134
rect 542222 398898 542404 399134
rect 541804 363454 542404 398898
rect 541804 363218 541986 363454
rect 542222 363218 542404 363454
rect 541804 363134 542404 363218
rect 541804 362898 541986 363134
rect 542222 362898 542404 363134
rect 541804 327454 542404 362898
rect 541804 327218 541986 327454
rect 542222 327218 542404 327454
rect 541804 327134 542404 327218
rect 541804 326898 541986 327134
rect 542222 326898 542404 327134
rect 541804 291454 542404 326898
rect 541804 291218 541986 291454
rect 542222 291218 542404 291454
rect 541804 291134 542404 291218
rect 541804 290898 541986 291134
rect 542222 290898 542404 291134
rect 541804 255454 542404 290898
rect 541804 255218 541986 255454
rect 542222 255218 542404 255454
rect 541804 255134 542404 255218
rect 541804 254898 541986 255134
rect 542222 254898 542404 255134
rect 541804 219454 542404 254898
rect 541804 219218 541986 219454
rect 542222 219218 542404 219454
rect 541804 219134 542404 219218
rect 541804 218898 541986 219134
rect 542222 218898 542404 219134
rect 541804 183454 542404 218898
rect 541804 183218 541986 183454
rect 542222 183218 542404 183454
rect 541804 183134 542404 183218
rect 541804 182898 541986 183134
rect 542222 182898 542404 183134
rect 541804 147454 542404 182898
rect 541804 147218 541986 147454
rect 542222 147218 542404 147454
rect 541804 147134 542404 147218
rect 541804 146898 541986 147134
rect 542222 146898 542404 147134
rect 541804 111454 542404 146898
rect 541804 111218 541986 111454
rect 542222 111218 542404 111454
rect 541804 111134 542404 111218
rect 541804 110898 541986 111134
rect 542222 110898 542404 111134
rect 541804 75454 542404 110898
rect 541804 75218 541986 75454
rect 542222 75218 542404 75454
rect 541804 75134 542404 75218
rect 541804 74898 541986 75134
rect 542222 74898 542404 75134
rect 541804 39454 542404 74898
rect 541804 39218 541986 39454
rect 542222 39218 542404 39454
rect 541804 39134 542404 39218
rect 541804 38898 541986 39134
rect 542222 38898 542404 39134
rect 541804 3454 542404 38898
rect 541804 3218 541986 3454
rect 542222 3218 542404 3454
rect 541804 3134 542404 3218
rect 541804 2898 541986 3134
rect 542222 2898 542404 3134
rect 541804 -346 542404 2898
rect 541804 -582 541986 -346
rect 542222 -582 542404 -346
rect 541804 -666 542404 -582
rect 541804 -902 541986 -666
rect 542222 -902 542404 -666
rect 541804 -1864 542404 -902
rect 545404 691054 546004 706162
rect 545404 690818 545586 691054
rect 545822 690818 546004 691054
rect 545404 690734 546004 690818
rect 545404 690498 545586 690734
rect 545822 690498 546004 690734
rect 545404 655054 546004 690498
rect 545404 654818 545586 655054
rect 545822 654818 546004 655054
rect 545404 654734 546004 654818
rect 545404 654498 545586 654734
rect 545822 654498 546004 654734
rect 545404 619054 546004 654498
rect 545404 618818 545586 619054
rect 545822 618818 546004 619054
rect 545404 618734 546004 618818
rect 545404 618498 545586 618734
rect 545822 618498 546004 618734
rect 545404 583054 546004 618498
rect 545404 582818 545586 583054
rect 545822 582818 546004 583054
rect 545404 582734 546004 582818
rect 545404 582498 545586 582734
rect 545822 582498 546004 582734
rect 545404 547054 546004 582498
rect 545404 546818 545586 547054
rect 545822 546818 546004 547054
rect 545404 546734 546004 546818
rect 545404 546498 545586 546734
rect 545822 546498 546004 546734
rect 545404 511054 546004 546498
rect 545404 510818 545586 511054
rect 545822 510818 546004 511054
rect 545404 510734 546004 510818
rect 545404 510498 545586 510734
rect 545822 510498 546004 510734
rect 545404 475054 546004 510498
rect 545404 474818 545586 475054
rect 545822 474818 546004 475054
rect 545404 474734 546004 474818
rect 545404 474498 545586 474734
rect 545822 474498 546004 474734
rect 545404 439054 546004 474498
rect 545404 438818 545586 439054
rect 545822 438818 546004 439054
rect 545404 438734 546004 438818
rect 545404 438498 545586 438734
rect 545822 438498 546004 438734
rect 545404 403054 546004 438498
rect 545404 402818 545586 403054
rect 545822 402818 546004 403054
rect 545404 402734 546004 402818
rect 545404 402498 545586 402734
rect 545822 402498 546004 402734
rect 545404 367054 546004 402498
rect 545404 366818 545586 367054
rect 545822 366818 546004 367054
rect 545404 366734 546004 366818
rect 545404 366498 545586 366734
rect 545822 366498 546004 366734
rect 545404 331054 546004 366498
rect 545404 330818 545586 331054
rect 545822 330818 546004 331054
rect 545404 330734 546004 330818
rect 545404 330498 545586 330734
rect 545822 330498 546004 330734
rect 545404 295054 546004 330498
rect 545404 294818 545586 295054
rect 545822 294818 546004 295054
rect 545404 294734 546004 294818
rect 545404 294498 545586 294734
rect 545822 294498 546004 294734
rect 545404 259054 546004 294498
rect 545404 258818 545586 259054
rect 545822 258818 546004 259054
rect 545404 258734 546004 258818
rect 545404 258498 545586 258734
rect 545822 258498 546004 258734
rect 545404 223054 546004 258498
rect 545404 222818 545586 223054
rect 545822 222818 546004 223054
rect 545404 222734 546004 222818
rect 545404 222498 545586 222734
rect 545822 222498 546004 222734
rect 545404 187054 546004 222498
rect 545404 186818 545586 187054
rect 545822 186818 546004 187054
rect 545404 186734 546004 186818
rect 545404 186498 545586 186734
rect 545822 186498 546004 186734
rect 545404 151054 546004 186498
rect 545404 150818 545586 151054
rect 545822 150818 546004 151054
rect 545404 150734 546004 150818
rect 545404 150498 545586 150734
rect 545822 150498 546004 150734
rect 545404 115054 546004 150498
rect 545404 114818 545586 115054
rect 545822 114818 546004 115054
rect 545404 114734 546004 114818
rect 545404 114498 545586 114734
rect 545822 114498 546004 114734
rect 545404 79054 546004 114498
rect 545404 78818 545586 79054
rect 545822 78818 546004 79054
rect 545404 78734 546004 78818
rect 545404 78498 545586 78734
rect 545822 78498 546004 78734
rect 545404 43054 546004 78498
rect 545404 42818 545586 43054
rect 545822 42818 546004 43054
rect 545404 42734 546004 42818
rect 545404 42498 545586 42734
rect 545822 42498 546004 42734
rect 545404 7054 546004 42498
rect 545404 6818 545586 7054
rect 545822 6818 546004 7054
rect 545404 6734 546004 6818
rect 545404 6498 545586 6734
rect 545822 6498 546004 6734
rect 545404 -2226 546004 6498
rect 545404 -2462 545586 -2226
rect 545822 -2462 546004 -2226
rect 545404 -2546 546004 -2462
rect 545404 -2782 545586 -2546
rect 545822 -2782 546004 -2546
rect 545404 -3744 546004 -2782
rect 549004 694654 549604 708042
rect 549004 694418 549186 694654
rect 549422 694418 549604 694654
rect 549004 694334 549604 694418
rect 549004 694098 549186 694334
rect 549422 694098 549604 694334
rect 549004 658654 549604 694098
rect 549004 658418 549186 658654
rect 549422 658418 549604 658654
rect 549004 658334 549604 658418
rect 549004 658098 549186 658334
rect 549422 658098 549604 658334
rect 549004 622654 549604 658098
rect 549004 622418 549186 622654
rect 549422 622418 549604 622654
rect 549004 622334 549604 622418
rect 549004 622098 549186 622334
rect 549422 622098 549604 622334
rect 549004 586654 549604 622098
rect 549004 586418 549186 586654
rect 549422 586418 549604 586654
rect 549004 586334 549604 586418
rect 549004 586098 549186 586334
rect 549422 586098 549604 586334
rect 549004 550654 549604 586098
rect 549004 550418 549186 550654
rect 549422 550418 549604 550654
rect 549004 550334 549604 550418
rect 549004 550098 549186 550334
rect 549422 550098 549604 550334
rect 549004 514654 549604 550098
rect 549004 514418 549186 514654
rect 549422 514418 549604 514654
rect 549004 514334 549604 514418
rect 549004 514098 549186 514334
rect 549422 514098 549604 514334
rect 549004 478654 549604 514098
rect 549004 478418 549186 478654
rect 549422 478418 549604 478654
rect 549004 478334 549604 478418
rect 549004 478098 549186 478334
rect 549422 478098 549604 478334
rect 549004 442654 549604 478098
rect 549004 442418 549186 442654
rect 549422 442418 549604 442654
rect 549004 442334 549604 442418
rect 549004 442098 549186 442334
rect 549422 442098 549604 442334
rect 549004 406654 549604 442098
rect 549004 406418 549186 406654
rect 549422 406418 549604 406654
rect 549004 406334 549604 406418
rect 549004 406098 549186 406334
rect 549422 406098 549604 406334
rect 549004 370654 549604 406098
rect 549004 370418 549186 370654
rect 549422 370418 549604 370654
rect 549004 370334 549604 370418
rect 549004 370098 549186 370334
rect 549422 370098 549604 370334
rect 549004 334654 549604 370098
rect 549004 334418 549186 334654
rect 549422 334418 549604 334654
rect 549004 334334 549604 334418
rect 549004 334098 549186 334334
rect 549422 334098 549604 334334
rect 549004 298654 549604 334098
rect 549004 298418 549186 298654
rect 549422 298418 549604 298654
rect 549004 298334 549604 298418
rect 549004 298098 549186 298334
rect 549422 298098 549604 298334
rect 549004 262654 549604 298098
rect 549004 262418 549186 262654
rect 549422 262418 549604 262654
rect 549004 262334 549604 262418
rect 549004 262098 549186 262334
rect 549422 262098 549604 262334
rect 549004 226654 549604 262098
rect 549004 226418 549186 226654
rect 549422 226418 549604 226654
rect 549004 226334 549604 226418
rect 549004 226098 549186 226334
rect 549422 226098 549604 226334
rect 549004 190654 549604 226098
rect 549004 190418 549186 190654
rect 549422 190418 549604 190654
rect 549004 190334 549604 190418
rect 549004 190098 549186 190334
rect 549422 190098 549604 190334
rect 549004 154654 549604 190098
rect 549004 154418 549186 154654
rect 549422 154418 549604 154654
rect 549004 154334 549604 154418
rect 549004 154098 549186 154334
rect 549422 154098 549604 154334
rect 549004 118654 549604 154098
rect 549004 118418 549186 118654
rect 549422 118418 549604 118654
rect 549004 118334 549604 118418
rect 549004 118098 549186 118334
rect 549422 118098 549604 118334
rect 549004 82654 549604 118098
rect 549004 82418 549186 82654
rect 549422 82418 549604 82654
rect 549004 82334 549604 82418
rect 549004 82098 549186 82334
rect 549422 82098 549604 82334
rect 549004 46654 549604 82098
rect 549004 46418 549186 46654
rect 549422 46418 549604 46654
rect 549004 46334 549604 46418
rect 549004 46098 549186 46334
rect 549422 46098 549604 46334
rect 549004 10654 549604 46098
rect 549004 10418 549186 10654
rect 549422 10418 549604 10654
rect 549004 10334 549604 10418
rect 549004 10098 549186 10334
rect 549422 10098 549604 10334
rect 549004 -4106 549604 10098
rect 549004 -4342 549186 -4106
rect 549422 -4342 549604 -4106
rect 549004 -4426 549604 -4342
rect 549004 -4662 549186 -4426
rect 549422 -4662 549604 -4426
rect 549004 -5624 549604 -4662
rect 552604 698254 553204 709922
rect 570604 711418 571204 711440
rect 570604 711182 570786 711418
rect 571022 711182 571204 711418
rect 570604 711098 571204 711182
rect 570604 710862 570786 711098
rect 571022 710862 571204 711098
rect 567004 709538 567604 709560
rect 567004 709302 567186 709538
rect 567422 709302 567604 709538
rect 567004 709218 567604 709302
rect 567004 708982 567186 709218
rect 567422 708982 567604 709218
rect 563404 707658 564004 707680
rect 563404 707422 563586 707658
rect 563822 707422 564004 707658
rect 563404 707338 564004 707422
rect 563404 707102 563586 707338
rect 563822 707102 564004 707338
rect 552604 698018 552786 698254
rect 553022 698018 553204 698254
rect 552604 697934 553204 698018
rect 552604 697698 552786 697934
rect 553022 697698 553204 697934
rect 552604 662254 553204 697698
rect 552604 662018 552786 662254
rect 553022 662018 553204 662254
rect 552604 661934 553204 662018
rect 552604 661698 552786 661934
rect 553022 661698 553204 661934
rect 552604 626254 553204 661698
rect 552604 626018 552786 626254
rect 553022 626018 553204 626254
rect 552604 625934 553204 626018
rect 552604 625698 552786 625934
rect 553022 625698 553204 625934
rect 552604 590254 553204 625698
rect 552604 590018 552786 590254
rect 553022 590018 553204 590254
rect 552604 589934 553204 590018
rect 552604 589698 552786 589934
rect 553022 589698 553204 589934
rect 552604 554254 553204 589698
rect 552604 554018 552786 554254
rect 553022 554018 553204 554254
rect 552604 553934 553204 554018
rect 552604 553698 552786 553934
rect 553022 553698 553204 553934
rect 552604 518254 553204 553698
rect 552604 518018 552786 518254
rect 553022 518018 553204 518254
rect 552604 517934 553204 518018
rect 552604 517698 552786 517934
rect 553022 517698 553204 517934
rect 552604 482254 553204 517698
rect 552604 482018 552786 482254
rect 553022 482018 553204 482254
rect 552604 481934 553204 482018
rect 552604 481698 552786 481934
rect 553022 481698 553204 481934
rect 552604 446254 553204 481698
rect 552604 446018 552786 446254
rect 553022 446018 553204 446254
rect 552604 445934 553204 446018
rect 552604 445698 552786 445934
rect 553022 445698 553204 445934
rect 552604 410254 553204 445698
rect 552604 410018 552786 410254
rect 553022 410018 553204 410254
rect 552604 409934 553204 410018
rect 552604 409698 552786 409934
rect 553022 409698 553204 409934
rect 552604 374254 553204 409698
rect 552604 374018 552786 374254
rect 553022 374018 553204 374254
rect 552604 373934 553204 374018
rect 552604 373698 552786 373934
rect 553022 373698 553204 373934
rect 552604 338254 553204 373698
rect 552604 338018 552786 338254
rect 553022 338018 553204 338254
rect 552604 337934 553204 338018
rect 552604 337698 552786 337934
rect 553022 337698 553204 337934
rect 552604 302254 553204 337698
rect 552604 302018 552786 302254
rect 553022 302018 553204 302254
rect 552604 301934 553204 302018
rect 552604 301698 552786 301934
rect 553022 301698 553204 301934
rect 552604 266254 553204 301698
rect 552604 266018 552786 266254
rect 553022 266018 553204 266254
rect 552604 265934 553204 266018
rect 552604 265698 552786 265934
rect 553022 265698 553204 265934
rect 552604 230254 553204 265698
rect 552604 230018 552786 230254
rect 553022 230018 553204 230254
rect 552604 229934 553204 230018
rect 552604 229698 552786 229934
rect 553022 229698 553204 229934
rect 552604 194254 553204 229698
rect 552604 194018 552786 194254
rect 553022 194018 553204 194254
rect 552604 193934 553204 194018
rect 552604 193698 552786 193934
rect 553022 193698 553204 193934
rect 552604 158254 553204 193698
rect 552604 158018 552786 158254
rect 553022 158018 553204 158254
rect 552604 157934 553204 158018
rect 552604 157698 552786 157934
rect 553022 157698 553204 157934
rect 552604 122254 553204 157698
rect 552604 122018 552786 122254
rect 553022 122018 553204 122254
rect 552604 121934 553204 122018
rect 552604 121698 552786 121934
rect 553022 121698 553204 121934
rect 552604 86254 553204 121698
rect 552604 86018 552786 86254
rect 553022 86018 553204 86254
rect 552604 85934 553204 86018
rect 552604 85698 552786 85934
rect 553022 85698 553204 85934
rect 552604 50254 553204 85698
rect 552604 50018 552786 50254
rect 553022 50018 553204 50254
rect 552604 49934 553204 50018
rect 552604 49698 552786 49934
rect 553022 49698 553204 49934
rect 552604 14254 553204 49698
rect 552604 14018 552786 14254
rect 553022 14018 553204 14254
rect 552604 13934 553204 14018
rect 552604 13698 552786 13934
rect 553022 13698 553204 13934
rect 534604 -7162 534786 -6926
rect 535022 -7162 535204 -6926
rect 534604 -7246 535204 -7162
rect 534604 -7482 534786 -7246
rect 535022 -7482 535204 -7246
rect 534604 -7504 535204 -7482
rect 552604 -5986 553204 13698
rect 559804 705778 560404 705800
rect 559804 705542 559986 705778
rect 560222 705542 560404 705778
rect 559804 705458 560404 705542
rect 559804 705222 559986 705458
rect 560222 705222 560404 705458
rect 559804 669454 560404 705222
rect 559804 669218 559986 669454
rect 560222 669218 560404 669454
rect 559804 669134 560404 669218
rect 559804 668898 559986 669134
rect 560222 668898 560404 669134
rect 559804 633454 560404 668898
rect 559804 633218 559986 633454
rect 560222 633218 560404 633454
rect 559804 633134 560404 633218
rect 559804 632898 559986 633134
rect 560222 632898 560404 633134
rect 559804 597454 560404 632898
rect 559804 597218 559986 597454
rect 560222 597218 560404 597454
rect 559804 597134 560404 597218
rect 559804 596898 559986 597134
rect 560222 596898 560404 597134
rect 559804 561454 560404 596898
rect 559804 561218 559986 561454
rect 560222 561218 560404 561454
rect 559804 561134 560404 561218
rect 559804 560898 559986 561134
rect 560222 560898 560404 561134
rect 559804 525454 560404 560898
rect 559804 525218 559986 525454
rect 560222 525218 560404 525454
rect 559804 525134 560404 525218
rect 559804 524898 559986 525134
rect 560222 524898 560404 525134
rect 559804 489454 560404 524898
rect 559804 489218 559986 489454
rect 560222 489218 560404 489454
rect 559804 489134 560404 489218
rect 559804 488898 559986 489134
rect 560222 488898 560404 489134
rect 559804 453454 560404 488898
rect 559804 453218 559986 453454
rect 560222 453218 560404 453454
rect 559804 453134 560404 453218
rect 559804 452898 559986 453134
rect 560222 452898 560404 453134
rect 559804 417454 560404 452898
rect 559804 417218 559986 417454
rect 560222 417218 560404 417454
rect 559804 417134 560404 417218
rect 559804 416898 559986 417134
rect 560222 416898 560404 417134
rect 559804 381454 560404 416898
rect 559804 381218 559986 381454
rect 560222 381218 560404 381454
rect 559804 381134 560404 381218
rect 559804 380898 559986 381134
rect 560222 380898 560404 381134
rect 559804 345454 560404 380898
rect 559804 345218 559986 345454
rect 560222 345218 560404 345454
rect 559804 345134 560404 345218
rect 559804 344898 559986 345134
rect 560222 344898 560404 345134
rect 559804 309454 560404 344898
rect 559804 309218 559986 309454
rect 560222 309218 560404 309454
rect 559804 309134 560404 309218
rect 559804 308898 559986 309134
rect 560222 308898 560404 309134
rect 559804 273454 560404 308898
rect 559804 273218 559986 273454
rect 560222 273218 560404 273454
rect 559804 273134 560404 273218
rect 559804 272898 559986 273134
rect 560222 272898 560404 273134
rect 559804 237454 560404 272898
rect 559804 237218 559986 237454
rect 560222 237218 560404 237454
rect 559804 237134 560404 237218
rect 559804 236898 559986 237134
rect 560222 236898 560404 237134
rect 559804 201454 560404 236898
rect 559804 201218 559986 201454
rect 560222 201218 560404 201454
rect 559804 201134 560404 201218
rect 559804 200898 559986 201134
rect 560222 200898 560404 201134
rect 559804 165454 560404 200898
rect 559804 165218 559986 165454
rect 560222 165218 560404 165454
rect 559804 165134 560404 165218
rect 559804 164898 559986 165134
rect 560222 164898 560404 165134
rect 559804 129454 560404 164898
rect 559804 129218 559986 129454
rect 560222 129218 560404 129454
rect 559804 129134 560404 129218
rect 559804 128898 559986 129134
rect 560222 128898 560404 129134
rect 559804 93454 560404 128898
rect 559804 93218 559986 93454
rect 560222 93218 560404 93454
rect 559804 93134 560404 93218
rect 559804 92898 559986 93134
rect 560222 92898 560404 93134
rect 559804 57454 560404 92898
rect 559804 57218 559986 57454
rect 560222 57218 560404 57454
rect 559804 57134 560404 57218
rect 559804 56898 559986 57134
rect 560222 56898 560404 57134
rect 559804 21454 560404 56898
rect 559804 21218 559986 21454
rect 560222 21218 560404 21454
rect 559804 21134 560404 21218
rect 559804 20898 559986 21134
rect 560222 20898 560404 21134
rect 559804 -1286 560404 20898
rect 559804 -1522 559986 -1286
rect 560222 -1522 560404 -1286
rect 559804 -1606 560404 -1522
rect 559804 -1842 559986 -1606
rect 560222 -1842 560404 -1606
rect 559804 -1864 560404 -1842
rect 563404 673054 564004 707102
rect 563404 672818 563586 673054
rect 563822 672818 564004 673054
rect 563404 672734 564004 672818
rect 563404 672498 563586 672734
rect 563822 672498 564004 672734
rect 563404 637054 564004 672498
rect 563404 636818 563586 637054
rect 563822 636818 564004 637054
rect 563404 636734 564004 636818
rect 563404 636498 563586 636734
rect 563822 636498 564004 636734
rect 563404 601054 564004 636498
rect 563404 600818 563586 601054
rect 563822 600818 564004 601054
rect 563404 600734 564004 600818
rect 563404 600498 563586 600734
rect 563822 600498 564004 600734
rect 563404 565054 564004 600498
rect 563404 564818 563586 565054
rect 563822 564818 564004 565054
rect 563404 564734 564004 564818
rect 563404 564498 563586 564734
rect 563822 564498 564004 564734
rect 563404 529054 564004 564498
rect 563404 528818 563586 529054
rect 563822 528818 564004 529054
rect 563404 528734 564004 528818
rect 563404 528498 563586 528734
rect 563822 528498 564004 528734
rect 563404 493054 564004 528498
rect 563404 492818 563586 493054
rect 563822 492818 564004 493054
rect 563404 492734 564004 492818
rect 563404 492498 563586 492734
rect 563822 492498 564004 492734
rect 563404 457054 564004 492498
rect 563404 456818 563586 457054
rect 563822 456818 564004 457054
rect 563404 456734 564004 456818
rect 563404 456498 563586 456734
rect 563822 456498 564004 456734
rect 563404 421054 564004 456498
rect 563404 420818 563586 421054
rect 563822 420818 564004 421054
rect 563404 420734 564004 420818
rect 563404 420498 563586 420734
rect 563822 420498 564004 420734
rect 563404 385054 564004 420498
rect 563404 384818 563586 385054
rect 563822 384818 564004 385054
rect 563404 384734 564004 384818
rect 563404 384498 563586 384734
rect 563822 384498 564004 384734
rect 563404 349054 564004 384498
rect 563404 348818 563586 349054
rect 563822 348818 564004 349054
rect 563404 348734 564004 348818
rect 563404 348498 563586 348734
rect 563822 348498 564004 348734
rect 563404 313054 564004 348498
rect 563404 312818 563586 313054
rect 563822 312818 564004 313054
rect 563404 312734 564004 312818
rect 563404 312498 563586 312734
rect 563822 312498 564004 312734
rect 563404 277054 564004 312498
rect 563404 276818 563586 277054
rect 563822 276818 564004 277054
rect 563404 276734 564004 276818
rect 563404 276498 563586 276734
rect 563822 276498 564004 276734
rect 563404 241054 564004 276498
rect 563404 240818 563586 241054
rect 563822 240818 564004 241054
rect 563404 240734 564004 240818
rect 563404 240498 563586 240734
rect 563822 240498 564004 240734
rect 563404 205054 564004 240498
rect 563404 204818 563586 205054
rect 563822 204818 564004 205054
rect 563404 204734 564004 204818
rect 563404 204498 563586 204734
rect 563822 204498 564004 204734
rect 563404 169054 564004 204498
rect 563404 168818 563586 169054
rect 563822 168818 564004 169054
rect 563404 168734 564004 168818
rect 563404 168498 563586 168734
rect 563822 168498 564004 168734
rect 563404 133054 564004 168498
rect 563404 132818 563586 133054
rect 563822 132818 564004 133054
rect 563404 132734 564004 132818
rect 563404 132498 563586 132734
rect 563822 132498 564004 132734
rect 563404 97054 564004 132498
rect 563404 96818 563586 97054
rect 563822 96818 564004 97054
rect 563404 96734 564004 96818
rect 563404 96498 563586 96734
rect 563822 96498 564004 96734
rect 563404 61054 564004 96498
rect 563404 60818 563586 61054
rect 563822 60818 564004 61054
rect 563404 60734 564004 60818
rect 563404 60498 563586 60734
rect 563822 60498 564004 60734
rect 563404 25054 564004 60498
rect 563404 24818 563586 25054
rect 563822 24818 564004 25054
rect 563404 24734 564004 24818
rect 563404 24498 563586 24734
rect 563822 24498 564004 24734
rect 563404 -3166 564004 24498
rect 563404 -3402 563586 -3166
rect 563822 -3402 564004 -3166
rect 563404 -3486 564004 -3402
rect 563404 -3722 563586 -3486
rect 563822 -3722 564004 -3486
rect 563404 -3744 564004 -3722
rect 567004 676654 567604 708982
rect 567004 676418 567186 676654
rect 567422 676418 567604 676654
rect 567004 676334 567604 676418
rect 567004 676098 567186 676334
rect 567422 676098 567604 676334
rect 567004 640654 567604 676098
rect 567004 640418 567186 640654
rect 567422 640418 567604 640654
rect 567004 640334 567604 640418
rect 567004 640098 567186 640334
rect 567422 640098 567604 640334
rect 567004 604654 567604 640098
rect 567004 604418 567186 604654
rect 567422 604418 567604 604654
rect 567004 604334 567604 604418
rect 567004 604098 567186 604334
rect 567422 604098 567604 604334
rect 567004 568654 567604 604098
rect 567004 568418 567186 568654
rect 567422 568418 567604 568654
rect 567004 568334 567604 568418
rect 567004 568098 567186 568334
rect 567422 568098 567604 568334
rect 567004 532654 567604 568098
rect 567004 532418 567186 532654
rect 567422 532418 567604 532654
rect 567004 532334 567604 532418
rect 567004 532098 567186 532334
rect 567422 532098 567604 532334
rect 567004 496654 567604 532098
rect 567004 496418 567186 496654
rect 567422 496418 567604 496654
rect 567004 496334 567604 496418
rect 567004 496098 567186 496334
rect 567422 496098 567604 496334
rect 567004 460654 567604 496098
rect 567004 460418 567186 460654
rect 567422 460418 567604 460654
rect 567004 460334 567604 460418
rect 567004 460098 567186 460334
rect 567422 460098 567604 460334
rect 567004 424654 567604 460098
rect 567004 424418 567186 424654
rect 567422 424418 567604 424654
rect 567004 424334 567604 424418
rect 567004 424098 567186 424334
rect 567422 424098 567604 424334
rect 567004 388654 567604 424098
rect 567004 388418 567186 388654
rect 567422 388418 567604 388654
rect 567004 388334 567604 388418
rect 567004 388098 567186 388334
rect 567422 388098 567604 388334
rect 567004 352654 567604 388098
rect 567004 352418 567186 352654
rect 567422 352418 567604 352654
rect 567004 352334 567604 352418
rect 567004 352098 567186 352334
rect 567422 352098 567604 352334
rect 567004 316654 567604 352098
rect 567004 316418 567186 316654
rect 567422 316418 567604 316654
rect 567004 316334 567604 316418
rect 567004 316098 567186 316334
rect 567422 316098 567604 316334
rect 567004 280654 567604 316098
rect 567004 280418 567186 280654
rect 567422 280418 567604 280654
rect 567004 280334 567604 280418
rect 567004 280098 567186 280334
rect 567422 280098 567604 280334
rect 567004 244654 567604 280098
rect 567004 244418 567186 244654
rect 567422 244418 567604 244654
rect 567004 244334 567604 244418
rect 567004 244098 567186 244334
rect 567422 244098 567604 244334
rect 567004 208654 567604 244098
rect 567004 208418 567186 208654
rect 567422 208418 567604 208654
rect 567004 208334 567604 208418
rect 567004 208098 567186 208334
rect 567422 208098 567604 208334
rect 567004 172654 567604 208098
rect 567004 172418 567186 172654
rect 567422 172418 567604 172654
rect 567004 172334 567604 172418
rect 567004 172098 567186 172334
rect 567422 172098 567604 172334
rect 567004 136654 567604 172098
rect 567004 136418 567186 136654
rect 567422 136418 567604 136654
rect 567004 136334 567604 136418
rect 567004 136098 567186 136334
rect 567422 136098 567604 136334
rect 567004 100654 567604 136098
rect 567004 100418 567186 100654
rect 567422 100418 567604 100654
rect 567004 100334 567604 100418
rect 567004 100098 567186 100334
rect 567422 100098 567604 100334
rect 567004 64654 567604 100098
rect 567004 64418 567186 64654
rect 567422 64418 567604 64654
rect 567004 64334 567604 64418
rect 567004 64098 567186 64334
rect 567422 64098 567604 64334
rect 567004 28654 567604 64098
rect 567004 28418 567186 28654
rect 567422 28418 567604 28654
rect 567004 28334 567604 28418
rect 567004 28098 567186 28334
rect 567422 28098 567604 28334
rect 567004 -5046 567604 28098
rect 567004 -5282 567186 -5046
rect 567422 -5282 567604 -5046
rect 567004 -5366 567604 -5282
rect 567004 -5602 567186 -5366
rect 567422 -5602 567604 -5366
rect 567004 -5624 567604 -5602
rect 570604 680254 571204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 581404 706718 582004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 581404 706482 581586 706718
rect 581822 706482 582004 706718
rect 581404 706398 582004 706482
rect 581404 706162 581586 706398
rect 581822 706162 582004 706398
rect 570604 680018 570786 680254
rect 571022 680018 571204 680254
rect 570604 679934 571204 680018
rect 570604 679698 570786 679934
rect 571022 679698 571204 679934
rect 570604 644254 571204 679698
rect 570604 644018 570786 644254
rect 571022 644018 571204 644254
rect 570604 643934 571204 644018
rect 570604 643698 570786 643934
rect 571022 643698 571204 643934
rect 570604 608254 571204 643698
rect 570604 608018 570786 608254
rect 571022 608018 571204 608254
rect 570604 607934 571204 608018
rect 570604 607698 570786 607934
rect 571022 607698 571204 607934
rect 570604 572254 571204 607698
rect 570604 572018 570786 572254
rect 571022 572018 571204 572254
rect 570604 571934 571204 572018
rect 570604 571698 570786 571934
rect 571022 571698 571204 571934
rect 570604 536254 571204 571698
rect 570604 536018 570786 536254
rect 571022 536018 571204 536254
rect 570604 535934 571204 536018
rect 570604 535698 570786 535934
rect 571022 535698 571204 535934
rect 570604 500254 571204 535698
rect 570604 500018 570786 500254
rect 571022 500018 571204 500254
rect 570604 499934 571204 500018
rect 570604 499698 570786 499934
rect 571022 499698 571204 499934
rect 570604 464254 571204 499698
rect 570604 464018 570786 464254
rect 571022 464018 571204 464254
rect 570604 463934 571204 464018
rect 570604 463698 570786 463934
rect 571022 463698 571204 463934
rect 570604 428254 571204 463698
rect 570604 428018 570786 428254
rect 571022 428018 571204 428254
rect 570604 427934 571204 428018
rect 570604 427698 570786 427934
rect 571022 427698 571204 427934
rect 570604 392254 571204 427698
rect 570604 392018 570786 392254
rect 571022 392018 571204 392254
rect 570604 391934 571204 392018
rect 570604 391698 570786 391934
rect 571022 391698 571204 391934
rect 570604 356254 571204 391698
rect 570604 356018 570786 356254
rect 571022 356018 571204 356254
rect 570604 355934 571204 356018
rect 570604 355698 570786 355934
rect 571022 355698 571204 355934
rect 570604 320254 571204 355698
rect 570604 320018 570786 320254
rect 571022 320018 571204 320254
rect 570604 319934 571204 320018
rect 570604 319698 570786 319934
rect 571022 319698 571204 319934
rect 570604 284254 571204 319698
rect 570604 284018 570786 284254
rect 571022 284018 571204 284254
rect 570604 283934 571204 284018
rect 570604 283698 570786 283934
rect 571022 283698 571204 283934
rect 570604 248254 571204 283698
rect 570604 248018 570786 248254
rect 571022 248018 571204 248254
rect 570604 247934 571204 248018
rect 570604 247698 570786 247934
rect 571022 247698 571204 247934
rect 570604 212254 571204 247698
rect 570604 212018 570786 212254
rect 571022 212018 571204 212254
rect 570604 211934 571204 212018
rect 570604 211698 570786 211934
rect 571022 211698 571204 211934
rect 570604 176254 571204 211698
rect 570604 176018 570786 176254
rect 571022 176018 571204 176254
rect 570604 175934 571204 176018
rect 570604 175698 570786 175934
rect 571022 175698 571204 175934
rect 570604 140254 571204 175698
rect 570604 140018 570786 140254
rect 571022 140018 571204 140254
rect 570604 139934 571204 140018
rect 570604 139698 570786 139934
rect 571022 139698 571204 139934
rect 570604 104254 571204 139698
rect 570604 104018 570786 104254
rect 571022 104018 571204 104254
rect 570604 103934 571204 104018
rect 570604 103698 570786 103934
rect 571022 103698 571204 103934
rect 570604 68254 571204 103698
rect 570604 68018 570786 68254
rect 571022 68018 571204 68254
rect 570604 67934 571204 68018
rect 570604 67698 570786 67934
rect 571022 67698 571204 67934
rect 570604 32254 571204 67698
rect 570604 32018 570786 32254
rect 571022 32018 571204 32254
rect 570604 31934 571204 32018
rect 570604 31698 570786 31934
rect 571022 31698 571204 31934
rect 552604 -6222 552786 -5986
rect 553022 -6222 553204 -5986
rect 552604 -6306 553204 -6222
rect 552604 -6542 552786 -6306
rect 553022 -6542 553204 -6306
rect 552604 -7504 553204 -6542
rect 570604 -6926 571204 31698
rect 577804 704838 578404 705800
rect 577804 704602 577986 704838
rect 578222 704602 578404 704838
rect 577804 704518 578404 704602
rect 577804 704282 577986 704518
rect 578222 704282 578404 704518
rect 577804 687454 578404 704282
rect 577804 687218 577986 687454
rect 578222 687218 578404 687454
rect 577804 687134 578404 687218
rect 577804 686898 577986 687134
rect 578222 686898 578404 687134
rect 577804 651454 578404 686898
rect 577804 651218 577986 651454
rect 578222 651218 578404 651454
rect 577804 651134 578404 651218
rect 577804 650898 577986 651134
rect 578222 650898 578404 651134
rect 577804 615454 578404 650898
rect 577804 615218 577986 615454
rect 578222 615218 578404 615454
rect 577804 615134 578404 615218
rect 577804 614898 577986 615134
rect 578222 614898 578404 615134
rect 577804 579454 578404 614898
rect 577804 579218 577986 579454
rect 578222 579218 578404 579454
rect 577804 579134 578404 579218
rect 577804 578898 577986 579134
rect 578222 578898 578404 579134
rect 577804 543454 578404 578898
rect 577804 543218 577986 543454
rect 578222 543218 578404 543454
rect 577804 543134 578404 543218
rect 577804 542898 577986 543134
rect 578222 542898 578404 543134
rect 577804 507454 578404 542898
rect 577804 507218 577986 507454
rect 578222 507218 578404 507454
rect 577804 507134 578404 507218
rect 577804 506898 577986 507134
rect 578222 506898 578404 507134
rect 577804 471454 578404 506898
rect 577804 471218 577986 471454
rect 578222 471218 578404 471454
rect 577804 471134 578404 471218
rect 577804 470898 577986 471134
rect 578222 470898 578404 471134
rect 577804 435454 578404 470898
rect 577804 435218 577986 435454
rect 578222 435218 578404 435454
rect 577804 435134 578404 435218
rect 577804 434898 577986 435134
rect 578222 434898 578404 435134
rect 577804 399454 578404 434898
rect 577804 399218 577986 399454
rect 578222 399218 578404 399454
rect 577804 399134 578404 399218
rect 577804 398898 577986 399134
rect 578222 398898 578404 399134
rect 577804 363454 578404 398898
rect 577804 363218 577986 363454
rect 578222 363218 578404 363454
rect 577804 363134 578404 363218
rect 577804 362898 577986 363134
rect 578222 362898 578404 363134
rect 577804 327454 578404 362898
rect 577804 327218 577986 327454
rect 578222 327218 578404 327454
rect 577804 327134 578404 327218
rect 577804 326898 577986 327134
rect 578222 326898 578404 327134
rect 577804 291454 578404 326898
rect 577804 291218 577986 291454
rect 578222 291218 578404 291454
rect 577804 291134 578404 291218
rect 577804 290898 577986 291134
rect 578222 290898 578404 291134
rect 577804 255454 578404 290898
rect 577804 255218 577986 255454
rect 578222 255218 578404 255454
rect 577804 255134 578404 255218
rect 577804 254898 577986 255134
rect 578222 254898 578404 255134
rect 577804 219454 578404 254898
rect 577804 219218 577986 219454
rect 578222 219218 578404 219454
rect 577804 219134 578404 219218
rect 577804 218898 577986 219134
rect 578222 218898 578404 219134
rect 577804 183454 578404 218898
rect 577804 183218 577986 183454
rect 578222 183218 578404 183454
rect 577804 183134 578404 183218
rect 577804 182898 577986 183134
rect 578222 182898 578404 183134
rect 577804 147454 578404 182898
rect 577804 147218 577986 147454
rect 578222 147218 578404 147454
rect 577804 147134 578404 147218
rect 577804 146898 577986 147134
rect 578222 146898 578404 147134
rect 577804 111454 578404 146898
rect 577804 111218 577986 111454
rect 578222 111218 578404 111454
rect 577804 111134 578404 111218
rect 577804 110898 577986 111134
rect 578222 110898 578404 111134
rect 577804 75454 578404 110898
rect 577804 75218 577986 75454
rect 578222 75218 578404 75454
rect 577804 75134 578404 75218
rect 577804 74898 577986 75134
rect 578222 74898 578404 75134
rect 577804 39454 578404 74898
rect 577804 39218 577986 39454
rect 578222 39218 578404 39454
rect 577804 39134 578404 39218
rect 577804 38898 577986 39134
rect 578222 38898 578404 39134
rect 577804 3454 578404 38898
rect 577804 3218 577986 3454
rect 578222 3218 578404 3454
rect 577804 3134 578404 3218
rect 577804 2898 577986 3134
rect 578222 2898 578404 3134
rect 577804 -346 578404 2898
rect 577804 -582 577986 -346
rect 578222 -582 578404 -346
rect 577804 -666 578404 -582
rect 577804 -902 577986 -666
rect 578222 -902 578404 -666
rect 577804 -1864 578404 -902
rect 581404 691054 582004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 581404 690818 581586 691054
rect 581822 690818 582004 691054
rect 581404 690734 582004 690818
rect 581404 690498 581586 690734
rect 581822 690498 582004 690734
rect 581404 655054 582004 690498
rect 581404 654818 581586 655054
rect 581822 654818 582004 655054
rect 581404 654734 582004 654818
rect 581404 654498 581586 654734
rect 581822 654498 582004 654734
rect 581404 619054 582004 654498
rect 581404 618818 581586 619054
rect 581822 618818 582004 619054
rect 581404 618734 582004 618818
rect 581404 618498 581586 618734
rect 581822 618498 582004 618734
rect 581404 583054 582004 618498
rect 581404 582818 581586 583054
rect 581822 582818 582004 583054
rect 581404 582734 582004 582818
rect 581404 582498 581586 582734
rect 581822 582498 582004 582734
rect 581404 547054 582004 582498
rect 581404 546818 581586 547054
rect 581822 546818 582004 547054
rect 581404 546734 582004 546818
rect 581404 546498 581586 546734
rect 581822 546498 582004 546734
rect 581404 511054 582004 546498
rect 581404 510818 581586 511054
rect 581822 510818 582004 511054
rect 581404 510734 582004 510818
rect 581404 510498 581586 510734
rect 581822 510498 582004 510734
rect 581404 475054 582004 510498
rect 581404 474818 581586 475054
rect 581822 474818 582004 475054
rect 581404 474734 582004 474818
rect 581404 474498 581586 474734
rect 581822 474498 582004 474734
rect 581404 439054 582004 474498
rect 581404 438818 581586 439054
rect 581822 438818 582004 439054
rect 581404 438734 582004 438818
rect 581404 438498 581586 438734
rect 581822 438498 582004 438734
rect 581404 403054 582004 438498
rect 581404 402818 581586 403054
rect 581822 402818 582004 403054
rect 581404 402734 582004 402818
rect 581404 402498 581586 402734
rect 581822 402498 582004 402734
rect 581404 367054 582004 402498
rect 581404 366818 581586 367054
rect 581822 366818 582004 367054
rect 581404 366734 582004 366818
rect 581404 366498 581586 366734
rect 581822 366498 582004 366734
rect 581404 331054 582004 366498
rect 581404 330818 581586 331054
rect 581822 330818 582004 331054
rect 581404 330734 582004 330818
rect 581404 330498 581586 330734
rect 581822 330498 582004 330734
rect 581404 295054 582004 330498
rect 581404 294818 581586 295054
rect 581822 294818 582004 295054
rect 581404 294734 582004 294818
rect 581404 294498 581586 294734
rect 581822 294498 582004 294734
rect 581404 259054 582004 294498
rect 581404 258818 581586 259054
rect 581822 258818 582004 259054
rect 581404 258734 582004 258818
rect 581404 258498 581586 258734
rect 581822 258498 582004 258734
rect 581404 223054 582004 258498
rect 581404 222818 581586 223054
rect 581822 222818 582004 223054
rect 581404 222734 582004 222818
rect 581404 222498 581586 222734
rect 581822 222498 582004 222734
rect 581404 187054 582004 222498
rect 581404 186818 581586 187054
rect 581822 186818 582004 187054
rect 581404 186734 582004 186818
rect 581404 186498 581586 186734
rect 581822 186498 582004 186734
rect 581404 151054 582004 186498
rect 581404 150818 581586 151054
rect 581822 150818 582004 151054
rect 581404 150734 582004 150818
rect 581404 150498 581586 150734
rect 581822 150498 582004 150734
rect 581404 115054 582004 150498
rect 581404 114818 581586 115054
rect 581822 114818 582004 115054
rect 581404 114734 582004 114818
rect 581404 114498 581586 114734
rect 581822 114498 582004 114734
rect 581404 79054 582004 114498
rect 581404 78818 581586 79054
rect 581822 78818 582004 79054
rect 581404 78734 582004 78818
rect 581404 78498 581586 78734
rect 581822 78498 582004 78734
rect 581404 43054 582004 78498
rect 581404 42818 581586 43054
rect 581822 42818 582004 43054
rect 581404 42734 582004 42818
rect 581404 42498 581586 42734
rect 581822 42498 582004 42734
rect 581404 7054 582004 42498
rect 581404 6818 581586 7054
rect 581822 6818 582004 7054
rect 581404 6734 582004 6818
rect 581404 6498 581586 6734
rect 581822 6498 582004 6734
rect 581404 -2226 582004 6498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 687454 585920 704282
rect 585320 687218 585502 687454
rect 585738 687218 585920 687454
rect 585320 687134 585920 687218
rect 585320 686898 585502 687134
rect 585738 686898 585920 687134
rect 585320 651454 585920 686898
rect 585320 651218 585502 651454
rect 585738 651218 585920 651454
rect 585320 651134 585920 651218
rect 585320 650898 585502 651134
rect 585738 650898 585920 651134
rect 585320 615454 585920 650898
rect 585320 615218 585502 615454
rect 585738 615218 585920 615454
rect 585320 615134 585920 615218
rect 585320 614898 585502 615134
rect 585738 614898 585920 615134
rect 585320 579454 585920 614898
rect 585320 579218 585502 579454
rect 585738 579218 585920 579454
rect 585320 579134 585920 579218
rect 585320 578898 585502 579134
rect 585738 578898 585920 579134
rect 585320 543454 585920 578898
rect 585320 543218 585502 543454
rect 585738 543218 585920 543454
rect 585320 543134 585920 543218
rect 585320 542898 585502 543134
rect 585738 542898 585920 543134
rect 585320 507454 585920 542898
rect 585320 507218 585502 507454
rect 585738 507218 585920 507454
rect 585320 507134 585920 507218
rect 585320 506898 585502 507134
rect 585738 506898 585920 507134
rect 585320 471454 585920 506898
rect 585320 471218 585502 471454
rect 585738 471218 585920 471454
rect 585320 471134 585920 471218
rect 585320 470898 585502 471134
rect 585738 470898 585920 471134
rect 585320 435454 585920 470898
rect 585320 435218 585502 435454
rect 585738 435218 585920 435454
rect 585320 435134 585920 435218
rect 585320 434898 585502 435134
rect 585738 434898 585920 435134
rect 585320 399454 585920 434898
rect 585320 399218 585502 399454
rect 585738 399218 585920 399454
rect 585320 399134 585920 399218
rect 585320 398898 585502 399134
rect 585738 398898 585920 399134
rect 585320 363454 585920 398898
rect 585320 363218 585502 363454
rect 585738 363218 585920 363454
rect 585320 363134 585920 363218
rect 585320 362898 585502 363134
rect 585738 362898 585920 363134
rect 585320 327454 585920 362898
rect 585320 327218 585502 327454
rect 585738 327218 585920 327454
rect 585320 327134 585920 327218
rect 585320 326898 585502 327134
rect 585738 326898 585920 327134
rect 585320 291454 585920 326898
rect 585320 291218 585502 291454
rect 585738 291218 585920 291454
rect 585320 291134 585920 291218
rect 585320 290898 585502 291134
rect 585738 290898 585920 291134
rect 585320 255454 585920 290898
rect 585320 255218 585502 255454
rect 585738 255218 585920 255454
rect 585320 255134 585920 255218
rect 585320 254898 585502 255134
rect 585738 254898 585920 255134
rect 585320 219454 585920 254898
rect 585320 219218 585502 219454
rect 585738 219218 585920 219454
rect 585320 219134 585920 219218
rect 585320 218898 585502 219134
rect 585738 218898 585920 219134
rect 585320 183454 585920 218898
rect 585320 183218 585502 183454
rect 585738 183218 585920 183454
rect 585320 183134 585920 183218
rect 585320 182898 585502 183134
rect 585738 182898 585920 183134
rect 585320 147454 585920 182898
rect 585320 147218 585502 147454
rect 585738 147218 585920 147454
rect 585320 147134 585920 147218
rect 585320 146898 585502 147134
rect 585738 146898 585920 147134
rect 585320 111454 585920 146898
rect 585320 111218 585502 111454
rect 585738 111218 585920 111454
rect 585320 111134 585920 111218
rect 585320 110898 585502 111134
rect 585738 110898 585920 111134
rect 585320 75454 585920 110898
rect 585320 75218 585502 75454
rect 585738 75218 585920 75454
rect 585320 75134 585920 75218
rect 585320 74898 585502 75134
rect 585738 74898 585920 75134
rect 585320 39454 585920 74898
rect 585320 39218 585502 39454
rect 585738 39218 585920 39454
rect 585320 39134 585920 39218
rect 585320 38898 585502 39134
rect 585738 38898 585920 39134
rect 585320 3454 585920 38898
rect 585320 3218 585502 3454
rect 585738 3218 585920 3454
rect 585320 3134 585920 3218
rect 585320 2898 585502 3134
rect 585738 2898 585920 3134
rect 585320 -346 585920 2898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 669454 586860 705222
rect 586260 669218 586442 669454
rect 586678 669218 586860 669454
rect 586260 669134 586860 669218
rect 586260 668898 586442 669134
rect 586678 668898 586860 669134
rect 586260 633454 586860 668898
rect 586260 633218 586442 633454
rect 586678 633218 586860 633454
rect 586260 633134 586860 633218
rect 586260 632898 586442 633134
rect 586678 632898 586860 633134
rect 586260 597454 586860 632898
rect 586260 597218 586442 597454
rect 586678 597218 586860 597454
rect 586260 597134 586860 597218
rect 586260 596898 586442 597134
rect 586678 596898 586860 597134
rect 586260 561454 586860 596898
rect 586260 561218 586442 561454
rect 586678 561218 586860 561454
rect 586260 561134 586860 561218
rect 586260 560898 586442 561134
rect 586678 560898 586860 561134
rect 586260 525454 586860 560898
rect 586260 525218 586442 525454
rect 586678 525218 586860 525454
rect 586260 525134 586860 525218
rect 586260 524898 586442 525134
rect 586678 524898 586860 525134
rect 586260 489454 586860 524898
rect 586260 489218 586442 489454
rect 586678 489218 586860 489454
rect 586260 489134 586860 489218
rect 586260 488898 586442 489134
rect 586678 488898 586860 489134
rect 586260 453454 586860 488898
rect 586260 453218 586442 453454
rect 586678 453218 586860 453454
rect 586260 453134 586860 453218
rect 586260 452898 586442 453134
rect 586678 452898 586860 453134
rect 586260 417454 586860 452898
rect 586260 417218 586442 417454
rect 586678 417218 586860 417454
rect 586260 417134 586860 417218
rect 586260 416898 586442 417134
rect 586678 416898 586860 417134
rect 586260 381454 586860 416898
rect 586260 381218 586442 381454
rect 586678 381218 586860 381454
rect 586260 381134 586860 381218
rect 586260 380898 586442 381134
rect 586678 380898 586860 381134
rect 586260 345454 586860 380898
rect 586260 345218 586442 345454
rect 586678 345218 586860 345454
rect 586260 345134 586860 345218
rect 586260 344898 586442 345134
rect 586678 344898 586860 345134
rect 586260 309454 586860 344898
rect 586260 309218 586442 309454
rect 586678 309218 586860 309454
rect 586260 309134 586860 309218
rect 586260 308898 586442 309134
rect 586678 308898 586860 309134
rect 586260 273454 586860 308898
rect 586260 273218 586442 273454
rect 586678 273218 586860 273454
rect 586260 273134 586860 273218
rect 586260 272898 586442 273134
rect 586678 272898 586860 273134
rect 586260 237454 586860 272898
rect 586260 237218 586442 237454
rect 586678 237218 586860 237454
rect 586260 237134 586860 237218
rect 586260 236898 586442 237134
rect 586678 236898 586860 237134
rect 586260 201454 586860 236898
rect 586260 201218 586442 201454
rect 586678 201218 586860 201454
rect 586260 201134 586860 201218
rect 586260 200898 586442 201134
rect 586678 200898 586860 201134
rect 586260 165454 586860 200898
rect 586260 165218 586442 165454
rect 586678 165218 586860 165454
rect 586260 165134 586860 165218
rect 586260 164898 586442 165134
rect 586678 164898 586860 165134
rect 586260 129454 586860 164898
rect 586260 129218 586442 129454
rect 586678 129218 586860 129454
rect 586260 129134 586860 129218
rect 586260 128898 586442 129134
rect 586678 128898 586860 129134
rect 586260 93454 586860 128898
rect 586260 93218 586442 93454
rect 586678 93218 586860 93454
rect 586260 93134 586860 93218
rect 586260 92898 586442 93134
rect 586678 92898 586860 93134
rect 586260 57454 586860 92898
rect 586260 57218 586442 57454
rect 586678 57218 586860 57454
rect 586260 57134 586860 57218
rect 586260 56898 586442 57134
rect 586678 56898 586860 57134
rect 586260 21454 586860 56898
rect 586260 21218 586442 21454
rect 586678 21218 586860 21454
rect 586260 21134 586860 21218
rect 586260 20898 586442 21134
rect 586678 20898 586860 21134
rect 586260 -1286 586860 20898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 691054 587800 706162
rect 587200 690818 587382 691054
rect 587618 690818 587800 691054
rect 587200 690734 587800 690818
rect 587200 690498 587382 690734
rect 587618 690498 587800 690734
rect 587200 655054 587800 690498
rect 587200 654818 587382 655054
rect 587618 654818 587800 655054
rect 587200 654734 587800 654818
rect 587200 654498 587382 654734
rect 587618 654498 587800 654734
rect 587200 619054 587800 654498
rect 587200 618818 587382 619054
rect 587618 618818 587800 619054
rect 587200 618734 587800 618818
rect 587200 618498 587382 618734
rect 587618 618498 587800 618734
rect 587200 583054 587800 618498
rect 587200 582818 587382 583054
rect 587618 582818 587800 583054
rect 587200 582734 587800 582818
rect 587200 582498 587382 582734
rect 587618 582498 587800 582734
rect 587200 547054 587800 582498
rect 587200 546818 587382 547054
rect 587618 546818 587800 547054
rect 587200 546734 587800 546818
rect 587200 546498 587382 546734
rect 587618 546498 587800 546734
rect 587200 511054 587800 546498
rect 587200 510818 587382 511054
rect 587618 510818 587800 511054
rect 587200 510734 587800 510818
rect 587200 510498 587382 510734
rect 587618 510498 587800 510734
rect 587200 475054 587800 510498
rect 587200 474818 587382 475054
rect 587618 474818 587800 475054
rect 587200 474734 587800 474818
rect 587200 474498 587382 474734
rect 587618 474498 587800 474734
rect 587200 439054 587800 474498
rect 587200 438818 587382 439054
rect 587618 438818 587800 439054
rect 587200 438734 587800 438818
rect 587200 438498 587382 438734
rect 587618 438498 587800 438734
rect 587200 403054 587800 438498
rect 587200 402818 587382 403054
rect 587618 402818 587800 403054
rect 587200 402734 587800 402818
rect 587200 402498 587382 402734
rect 587618 402498 587800 402734
rect 587200 367054 587800 402498
rect 587200 366818 587382 367054
rect 587618 366818 587800 367054
rect 587200 366734 587800 366818
rect 587200 366498 587382 366734
rect 587618 366498 587800 366734
rect 587200 331054 587800 366498
rect 587200 330818 587382 331054
rect 587618 330818 587800 331054
rect 587200 330734 587800 330818
rect 587200 330498 587382 330734
rect 587618 330498 587800 330734
rect 587200 295054 587800 330498
rect 587200 294818 587382 295054
rect 587618 294818 587800 295054
rect 587200 294734 587800 294818
rect 587200 294498 587382 294734
rect 587618 294498 587800 294734
rect 587200 259054 587800 294498
rect 587200 258818 587382 259054
rect 587618 258818 587800 259054
rect 587200 258734 587800 258818
rect 587200 258498 587382 258734
rect 587618 258498 587800 258734
rect 587200 223054 587800 258498
rect 587200 222818 587382 223054
rect 587618 222818 587800 223054
rect 587200 222734 587800 222818
rect 587200 222498 587382 222734
rect 587618 222498 587800 222734
rect 587200 187054 587800 222498
rect 587200 186818 587382 187054
rect 587618 186818 587800 187054
rect 587200 186734 587800 186818
rect 587200 186498 587382 186734
rect 587618 186498 587800 186734
rect 587200 151054 587800 186498
rect 587200 150818 587382 151054
rect 587618 150818 587800 151054
rect 587200 150734 587800 150818
rect 587200 150498 587382 150734
rect 587618 150498 587800 150734
rect 587200 115054 587800 150498
rect 587200 114818 587382 115054
rect 587618 114818 587800 115054
rect 587200 114734 587800 114818
rect 587200 114498 587382 114734
rect 587618 114498 587800 114734
rect 587200 79054 587800 114498
rect 587200 78818 587382 79054
rect 587618 78818 587800 79054
rect 587200 78734 587800 78818
rect 587200 78498 587382 78734
rect 587618 78498 587800 78734
rect 587200 43054 587800 78498
rect 587200 42818 587382 43054
rect 587618 42818 587800 43054
rect 587200 42734 587800 42818
rect 587200 42498 587382 42734
rect 587618 42498 587800 42734
rect 587200 7054 587800 42498
rect 587200 6818 587382 7054
rect 587618 6818 587800 7054
rect 587200 6734 587800 6818
rect 587200 6498 587382 6734
rect 587618 6498 587800 6734
rect 581404 -2462 581586 -2226
rect 581822 -2462 582004 -2226
rect 581404 -2546 582004 -2462
rect 581404 -2782 581586 -2546
rect 581822 -2782 582004 -2546
rect 581404 -3744 582004 -2782
rect 587200 -2226 587800 6498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 673054 588740 707102
rect 588140 672818 588322 673054
rect 588558 672818 588740 673054
rect 588140 672734 588740 672818
rect 588140 672498 588322 672734
rect 588558 672498 588740 672734
rect 588140 637054 588740 672498
rect 588140 636818 588322 637054
rect 588558 636818 588740 637054
rect 588140 636734 588740 636818
rect 588140 636498 588322 636734
rect 588558 636498 588740 636734
rect 588140 601054 588740 636498
rect 588140 600818 588322 601054
rect 588558 600818 588740 601054
rect 588140 600734 588740 600818
rect 588140 600498 588322 600734
rect 588558 600498 588740 600734
rect 588140 565054 588740 600498
rect 588140 564818 588322 565054
rect 588558 564818 588740 565054
rect 588140 564734 588740 564818
rect 588140 564498 588322 564734
rect 588558 564498 588740 564734
rect 588140 529054 588740 564498
rect 588140 528818 588322 529054
rect 588558 528818 588740 529054
rect 588140 528734 588740 528818
rect 588140 528498 588322 528734
rect 588558 528498 588740 528734
rect 588140 493054 588740 528498
rect 588140 492818 588322 493054
rect 588558 492818 588740 493054
rect 588140 492734 588740 492818
rect 588140 492498 588322 492734
rect 588558 492498 588740 492734
rect 588140 457054 588740 492498
rect 588140 456818 588322 457054
rect 588558 456818 588740 457054
rect 588140 456734 588740 456818
rect 588140 456498 588322 456734
rect 588558 456498 588740 456734
rect 588140 421054 588740 456498
rect 588140 420818 588322 421054
rect 588558 420818 588740 421054
rect 588140 420734 588740 420818
rect 588140 420498 588322 420734
rect 588558 420498 588740 420734
rect 588140 385054 588740 420498
rect 588140 384818 588322 385054
rect 588558 384818 588740 385054
rect 588140 384734 588740 384818
rect 588140 384498 588322 384734
rect 588558 384498 588740 384734
rect 588140 349054 588740 384498
rect 588140 348818 588322 349054
rect 588558 348818 588740 349054
rect 588140 348734 588740 348818
rect 588140 348498 588322 348734
rect 588558 348498 588740 348734
rect 588140 313054 588740 348498
rect 588140 312818 588322 313054
rect 588558 312818 588740 313054
rect 588140 312734 588740 312818
rect 588140 312498 588322 312734
rect 588558 312498 588740 312734
rect 588140 277054 588740 312498
rect 588140 276818 588322 277054
rect 588558 276818 588740 277054
rect 588140 276734 588740 276818
rect 588140 276498 588322 276734
rect 588558 276498 588740 276734
rect 588140 241054 588740 276498
rect 588140 240818 588322 241054
rect 588558 240818 588740 241054
rect 588140 240734 588740 240818
rect 588140 240498 588322 240734
rect 588558 240498 588740 240734
rect 588140 205054 588740 240498
rect 588140 204818 588322 205054
rect 588558 204818 588740 205054
rect 588140 204734 588740 204818
rect 588140 204498 588322 204734
rect 588558 204498 588740 204734
rect 588140 169054 588740 204498
rect 588140 168818 588322 169054
rect 588558 168818 588740 169054
rect 588140 168734 588740 168818
rect 588140 168498 588322 168734
rect 588558 168498 588740 168734
rect 588140 133054 588740 168498
rect 588140 132818 588322 133054
rect 588558 132818 588740 133054
rect 588140 132734 588740 132818
rect 588140 132498 588322 132734
rect 588558 132498 588740 132734
rect 588140 97054 588740 132498
rect 588140 96818 588322 97054
rect 588558 96818 588740 97054
rect 588140 96734 588740 96818
rect 588140 96498 588322 96734
rect 588558 96498 588740 96734
rect 588140 61054 588740 96498
rect 588140 60818 588322 61054
rect 588558 60818 588740 61054
rect 588140 60734 588740 60818
rect 588140 60498 588322 60734
rect 588558 60498 588740 60734
rect 588140 25054 588740 60498
rect 588140 24818 588322 25054
rect 588558 24818 588740 25054
rect 588140 24734 588740 24818
rect 588140 24498 588322 24734
rect 588558 24498 588740 24734
rect 588140 -3166 588740 24498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 694654 589680 708042
rect 589080 694418 589262 694654
rect 589498 694418 589680 694654
rect 589080 694334 589680 694418
rect 589080 694098 589262 694334
rect 589498 694098 589680 694334
rect 589080 658654 589680 694098
rect 589080 658418 589262 658654
rect 589498 658418 589680 658654
rect 589080 658334 589680 658418
rect 589080 658098 589262 658334
rect 589498 658098 589680 658334
rect 589080 622654 589680 658098
rect 589080 622418 589262 622654
rect 589498 622418 589680 622654
rect 589080 622334 589680 622418
rect 589080 622098 589262 622334
rect 589498 622098 589680 622334
rect 589080 586654 589680 622098
rect 589080 586418 589262 586654
rect 589498 586418 589680 586654
rect 589080 586334 589680 586418
rect 589080 586098 589262 586334
rect 589498 586098 589680 586334
rect 589080 550654 589680 586098
rect 589080 550418 589262 550654
rect 589498 550418 589680 550654
rect 589080 550334 589680 550418
rect 589080 550098 589262 550334
rect 589498 550098 589680 550334
rect 589080 514654 589680 550098
rect 589080 514418 589262 514654
rect 589498 514418 589680 514654
rect 589080 514334 589680 514418
rect 589080 514098 589262 514334
rect 589498 514098 589680 514334
rect 589080 478654 589680 514098
rect 589080 478418 589262 478654
rect 589498 478418 589680 478654
rect 589080 478334 589680 478418
rect 589080 478098 589262 478334
rect 589498 478098 589680 478334
rect 589080 442654 589680 478098
rect 589080 442418 589262 442654
rect 589498 442418 589680 442654
rect 589080 442334 589680 442418
rect 589080 442098 589262 442334
rect 589498 442098 589680 442334
rect 589080 406654 589680 442098
rect 589080 406418 589262 406654
rect 589498 406418 589680 406654
rect 589080 406334 589680 406418
rect 589080 406098 589262 406334
rect 589498 406098 589680 406334
rect 589080 370654 589680 406098
rect 589080 370418 589262 370654
rect 589498 370418 589680 370654
rect 589080 370334 589680 370418
rect 589080 370098 589262 370334
rect 589498 370098 589680 370334
rect 589080 334654 589680 370098
rect 589080 334418 589262 334654
rect 589498 334418 589680 334654
rect 589080 334334 589680 334418
rect 589080 334098 589262 334334
rect 589498 334098 589680 334334
rect 589080 298654 589680 334098
rect 589080 298418 589262 298654
rect 589498 298418 589680 298654
rect 589080 298334 589680 298418
rect 589080 298098 589262 298334
rect 589498 298098 589680 298334
rect 589080 262654 589680 298098
rect 589080 262418 589262 262654
rect 589498 262418 589680 262654
rect 589080 262334 589680 262418
rect 589080 262098 589262 262334
rect 589498 262098 589680 262334
rect 589080 226654 589680 262098
rect 589080 226418 589262 226654
rect 589498 226418 589680 226654
rect 589080 226334 589680 226418
rect 589080 226098 589262 226334
rect 589498 226098 589680 226334
rect 589080 190654 589680 226098
rect 589080 190418 589262 190654
rect 589498 190418 589680 190654
rect 589080 190334 589680 190418
rect 589080 190098 589262 190334
rect 589498 190098 589680 190334
rect 589080 154654 589680 190098
rect 589080 154418 589262 154654
rect 589498 154418 589680 154654
rect 589080 154334 589680 154418
rect 589080 154098 589262 154334
rect 589498 154098 589680 154334
rect 589080 118654 589680 154098
rect 589080 118418 589262 118654
rect 589498 118418 589680 118654
rect 589080 118334 589680 118418
rect 589080 118098 589262 118334
rect 589498 118098 589680 118334
rect 589080 82654 589680 118098
rect 589080 82418 589262 82654
rect 589498 82418 589680 82654
rect 589080 82334 589680 82418
rect 589080 82098 589262 82334
rect 589498 82098 589680 82334
rect 589080 46654 589680 82098
rect 589080 46418 589262 46654
rect 589498 46418 589680 46654
rect 589080 46334 589680 46418
rect 589080 46098 589262 46334
rect 589498 46098 589680 46334
rect 589080 10654 589680 46098
rect 589080 10418 589262 10654
rect 589498 10418 589680 10654
rect 589080 10334 589680 10418
rect 589080 10098 589262 10334
rect 589498 10098 589680 10334
rect 589080 -4106 589680 10098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 676654 590620 708982
rect 590020 676418 590202 676654
rect 590438 676418 590620 676654
rect 590020 676334 590620 676418
rect 590020 676098 590202 676334
rect 590438 676098 590620 676334
rect 590020 640654 590620 676098
rect 590020 640418 590202 640654
rect 590438 640418 590620 640654
rect 590020 640334 590620 640418
rect 590020 640098 590202 640334
rect 590438 640098 590620 640334
rect 590020 604654 590620 640098
rect 590020 604418 590202 604654
rect 590438 604418 590620 604654
rect 590020 604334 590620 604418
rect 590020 604098 590202 604334
rect 590438 604098 590620 604334
rect 590020 568654 590620 604098
rect 590020 568418 590202 568654
rect 590438 568418 590620 568654
rect 590020 568334 590620 568418
rect 590020 568098 590202 568334
rect 590438 568098 590620 568334
rect 590020 532654 590620 568098
rect 590020 532418 590202 532654
rect 590438 532418 590620 532654
rect 590020 532334 590620 532418
rect 590020 532098 590202 532334
rect 590438 532098 590620 532334
rect 590020 496654 590620 532098
rect 590020 496418 590202 496654
rect 590438 496418 590620 496654
rect 590020 496334 590620 496418
rect 590020 496098 590202 496334
rect 590438 496098 590620 496334
rect 590020 460654 590620 496098
rect 590020 460418 590202 460654
rect 590438 460418 590620 460654
rect 590020 460334 590620 460418
rect 590020 460098 590202 460334
rect 590438 460098 590620 460334
rect 590020 424654 590620 460098
rect 590020 424418 590202 424654
rect 590438 424418 590620 424654
rect 590020 424334 590620 424418
rect 590020 424098 590202 424334
rect 590438 424098 590620 424334
rect 590020 388654 590620 424098
rect 590020 388418 590202 388654
rect 590438 388418 590620 388654
rect 590020 388334 590620 388418
rect 590020 388098 590202 388334
rect 590438 388098 590620 388334
rect 590020 352654 590620 388098
rect 590020 352418 590202 352654
rect 590438 352418 590620 352654
rect 590020 352334 590620 352418
rect 590020 352098 590202 352334
rect 590438 352098 590620 352334
rect 590020 316654 590620 352098
rect 590020 316418 590202 316654
rect 590438 316418 590620 316654
rect 590020 316334 590620 316418
rect 590020 316098 590202 316334
rect 590438 316098 590620 316334
rect 590020 280654 590620 316098
rect 590020 280418 590202 280654
rect 590438 280418 590620 280654
rect 590020 280334 590620 280418
rect 590020 280098 590202 280334
rect 590438 280098 590620 280334
rect 590020 244654 590620 280098
rect 590020 244418 590202 244654
rect 590438 244418 590620 244654
rect 590020 244334 590620 244418
rect 590020 244098 590202 244334
rect 590438 244098 590620 244334
rect 590020 208654 590620 244098
rect 590020 208418 590202 208654
rect 590438 208418 590620 208654
rect 590020 208334 590620 208418
rect 590020 208098 590202 208334
rect 590438 208098 590620 208334
rect 590020 172654 590620 208098
rect 590020 172418 590202 172654
rect 590438 172418 590620 172654
rect 590020 172334 590620 172418
rect 590020 172098 590202 172334
rect 590438 172098 590620 172334
rect 590020 136654 590620 172098
rect 590020 136418 590202 136654
rect 590438 136418 590620 136654
rect 590020 136334 590620 136418
rect 590020 136098 590202 136334
rect 590438 136098 590620 136334
rect 590020 100654 590620 136098
rect 590020 100418 590202 100654
rect 590438 100418 590620 100654
rect 590020 100334 590620 100418
rect 590020 100098 590202 100334
rect 590438 100098 590620 100334
rect 590020 64654 590620 100098
rect 590020 64418 590202 64654
rect 590438 64418 590620 64654
rect 590020 64334 590620 64418
rect 590020 64098 590202 64334
rect 590438 64098 590620 64334
rect 590020 28654 590620 64098
rect 590020 28418 590202 28654
rect 590438 28418 590620 28654
rect 590020 28334 590620 28418
rect 590020 28098 590202 28334
rect 590438 28098 590620 28334
rect 590020 -5046 590620 28098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 698254 591560 709922
rect 590960 698018 591142 698254
rect 591378 698018 591560 698254
rect 590960 697934 591560 698018
rect 590960 697698 591142 697934
rect 591378 697698 591560 697934
rect 590960 662254 591560 697698
rect 590960 662018 591142 662254
rect 591378 662018 591560 662254
rect 590960 661934 591560 662018
rect 590960 661698 591142 661934
rect 591378 661698 591560 661934
rect 590960 626254 591560 661698
rect 590960 626018 591142 626254
rect 591378 626018 591560 626254
rect 590960 625934 591560 626018
rect 590960 625698 591142 625934
rect 591378 625698 591560 625934
rect 590960 590254 591560 625698
rect 590960 590018 591142 590254
rect 591378 590018 591560 590254
rect 590960 589934 591560 590018
rect 590960 589698 591142 589934
rect 591378 589698 591560 589934
rect 590960 554254 591560 589698
rect 590960 554018 591142 554254
rect 591378 554018 591560 554254
rect 590960 553934 591560 554018
rect 590960 553698 591142 553934
rect 591378 553698 591560 553934
rect 590960 518254 591560 553698
rect 590960 518018 591142 518254
rect 591378 518018 591560 518254
rect 590960 517934 591560 518018
rect 590960 517698 591142 517934
rect 591378 517698 591560 517934
rect 590960 482254 591560 517698
rect 590960 482018 591142 482254
rect 591378 482018 591560 482254
rect 590960 481934 591560 482018
rect 590960 481698 591142 481934
rect 591378 481698 591560 481934
rect 590960 446254 591560 481698
rect 590960 446018 591142 446254
rect 591378 446018 591560 446254
rect 590960 445934 591560 446018
rect 590960 445698 591142 445934
rect 591378 445698 591560 445934
rect 590960 410254 591560 445698
rect 590960 410018 591142 410254
rect 591378 410018 591560 410254
rect 590960 409934 591560 410018
rect 590960 409698 591142 409934
rect 591378 409698 591560 409934
rect 590960 374254 591560 409698
rect 590960 374018 591142 374254
rect 591378 374018 591560 374254
rect 590960 373934 591560 374018
rect 590960 373698 591142 373934
rect 591378 373698 591560 373934
rect 590960 338254 591560 373698
rect 590960 338018 591142 338254
rect 591378 338018 591560 338254
rect 590960 337934 591560 338018
rect 590960 337698 591142 337934
rect 591378 337698 591560 337934
rect 590960 302254 591560 337698
rect 590960 302018 591142 302254
rect 591378 302018 591560 302254
rect 590960 301934 591560 302018
rect 590960 301698 591142 301934
rect 591378 301698 591560 301934
rect 590960 266254 591560 301698
rect 590960 266018 591142 266254
rect 591378 266018 591560 266254
rect 590960 265934 591560 266018
rect 590960 265698 591142 265934
rect 591378 265698 591560 265934
rect 590960 230254 591560 265698
rect 590960 230018 591142 230254
rect 591378 230018 591560 230254
rect 590960 229934 591560 230018
rect 590960 229698 591142 229934
rect 591378 229698 591560 229934
rect 590960 194254 591560 229698
rect 590960 194018 591142 194254
rect 591378 194018 591560 194254
rect 590960 193934 591560 194018
rect 590960 193698 591142 193934
rect 591378 193698 591560 193934
rect 590960 158254 591560 193698
rect 590960 158018 591142 158254
rect 591378 158018 591560 158254
rect 590960 157934 591560 158018
rect 590960 157698 591142 157934
rect 591378 157698 591560 157934
rect 590960 122254 591560 157698
rect 590960 122018 591142 122254
rect 591378 122018 591560 122254
rect 590960 121934 591560 122018
rect 590960 121698 591142 121934
rect 591378 121698 591560 121934
rect 590960 86254 591560 121698
rect 590960 86018 591142 86254
rect 591378 86018 591560 86254
rect 590960 85934 591560 86018
rect 590960 85698 591142 85934
rect 591378 85698 591560 85934
rect 590960 50254 591560 85698
rect 590960 50018 591142 50254
rect 591378 50018 591560 50254
rect 590960 49934 591560 50018
rect 590960 49698 591142 49934
rect 591378 49698 591560 49934
rect 590960 14254 591560 49698
rect 590960 14018 591142 14254
rect 591378 14018 591560 14254
rect 590960 13934 591560 14018
rect 590960 13698 591142 13934
rect 591378 13698 591560 13934
rect 590960 -5986 591560 13698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 680254 592500 710862
rect 591900 680018 592082 680254
rect 592318 680018 592500 680254
rect 591900 679934 592500 680018
rect 591900 679698 592082 679934
rect 592318 679698 592500 679934
rect 591900 644254 592500 679698
rect 591900 644018 592082 644254
rect 592318 644018 592500 644254
rect 591900 643934 592500 644018
rect 591900 643698 592082 643934
rect 592318 643698 592500 643934
rect 591900 608254 592500 643698
rect 591900 608018 592082 608254
rect 592318 608018 592500 608254
rect 591900 607934 592500 608018
rect 591900 607698 592082 607934
rect 592318 607698 592500 607934
rect 591900 572254 592500 607698
rect 591900 572018 592082 572254
rect 592318 572018 592500 572254
rect 591900 571934 592500 572018
rect 591900 571698 592082 571934
rect 592318 571698 592500 571934
rect 591900 536254 592500 571698
rect 591900 536018 592082 536254
rect 592318 536018 592500 536254
rect 591900 535934 592500 536018
rect 591900 535698 592082 535934
rect 592318 535698 592500 535934
rect 591900 500254 592500 535698
rect 591900 500018 592082 500254
rect 592318 500018 592500 500254
rect 591900 499934 592500 500018
rect 591900 499698 592082 499934
rect 592318 499698 592500 499934
rect 591900 464254 592500 499698
rect 591900 464018 592082 464254
rect 592318 464018 592500 464254
rect 591900 463934 592500 464018
rect 591900 463698 592082 463934
rect 592318 463698 592500 463934
rect 591900 428254 592500 463698
rect 591900 428018 592082 428254
rect 592318 428018 592500 428254
rect 591900 427934 592500 428018
rect 591900 427698 592082 427934
rect 592318 427698 592500 427934
rect 591900 392254 592500 427698
rect 591900 392018 592082 392254
rect 592318 392018 592500 392254
rect 591900 391934 592500 392018
rect 591900 391698 592082 391934
rect 592318 391698 592500 391934
rect 591900 356254 592500 391698
rect 591900 356018 592082 356254
rect 592318 356018 592500 356254
rect 591900 355934 592500 356018
rect 591900 355698 592082 355934
rect 592318 355698 592500 355934
rect 591900 320254 592500 355698
rect 591900 320018 592082 320254
rect 592318 320018 592500 320254
rect 591900 319934 592500 320018
rect 591900 319698 592082 319934
rect 592318 319698 592500 319934
rect 591900 284254 592500 319698
rect 591900 284018 592082 284254
rect 592318 284018 592500 284254
rect 591900 283934 592500 284018
rect 591900 283698 592082 283934
rect 592318 283698 592500 283934
rect 591900 248254 592500 283698
rect 591900 248018 592082 248254
rect 592318 248018 592500 248254
rect 591900 247934 592500 248018
rect 591900 247698 592082 247934
rect 592318 247698 592500 247934
rect 591900 212254 592500 247698
rect 591900 212018 592082 212254
rect 592318 212018 592500 212254
rect 591900 211934 592500 212018
rect 591900 211698 592082 211934
rect 592318 211698 592500 211934
rect 591900 176254 592500 211698
rect 591900 176018 592082 176254
rect 592318 176018 592500 176254
rect 591900 175934 592500 176018
rect 591900 175698 592082 175934
rect 592318 175698 592500 175934
rect 591900 140254 592500 175698
rect 591900 140018 592082 140254
rect 592318 140018 592500 140254
rect 591900 139934 592500 140018
rect 591900 139698 592082 139934
rect 592318 139698 592500 139934
rect 591900 104254 592500 139698
rect 591900 104018 592082 104254
rect 592318 104018 592500 104254
rect 591900 103934 592500 104018
rect 591900 103698 592082 103934
rect 592318 103698 592500 103934
rect 591900 68254 592500 103698
rect 591900 68018 592082 68254
rect 592318 68018 592500 68254
rect 591900 67934 592500 68018
rect 591900 67698 592082 67934
rect 592318 67698 592500 67934
rect 591900 32254 592500 67698
rect 591900 32018 592082 32254
rect 592318 32018 592500 32254
rect 591900 31934 592500 32018
rect 591900 31698 592082 31934
rect 592318 31698 592500 31934
rect 570604 -7162 570786 -6926
rect 571022 -7162 571204 -6926
rect 570604 -7246 571204 -7162
rect 570604 -7482 570786 -7246
rect 571022 -7482 571204 -7246
rect 570604 -7504 571204 -7482
rect 591900 -6926 592500 31698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 680018 -8158 680254
rect -8394 679698 -8158 679934
rect -8394 644018 -8158 644254
rect -8394 643698 -8158 643934
rect -8394 608018 -8158 608254
rect -8394 607698 -8158 607934
rect -8394 572018 -8158 572254
rect -8394 571698 -8158 571934
rect -8394 536018 -8158 536254
rect -8394 535698 -8158 535934
rect -8394 500018 -8158 500254
rect -8394 499698 -8158 499934
rect -8394 464018 -8158 464254
rect -8394 463698 -8158 463934
rect -8394 428018 -8158 428254
rect -8394 427698 -8158 427934
rect -8394 392018 -8158 392254
rect -8394 391698 -8158 391934
rect -8394 356018 -8158 356254
rect -8394 355698 -8158 355934
rect -8394 320018 -8158 320254
rect -8394 319698 -8158 319934
rect -8394 284018 -8158 284254
rect -8394 283698 -8158 283934
rect -8394 248018 -8158 248254
rect -8394 247698 -8158 247934
rect -8394 212018 -8158 212254
rect -8394 211698 -8158 211934
rect -8394 176018 -8158 176254
rect -8394 175698 -8158 175934
rect -8394 140018 -8158 140254
rect -8394 139698 -8158 139934
rect -8394 104018 -8158 104254
rect -8394 103698 -8158 103934
rect -8394 68018 -8158 68254
rect -8394 67698 -8158 67934
rect -8394 32018 -8158 32254
rect -8394 31698 -8158 31934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 12786 710242 13022 710478
rect 12786 709922 13022 710158
rect -7454 698018 -7218 698254
rect -7454 697698 -7218 697934
rect -7454 662018 -7218 662254
rect -7454 661698 -7218 661934
rect -7454 626018 -7218 626254
rect -7454 625698 -7218 625934
rect -7454 590018 -7218 590254
rect -7454 589698 -7218 589934
rect -7454 554018 -7218 554254
rect -7454 553698 -7218 553934
rect -7454 518018 -7218 518254
rect -7454 517698 -7218 517934
rect -7454 482018 -7218 482254
rect -7454 481698 -7218 481934
rect -7454 446018 -7218 446254
rect -7454 445698 -7218 445934
rect -7454 410018 -7218 410254
rect -7454 409698 -7218 409934
rect -7454 374018 -7218 374254
rect -7454 373698 -7218 373934
rect -7454 338018 -7218 338254
rect -7454 337698 -7218 337934
rect -7454 302018 -7218 302254
rect -7454 301698 -7218 301934
rect -7454 266018 -7218 266254
rect -7454 265698 -7218 265934
rect -7454 230018 -7218 230254
rect -7454 229698 -7218 229934
rect -7454 194018 -7218 194254
rect -7454 193698 -7218 193934
rect -7454 158018 -7218 158254
rect -7454 157698 -7218 157934
rect -7454 122018 -7218 122254
rect -7454 121698 -7218 121934
rect -7454 86018 -7218 86254
rect -7454 85698 -7218 85934
rect -7454 50018 -7218 50254
rect -7454 49698 -7218 49934
rect -7454 14018 -7218 14254
rect -7454 13698 -7218 13934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 676418 -6278 676654
rect -6514 676098 -6278 676334
rect -6514 640418 -6278 640654
rect -6514 640098 -6278 640334
rect -6514 604418 -6278 604654
rect -6514 604098 -6278 604334
rect -6514 568418 -6278 568654
rect -6514 568098 -6278 568334
rect -6514 532418 -6278 532654
rect -6514 532098 -6278 532334
rect -6514 496418 -6278 496654
rect -6514 496098 -6278 496334
rect -6514 460418 -6278 460654
rect -6514 460098 -6278 460334
rect -6514 424418 -6278 424654
rect -6514 424098 -6278 424334
rect -6514 388418 -6278 388654
rect -6514 388098 -6278 388334
rect -6514 352418 -6278 352654
rect -6514 352098 -6278 352334
rect -6514 316418 -6278 316654
rect -6514 316098 -6278 316334
rect -6514 280418 -6278 280654
rect -6514 280098 -6278 280334
rect -6514 244418 -6278 244654
rect -6514 244098 -6278 244334
rect -6514 208418 -6278 208654
rect -6514 208098 -6278 208334
rect -6514 172418 -6278 172654
rect -6514 172098 -6278 172334
rect -6514 136418 -6278 136654
rect -6514 136098 -6278 136334
rect -6514 100418 -6278 100654
rect -6514 100098 -6278 100334
rect -6514 64418 -6278 64654
rect -6514 64098 -6278 64334
rect -6514 28418 -6278 28654
rect -6514 28098 -6278 28334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 9186 708362 9422 708598
rect 9186 708042 9422 708278
rect -5574 694418 -5338 694654
rect -5574 694098 -5338 694334
rect -5574 658418 -5338 658654
rect -5574 658098 -5338 658334
rect -5574 622418 -5338 622654
rect -5574 622098 -5338 622334
rect -5574 586418 -5338 586654
rect -5574 586098 -5338 586334
rect -5574 550418 -5338 550654
rect -5574 550098 -5338 550334
rect -5574 514418 -5338 514654
rect -5574 514098 -5338 514334
rect -5574 478418 -5338 478654
rect -5574 478098 -5338 478334
rect -5574 442418 -5338 442654
rect -5574 442098 -5338 442334
rect -5574 406418 -5338 406654
rect -5574 406098 -5338 406334
rect -5574 370418 -5338 370654
rect -5574 370098 -5338 370334
rect -5574 334418 -5338 334654
rect -5574 334098 -5338 334334
rect -5574 298418 -5338 298654
rect -5574 298098 -5338 298334
rect -5574 262418 -5338 262654
rect -5574 262098 -5338 262334
rect -5574 226418 -5338 226654
rect -5574 226098 -5338 226334
rect -5574 190418 -5338 190654
rect -5574 190098 -5338 190334
rect -5574 154418 -5338 154654
rect -5574 154098 -5338 154334
rect -5574 118418 -5338 118654
rect -5574 118098 -5338 118334
rect -5574 82418 -5338 82654
rect -5574 82098 -5338 82334
rect -5574 46418 -5338 46654
rect -5574 46098 -5338 46334
rect -5574 10418 -5338 10654
rect -5574 10098 -5338 10334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 672818 -4398 673054
rect -4634 672498 -4398 672734
rect -4634 636818 -4398 637054
rect -4634 636498 -4398 636734
rect -4634 600818 -4398 601054
rect -4634 600498 -4398 600734
rect -4634 564818 -4398 565054
rect -4634 564498 -4398 564734
rect -4634 528818 -4398 529054
rect -4634 528498 -4398 528734
rect -4634 492818 -4398 493054
rect -4634 492498 -4398 492734
rect -4634 456818 -4398 457054
rect -4634 456498 -4398 456734
rect -4634 420818 -4398 421054
rect -4634 420498 -4398 420734
rect -4634 384818 -4398 385054
rect -4634 384498 -4398 384734
rect -4634 348818 -4398 349054
rect -4634 348498 -4398 348734
rect -4634 312818 -4398 313054
rect -4634 312498 -4398 312734
rect -4634 276818 -4398 277054
rect -4634 276498 -4398 276734
rect -4634 240818 -4398 241054
rect -4634 240498 -4398 240734
rect -4634 204818 -4398 205054
rect -4634 204498 -4398 204734
rect -4634 168818 -4398 169054
rect -4634 168498 -4398 168734
rect -4634 132818 -4398 133054
rect -4634 132498 -4398 132734
rect -4634 96818 -4398 97054
rect -4634 96498 -4398 96734
rect -4634 60818 -4398 61054
rect -4634 60498 -4398 60734
rect -4634 24818 -4398 25054
rect -4634 24498 -4398 24734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 5586 706482 5822 706718
rect 5586 706162 5822 706398
rect -3694 690818 -3458 691054
rect -3694 690498 -3458 690734
rect -3694 654818 -3458 655054
rect -3694 654498 -3458 654734
rect -3694 618818 -3458 619054
rect -3694 618498 -3458 618734
rect -3694 582818 -3458 583054
rect -3694 582498 -3458 582734
rect -3694 546818 -3458 547054
rect -3694 546498 -3458 546734
rect -3694 510818 -3458 511054
rect -3694 510498 -3458 510734
rect -3694 474818 -3458 475054
rect -3694 474498 -3458 474734
rect -3694 438818 -3458 439054
rect -3694 438498 -3458 438734
rect -3694 402818 -3458 403054
rect -3694 402498 -3458 402734
rect -3694 366818 -3458 367054
rect -3694 366498 -3458 366734
rect -3694 330818 -3458 331054
rect -3694 330498 -3458 330734
rect -3694 294818 -3458 295054
rect -3694 294498 -3458 294734
rect -3694 258818 -3458 259054
rect -3694 258498 -3458 258734
rect -3694 222818 -3458 223054
rect -3694 222498 -3458 222734
rect -3694 186818 -3458 187054
rect -3694 186498 -3458 186734
rect -3694 150818 -3458 151054
rect -3694 150498 -3458 150734
rect -3694 114818 -3458 115054
rect -3694 114498 -3458 114734
rect -3694 78818 -3458 79054
rect -3694 78498 -3458 78734
rect -3694 42818 -3458 43054
rect -3694 42498 -3458 42734
rect -3694 6818 -3458 7054
rect -3694 6498 -3458 6734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 669218 -2518 669454
rect -2754 668898 -2518 669134
rect -2754 633218 -2518 633454
rect -2754 632898 -2518 633134
rect -2754 597218 -2518 597454
rect -2754 596898 -2518 597134
rect -2754 561218 -2518 561454
rect -2754 560898 -2518 561134
rect -2754 525218 -2518 525454
rect -2754 524898 -2518 525134
rect -2754 489218 -2518 489454
rect -2754 488898 -2518 489134
rect -2754 453218 -2518 453454
rect -2754 452898 -2518 453134
rect -2754 417218 -2518 417454
rect -2754 416898 -2518 417134
rect -2754 381218 -2518 381454
rect -2754 380898 -2518 381134
rect -2754 345218 -2518 345454
rect -2754 344898 -2518 345134
rect -2754 309218 -2518 309454
rect -2754 308898 -2518 309134
rect -2754 273218 -2518 273454
rect -2754 272898 -2518 273134
rect -2754 237218 -2518 237454
rect -2754 236898 -2518 237134
rect -2754 201218 -2518 201454
rect -2754 200898 -2518 201134
rect -2754 165218 -2518 165454
rect -2754 164898 -2518 165134
rect -2754 129218 -2518 129454
rect -2754 128898 -2518 129134
rect -2754 93218 -2518 93454
rect -2754 92898 -2518 93134
rect -2754 57218 -2518 57454
rect -2754 56898 -2518 57134
rect -2754 21218 -2518 21454
rect -2754 20898 -2518 21134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 687218 -1578 687454
rect -1814 686898 -1578 687134
rect -1814 651218 -1578 651454
rect -1814 650898 -1578 651134
rect -1814 615218 -1578 615454
rect -1814 614898 -1578 615134
rect -1814 579218 -1578 579454
rect -1814 578898 -1578 579134
rect -1814 543218 -1578 543454
rect -1814 542898 -1578 543134
rect -1814 507218 -1578 507454
rect -1814 506898 -1578 507134
rect -1814 471218 -1578 471454
rect -1814 470898 -1578 471134
rect -1814 435218 -1578 435454
rect -1814 434898 -1578 435134
rect -1814 399218 -1578 399454
rect -1814 398898 -1578 399134
rect -1814 363218 -1578 363454
rect -1814 362898 -1578 363134
rect -1814 327218 -1578 327454
rect -1814 326898 -1578 327134
rect -1814 291218 -1578 291454
rect -1814 290898 -1578 291134
rect -1814 255218 -1578 255454
rect -1814 254898 -1578 255134
rect -1814 219218 -1578 219454
rect -1814 218898 -1578 219134
rect -1814 183218 -1578 183454
rect -1814 182898 -1578 183134
rect -1814 147218 -1578 147454
rect -1814 146898 -1578 147134
rect -1814 111218 -1578 111454
rect -1814 110898 -1578 111134
rect -1814 75218 -1578 75454
rect -1814 74898 -1578 75134
rect -1814 39218 -1578 39454
rect -1814 38898 -1578 39134
rect -1814 3218 -1578 3454
rect -1814 2898 -1578 3134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 1986 704602 2222 704838
rect 1986 704282 2222 704518
rect 1986 687218 2222 687454
rect 1986 686898 2222 687134
rect 5586 690818 5822 691054
rect 5586 690498 5822 690734
rect 1986 651218 2222 651454
rect 1986 650898 2222 651134
rect 1986 615218 2222 615454
rect 1986 614898 2222 615134
rect 1986 579218 2222 579454
rect 1986 578898 2222 579134
rect 1986 543218 2222 543454
rect 1986 542898 2222 543134
rect 1986 507218 2222 507454
rect 1986 506898 2222 507134
rect 5586 654818 5822 655054
rect 5586 654498 5822 654734
rect 5586 618818 5822 619054
rect 5586 618498 5822 618734
rect 5586 582818 5822 583054
rect 5586 582498 5822 582734
rect 5586 546818 5822 547054
rect 5586 546498 5822 546734
rect 5586 510818 5822 511054
rect 5586 510498 5822 510734
rect 5586 474818 5822 475054
rect 5586 474498 5822 474734
rect 1986 471218 2222 471454
rect 1986 470898 2222 471134
rect 1986 435218 2222 435454
rect 1986 434898 2222 435134
rect 1986 399218 2222 399454
rect 1986 398898 2222 399134
rect 1986 363218 2222 363454
rect 1986 362898 2222 363134
rect 1986 327218 2222 327454
rect 1986 326898 2222 327134
rect 1986 291218 2222 291454
rect 1986 290898 2222 291134
rect 1986 255218 2222 255454
rect 1986 254898 2222 255134
rect 1986 219218 2222 219454
rect 1986 218898 2222 219134
rect 1986 183218 2222 183454
rect 1986 182898 2222 183134
rect 1986 147218 2222 147454
rect 1986 146898 2222 147134
rect 1986 111218 2222 111454
rect 1986 110898 2222 111134
rect 1986 75218 2222 75454
rect 1986 74898 2222 75134
rect 1986 39218 2222 39454
rect 1986 38898 2222 39134
rect 1986 3218 2222 3454
rect 1986 2898 2222 3134
rect 1986 -582 2222 -346
rect 1986 -902 2222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 5586 438818 5822 439054
rect 5586 438498 5822 438734
rect 5586 402818 5822 403054
rect 5586 402498 5822 402734
rect 5586 366818 5822 367054
rect 5586 366498 5822 366734
rect 5586 330818 5822 331054
rect 5586 330498 5822 330734
rect 5586 294818 5822 295054
rect 5586 294498 5822 294734
rect 5586 258818 5822 259054
rect 5586 258498 5822 258734
rect 5586 222818 5822 223054
rect 5586 222498 5822 222734
rect 5586 186818 5822 187054
rect 5586 186498 5822 186734
rect 5586 150818 5822 151054
rect 5586 150498 5822 150734
rect 5586 114818 5822 115054
rect 5586 114498 5822 114734
rect 5586 78818 5822 79054
rect 5586 78498 5822 78734
rect 5586 42818 5822 43054
rect 5586 42498 5822 42734
rect 5586 6818 5822 7054
rect 5586 6498 5822 6734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 5586 -2462 5822 -2226
rect 5586 -2782 5822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 9186 694418 9422 694654
rect 9186 694098 9422 694334
rect 9186 658418 9422 658654
rect 9186 658098 9422 658334
rect 9186 622418 9422 622654
rect 9186 622098 9422 622334
rect 9186 586418 9422 586654
rect 9186 586098 9422 586334
rect 9186 550418 9422 550654
rect 9186 550098 9422 550334
rect 9186 514418 9422 514654
rect 9186 514098 9422 514334
rect 9186 478418 9422 478654
rect 9186 478098 9422 478334
rect 9186 442418 9422 442654
rect 9186 442098 9422 442334
rect 9186 406418 9422 406654
rect 9186 406098 9422 406334
rect 9186 370418 9422 370654
rect 9186 370098 9422 370334
rect 9186 334418 9422 334654
rect 9186 334098 9422 334334
rect 9186 298418 9422 298654
rect 9186 298098 9422 298334
rect 9186 262418 9422 262654
rect 9186 262098 9422 262334
rect 9186 226418 9422 226654
rect 9186 226098 9422 226334
rect 9186 190418 9422 190654
rect 9186 190098 9422 190334
rect 9186 154418 9422 154654
rect 9186 154098 9422 154334
rect 9186 118418 9422 118654
rect 9186 118098 9422 118334
rect 9186 82418 9422 82654
rect 9186 82098 9422 82334
rect 9186 46418 9422 46654
rect 9186 46098 9422 46334
rect 9186 10418 9422 10654
rect 9186 10098 9422 10334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 9186 -4342 9422 -4106
rect 9186 -4662 9422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 30786 711182 31022 711418
rect 30786 710862 31022 711098
rect 27186 709302 27422 709538
rect 27186 708982 27422 709218
rect 23586 707422 23822 707658
rect 23586 707102 23822 707338
rect 12786 698018 13022 698254
rect 12786 697698 13022 697934
rect 12786 662018 13022 662254
rect 12786 661698 13022 661934
rect 12786 626018 13022 626254
rect 12786 625698 13022 625934
rect 12786 590018 13022 590254
rect 12786 589698 13022 589934
rect 12786 554018 13022 554254
rect 12786 553698 13022 553934
rect 12786 518018 13022 518254
rect 12786 517698 13022 517934
rect 12786 482018 13022 482254
rect 12786 481698 13022 481934
rect 12786 446018 13022 446254
rect 12786 445698 13022 445934
rect 12786 410018 13022 410254
rect 12786 409698 13022 409934
rect 12786 374018 13022 374254
rect 12786 373698 13022 373934
rect 12786 338018 13022 338254
rect 12786 337698 13022 337934
rect 12786 302018 13022 302254
rect 12786 301698 13022 301934
rect 12786 266018 13022 266254
rect 12786 265698 13022 265934
rect 12786 230018 13022 230254
rect 12786 229698 13022 229934
rect 12786 194018 13022 194254
rect 12786 193698 13022 193934
rect 12786 158018 13022 158254
rect 12786 157698 13022 157934
rect 12786 122018 13022 122254
rect 12786 121698 13022 121934
rect 12786 86018 13022 86254
rect 12786 85698 13022 85934
rect 12786 50018 13022 50254
rect 12786 49698 13022 49934
rect 12786 14018 13022 14254
rect 12786 13698 13022 13934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 19986 705542 20222 705778
rect 19986 705222 20222 705458
rect 19986 669218 20222 669454
rect 19986 668898 20222 669134
rect 19986 633218 20222 633454
rect 19986 632898 20222 633134
rect 19986 597218 20222 597454
rect 19986 596898 20222 597134
rect 19986 561218 20222 561454
rect 19986 560898 20222 561134
rect 19986 525218 20222 525454
rect 19986 524898 20222 525134
rect 19986 489218 20222 489454
rect 19986 488898 20222 489134
rect 19986 453218 20222 453454
rect 19986 452898 20222 453134
rect 19986 417218 20222 417454
rect 19986 416898 20222 417134
rect 19986 381218 20222 381454
rect 19986 380898 20222 381134
rect 19986 345218 20222 345454
rect 19986 344898 20222 345134
rect 19986 309218 20222 309454
rect 19986 308898 20222 309134
rect 19986 273218 20222 273454
rect 19986 272898 20222 273134
rect 19986 237218 20222 237454
rect 19986 236898 20222 237134
rect 19986 201218 20222 201454
rect 19986 200898 20222 201134
rect 19986 165218 20222 165454
rect 19986 164898 20222 165134
rect 19986 129218 20222 129454
rect 19986 128898 20222 129134
rect 19986 93218 20222 93454
rect 19986 92898 20222 93134
rect 19986 57218 20222 57454
rect 19986 56898 20222 57134
rect 19986 21218 20222 21454
rect 19986 20898 20222 21134
rect 19986 -1522 20222 -1286
rect 19986 -1842 20222 -1606
rect 23586 672818 23822 673054
rect 23586 672498 23822 672734
rect 23586 636818 23822 637054
rect 23586 636498 23822 636734
rect 23586 600818 23822 601054
rect 23586 600498 23822 600734
rect 23586 564818 23822 565054
rect 23586 564498 23822 564734
rect 23586 528818 23822 529054
rect 23586 528498 23822 528734
rect 23586 492818 23822 493054
rect 23586 492498 23822 492734
rect 23586 456818 23822 457054
rect 23586 456498 23822 456734
rect 23586 420818 23822 421054
rect 23586 420498 23822 420734
rect 23586 384818 23822 385054
rect 23586 384498 23822 384734
rect 23586 348818 23822 349054
rect 23586 348498 23822 348734
rect 23586 312818 23822 313054
rect 23586 312498 23822 312734
rect 23586 276818 23822 277054
rect 23586 276498 23822 276734
rect 23586 240818 23822 241054
rect 23586 240498 23822 240734
rect 23586 204818 23822 205054
rect 23586 204498 23822 204734
rect 23586 168818 23822 169054
rect 23586 168498 23822 168734
rect 23586 132818 23822 133054
rect 23586 132498 23822 132734
rect 23586 96818 23822 97054
rect 23586 96498 23822 96734
rect 23586 60818 23822 61054
rect 23586 60498 23822 60734
rect 23586 24818 23822 25054
rect 23586 24498 23822 24734
rect 23586 -3402 23822 -3166
rect 23586 -3722 23822 -3486
rect 27186 676418 27422 676654
rect 27186 676098 27422 676334
rect 27186 640418 27422 640654
rect 27186 640098 27422 640334
rect 27186 604418 27422 604654
rect 27186 604098 27422 604334
rect 27186 568418 27422 568654
rect 27186 568098 27422 568334
rect 27186 532418 27422 532654
rect 27186 532098 27422 532334
rect 27186 496418 27422 496654
rect 27186 496098 27422 496334
rect 27186 460418 27422 460654
rect 27186 460098 27422 460334
rect 27186 424418 27422 424654
rect 27186 424098 27422 424334
rect 27186 388418 27422 388654
rect 27186 388098 27422 388334
rect 27186 352418 27422 352654
rect 27186 352098 27422 352334
rect 27186 316418 27422 316654
rect 27186 316098 27422 316334
rect 27186 280418 27422 280654
rect 27186 280098 27422 280334
rect 27186 244418 27422 244654
rect 27186 244098 27422 244334
rect 27186 208418 27422 208654
rect 27186 208098 27422 208334
rect 27186 172418 27422 172654
rect 27186 172098 27422 172334
rect 27186 136418 27422 136654
rect 27186 136098 27422 136334
rect 27186 100418 27422 100654
rect 27186 100098 27422 100334
rect 27186 64418 27422 64654
rect 27186 64098 27422 64334
rect 27186 28418 27422 28654
rect 27186 28098 27422 28334
rect 27186 -5282 27422 -5046
rect 27186 -5602 27422 -5366
rect 48786 710242 49022 710478
rect 48786 709922 49022 710158
rect 45186 708362 45422 708598
rect 45186 708042 45422 708278
rect 41586 706482 41822 706718
rect 41586 706162 41822 706398
rect 30786 680018 31022 680254
rect 30786 679698 31022 679934
rect 30786 644018 31022 644254
rect 30786 643698 31022 643934
rect 30786 608018 31022 608254
rect 30786 607698 31022 607934
rect 30786 572018 31022 572254
rect 30786 571698 31022 571934
rect 30786 536018 31022 536254
rect 30786 535698 31022 535934
rect 30786 500018 31022 500254
rect 30786 499698 31022 499934
rect 30786 464018 31022 464254
rect 30786 463698 31022 463934
rect 30786 428018 31022 428254
rect 30786 427698 31022 427934
rect 30786 392018 31022 392254
rect 30786 391698 31022 391934
rect 30786 356018 31022 356254
rect 30786 355698 31022 355934
rect 30786 320018 31022 320254
rect 30786 319698 31022 319934
rect 30786 284018 31022 284254
rect 30786 283698 31022 283934
rect 30786 248018 31022 248254
rect 30786 247698 31022 247934
rect 30786 212018 31022 212254
rect 30786 211698 31022 211934
rect 30786 176018 31022 176254
rect 30786 175698 31022 175934
rect 30786 140018 31022 140254
rect 30786 139698 31022 139934
rect 30786 104018 31022 104254
rect 30786 103698 31022 103934
rect 30786 68018 31022 68254
rect 30786 67698 31022 67934
rect 30786 32018 31022 32254
rect 30786 31698 31022 31934
rect 12786 -6222 13022 -5986
rect 12786 -6542 13022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 37986 704602 38222 704838
rect 37986 704282 38222 704518
rect 37986 687218 38222 687454
rect 37986 686898 38222 687134
rect 37986 651218 38222 651454
rect 37986 650898 38222 651134
rect 37986 615218 38222 615454
rect 37986 614898 38222 615134
rect 37986 579218 38222 579454
rect 37986 578898 38222 579134
rect 37986 543218 38222 543454
rect 37986 542898 38222 543134
rect 37986 507218 38222 507454
rect 37986 506898 38222 507134
rect 37986 471218 38222 471454
rect 37986 470898 38222 471134
rect 37986 435218 38222 435454
rect 37986 434898 38222 435134
rect 37986 399218 38222 399454
rect 37986 398898 38222 399134
rect 37986 363218 38222 363454
rect 37986 362898 38222 363134
rect 37986 327218 38222 327454
rect 37986 326898 38222 327134
rect 37986 291218 38222 291454
rect 37986 290898 38222 291134
rect 37986 255218 38222 255454
rect 37986 254898 38222 255134
rect 37986 219218 38222 219454
rect 37986 218898 38222 219134
rect 37986 183218 38222 183454
rect 37986 182898 38222 183134
rect 37986 147218 38222 147454
rect 37986 146898 38222 147134
rect 37986 111218 38222 111454
rect 37986 110898 38222 111134
rect 37986 75218 38222 75454
rect 37986 74898 38222 75134
rect 37986 39218 38222 39454
rect 37986 38898 38222 39134
rect 37986 3218 38222 3454
rect 37986 2898 38222 3134
rect 37986 -582 38222 -346
rect 37986 -902 38222 -666
rect 41586 690818 41822 691054
rect 41586 690498 41822 690734
rect 41586 654818 41822 655054
rect 41586 654498 41822 654734
rect 41586 618818 41822 619054
rect 41586 618498 41822 618734
rect 41586 582818 41822 583054
rect 41586 582498 41822 582734
rect 41586 546818 41822 547054
rect 41586 546498 41822 546734
rect 41586 510818 41822 511054
rect 41586 510498 41822 510734
rect 41586 474818 41822 475054
rect 41586 474498 41822 474734
rect 41586 438818 41822 439054
rect 41586 438498 41822 438734
rect 41586 402818 41822 403054
rect 41586 402498 41822 402734
rect 41586 366818 41822 367054
rect 41586 366498 41822 366734
rect 41586 330818 41822 331054
rect 41586 330498 41822 330734
rect 41586 294818 41822 295054
rect 41586 294498 41822 294734
rect 41586 258818 41822 259054
rect 41586 258498 41822 258734
rect 41586 222818 41822 223054
rect 41586 222498 41822 222734
rect 41586 186818 41822 187054
rect 41586 186498 41822 186734
rect 41586 150818 41822 151054
rect 41586 150498 41822 150734
rect 41586 114818 41822 115054
rect 41586 114498 41822 114734
rect 41586 78818 41822 79054
rect 41586 78498 41822 78734
rect 41586 42818 41822 43054
rect 41586 42498 41822 42734
rect 41586 6818 41822 7054
rect 41586 6498 41822 6734
rect 41586 -2462 41822 -2226
rect 41586 -2782 41822 -2546
rect 45186 694418 45422 694654
rect 45186 694098 45422 694334
rect 45186 658418 45422 658654
rect 45186 658098 45422 658334
rect 45186 622418 45422 622654
rect 45186 622098 45422 622334
rect 45186 586418 45422 586654
rect 45186 586098 45422 586334
rect 45186 550418 45422 550654
rect 45186 550098 45422 550334
rect 45186 514418 45422 514654
rect 45186 514098 45422 514334
rect 45186 478418 45422 478654
rect 45186 478098 45422 478334
rect 45186 442418 45422 442654
rect 45186 442098 45422 442334
rect 45186 406418 45422 406654
rect 45186 406098 45422 406334
rect 45186 370418 45422 370654
rect 45186 370098 45422 370334
rect 45186 334418 45422 334654
rect 45186 334098 45422 334334
rect 45186 298418 45422 298654
rect 45186 298098 45422 298334
rect 45186 262418 45422 262654
rect 45186 262098 45422 262334
rect 45186 226418 45422 226654
rect 45186 226098 45422 226334
rect 45186 190418 45422 190654
rect 45186 190098 45422 190334
rect 45186 154418 45422 154654
rect 45186 154098 45422 154334
rect 45186 118418 45422 118654
rect 45186 118098 45422 118334
rect 45186 82418 45422 82654
rect 45186 82098 45422 82334
rect 45186 46418 45422 46654
rect 45186 46098 45422 46334
rect 45186 10418 45422 10654
rect 45186 10098 45422 10334
rect 45186 -4342 45422 -4106
rect 45186 -4662 45422 -4426
rect 66786 711182 67022 711418
rect 66786 710862 67022 711098
rect 63186 709302 63422 709538
rect 63186 708982 63422 709218
rect 59586 707422 59822 707658
rect 59586 707102 59822 707338
rect 48786 698018 49022 698254
rect 48786 697698 49022 697934
rect 48786 662018 49022 662254
rect 48786 661698 49022 661934
rect 48786 626018 49022 626254
rect 48786 625698 49022 625934
rect 48786 590018 49022 590254
rect 48786 589698 49022 589934
rect 48786 554018 49022 554254
rect 48786 553698 49022 553934
rect 48786 518018 49022 518254
rect 48786 517698 49022 517934
rect 48786 482018 49022 482254
rect 48786 481698 49022 481934
rect 48786 446018 49022 446254
rect 48786 445698 49022 445934
rect 48786 410018 49022 410254
rect 48786 409698 49022 409934
rect 48786 374018 49022 374254
rect 48786 373698 49022 373934
rect 48786 338018 49022 338254
rect 48786 337698 49022 337934
rect 48786 302018 49022 302254
rect 48786 301698 49022 301934
rect 48786 266018 49022 266254
rect 48786 265698 49022 265934
rect 48786 230018 49022 230254
rect 48786 229698 49022 229934
rect 48786 194018 49022 194254
rect 48786 193698 49022 193934
rect 48786 158018 49022 158254
rect 48786 157698 49022 157934
rect 48786 122018 49022 122254
rect 48786 121698 49022 121934
rect 48786 86018 49022 86254
rect 48786 85698 49022 85934
rect 48786 50018 49022 50254
rect 48786 49698 49022 49934
rect 48786 14018 49022 14254
rect 48786 13698 49022 13934
rect 30786 -7162 31022 -6926
rect 30786 -7482 31022 -7246
rect 55986 705542 56222 705778
rect 55986 705222 56222 705458
rect 55986 669218 56222 669454
rect 55986 668898 56222 669134
rect 55986 633218 56222 633454
rect 55986 632898 56222 633134
rect 55986 597218 56222 597454
rect 55986 596898 56222 597134
rect 55986 561218 56222 561454
rect 55986 560898 56222 561134
rect 55986 525218 56222 525454
rect 55986 524898 56222 525134
rect 55986 489218 56222 489454
rect 55986 488898 56222 489134
rect 55986 453218 56222 453454
rect 55986 452898 56222 453134
rect 55986 417218 56222 417454
rect 55986 416898 56222 417134
rect 55986 381218 56222 381454
rect 55986 380898 56222 381134
rect 55986 345218 56222 345454
rect 55986 344898 56222 345134
rect 55986 309218 56222 309454
rect 55986 308898 56222 309134
rect 55986 273218 56222 273454
rect 55986 272898 56222 273134
rect 55986 237218 56222 237454
rect 55986 236898 56222 237134
rect 55986 201218 56222 201454
rect 55986 200898 56222 201134
rect 55986 165218 56222 165454
rect 55986 164898 56222 165134
rect 55986 129218 56222 129454
rect 55986 128898 56222 129134
rect 55986 93218 56222 93454
rect 55986 92898 56222 93134
rect 55986 57218 56222 57454
rect 55986 56898 56222 57134
rect 55986 21218 56222 21454
rect 55986 20898 56222 21134
rect 55986 -1522 56222 -1286
rect 55986 -1842 56222 -1606
rect 59586 672818 59822 673054
rect 59586 672498 59822 672734
rect 59586 636818 59822 637054
rect 59586 636498 59822 636734
rect 59586 600818 59822 601054
rect 59586 600498 59822 600734
rect 59586 564818 59822 565054
rect 59586 564498 59822 564734
rect 59586 528818 59822 529054
rect 59586 528498 59822 528734
rect 59586 492818 59822 493054
rect 59586 492498 59822 492734
rect 59586 456818 59822 457054
rect 59586 456498 59822 456734
rect 59586 420818 59822 421054
rect 59586 420498 59822 420734
rect 59586 384818 59822 385054
rect 59586 384498 59822 384734
rect 59586 348818 59822 349054
rect 59586 348498 59822 348734
rect 59586 312818 59822 313054
rect 59586 312498 59822 312734
rect 59586 276818 59822 277054
rect 59586 276498 59822 276734
rect 59586 240818 59822 241054
rect 59586 240498 59822 240734
rect 59586 204818 59822 205054
rect 59586 204498 59822 204734
rect 59586 168818 59822 169054
rect 59586 168498 59822 168734
rect 59586 132818 59822 133054
rect 59586 132498 59822 132734
rect 59586 96818 59822 97054
rect 59586 96498 59822 96734
rect 59586 60818 59822 61054
rect 59586 60498 59822 60734
rect 59586 24818 59822 25054
rect 59586 24498 59822 24734
rect 59586 -3402 59822 -3166
rect 59586 -3722 59822 -3486
rect 63186 676418 63422 676654
rect 63186 676098 63422 676334
rect 63186 640418 63422 640654
rect 63186 640098 63422 640334
rect 63186 604418 63422 604654
rect 63186 604098 63422 604334
rect 63186 568418 63422 568654
rect 63186 568098 63422 568334
rect 63186 532418 63422 532654
rect 63186 532098 63422 532334
rect 63186 496418 63422 496654
rect 63186 496098 63422 496334
rect 63186 460418 63422 460654
rect 63186 460098 63422 460334
rect 63186 424418 63422 424654
rect 63186 424098 63422 424334
rect 63186 388418 63422 388654
rect 63186 388098 63422 388334
rect 63186 352418 63422 352654
rect 63186 352098 63422 352334
rect 63186 316418 63422 316654
rect 63186 316098 63422 316334
rect 63186 280418 63422 280654
rect 63186 280098 63422 280334
rect 63186 244418 63422 244654
rect 63186 244098 63422 244334
rect 63186 208418 63422 208654
rect 63186 208098 63422 208334
rect 63186 172418 63422 172654
rect 63186 172098 63422 172334
rect 63186 136418 63422 136654
rect 63186 136098 63422 136334
rect 63186 100418 63422 100654
rect 63186 100098 63422 100334
rect 63186 64418 63422 64654
rect 63186 64098 63422 64334
rect 63186 28418 63422 28654
rect 63186 28098 63422 28334
rect 63186 -5282 63422 -5046
rect 63186 -5602 63422 -5366
rect 84786 710242 85022 710478
rect 84786 709922 85022 710158
rect 81186 708362 81422 708598
rect 81186 708042 81422 708278
rect 77586 706482 77822 706718
rect 77586 706162 77822 706398
rect 66786 680018 67022 680254
rect 66786 679698 67022 679934
rect 66786 644018 67022 644254
rect 66786 643698 67022 643934
rect 66786 608018 67022 608254
rect 66786 607698 67022 607934
rect 66786 572018 67022 572254
rect 66786 571698 67022 571934
rect 66786 536018 67022 536254
rect 66786 535698 67022 535934
rect 66786 500018 67022 500254
rect 66786 499698 67022 499934
rect 66786 464018 67022 464254
rect 66786 463698 67022 463934
rect 66786 428018 67022 428254
rect 66786 427698 67022 427934
rect 66786 392018 67022 392254
rect 66786 391698 67022 391934
rect 66786 356018 67022 356254
rect 66786 355698 67022 355934
rect 66786 320018 67022 320254
rect 66786 319698 67022 319934
rect 66786 284018 67022 284254
rect 66786 283698 67022 283934
rect 66786 248018 67022 248254
rect 66786 247698 67022 247934
rect 66786 212018 67022 212254
rect 66786 211698 67022 211934
rect 66786 176018 67022 176254
rect 66786 175698 67022 175934
rect 66786 140018 67022 140254
rect 66786 139698 67022 139934
rect 66786 104018 67022 104254
rect 66786 103698 67022 103934
rect 66786 68018 67022 68254
rect 66786 67698 67022 67934
rect 66786 32018 67022 32254
rect 66786 31698 67022 31934
rect 48786 -6222 49022 -5986
rect 48786 -6542 49022 -6306
rect 73986 704602 74222 704838
rect 73986 704282 74222 704518
rect 73986 687218 74222 687454
rect 73986 686898 74222 687134
rect 73986 651218 74222 651454
rect 73986 650898 74222 651134
rect 73986 615218 74222 615454
rect 73986 614898 74222 615134
rect 73986 579218 74222 579454
rect 73986 578898 74222 579134
rect 73986 543218 74222 543454
rect 73986 542898 74222 543134
rect 73986 507218 74222 507454
rect 73986 506898 74222 507134
rect 73986 471218 74222 471454
rect 73986 470898 74222 471134
rect 73986 435218 74222 435454
rect 73986 434898 74222 435134
rect 73986 399218 74222 399454
rect 73986 398898 74222 399134
rect 73986 363218 74222 363454
rect 73986 362898 74222 363134
rect 73986 327218 74222 327454
rect 73986 326898 74222 327134
rect 73986 291218 74222 291454
rect 73986 290898 74222 291134
rect 73986 255218 74222 255454
rect 73986 254898 74222 255134
rect 73986 219218 74222 219454
rect 73986 218898 74222 219134
rect 73986 183218 74222 183454
rect 73986 182898 74222 183134
rect 73986 147218 74222 147454
rect 73986 146898 74222 147134
rect 73986 111218 74222 111454
rect 73986 110898 74222 111134
rect 73986 75218 74222 75454
rect 73986 74898 74222 75134
rect 73986 39218 74222 39454
rect 73986 38898 74222 39134
rect 73986 3218 74222 3454
rect 73986 2898 74222 3134
rect 73986 -582 74222 -346
rect 73986 -902 74222 -666
rect 77586 690818 77822 691054
rect 77586 690498 77822 690734
rect 77586 654818 77822 655054
rect 77586 654498 77822 654734
rect 77586 618818 77822 619054
rect 77586 618498 77822 618734
rect 77586 582818 77822 583054
rect 77586 582498 77822 582734
rect 77586 546818 77822 547054
rect 77586 546498 77822 546734
rect 77586 510818 77822 511054
rect 77586 510498 77822 510734
rect 77586 474818 77822 475054
rect 77586 474498 77822 474734
rect 77586 438818 77822 439054
rect 77586 438498 77822 438734
rect 77586 402818 77822 403054
rect 77586 402498 77822 402734
rect 77586 366818 77822 367054
rect 77586 366498 77822 366734
rect 77586 330818 77822 331054
rect 77586 330498 77822 330734
rect 77586 294818 77822 295054
rect 77586 294498 77822 294734
rect 77586 258818 77822 259054
rect 77586 258498 77822 258734
rect 77586 222818 77822 223054
rect 77586 222498 77822 222734
rect 77586 186818 77822 187054
rect 77586 186498 77822 186734
rect 77586 150818 77822 151054
rect 77586 150498 77822 150734
rect 77586 114818 77822 115054
rect 77586 114498 77822 114734
rect 77586 78818 77822 79054
rect 77586 78498 77822 78734
rect 77586 42818 77822 43054
rect 77586 42498 77822 42734
rect 77586 6818 77822 7054
rect 77586 6498 77822 6734
rect 77586 -2462 77822 -2226
rect 77586 -2782 77822 -2546
rect 81186 694418 81422 694654
rect 81186 694098 81422 694334
rect 81186 658418 81422 658654
rect 81186 658098 81422 658334
rect 81186 622418 81422 622654
rect 81186 622098 81422 622334
rect 81186 586418 81422 586654
rect 81186 586098 81422 586334
rect 81186 550418 81422 550654
rect 81186 550098 81422 550334
rect 81186 514418 81422 514654
rect 81186 514098 81422 514334
rect 81186 478418 81422 478654
rect 81186 478098 81422 478334
rect 81186 442418 81422 442654
rect 81186 442098 81422 442334
rect 81186 406418 81422 406654
rect 81186 406098 81422 406334
rect 81186 370418 81422 370654
rect 81186 370098 81422 370334
rect 81186 334418 81422 334654
rect 81186 334098 81422 334334
rect 81186 298418 81422 298654
rect 81186 298098 81422 298334
rect 81186 262418 81422 262654
rect 81186 262098 81422 262334
rect 81186 226418 81422 226654
rect 81186 226098 81422 226334
rect 81186 190418 81422 190654
rect 81186 190098 81422 190334
rect 81186 154418 81422 154654
rect 81186 154098 81422 154334
rect 81186 118418 81422 118654
rect 81186 118098 81422 118334
rect 81186 82418 81422 82654
rect 81186 82098 81422 82334
rect 81186 46418 81422 46654
rect 81186 46098 81422 46334
rect 81186 10418 81422 10654
rect 81186 10098 81422 10334
rect 81186 -4342 81422 -4106
rect 81186 -4662 81422 -4426
rect 102786 711182 103022 711418
rect 102786 710862 103022 711098
rect 99186 709302 99422 709538
rect 99186 708982 99422 709218
rect 95586 707422 95822 707658
rect 95586 707102 95822 707338
rect 84786 698018 85022 698254
rect 84786 697698 85022 697934
rect 84786 662018 85022 662254
rect 84786 661698 85022 661934
rect 84786 626018 85022 626254
rect 84786 625698 85022 625934
rect 84786 590018 85022 590254
rect 84786 589698 85022 589934
rect 84786 554018 85022 554254
rect 84786 553698 85022 553934
rect 84786 518018 85022 518254
rect 84786 517698 85022 517934
rect 84786 482018 85022 482254
rect 84786 481698 85022 481934
rect 84786 446018 85022 446254
rect 84786 445698 85022 445934
rect 84786 410018 85022 410254
rect 84786 409698 85022 409934
rect 84786 374018 85022 374254
rect 84786 373698 85022 373934
rect 84786 338018 85022 338254
rect 84786 337698 85022 337934
rect 84786 302018 85022 302254
rect 84786 301698 85022 301934
rect 84786 266018 85022 266254
rect 84786 265698 85022 265934
rect 84786 230018 85022 230254
rect 84786 229698 85022 229934
rect 84786 194018 85022 194254
rect 84786 193698 85022 193934
rect 84786 158018 85022 158254
rect 84786 157698 85022 157934
rect 84786 122018 85022 122254
rect 84786 121698 85022 121934
rect 84786 86018 85022 86254
rect 84786 85698 85022 85934
rect 84786 50018 85022 50254
rect 84786 49698 85022 49934
rect 84786 14018 85022 14254
rect 84786 13698 85022 13934
rect 66786 -7162 67022 -6926
rect 66786 -7482 67022 -7246
rect 91986 705542 92222 705778
rect 91986 705222 92222 705458
rect 91986 669218 92222 669454
rect 91986 668898 92222 669134
rect 91986 633218 92222 633454
rect 91986 632898 92222 633134
rect 91986 597218 92222 597454
rect 91986 596898 92222 597134
rect 91986 561218 92222 561454
rect 91986 560898 92222 561134
rect 91986 525218 92222 525454
rect 91986 524898 92222 525134
rect 91986 489218 92222 489454
rect 91986 488898 92222 489134
rect 91986 453218 92222 453454
rect 91986 452898 92222 453134
rect 91986 417218 92222 417454
rect 91986 416898 92222 417134
rect 91986 381218 92222 381454
rect 91986 380898 92222 381134
rect 91986 345218 92222 345454
rect 91986 344898 92222 345134
rect 91986 309218 92222 309454
rect 91986 308898 92222 309134
rect 91986 273218 92222 273454
rect 91986 272898 92222 273134
rect 91986 237218 92222 237454
rect 91986 236898 92222 237134
rect 91986 201218 92222 201454
rect 91986 200898 92222 201134
rect 91986 165218 92222 165454
rect 91986 164898 92222 165134
rect 91986 129218 92222 129454
rect 91986 128898 92222 129134
rect 91986 93218 92222 93454
rect 91986 92898 92222 93134
rect 91986 57218 92222 57454
rect 91986 56898 92222 57134
rect 91986 21218 92222 21454
rect 91986 20898 92222 21134
rect 91986 -1522 92222 -1286
rect 91986 -1842 92222 -1606
rect 95586 672818 95822 673054
rect 95586 672498 95822 672734
rect 95586 636818 95822 637054
rect 95586 636498 95822 636734
rect 95586 600818 95822 601054
rect 95586 600498 95822 600734
rect 95586 564818 95822 565054
rect 95586 564498 95822 564734
rect 95586 528818 95822 529054
rect 95586 528498 95822 528734
rect 95586 492818 95822 493054
rect 95586 492498 95822 492734
rect 95586 456818 95822 457054
rect 95586 456498 95822 456734
rect 95586 420818 95822 421054
rect 95586 420498 95822 420734
rect 95586 384818 95822 385054
rect 95586 384498 95822 384734
rect 95586 348818 95822 349054
rect 95586 348498 95822 348734
rect 95586 312818 95822 313054
rect 95586 312498 95822 312734
rect 95586 276818 95822 277054
rect 95586 276498 95822 276734
rect 95586 240818 95822 241054
rect 95586 240498 95822 240734
rect 95586 204818 95822 205054
rect 95586 204498 95822 204734
rect 95586 168818 95822 169054
rect 95586 168498 95822 168734
rect 95586 132818 95822 133054
rect 95586 132498 95822 132734
rect 95586 96818 95822 97054
rect 95586 96498 95822 96734
rect 95586 60818 95822 61054
rect 95586 60498 95822 60734
rect 95586 24818 95822 25054
rect 95586 24498 95822 24734
rect 95586 -3402 95822 -3166
rect 95586 -3722 95822 -3486
rect 99186 676418 99422 676654
rect 99186 676098 99422 676334
rect 99186 640418 99422 640654
rect 99186 640098 99422 640334
rect 99186 604418 99422 604654
rect 99186 604098 99422 604334
rect 99186 568418 99422 568654
rect 99186 568098 99422 568334
rect 99186 532418 99422 532654
rect 99186 532098 99422 532334
rect 99186 496418 99422 496654
rect 99186 496098 99422 496334
rect 99186 460418 99422 460654
rect 99186 460098 99422 460334
rect 99186 424418 99422 424654
rect 99186 424098 99422 424334
rect 99186 388418 99422 388654
rect 99186 388098 99422 388334
rect 99186 352418 99422 352654
rect 99186 352098 99422 352334
rect 99186 316418 99422 316654
rect 99186 316098 99422 316334
rect 99186 280418 99422 280654
rect 99186 280098 99422 280334
rect 99186 244418 99422 244654
rect 99186 244098 99422 244334
rect 99186 208418 99422 208654
rect 99186 208098 99422 208334
rect 99186 172418 99422 172654
rect 99186 172098 99422 172334
rect 99186 136418 99422 136654
rect 99186 136098 99422 136334
rect 99186 100418 99422 100654
rect 99186 100098 99422 100334
rect 99186 64418 99422 64654
rect 99186 64098 99422 64334
rect 99186 28418 99422 28654
rect 99186 28098 99422 28334
rect 99186 -5282 99422 -5046
rect 99186 -5602 99422 -5366
rect 120786 710242 121022 710478
rect 120786 709922 121022 710158
rect 117186 708362 117422 708598
rect 117186 708042 117422 708278
rect 113586 706482 113822 706718
rect 113586 706162 113822 706398
rect 102786 680018 103022 680254
rect 102786 679698 103022 679934
rect 102786 644018 103022 644254
rect 102786 643698 103022 643934
rect 102786 608018 103022 608254
rect 102786 607698 103022 607934
rect 109986 704602 110222 704838
rect 109986 704282 110222 704518
rect 109986 687218 110222 687454
rect 109986 686898 110222 687134
rect 109986 651218 110222 651454
rect 109986 650898 110222 651134
rect 109986 615218 110222 615454
rect 109986 614898 110222 615134
rect 113586 690818 113822 691054
rect 113586 690498 113822 690734
rect 113586 654818 113822 655054
rect 113586 654498 113822 654734
rect 113586 618818 113822 619054
rect 113586 618498 113822 618734
rect 117186 694418 117422 694654
rect 117186 694098 117422 694334
rect 117186 658418 117422 658654
rect 117186 658098 117422 658334
rect 117186 622418 117422 622654
rect 117186 622098 117422 622334
rect 138786 711182 139022 711418
rect 138786 710862 139022 711098
rect 135186 709302 135422 709538
rect 135186 708982 135422 709218
rect 131586 707422 131822 707658
rect 131586 707102 131822 707338
rect 120786 698018 121022 698254
rect 120786 697698 121022 697934
rect 120786 662018 121022 662254
rect 120786 661698 121022 661934
rect 120786 626018 121022 626254
rect 120786 625698 121022 625934
rect 127986 705542 128222 705778
rect 127986 705222 128222 705458
rect 127986 669218 128222 669454
rect 127986 668898 128222 669134
rect 127986 633218 128222 633454
rect 127986 632898 128222 633134
rect 131586 672818 131822 673054
rect 131586 672498 131822 672734
rect 131586 636818 131822 637054
rect 131586 636498 131822 636734
rect 131586 600818 131822 601054
rect 131586 600498 131822 600734
rect 135186 676418 135422 676654
rect 135186 676098 135422 676334
rect 135186 640418 135422 640654
rect 135186 640098 135422 640334
rect 135186 604418 135422 604654
rect 135186 604098 135422 604334
rect 156786 710242 157022 710478
rect 156786 709922 157022 710158
rect 153186 708362 153422 708598
rect 153186 708042 153422 708278
rect 149586 706482 149822 706718
rect 149586 706162 149822 706398
rect 138786 680018 139022 680254
rect 138786 679698 139022 679934
rect 138786 644018 139022 644254
rect 138786 643698 139022 643934
rect 138786 608018 139022 608254
rect 138786 607698 139022 607934
rect 145986 704602 146222 704838
rect 145986 704282 146222 704518
rect 145986 687218 146222 687454
rect 145986 686898 146222 687134
rect 145986 651218 146222 651454
rect 145986 650898 146222 651134
rect 145986 615218 146222 615454
rect 145986 614898 146222 615134
rect 149586 690818 149822 691054
rect 149586 690498 149822 690734
rect 149586 654818 149822 655054
rect 149586 654498 149822 654734
rect 149586 618818 149822 619054
rect 149586 618498 149822 618734
rect 153186 694418 153422 694654
rect 153186 694098 153422 694334
rect 153186 658418 153422 658654
rect 153186 658098 153422 658334
rect 153186 622418 153422 622654
rect 153186 622098 153422 622334
rect 174786 711182 175022 711418
rect 174786 710862 175022 711098
rect 171186 709302 171422 709538
rect 171186 708982 171422 709218
rect 167586 707422 167822 707658
rect 167586 707102 167822 707338
rect 156786 698018 157022 698254
rect 156786 697698 157022 697934
rect 156786 662018 157022 662254
rect 156786 661698 157022 661934
rect 156786 626018 157022 626254
rect 156786 625698 157022 625934
rect 163986 705542 164222 705778
rect 163986 705222 164222 705458
rect 163986 669218 164222 669454
rect 163986 668898 164222 669134
rect 163986 633218 164222 633454
rect 163986 632898 164222 633134
rect 167586 672818 167822 673054
rect 167586 672498 167822 672734
rect 167586 636818 167822 637054
rect 167586 636498 167822 636734
rect 167586 600818 167822 601054
rect 167586 600498 167822 600734
rect 171186 676418 171422 676654
rect 171186 676098 171422 676334
rect 171186 640418 171422 640654
rect 171186 640098 171422 640334
rect 171186 604418 171422 604654
rect 171186 604098 171422 604334
rect 192786 710242 193022 710478
rect 192786 709922 193022 710158
rect 189186 708362 189422 708598
rect 189186 708042 189422 708278
rect 185586 706482 185822 706718
rect 185586 706162 185822 706398
rect 174786 680018 175022 680254
rect 174786 679698 175022 679934
rect 174786 644018 175022 644254
rect 174786 643698 175022 643934
rect 174786 608018 175022 608254
rect 174786 607698 175022 607934
rect 181986 704602 182222 704838
rect 181986 704282 182222 704518
rect 181986 687218 182222 687454
rect 181986 686898 182222 687134
rect 181986 651218 182222 651454
rect 181986 650898 182222 651134
rect 181986 615218 182222 615454
rect 181986 614898 182222 615134
rect 185586 690818 185822 691054
rect 185586 690498 185822 690734
rect 185586 654818 185822 655054
rect 185586 654498 185822 654734
rect 185586 618818 185822 619054
rect 185586 618498 185822 618734
rect 189186 694418 189422 694654
rect 189186 694098 189422 694334
rect 189186 658418 189422 658654
rect 189186 658098 189422 658334
rect 189186 622418 189422 622654
rect 189186 622098 189422 622334
rect 210786 711182 211022 711418
rect 210786 710862 211022 711098
rect 207186 709302 207422 709538
rect 207186 708982 207422 709218
rect 203586 707422 203822 707658
rect 203586 707102 203822 707338
rect 192786 698018 193022 698254
rect 192786 697698 193022 697934
rect 192786 662018 193022 662254
rect 192786 661698 193022 661934
rect 192786 626018 193022 626254
rect 192786 625698 193022 625934
rect 199986 705542 200222 705778
rect 199986 705222 200222 705458
rect 199986 669218 200222 669454
rect 199986 668898 200222 669134
rect 199986 633218 200222 633454
rect 199986 632898 200222 633134
rect 203586 672818 203822 673054
rect 203586 672498 203822 672734
rect 203586 636818 203822 637054
rect 203586 636498 203822 636734
rect 203586 600818 203822 601054
rect 203586 600498 203822 600734
rect 207186 676418 207422 676654
rect 207186 676098 207422 676334
rect 207186 640418 207422 640654
rect 207186 640098 207422 640334
rect 207186 604418 207422 604654
rect 207186 604098 207422 604334
rect 228786 710242 229022 710478
rect 228786 709922 229022 710158
rect 225186 708362 225422 708598
rect 225186 708042 225422 708278
rect 221586 706482 221822 706718
rect 221586 706162 221822 706398
rect 210786 680018 211022 680254
rect 210786 679698 211022 679934
rect 210786 644018 211022 644254
rect 210786 643698 211022 643934
rect 210786 608018 211022 608254
rect 210786 607698 211022 607934
rect 217986 704602 218222 704838
rect 217986 704282 218222 704518
rect 217986 687218 218222 687454
rect 217986 686898 218222 687134
rect 217986 651218 218222 651454
rect 217986 650898 218222 651134
rect 217986 615218 218222 615454
rect 217986 614898 218222 615134
rect 221586 690818 221822 691054
rect 221586 690498 221822 690734
rect 221586 654818 221822 655054
rect 221586 654498 221822 654734
rect 221586 618818 221822 619054
rect 221586 618498 221822 618734
rect 225186 694418 225422 694654
rect 225186 694098 225422 694334
rect 225186 658418 225422 658654
rect 225186 658098 225422 658334
rect 225186 622418 225422 622654
rect 225186 622098 225422 622334
rect 246786 711182 247022 711418
rect 246786 710862 247022 711098
rect 243186 709302 243422 709538
rect 243186 708982 243422 709218
rect 239586 707422 239822 707658
rect 239586 707102 239822 707338
rect 228786 698018 229022 698254
rect 228786 697698 229022 697934
rect 228786 662018 229022 662254
rect 228786 661698 229022 661934
rect 228786 626018 229022 626254
rect 228786 625698 229022 625934
rect 235986 705542 236222 705778
rect 235986 705222 236222 705458
rect 235986 669218 236222 669454
rect 235986 668898 236222 669134
rect 235986 633218 236222 633454
rect 235986 632898 236222 633134
rect 239586 672818 239822 673054
rect 239586 672498 239822 672734
rect 239586 636818 239822 637054
rect 239586 636498 239822 636734
rect 239586 600818 239822 601054
rect 239586 600498 239822 600734
rect 243186 676418 243422 676654
rect 243186 676098 243422 676334
rect 243186 640418 243422 640654
rect 243186 640098 243422 640334
rect 243186 604418 243422 604654
rect 243186 604098 243422 604334
rect 264786 710242 265022 710478
rect 264786 709922 265022 710158
rect 261186 708362 261422 708598
rect 261186 708042 261422 708278
rect 257586 706482 257822 706718
rect 257586 706162 257822 706398
rect 246786 680018 247022 680254
rect 246786 679698 247022 679934
rect 246786 644018 247022 644254
rect 246786 643698 247022 643934
rect 246786 608018 247022 608254
rect 246786 607698 247022 607934
rect 253986 704602 254222 704838
rect 253986 704282 254222 704518
rect 253986 687218 254222 687454
rect 253986 686898 254222 687134
rect 253986 651218 254222 651454
rect 253986 650898 254222 651134
rect 253986 615218 254222 615454
rect 253986 614898 254222 615134
rect 257586 690818 257822 691054
rect 257586 690498 257822 690734
rect 257586 654818 257822 655054
rect 257586 654498 257822 654734
rect 257586 618818 257822 619054
rect 257586 618498 257822 618734
rect 261186 694418 261422 694654
rect 261186 694098 261422 694334
rect 261186 658418 261422 658654
rect 261186 658098 261422 658334
rect 261186 622418 261422 622654
rect 261186 622098 261422 622334
rect 282786 711182 283022 711418
rect 282786 710862 283022 711098
rect 279186 709302 279422 709538
rect 279186 708982 279422 709218
rect 275586 707422 275822 707658
rect 275586 707102 275822 707338
rect 264786 698018 265022 698254
rect 264786 697698 265022 697934
rect 264786 662018 265022 662254
rect 264786 661698 265022 661934
rect 264786 626018 265022 626254
rect 264786 625698 265022 625934
rect 271986 705542 272222 705778
rect 271986 705222 272222 705458
rect 271986 669218 272222 669454
rect 271986 668898 272222 669134
rect 271986 633218 272222 633454
rect 271986 632898 272222 633134
rect 275586 672818 275822 673054
rect 275586 672498 275822 672734
rect 275586 636818 275822 637054
rect 275586 636498 275822 636734
rect 275586 600818 275822 601054
rect 275586 600498 275822 600734
rect 279186 676418 279422 676654
rect 279186 676098 279422 676334
rect 279186 640418 279422 640654
rect 279186 640098 279422 640334
rect 279186 604418 279422 604654
rect 279186 604098 279422 604334
rect 300786 710242 301022 710478
rect 300786 709922 301022 710158
rect 297186 708362 297422 708598
rect 297186 708042 297422 708278
rect 293586 706482 293822 706718
rect 293586 706162 293822 706398
rect 282786 680018 283022 680254
rect 282786 679698 283022 679934
rect 282786 644018 283022 644254
rect 282786 643698 283022 643934
rect 282786 608018 283022 608254
rect 282786 607698 283022 607934
rect 289986 704602 290222 704838
rect 289986 704282 290222 704518
rect 289986 687218 290222 687454
rect 289986 686898 290222 687134
rect 289986 651218 290222 651454
rect 289986 650898 290222 651134
rect 289986 615218 290222 615454
rect 289986 614898 290222 615134
rect 293586 690818 293822 691054
rect 293586 690498 293822 690734
rect 293586 654818 293822 655054
rect 293586 654498 293822 654734
rect 293586 618818 293822 619054
rect 293586 618498 293822 618734
rect 297186 694418 297422 694654
rect 297186 694098 297422 694334
rect 297186 658418 297422 658654
rect 297186 658098 297422 658334
rect 297186 622418 297422 622654
rect 297186 622098 297422 622334
rect 318786 711182 319022 711418
rect 318786 710862 319022 711098
rect 315186 709302 315422 709538
rect 315186 708982 315422 709218
rect 311586 707422 311822 707658
rect 311586 707102 311822 707338
rect 300786 698018 301022 698254
rect 300786 697698 301022 697934
rect 300786 662018 301022 662254
rect 300786 661698 301022 661934
rect 300786 626018 301022 626254
rect 300786 625698 301022 625934
rect 307986 705542 308222 705778
rect 307986 705222 308222 705458
rect 307986 669218 308222 669454
rect 307986 668898 308222 669134
rect 307986 633218 308222 633454
rect 307986 632898 308222 633134
rect 311586 672818 311822 673054
rect 311586 672498 311822 672734
rect 311586 636818 311822 637054
rect 311586 636498 311822 636734
rect 311586 600818 311822 601054
rect 311586 600498 311822 600734
rect 315186 676418 315422 676654
rect 315186 676098 315422 676334
rect 315186 640418 315422 640654
rect 315186 640098 315422 640334
rect 315186 604418 315422 604654
rect 315186 604098 315422 604334
rect 336786 710242 337022 710478
rect 336786 709922 337022 710158
rect 333186 708362 333422 708598
rect 333186 708042 333422 708278
rect 329586 706482 329822 706718
rect 329586 706162 329822 706398
rect 318786 680018 319022 680254
rect 318786 679698 319022 679934
rect 318786 644018 319022 644254
rect 318786 643698 319022 643934
rect 318786 608018 319022 608254
rect 318786 607698 319022 607934
rect 325986 704602 326222 704838
rect 325986 704282 326222 704518
rect 325986 687218 326222 687454
rect 325986 686898 326222 687134
rect 325986 651218 326222 651454
rect 325986 650898 326222 651134
rect 325986 615218 326222 615454
rect 325986 614898 326222 615134
rect 329586 690818 329822 691054
rect 329586 690498 329822 690734
rect 329586 654818 329822 655054
rect 329586 654498 329822 654734
rect 329586 618818 329822 619054
rect 329586 618498 329822 618734
rect 333186 694418 333422 694654
rect 333186 694098 333422 694334
rect 333186 658418 333422 658654
rect 333186 658098 333422 658334
rect 333186 622418 333422 622654
rect 333186 622098 333422 622334
rect 354786 711182 355022 711418
rect 354786 710862 355022 711098
rect 351186 709302 351422 709538
rect 351186 708982 351422 709218
rect 347586 707422 347822 707658
rect 347586 707102 347822 707338
rect 336786 698018 337022 698254
rect 336786 697698 337022 697934
rect 336786 662018 337022 662254
rect 336786 661698 337022 661934
rect 336786 626018 337022 626254
rect 336786 625698 337022 625934
rect 343986 705542 344222 705778
rect 343986 705222 344222 705458
rect 343986 669218 344222 669454
rect 343986 668898 344222 669134
rect 343986 633218 344222 633454
rect 343986 632898 344222 633134
rect 347586 672818 347822 673054
rect 347586 672498 347822 672734
rect 347586 636818 347822 637054
rect 347586 636498 347822 636734
rect 347586 600818 347822 601054
rect 347586 600498 347822 600734
rect 351186 676418 351422 676654
rect 351186 676098 351422 676334
rect 351186 640418 351422 640654
rect 351186 640098 351422 640334
rect 351186 604418 351422 604654
rect 351186 604098 351422 604334
rect 372786 710242 373022 710478
rect 372786 709922 373022 710158
rect 369186 708362 369422 708598
rect 369186 708042 369422 708278
rect 365586 706482 365822 706718
rect 365586 706162 365822 706398
rect 354786 680018 355022 680254
rect 354786 679698 355022 679934
rect 354786 644018 355022 644254
rect 354786 643698 355022 643934
rect 354786 608018 355022 608254
rect 354786 607698 355022 607934
rect 361986 704602 362222 704838
rect 361986 704282 362222 704518
rect 361986 687218 362222 687454
rect 361986 686898 362222 687134
rect 361986 651218 362222 651454
rect 361986 650898 362222 651134
rect 361986 615218 362222 615454
rect 361986 614898 362222 615134
rect 365586 690818 365822 691054
rect 365586 690498 365822 690734
rect 365586 654818 365822 655054
rect 365586 654498 365822 654734
rect 365586 618818 365822 619054
rect 365586 618498 365822 618734
rect 369186 694418 369422 694654
rect 369186 694098 369422 694334
rect 369186 658418 369422 658654
rect 369186 658098 369422 658334
rect 369186 622418 369422 622654
rect 369186 622098 369422 622334
rect 390786 711182 391022 711418
rect 390786 710862 391022 711098
rect 387186 709302 387422 709538
rect 387186 708982 387422 709218
rect 383586 707422 383822 707658
rect 383586 707102 383822 707338
rect 372786 698018 373022 698254
rect 372786 697698 373022 697934
rect 372786 662018 373022 662254
rect 372786 661698 373022 661934
rect 372786 626018 373022 626254
rect 372786 625698 373022 625934
rect 379986 705542 380222 705778
rect 379986 705222 380222 705458
rect 379986 669218 380222 669454
rect 379986 668898 380222 669134
rect 379986 633218 380222 633454
rect 379986 632898 380222 633134
rect 383586 672818 383822 673054
rect 383586 672498 383822 672734
rect 383586 636818 383822 637054
rect 383586 636498 383822 636734
rect 383586 600818 383822 601054
rect 383586 600498 383822 600734
rect 387186 676418 387422 676654
rect 387186 676098 387422 676334
rect 387186 640418 387422 640654
rect 387186 640098 387422 640334
rect 387186 604418 387422 604654
rect 387186 604098 387422 604334
rect 408786 710242 409022 710478
rect 408786 709922 409022 710158
rect 405186 708362 405422 708598
rect 405186 708042 405422 708278
rect 401586 706482 401822 706718
rect 401586 706162 401822 706398
rect 390786 680018 391022 680254
rect 390786 679698 391022 679934
rect 390786 644018 391022 644254
rect 390786 643698 391022 643934
rect 390786 608018 391022 608254
rect 390786 607698 391022 607934
rect 397986 704602 398222 704838
rect 397986 704282 398222 704518
rect 397986 687218 398222 687454
rect 397986 686898 398222 687134
rect 397986 651218 398222 651454
rect 397986 650898 398222 651134
rect 397986 615218 398222 615454
rect 397986 614898 398222 615134
rect 401586 690818 401822 691054
rect 401586 690498 401822 690734
rect 401586 654818 401822 655054
rect 401586 654498 401822 654734
rect 401586 618818 401822 619054
rect 401586 618498 401822 618734
rect 405186 694418 405422 694654
rect 405186 694098 405422 694334
rect 405186 658418 405422 658654
rect 405186 658098 405422 658334
rect 405186 622418 405422 622654
rect 405186 622098 405422 622334
rect 426786 711182 427022 711418
rect 426786 710862 427022 711098
rect 423186 709302 423422 709538
rect 423186 708982 423422 709218
rect 419586 707422 419822 707658
rect 419586 707102 419822 707338
rect 408786 698018 409022 698254
rect 408786 697698 409022 697934
rect 408786 662018 409022 662254
rect 408786 661698 409022 661934
rect 408786 626018 409022 626254
rect 408786 625698 409022 625934
rect 415986 705542 416222 705778
rect 415986 705222 416222 705458
rect 415986 669218 416222 669454
rect 415986 668898 416222 669134
rect 415986 633218 416222 633454
rect 415986 632898 416222 633134
rect 419586 672818 419822 673054
rect 419586 672498 419822 672734
rect 419586 636818 419822 637054
rect 419586 636498 419822 636734
rect 419586 600818 419822 601054
rect 419586 600498 419822 600734
rect 423186 676418 423422 676654
rect 423186 676098 423422 676334
rect 423186 640418 423422 640654
rect 423186 640098 423422 640334
rect 423186 604418 423422 604654
rect 423186 604098 423422 604334
rect 444786 710242 445022 710478
rect 444786 709922 445022 710158
rect 441186 708362 441422 708598
rect 441186 708042 441422 708278
rect 437586 706482 437822 706718
rect 437586 706162 437822 706398
rect 426786 680018 427022 680254
rect 426786 679698 427022 679934
rect 426786 644018 427022 644254
rect 426786 643698 427022 643934
rect 426786 608018 427022 608254
rect 426786 607698 427022 607934
rect 433986 704602 434222 704838
rect 433986 704282 434222 704518
rect 433986 687218 434222 687454
rect 433986 686898 434222 687134
rect 433986 651218 434222 651454
rect 433986 650898 434222 651134
rect 433986 615218 434222 615454
rect 433986 614898 434222 615134
rect 437586 690818 437822 691054
rect 437586 690498 437822 690734
rect 437586 654818 437822 655054
rect 437586 654498 437822 654734
rect 437586 618818 437822 619054
rect 437586 618498 437822 618734
rect 441186 694418 441422 694654
rect 441186 694098 441422 694334
rect 441186 658418 441422 658654
rect 441186 658098 441422 658334
rect 441186 622418 441422 622654
rect 441186 622098 441422 622334
rect 462786 711182 463022 711418
rect 462786 710862 463022 711098
rect 459186 709302 459422 709538
rect 459186 708982 459422 709218
rect 455586 707422 455822 707658
rect 455586 707102 455822 707338
rect 444786 698018 445022 698254
rect 444786 697698 445022 697934
rect 444786 662018 445022 662254
rect 444786 661698 445022 661934
rect 444786 626018 445022 626254
rect 444786 625698 445022 625934
rect 451986 705542 452222 705778
rect 451986 705222 452222 705458
rect 451986 669218 452222 669454
rect 451986 668898 452222 669134
rect 451986 633218 452222 633454
rect 451986 632898 452222 633134
rect 451986 597218 452222 597454
rect 451986 596898 452222 597134
rect 102786 572018 103022 572254
rect 102786 571698 103022 571934
rect 102786 536018 103022 536254
rect 102786 535698 103022 535934
rect 102786 500018 103022 500254
rect 102786 499698 103022 499934
rect 102786 464018 103022 464254
rect 102786 463698 103022 463934
rect 102786 428018 103022 428254
rect 102786 427698 103022 427934
rect 102786 392018 103022 392254
rect 102786 391698 103022 391934
rect 102786 356018 103022 356254
rect 102786 355698 103022 355934
rect 102786 320018 103022 320254
rect 102786 319698 103022 319934
rect 102786 284018 103022 284254
rect 102786 283698 103022 283934
rect 102786 248018 103022 248254
rect 102786 247698 103022 247934
rect 123186 582663 123422 582899
rect 123581 582677 123817 582913
rect 123901 582677 124137 582913
rect 124275 582677 124511 582913
rect 124595 582677 124831 582913
rect 124982 582692 125218 582928
rect 125302 582692 125538 582928
rect 125676 582692 125912 582928
rect 125996 582692 126232 582928
rect 126391 582706 126627 582942
rect 126711 582706 126947 582942
rect 127085 582706 127321 582942
rect 127405 582706 127641 582942
rect 127871 582721 128107 582957
rect 128191 582721 128427 582957
rect 128565 582721 128801 582957
rect 128885 582721 129121 582957
rect 129280 582735 129516 582971
rect 129600 582735 129836 582971
rect 129974 582735 130210 582971
rect 130294 582735 130530 582971
rect 130681 582750 130917 582986
rect 131001 582750 131237 582986
rect 131375 582750 131611 582986
rect 131695 582750 131931 582986
rect 132090 582764 132326 583000
rect 132410 582764 132646 583000
rect 132784 582764 133020 583000
rect 133104 582764 133340 583000
rect 123273 546639 123509 546875
rect 123668 546653 123904 546889
rect 123988 546653 124224 546889
rect 124362 546653 124598 546889
rect 124682 546653 124918 546889
rect 125069 546668 125305 546904
rect 125389 546668 125625 546904
rect 125763 546668 125999 546904
rect 126083 546668 126319 546904
rect 126478 546682 126714 546918
rect 126798 546682 127034 546918
rect 127172 546682 127408 546918
rect 127492 546682 127728 546918
rect 127958 546697 128194 546933
rect 128278 546697 128514 546933
rect 128652 546697 128888 546933
rect 128972 546697 129208 546933
rect 129367 546711 129603 546947
rect 129687 546711 129923 546947
rect 130061 546711 130297 546947
rect 130381 546711 130617 546947
rect 130768 546726 131004 546962
rect 131088 546726 131324 546962
rect 131462 546726 131698 546962
rect 131782 546726 132018 546962
rect 132177 546740 132413 546976
rect 132497 546740 132733 546976
rect 132871 546740 133107 546976
rect 133191 546740 133427 546976
rect 123233 510636 123469 510872
rect 123628 510650 123864 510886
rect 123948 510650 124184 510886
rect 124322 510650 124558 510886
rect 124642 510650 124878 510886
rect 125029 510665 125265 510901
rect 125349 510665 125585 510901
rect 125723 510665 125959 510901
rect 126043 510665 126279 510901
rect 126438 510679 126674 510915
rect 126758 510679 126994 510915
rect 127132 510679 127368 510915
rect 127452 510679 127688 510915
rect 127918 510694 128154 510930
rect 128238 510694 128474 510930
rect 128612 510694 128848 510930
rect 128932 510694 129168 510930
rect 129327 510708 129563 510944
rect 129647 510708 129883 510944
rect 130021 510708 130257 510944
rect 130341 510708 130577 510944
rect 130728 510723 130964 510959
rect 131048 510723 131284 510959
rect 131422 510723 131658 510959
rect 131742 510723 131978 510959
rect 132137 510737 132373 510973
rect 132457 510737 132693 510973
rect 132831 510737 133067 510973
rect 133151 510737 133387 510973
rect 123412 473270 123648 473506
rect 123412 472950 123648 473186
rect 123412 472630 123648 472866
rect 123807 472644 124363 473520
rect 124501 472644 125057 473520
rect 125208 472659 125764 473535
rect 125902 472659 126458 473535
rect 126617 472673 127173 473549
rect 127311 472673 127867 473549
rect 128097 472688 128653 473564
rect 128791 472688 129347 473564
rect 129506 472702 130062 473578
rect 130200 472702 130756 473578
rect 130907 472717 131463 473593
rect 131601 472717 132157 473593
rect 132316 472731 132872 473607
rect 133010 472731 133566 473607
rect 123477 465284 123713 465520
rect 123477 464964 123713 465200
rect 123477 464644 123713 464880
rect 123872 464658 124428 465534
rect 124566 464658 125122 465534
rect 125273 464673 125829 465549
rect 125967 464673 126523 465549
rect 126682 464687 127238 465563
rect 127376 464687 127932 465563
rect 128162 464702 128718 465578
rect 128856 464702 129412 465578
rect 129571 464716 130127 465592
rect 130265 464716 130821 465592
rect 130972 464731 131528 465607
rect 131666 464731 132222 465607
rect 132381 464745 132937 465621
rect 133075 464745 133631 465621
rect 123337 457338 123573 457574
rect 123337 457018 123573 457254
rect 123337 456698 123573 456934
rect 123732 456712 124288 457588
rect 124426 456712 124982 457588
rect 125133 456727 125689 457603
rect 125827 456727 126383 457603
rect 126542 456741 127098 457617
rect 127236 456741 127792 457617
rect 128022 456756 128578 457632
rect 128716 456756 129272 457632
rect 129431 456770 129987 457646
rect 130125 456770 130681 457646
rect 130832 456785 131388 457661
rect 131526 456785 132082 457661
rect 132241 456799 132797 457675
rect 132935 456799 133491 457675
rect 123392 449305 123628 449541
rect 123392 448985 123628 449221
rect 123392 448665 123628 448901
rect 123787 448679 124343 449555
rect 124481 448679 125037 449555
rect 125188 448694 125744 449570
rect 125882 448694 126438 449570
rect 126597 448708 127153 449584
rect 127291 448708 127847 449584
rect 128077 448723 128633 449599
rect 128771 448723 129327 449599
rect 129486 448737 130042 449613
rect 130180 448737 130736 449613
rect 130887 448752 131443 449628
rect 131581 448752 132137 449628
rect 132296 448766 132852 449642
rect 132990 448766 133546 449642
rect 123506 441317 123742 441553
rect 123506 440997 123742 441233
rect 123506 440677 123742 440913
rect 123901 440691 124457 441567
rect 124595 440691 125151 441567
rect 125302 440706 125858 441582
rect 125996 440706 126552 441582
rect 126711 440720 127267 441596
rect 127405 440720 127961 441596
rect 128191 440735 128747 441611
rect 128885 440735 129441 441611
rect 129600 440749 130156 441625
rect 130294 440749 130850 441625
rect 131001 440764 131557 441640
rect 131695 440764 132251 441640
rect 132410 440778 132966 441654
rect 133104 440778 133660 441654
rect 123436 433272 123672 433508
rect 123436 432952 123672 433188
rect 123436 432632 123672 432868
rect 123831 432646 124387 433522
rect 124525 432646 125081 433522
rect 125232 432661 125788 433537
rect 125926 432661 126482 433537
rect 126641 432675 127197 433551
rect 127335 432675 127891 433551
rect 128121 432690 128677 433566
rect 128815 432690 129371 433566
rect 129530 432704 130086 433580
rect 130224 432704 130780 433580
rect 130931 432719 131487 433595
rect 131625 432719 132181 433595
rect 132340 432733 132896 433609
rect 133034 432733 133590 433609
rect 123438 425328 123674 425564
rect 123438 425008 123674 425244
rect 123438 424688 123674 424924
rect 123833 424702 124389 425578
rect 124527 424702 125083 425578
rect 125234 424717 125790 425593
rect 125928 424717 126484 425593
rect 126643 424731 127199 425607
rect 127337 424731 127893 425607
rect 128123 424746 128679 425622
rect 128817 424746 129373 425622
rect 129532 424760 130088 425636
rect 130226 424760 130782 425636
rect 130933 424775 131489 425651
rect 131627 424775 132183 425651
rect 132342 424789 132898 425665
rect 133036 424789 133592 425665
rect 123409 417269 123645 417505
rect 123409 416949 123645 417185
rect 123409 416629 123645 416865
rect 123804 416643 124360 417519
rect 124498 416643 125054 417519
rect 125205 416658 125761 417534
rect 125899 416658 126455 417534
rect 126614 416672 127170 417548
rect 127308 416672 127864 417548
rect 128094 416687 128650 417563
rect 128788 416687 129344 417563
rect 129503 416701 130059 417577
rect 130197 416701 130753 417577
rect 130904 416716 131460 417592
rect 131598 416716 132154 417592
rect 132313 416730 132869 417606
rect 133007 416730 133563 417606
rect 123496 409301 123732 409537
rect 123496 408981 123732 409217
rect 123496 408661 123732 408897
rect 123891 408675 124447 409551
rect 124585 408675 125141 409551
rect 125292 408690 125848 409566
rect 125986 408690 126542 409566
rect 126701 408704 127257 409580
rect 127395 408704 127951 409580
rect 128181 408719 128737 409595
rect 128875 408719 129431 409595
rect 129590 408733 130146 409609
rect 130284 408733 130840 409609
rect 130991 408748 131547 409624
rect 131685 408748 132241 409624
rect 132400 408762 132956 409638
rect 133094 408762 133650 409638
rect 123430 401303 123666 401539
rect 123430 400983 123666 401219
rect 123430 400663 123666 400899
rect 123825 400677 124381 401553
rect 124519 400677 125075 401553
rect 125226 400692 125782 401568
rect 125920 400692 126476 401568
rect 126635 400706 127191 401582
rect 127329 400706 127885 401582
rect 128115 400721 128671 401597
rect 128809 400721 129365 401597
rect 129524 400735 130080 401611
rect 130218 400735 130774 401611
rect 130925 400750 131481 401626
rect 131619 400750 132175 401626
rect 132334 400764 132890 401640
rect 133028 400764 133584 401640
rect 123400 393303 123636 393539
rect 123400 392983 123636 393219
rect 123400 392663 123636 392899
rect 123795 392677 124351 393553
rect 124489 392677 125045 393553
rect 125196 392692 125752 393568
rect 125890 392692 126446 393568
rect 126605 392706 127161 393582
rect 127299 392706 127855 393582
rect 128085 392721 128641 393597
rect 128779 392721 129335 393597
rect 129494 392735 130050 393611
rect 130188 392735 130744 393611
rect 130895 392750 131451 393626
rect 131589 392750 132145 393626
rect 132304 392764 132860 393640
rect 132998 392764 133554 393640
rect 123481 385275 123717 385511
rect 123481 384955 123717 385191
rect 123481 384635 123717 384871
rect 123876 384649 124432 385525
rect 124570 384649 125126 385525
rect 125277 384664 125833 385540
rect 125971 384664 126527 385540
rect 126686 384678 127242 385554
rect 127380 384678 127936 385554
rect 128166 384693 128722 385569
rect 128860 384693 129416 385569
rect 129575 384707 130131 385583
rect 130269 384707 130825 385583
rect 130976 384722 131532 385598
rect 131670 384722 132226 385598
rect 132385 384736 132941 385612
rect 133079 384736 133635 385612
rect 123413 377317 123649 377553
rect 123413 376997 123649 377233
rect 123413 376677 123649 376913
rect 123808 376691 124364 377567
rect 124502 376691 125058 377567
rect 125209 376706 125765 377582
rect 125903 376706 126459 377582
rect 126618 376720 127174 377596
rect 127312 376720 127868 377596
rect 128098 376735 128654 377611
rect 128792 376735 129348 377611
rect 129507 376749 130063 377625
rect 130201 376749 130757 377625
rect 130908 376764 131464 377640
rect 131602 376764 132158 377640
rect 132317 376778 132873 377654
rect 133011 376778 133567 377654
rect 123342 369255 123578 369491
rect 123342 368935 123578 369171
rect 123342 368615 123578 368851
rect 123737 368629 124293 369505
rect 124431 368629 124987 369505
rect 125138 368644 125694 369520
rect 125832 368644 126388 369520
rect 126547 368658 127103 369534
rect 127241 368658 127797 369534
rect 128027 368673 128583 369549
rect 128721 368673 129277 369549
rect 129436 368687 129992 369563
rect 130130 368687 130686 369563
rect 130837 368702 131393 369578
rect 131531 368702 132087 369578
rect 132246 368716 132802 369592
rect 132940 368716 133496 369592
rect 123481 361303 123717 361539
rect 123481 360983 123717 361219
rect 123481 360663 123717 360899
rect 123876 360677 124432 361553
rect 124570 360677 125126 361553
rect 125277 360692 125833 361568
rect 125971 360692 126527 361568
rect 126686 360706 127242 361582
rect 127380 360706 127936 361582
rect 128166 360721 128722 361597
rect 128860 360721 129416 361597
rect 129575 360735 130131 361611
rect 130269 360735 130825 361611
rect 130976 360750 131532 361626
rect 131670 360750 132226 361626
rect 132385 360764 132941 361640
rect 133079 360764 133635 361640
rect 123410 353277 123646 353513
rect 123410 352957 123646 353193
rect 123410 352637 123646 352873
rect 123805 352651 124361 353527
rect 124499 352651 125055 353527
rect 125206 352666 125762 353542
rect 125900 352666 126456 353542
rect 126615 352680 127171 353556
rect 127309 352680 127865 353556
rect 128095 352695 128651 353571
rect 128789 352695 129345 353571
rect 129504 352709 130060 353585
rect 130198 352709 130754 353585
rect 130905 352724 131461 353600
rect 131599 352724 132155 353600
rect 132314 352738 132870 353614
rect 133008 352738 133564 353614
rect 123512 345297 123748 345533
rect 123512 344977 123748 345213
rect 123512 344657 123748 344893
rect 123907 344671 124463 345547
rect 124601 344671 125157 345547
rect 125308 344686 125864 345562
rect 126002 344686 126558 345562
rect 126717 344700 127273 345576
rect 127411 344700 127967 345576
rect 128197 344715 128753 345591
rect 128891 344715 129447 345591
rect 129606 344729 130162 345605
rect 130300 344729 130856 345605
rect 131007 344744 131563 345620
rect 131701 344744 132257 345620
rect 132416 344758 132972 345634
rect 133110 344758 133666 345634
rect 123455 330610 123691 330846
rect 123850 330624 124086 330860
rect 124170 330624 124406 330860
rect 124544 330624 124780 330860
rect 124864 330624 125100 330860
rect 125251 330639 125487 330875
rect 125571 330639 125807 330875
rect 125945 330639 126181 330875
rect 126265 330639 126501 330875
rect 126660 330653 126896 330889
rect 126980 330653 127216 330889
rect 127354 330653 127590 330889
rect 127674 330653 127910 330889
rect 128140 330668 128376 330904
rect 128460 330668 128696 330904
rect 128834 330668 129070 330904
rect 129154 330668 129390 330904
rect 129549 330682 129785 330918
rect 129869 330682 130105 330918
rect 130243 330682 130479 330918
rect 130563 330682 130799 330918
rect 130950 330697 131186 330933
rect 131270 330697 131506 330933
rect 131644 330697 131880 330933
rect 131964 330697 132200 330933
rect 132359 330711 132595 330947
rect 132679 330711 132915 330947
rect 133053 330711 133289 330947
rect 133373 330711 133609 330947
rect 123472 294607 123708 294843
rect 123867 294621 124103 294857
rect 124187 294621 124423 294857
rect 124561 294621 124797 294857
rect 124881 294621 125117 294857
rect 125268 294636 125504 294872
rect 125588 294636 125824 294872
rect 125962 294636 126198 294872
rect 126282 294636 126518 294872
rect 126677 294650 126913 294886
rect 126997 294650 127233 294886
rect 127371 294650 127607 294886
rect 127691 294650 127927 294886
rect 128157 294665 128393 294901
rect 128477 294665 128713 294901
rect 128851 294665 129087 294901
rect 129171 294665 129407 294901
rect 129566 294679 129802 294915
rect 129886 294679 130122 294915
rect 130260 294679 130496 294915
rect 130580 294679 130816 294915
rect 130967 294694 131203 294930
rect 131287 294694 131523 294930
rect 131661 294694 131897 294930
rect 131981 294694 132217 294930
rect 132376 294708 132612 294944
rect 132696 294708 132932 294944
rect 133070 294708 133306 294944
rect 133390 294708 133626 294944
rect 123238 258607 123474 258843
rect 123633 258621 123869 258857
rect 123953 258621 124189 258857
rect 124327 258621 124563 258857
rect 124647 258621 124883 258857
rect 125034 258636 125270 258872
rect 125354 258636 125590 258872
rect 125728 258636 125964 258872
rect 126048 258636 126284 258872
rect 126443 258650 126679 258886
rect 126763 258650 126999 258886
rect 127137 258650 127373 258886
rect 127457 258650 127693 258886
rect 127923 258665 128159 258901
rect 128243 258665 128479 258901
rect 128617 258665 128853 258901
rect 128937 258665 129173 258901
rect 129332 258679 129568 258915
rect 129652 258679 129888 258915
rect 130026 258679 130262 258915
rect 130346 258679 130582 258915
rect 130733 258694 130969 258930
rect 131053 258694 131289 258930
rect 131427 258694 131663 258930
rect 131747 258694 131983 258930
rect 132142 258708 132378 258944
rect 132462 258708 132698 258944
rect 132836 258708 133072 258944
rect 133156 258708 133392 258944
rect 140937 579057 141173 579293
rect 141332 579071 141568 579307
rect 141652 579071 141888 579307
rect 142026 579071 142262 579307
rect 142346 579071 142582 579307
rect 142733 579086 142969 579322
rect 143053 579086 143289 579322
rect 143427 579086 143663 579322
rect 143747 579086 143983 579322
rect 144142 579100 144378 579336
rect 144462 579100 144698 579336
rect 144836 579100 145072 579336
rect 145156 579100 145392 579336
rect 145622 579115 145858 579351
rect 145942 579115 146178 579351
rect 146316 579115 146552 579351
rect 146636 579115 146872 579351
rect 147031 579129 147267 579365
rect 147351 579129 147587 579365
rect 147725 579129 147961 579365
rect 148045 579129 148281 579365
rect 148432 579144 148668 579380
rect 148752 579144 148988 579380
rect 149126 579144 149362 579380
rect 149446 579144 149682 579380
rect 149841 579158 150077 579394
rect 150161 579158 150397 579394
rect 150535 579158 150771 579394
rect 150855 579158 151091 579394
rect 141064 543036 141300 543272
rect 141459 543050 141695 543286
rect 141779 543050 142015 543286
rect 142153 543050 142389 543286
rect 142473 543050 142709 543286
rect 142860 543065 143096 543301
rect 143180 543065 143416 543301
rect 143554 543065 143790 543301
rect 143874 543065 144110 543301
rect 144269 543079 144505 543315
rect 144589 543079 144825 543315
rect 144963 543079 145199 543315
rect 145283 543079 145519 543315
rect 145749 543094 145985 543330
rect 146069 543094 146305 543330
rect 146443 543094 146679 543330
rect 146763 543094 146999 543330
rect 147158 543108 147394 543344
rect 147478 543108 147714 543344
rect 147852 543108 148088 543344
rect 148172 543108 148408 543344
rect 148559 543123 148795 543359
rect 148879 543123 149115 543359
rect 149253 543123 149489 543359
rect 149573 543123 149809 543359
rect 149968 543137 150204 543373
rect 150288 543137 150524 543373
rect 150662 543137 150898 543373
rect 150982 543137 151218 543373
rect 141248 507069 141484 507305
rect 141643 507083 141879 507319
rect 141963 507083 142199 507319
rect 142337 507083 142573 507319
rect 142657 507083 142893 507319
rect 143044 507098 143280 507334
rect 143364 507098 143600 507334
rect 143738 507098 143974 507334
rect 144058 507098 144294 507334
rect 144453 507112 144689 507348
rect 144773 507112 145009 507348
rect 145147 507112 145383 507348
rect 145467 507112 145703 507348
rect 145933 507127 146169 507363
rect 146253 507127 146489 507363
rect 146627 507127 146863 507363
rect 146947 507127 147183 507363
rect 147342 507141 147578 507377
rect 147662 507141 147898 507377
rect 148036 507141 148272 507377
rect 148356 507141 148592 507377
rect 148743 507156 148979 507392
rect 149063 507156 149299 507392
rect 149437 507156 149673 507392
rect 149757 507156 149993 507392
rect 150152 507170 150388 507406
rect 150472 507170 150708 507406
rect 150846 507170 151082 507406
rect 151166 507170 151402 507406
rect 141065 471572 141301 471808
rect 141065 471252 141301 471488
rect 141065 470932 141301 471168
rect 141460 470946 142016 471822
rect 142154 470946 142710 471822
rect 142861 470961 143417 471837
rect 143555 470961 144111 471837
rect 144270 470975 144826 471851
rect 144964 470975 145520 471851
rect 145750 470990 146306 471866
rect 146444 470990 147000 471866
rect 147159 471004 147715 471880
rect 147853 471004 148409 471880
rect 148560 471019 149116 471895
rect 149254 471019 149810 471895
rect 149969 471033 150525 471909
rect 150663 471033 151219 471909
rect 140945 463615 141181 463851
rect 140945 463295 141181 463531
rect 140945 462975 141181 463211
rect 141340 462989 141896 463865
rect 142034 462989 142590 463865
rect 142741 463004 143297 463880
rect 143435 463004 143991 463880
rect 144150 463018 144706 463894
rect 144844 463018 145400 463894
rect 145630 463033 146186 463909
rect 146324 463033 146880 463909
rect 147039 463047 147595 463923
rect 147733 463047 148289 463923
rect 148440 463062 148996 463938
rect 149134 463062 149690 463938
rect 149849 463076 150405 463952
rect 150543 463076 151099 463952
rect 141056 455655 141292 455891
rect 141056 455335 141292 455571
rect 141056 455015 141292 455251
rect 141451 455029 142007 455905
rect 142145 455029 142701 455905
rect 142852 455044 143408 455920
rect 143546 455044 144102 455920
rect 144261 455058 144817 455934
rect 144955 455058 145511 455934
rect 145741 455073 146297 455949
rect 146435 455073 146991 455949
rect 147150 455087 147706 455963
rect 147844 455087 148400 455963
rect 148551 455102 149107 455978
rect 149245 455102 149801 455978
rect 149960 455116 150516 455992
rect 150654 455116 151210 455992
rect 141129 447649 141365 447885
rect 141129 447329 141365 447565
rect 141129 447009 141365 447245
rect 141524 447023 142080 447899
rect 142218 447023 142774 447899
rect 142925 447038 143481 447914
rect 143619 447038 144175 447914
rect 144334 447052 144890 447928
rect 145028 447052 145584 447928
rect 145814 447067 146370 447943
rect 146508 447067 147064 447943
rect 147223 447081 147779 447957
rect 147917 447081 148473 447957
rect 148624 447096 149180 447972
rect 149318 447096 149874 447972
rect 150033 447110 150589 447986
rect 150727 447110 151283 447986
rect 141102 439692 141338 439928
rect 141102 439372 141338 439608
rect 141102 439052 141338 439288
rect 141497 439066 142053 439942
rect 142191 439066 142747 439942
rect 142898 439081 143454 439957
rect 143592 439081 144148 439957
rect 144307 439095 144863 439971
rect 145001 439095 145557 439971
rect 145787 439110 146343 439986
rect 146481 439110 147037 439986
rect 147196 439124 147752 440000
rect 147890 439124 148446 440000
rect 148597 439139 149153 440015
rect 149291 439139 149847 440015
rect 150006 439153 150562 440029
rect 150700 439153 151256 440029
rect 141073 431602 141309 431838
rect 141073 431282 141309 431518
rect 141073 430962 141309 431198
rect 141468 430976 142024 431852
rect 142162 430976 142718 431852
rect 142869 430991 143425 431867
rect 143563 430991 144119 431867
rect 144278 431005 144834 431881
rect 144972 431005 145528 431881
rect 145758 431020 146314 431896
rect 146452 431020 147008 431896
rect 147167 431034 147723 431910
rect 147861 431034 148417 431910
rect 148568 431049 149124 431925
rect 149262 431049 149818 431925
rect 149977 431063 150533 431939
rect 150671 431063 151227 431939
rect 141100 423625 141336 423861
rect 141100 423305 141336 423541
rect 141100 422985 141336 423221
rect 141495 422999 142051 423875
rect 142189 422999 142745 423875
rect 142896 423014 143452 423890
rect 143590 423014 144146 423890
rect 144305 423028 144861 423904
rect 144999 423028 145555 423904
rect 145785 423043 146341 423919
rect 146479 423043 147035 423919
rect 147194 423057 147750 423933
rect 147888 423057 148444 423933
rect 148595 423072 149151 423948
rect 149289 423072 149845 423948
rect 150004 423086 150560 423962
rect 150698 423086 151254 423962
rect 141035 415677 141271 415913
rect 141035 415357 141271 415593
rect 141035 415037 141271 415273
rect 141430 415051 141986 415927
rect 142124 415051 142680 415927
rect 142831 415066 143387 415942
rect 143525 415066 144081 415942
rect 144240 415080 144796 415956
rect 144934 415080 145490 415956
rect 145720 415095 146276 415971
rect 146414 415095 146970 415971
rect 147129 415109 147685 415985
rect 147823 415109 148379 415985
rect 148530 415124 149086 416000
rect 149224 415124 149780 416000
rect 149939 415138 150495 416014
rect 150633 415138 151189 416014
rect 140958 407614 141194 407850
rect 140958 407294 141194 407530
rect 140958 406974 141194 407210
rect 141353 406988 141909 407864
rect 142047 406988 142603 407864
rect 142754 407003 143310 407879
rect 143448 407003 144004 407879
rect 144163 407017 144719 407893
rect 144857 407017 145413 407893
rect 145643 407032 146199 407908
rect 146337 407032 146893 407908
rect 147052 407046 147608 407922
rect 147746 407046 148302 407922
rect 148453 407061 149009 407937
rect 149147 407061 149703 407937
rect 149862 407075 150418 407951
rect 150556 407075 151112 407951
rect 141050 399610 141286 399846
rect 141050 399290 141286 399526
rect 141050 398970 141286 399206
rect 141445 398984 142001 399860
rect 142139 398984 142695 399860
rect 142846 398999 143402 399875
rect 143540 398999 144096 399875
rect 144255 399013 144811 399889
rect 144949 399013 145505 399889
rect 145735 399028 146291 399904
rect 146429 399028 146985 399904
rect 147144 399042 147700 399918
rect 147838 399042 148394 399918
rect 148545 399057 149101 399933
rect 149239 399057 149795 399933
rect 149954 399071 150510 399947
rect 150648 399071 151204 399947
rect 141064 391606 141300 391842
rect 141064 391286 141300 391522
rect 141064 390966 141300 391202
rect 141459 390980 142015 391856
rect 142153 390980 142709 391856
rect 142860 390995 143416 391871
rect 143554 390995 144110 391871
rect 144269 391009 144825 391885
rect 144963 391009 145519 391885
rect 145749 391024 146305 391900
rect 146443 391024 146999 391900
rect 147158 391038 147714 391914
rect 147852 391038 148408 391914
rect 148559 391053 149115 391929
rect 149253 391053 149809 391929
rect 149968 391067 150524 391943
rect 150662 391067 151218 391943
rect 141069 383622 141305 383858
rect 141069 383302 141305 383538
rect 141069 382982 141305 383218
rect 141464 382996 142020 383872
rect 142158 382996 142714 383872
rect 142865 383011 143421 383887
rect 143559 383011 144115 383887
rect 144274 383025 144830 383901
rect 144968 383025 145524 383901
rect 145754 383040 146310 383916
rect 146448 383040 147004 383916
rect 147163 383054 147719 383930
rect 147857 383054 148413 383930
rect 148564 383069 149120 383945
rect 149258 383069 149814 383945
rect 149973 383083 150529 383959
rect 150667 383083 151223 383959
rect 141062 375603 141298 375839
rect 141062 375283 141298 375519
rect 141062 374963 141298 375199
rect 141457 374977 142013 375853
rect 142151 374977 142707 375853
rect 142858 374992 143414 375868
rect 143552 374992 144108 375868
rect 144267 375006 144823 375882
rect 144961 375006 145517 375882
rect 145747 375021 146303 375897
rect 146441 375021 146997 375897
rect 147156 375035 147712 375911
rect 147850 375035 148406 375911
rect 148557 375050 149113 375926
rect 149251 375050 149807 375926
rect 149966 375064 150522 375940
rect 150660 375064 151216 375940
rect 141060 367664 141296 367900
rect 141060 367344 141296 367580
rect 141060 367024 141296 367260
rect 141455 367038 142011 367914
rect 142149 367038 142705 367914
rect 142856 367053 143412 367929
rect 143550 367053 144106 367929
rect 144265 367067 144821 367943
rect 144959 367067 145515 367943
rect 145745 367082 146301 367958
rect 146439 367082 146995 367958
rect 147154 367096 147710 367972
rect 147848 367096 148404 367972
rect 148555 367111 149111 367987
rect 149249 367111 149805 367987
rect 149964 367125 150520 368001
rect 150658 367125 151214 368001
rect 140964 359583 141200 359819
rect 140964 359263 141200 359499
rect 140964 358943 141200 359179
rect 141359 358957 141915 359833
rect 142053 358957 142609 359833
rect 142760 358972 143316 359848
rect 143454 358972 144010 359848
rect 144169 358986 144725 359862
rect 144863 358986 145419 359862
rect 145649 359001 146205 359877
rect 146343 359001 146899 359877
rect 147058 359015 147614 359891
rect 147752 359015 148308 359891
rect 148459 359030 149015 359906
rect 149153 359030 149709 359906
rect 149868 359044 150424 359920
rect 150562 359044 151118 359920
rect 141042 351606 141278 351842
rect 141042 351286 141278 351522
rect 141042 350966 141278 351202
rect 141437 350980 141993 351856
rect 142131 350980 142687 351856
rect 142838 350995 143394 351871
rect 143532 350995 144088 351871
rect 144247 351009 144803 351885
rect 144941 351009 145497 351885
rect 145727 351024 146283 351900
rect 146421 351024 146977 351900
rect 147136 351038 147692 351914
rect 147830 351038 148386 351914
rect 148537 351053 149093 351929
rect 149231 351053 149787 351929
rect 149946 351067 150502 351943
rect 150640 351067 151196 351943
rect 407908 564622 408144 564858
rect 408303 564636 408539 564872
rect 408623 564636 408859 564872
rect 408997 564636 409233 564872
rect 409317 564636 409553 564872
rect 409704 564651 409940 564887
rect 410024 564651 410260 564887
rect 410398 564651 410634 564887
rect 410718 564651 410954 564887
rect 411113 564665 411349 564901
rect 411433 564665 411669 564901
rect 411807 564665 412043 564901
rect 412127 564665 412363 564901
rect 412593 564680 412829 564916
rect 412913 564680 413149 564916
rect 413287 564680 413523 564916
rect 413607 564680 413843 564916
rect 414002 564694 414238 564930
rect 414322 564694 414558 564930
rect 414696 564694 414932 564930
rect 415016 564694 415252 564930
rect 415403 564709 415639 564945
rect 415723 564709 415959 564945
rect 416097 564709 416333 564945
rect 416417 564709 416653 564945
rect 416812 564723 417048 564959
rect 417132 564723 417368 564959
rect 417506 564723 417742 564959
rect 417826 564723 418062 564959
rect 407832 528661 408068 528897
rect 408227 528675 408463 528911
rect 408547 528675 408783 528911
rect 408921 528675 409157 528911
rect 409241 528675 409477 528911
rect 409628 528690 409864 528926
rect 409948 528690 410184 528926
rect 410322 528690 410558 528926
rect 410642 528690 410878 528926
rect 411037 528704 411273 528940
rect 411357 528704 411593 528940
rect 411731 528704 411967 528940
rect 412051 528704 412287 528940
rect 412517 528719 412753 528955
rect 412837 528719 413073 528955
rect 413211 528719 413447 528955
rect 413531 528719 413767 528955
rect 413926 528733 414162 528969
rect 414246 528733 414482 528969
rect 414620 528733 414856 528969
rect 414940 528733 415176 528969
rect 415327 528748 415563 528984
rect 415647 528748 415883 528984
rect 416021 528748 416257 528984
rect 416341 528748 416577 528984
rect 416736 528762 416972 528998
rect 417056 528762 417292 528998
rect 417430 528762 417666 528998
rect 417750 528762 417986 528998
rect 407812 492634 408048 492870
rect 408207 492648 408443 492884
rect 408527 492648 408763 492884
rect 408901 492648 409137 492884
rect 409221 492648 409457 492884
rect 409608 492663 409844 492899
rect 409928 492663 410164 492899
rect 410302 492663 410538 492899
rect 410622 492663 410858 492899
rect 411017 492677 411253 492913
rect 411337 492677 411573 492913
rect 411711 492677 411947 492913
rect 412031 492677 412267 492913
rect 412497 492692 412733 492928
rect 412817 492692 413053 492928
rect 413191 492692 413427 492928
rect 413511 492692 413747 492928
rect 413906 492706 414142 492942
rect 414226 492706 414462 492942
rect 414600 492706 414836 492942
rect 414920 492706 415156 492942
rect 415307 492721 415543 492957
rect 415627 492721 415863 492957
rect 416001 492721 416237 492957
rect 416321 492721 416557 492957
rect 416716 492735 416952 492971
rect 417036 492735 417272 492971
rect 417410 492735 417646 492971
rect 417730 492735 417966 492971
rect 407906 469285 408142 469521
rect 407906 468965 408142 469201
rect 407906 468645 408142 468881
rect 408301 468659 408857 469535
rect 408995 468659 409551 469535
rect 409702 468674 410258 469550
rect 410396 468674 410952 469550
rect 411111 468688 411667 469564
rect 411805 468688 412361 469564
rect 412591 468703 413147 469579
rect 413285 468703 413841 469579
rect 414000 468717 414556 469593
rect 414694 468717 415250 469593
rect 415401 468732 415957 469608
rect 416095 468732 416651 469608
rect 416810 468746 417366 469622
rect 417504 468746 418060 469622
rect 407909 461282 408145 461518
rect 407909 460962 408145 461198
rect 407909 460642 408145 460878
rect 408304 460656 408860 461532
rect 408998 460656 409554 461532
rect 409705 460671 410261 461547
rect 410399 460671 410955 461547
rect 411114 460685 411670 461561
rect 411808 460685 412364 461561
rect 412594 460700 413150 461576
rect 413288 460700 413844 461576
rect 414003 460714 414559 461590
rect 414697 460714 415253 461590
rect 415404 460729 415960 461605
rect 416098 460729 416654 461605
rect 416813 460743 417369 461619
rect 417507 460743 418063 461619
rect 407868 453286 408104 453522
rect 407868 452966 408104 453202
rect 407868 452646 408104 452882
rect 408263 452660 408819 453536
rect 408957 452660 409513 453536
rect 409664 452675 410220 453551
rect 410358 452675 410914 453551
rect 411073 452689 411629 453565
rect 411767 452689 412323 453565
rect 412553 452704 413109 453580
rect 413247 452704 413803 453580
rect 413962 452718 414518 453594
rect 414656 452718 415212 453594
rect 415363 452733 415919 453609
rect 416057 452733 416613 453609
rect 416772 452747 417328 453623
rect 417466 452747 418022 453623
rect 407859 445277 408095 445513
rect 407859 444957 408095 445193
rect 407859 444637 408095 444873
rect 408254 444651 408810 445527
rect 408948 444651 409504 445527
rect 409655 444666 410211 445542
rect 410349 444666 410905 445542
rect 411064 444680 411620 445556
rect 411758 444680 412314 445556
rect 412544 444695 413100 445571
rect 413238 444695 413794 445571
rect 413953 444709 414509 445585
rect 414647 444709 415203 445585
rect 415354 444724 415910 445600
rect 416048 444724 416604 445600
rect 416763 444738 417319 445614
rect 417457 444738 418013 445614
rect 407832 437291 408068 437527
rect 407832 436971 408068 437207
rect 407832 436651 408068 436887
rect 408227 436665 408783 437541
rect 408921 436665 409477 437541
rect 409628 436680 410184 437556
rect 410322 436680 410878 437556
rect 411037 436694 411593 437570
rect 411731 436694 412287 437570
rect 412517 436709 413073 437585
rect 413211 436709 413767 437585
rect 413926 436723 414482 437599
rect 414620 436723 415176 437599
rect 415327 436738 415883 437614
rect 416021 436738 416577 437614
rect 416736 436752 417292 437628
rect 417430 436752 417986 437628
rect 407856 429260 408092 429496
rect 407856 428940 408092 429176
rect 407856 428620 408092 428856
rect 408251 428634 408807 429510
rect 408945 428634 409501 429510
rect 409652 428649 410208 429525
rect 410346 428649 410902 429525
rect 411061 428663 411617 429539
rect 411755 428663 412311 429539
rect 412541 428678 413097 429554
rect 413235 428678 413791 429554
rect 413950 428692 414506 429568
rect 414644 428692 415200 429568
rect 415351 428707 415907 429583
rect 416045 428707 416601 429583
rect 416760 428721 417316 429597
rect 417454 428721 418010 429597
rect 407918 421329 408154 421565
rect 407918 421009 408154 421245
rect 407918 420689 408154 420925
rect 408313 420703 408869 421579
rect 409007 420703 409563 421579
rect 409714 420718 410270 421594
rect 410408 420718 410964 421594
rect 411123 420732 411679 421608
rect 411817 420732 412373 421608
rect 412603 420747 413159 421623
rect 413297 420747 413853 421623
rect 414012 420761 414568 421637
rect 414706 420761 415262 421637
rect 415413 420776 415969 421652
rect 416107 420776 416663 421652
rect 416822 420790 417378 421666
rect 417516 420790 418072 421666
rect 407934 413299 408170 413535
rect 407934 412979 408170 413215
rect 407934 412659 408170 412895
rect 408329 412673 408885 413549
rect 409023 412673 409579 413549
rect 409730 412688 410286 413564
rect 410424 412688 410980 413564
rect 411139 412702 411695 413578
rect 411833 412702 412389 413578
rect 412619 412717 413175 413593
rect 413313 412717 413869 413593
rect 414028 412731 414584 413607
rect 414722 412731 415278 413607
rect 415429 412746 415985 413622
rect 416123 412746 416679 413622
rect 416838 412760 417394 413636
rect 417532 412760 418088 413636
rect 407908 405291 408144 405527
rect 407908 404971 408144 405207
rect 407908 404651 408144 404887
rect 408303 404665 408859 405541
rect 408997 404665 409553 405541
rect 409704 404680 410260 405556
rect 410398 404680 410954 405556
rect 411113 404694 411669 405570
rect 411807 404694 412363 405570
rect 412593 404709 413149 405585
rect 413287 404709 413843 405585
rect 414002 404723 414558 405599
rect 414696 404723 415252 405599
rect 415403 404738 415959 405614
rect 416097 404738 416653 405614
rect 416812 404752 417368 405628
rect 417506 404752 418062 405628
rect 407882 397272 408118 397508
rect 407882 396952 408118 397188
rect 407882 396632 408118 396868
rect 408277 396646 408833 397522
rect 408971 396646 409527 397522
rect 409678 396661 410234 397537
rect 410372 396661 410928 397537
rect 411087 396675 411643 397551
rect 411781 396675 412337 397551
rect 412567 396690 413123 397566
rect 413261 396690 413817 397566
rect 413976 396704 414532 397580
rect 414670 396704 415226 397580
rect 415377 396719 415933 397595
rect 416071 396719 416627 397595
rect 416786 396733 417342 397609
rect 417480 396733 418036 397609
rect 407973 389269 408209 389505
rect 407973 388949 408209 389185
rect 407973 388629 408209 388865
rect 408368 388643 408924 389519
rect 409062 388643 409618 389519
rect 409769 388658 410325 389534
rect 410463 388658 411019 389534
rect 411178 388672 411734 389548
rect 411872 388672 412428 389548
rect 412658 388687 413214 389563
rect 413352 388687 413908 389563
rect 414067 388701 414623 389577
rect 414761 388701 415317 389577
rect 415468 388716 416024 389592
rect 416162 388716 416718 389592
rect 416877 388730 417433 389606
rect 417571 388730 418127 389606
rect 407894 381318 408130 381554
rect 407894 380998 408130 381234
rect 407894 380678 408130 380914
rect 408289 380692 408845 381568
rect 408983 380692 409539 381568
rect 409690 380707 410246 381583
rect 410384 380707 410940 381583
rect 411099 380721 411655 381597
rect 411793 380721 412349 381597
rect 412579 380736 413135 381612
rect 413273 380736 413829 381612
rect 413988 380750 414544 381626
rect 414682 380750 415238 381626
rect 415389 380765 415945 381641
rect 416083 380765 416639 381641
rect 416798 380779 417354 381655
rect 417492 380779 418048 381655
rect 407885 373290 408121 373526
rect 407885 372970 408121 373206
rect 407885 372650 408121 372886
rect 408280 372664 408836 373540
rect 408974 372664 409530 373540
rect 409681 372679 410237 373555
rect 410375 372679 410931 373555
rect 411090 372693 411646 373569
rect 411784 372693 412340 373569
rect 412570 372708 413126 373584
rect 413264 372708 413820 373584
rect 413979 372722 414535 373598
rect 414673 372722 415229 373598
rect 415380 372737 415936 373613
rect 416074 372737 416630 373613
rect 416789 372751 417345 373627
rect 417483 372751 418039 373627
rect 407877 365299 408113 365535
rect 407877 364979 408113 365215
rect 407877 364659 408113 364895
rect 408272 364673 408828 365549
rect 408966 364673 409522 365549
rect 409673 364688 410229 365564
rect 410367 364688 410923 365564
rect 411082 364702 411638 365578
rect 411776 364702 412332 365578
rect 412562 364717 413118 365593
rect 413256 364717 413812 365593
rect 413971 364731 414527 365607
rect 414665 364731 415221 365607
rect 415372 364746 415928 365622
rect 416066 364746 416622 365622
rect 416781 364760 417337 365636
rect 417475 364760 418031 365636
rect 407814 357309 408050 357545
rect 407814 356989 408050 357225
rect 407814 356669 408050 356905
rect 408209 356683 408765 357559
rect 408903 356683 409459 357559
rect 409610 356698 410166 357574
rect 410304 356698 410860 357574
rect 411019 356712 411575 357588
rect 411713 356712 412269 357588
rect 412499 356727 413055 357603
rect 413193 356727 413749 357603
rect 413908 356741 414464 357617
rect 414602 356741 415158 357617
rect 415309 356756 415865 357632
rect 416003 356756 416559 357632
rect 416718 356770 417274 357646
rect 417412 356770 417968 357646
rect 407901 349296 408137 349532
rect 407901 348976 408137 349212
rect 407901 348656 408137 348892
rect 408296 348670 408852 349546
rect 408990 348670 409546 349546
rect 409697 348685 410253 349561
rect 410391 348685 410947 349561
rect 411106 348699 411662 349575
rect 411800 348699 412356 349575
rect 412586 348714 413142 349590
rect 413280 348714 413836 349590
rect 413995 348728 414551 349604
rect 414689 348728 415245 349604
rect 415396 348743 415952 349619
rect 416090 348743 416646 349619
rect 416805 348757 417361 349633
rect 417499 348757 418055 349633
rect 141117 343640 141353 343876
rect 141117 343320 141353 343556
rect 141117 343000 141353 343236
rect 141512 343014 142068 343890
rect 142206 343014 142762 343890
rect 142913 343029 143469 343905
rect 143607 343029 144163 343905
rect 144322 343043 144878 343919
rect 145016 343043 145572 343919
rect 145802 343058 146358 343934
rect 146496 343058 147052 343934
rect 147211 343072 147767 343948
rect 147905 343072 148461 343948
rect 148612 343087 149168 343963
rect 149306 343087 149862 343963
rect 150021 343101 150577 343977
rect 150715 343101 151271 343977
rect 141144 327031 141380 327267
rect 141539 327045 141775 327281
rect 141859 327045 142095 327281
rect 142233 327045 142469 327281
rect 142553 327045 142789 327281
rect 142940 327060 143176 327296
rect 143260 327060 143496 327296
rect 143634 327060 143870 327296
rect 143954 327060 144190 327296
rect 144349 327074 144585 327310
rect 144669 327074 144905 327310
rect 145043 327074 145279 327310
rect 145363 327074 145599 327310
rect 145829 327089 146065 327325
rect 146149 327089 146385 327325
rect 146523 327089 146759 327325
rect 146843 327089 147079 327325
rect 147238 327103 147474 327339
rect 147558 327103 147794 327339
rect 147932 327103 148168 327339
rect 148252 327103 148488 327339
rect 148639 327118 148875 327354
rect 148959 327118 149195 327354
rect 149333 327118 149569 327354
rect 149653 327118 149889 327354
rect 150048 327132 150284 327368
rect 150368 327132 150604 327368
rect 150742 327132 150978 327368
rect 151062 327132 151298 327368
rect 141017 290998 141253 291234
rect 141412 291012 141648 291248
rect 141732 291012 141968 291248
rect 142106 291012 142342 291248
rect 142426 291012 142662 291248
rect 142813 291027 143049 291263
rect 143133 291027 143369 291263
rect 143507 291027 143743 291263
rect 143827 291027 144063 291263
rect 144222 291041 144458 291277
rect 144542 291041 144778 291277
rect 144916 291041 145152 291277
rect 145236 291041 145472 291277
rect 145702 291056 145938 291292
rect 146022 291056 146258 291292
rect 146396 291056 146632 291292
rect 146716 291056 146952 291292
rect 147111 291070 147347 291306
rect 147431 291070 147667 291306
rect 147805 291070 148041 291306
rect 148125 291070 148361 291306
rect 148512 291085 148748 291321
rect 148832 291085 149068 291321
rect 149206 291085 149442 291321
rect 149526 291085 149762 291321
rect 149921 291099 150157 291335
rect 150241 291099 150477 291335
rect 150615 291099 150851 291335
rect 150935 291099 151171 291335
rect 141045 254988 141281 255224
rect 141440 255002 141676 255238
rect 141760 255002 141996 255238
rect 142134 255002 142370 255238
rect 142454 255002 142690 255238
rect 142841 255017 143077 255253
rect 143161 255017 143397 255253
rect 143535 255017 143771 255253
rect 143855 255017 144091 255253
rect 144250 255031 144486 255267
rect 144570 255031 144806 255267
rect 144944 255031 145180 255267
rect 145264 255031 145500 255267
rect 145730 255046 145966 255282
rect 146050 255046 146286 255282
rect 146424 255046 146660 255282
rect 146744 255046 146980 255282
rect 147139 255060 147375 255296
rect 147459 255060 147695 255296
rect 147833 255060 148069 255296
rect 148153 255060 148389 255296
rect 148540 255075 148776 255311
rect 148860 255075 149096 255311
rect 149234 255075 149470 255311
rect 149554 255075 149790 255311
rect 149949 255089 150185 255325
rect 150269 255089 150505 255325
rect 150643 255089 150879 255325
rect 150963 255089 151199 255325
rect 102786 212018 103022 212254
rect 102786 211698 103022 211934
rect 102786 176018 103022 176254
rect 102786 175698 103022 175934
rect 102786 140018 103022 140254
rect 102786 139698 103022 139934
rect 102786 104018 103022 104254
rect 102786 103698 103022 103934
rect 102786 68018 103022 68254
rect 102786 67698 103022 67934
rect 102786 32018 103022 32254
rect 102786 31698 103022 31934
rect 84786 -6222 85022 -5986
rect 84786 -6542 85022 -6306
rect 109986 183218 110222 183454
rect 109986 182898 110222 183134
rect 109986 147218 110222 147454
rect 109986 146898 110222 147134
rect 109986 111218 110222 111454
rect 109986 110898 110222 111134
rect 109986 75218 110222 75454
rect 109986 74898 110222 75134
rect 109986 39218 110222 39454
rect 109986 38898 110222 39134
rect 109986 3218 110222 3454
rect 109986 2898 110222 3134
rect 109986 -582 110222 -346
rect 109986 -902 110222 -666
rect 113586 186818 113822 187054
rect 113586 186498 113822 186734
rect 113586 150818 113822 151054
rect 113586 150498 113822 150734
rect 113586 114818 113822 115054
rect 113586 114498 113822 114734
rect 113586 78818 113822 79054
rect 113586 78498 113822 78734
rect 113586 42818 113822 43054
rect 113586 42498 113822 42734
rect 113586 6818 113822 7054
rect 113586 6498 113822 6734
rect 113586 -2462 113822 -2226
rect 113586 -2782 113822 -2546
rect 117186 190418 117422 190654
rect 117186 190098 117422 190334
rect 117186 154418 117422 154654
rect 117186 154098 117422 154334
rect 117186 118418 117422 118654
rect 117186 118098 117422 118334
rect 117186 82418 117422 82654
rect 117186 82098 117422 82334
rect 117186 46418 117422 46654
rect 117186 46098 117422 46334
rect 117186 10418 117422 10654
rect 117186 10098 117422 10334
rect 117186 -4342 117422 -4106
rect 117186 -4662 117422 -4426
rect 120786 194018 121022 194254
rect 120786 193698 121022 193934
rect 120786 158018 121022 158254
rect 120786 157698 121022 157934
rect 120786 122018 121022 122254
rect 120786 121698 121022 121934
rect 120786 86018 121022 86254
rect 120786 85698 121022 85934
rect 120786 50018 121022 50254
rect 120786 49698 121022 49934
rect 120786 14018 121022 14254
rect 120786 13698 121022 13934
rect 102786 -7162 103022 -6926
rect 102786 -7482 103022 -7246
rect 127986 201218 128222 201454
rect 127986 200898 128222 201134
rect 127986 165218 128222 165454
rect 127986 164898 128222 165134
rect 127986 129218 128222 129454
rect 127986 128898 128222 129134
rect 127986 93218 128222 93454
rect 127986 92898 128222 93134
rect 127986 57218 128222 57454
rect 127986 56898 128222 57134
rect 127986 21218 128222 21454
rect 127986 20898 128222 21134
rect 127986 -1522 128222 -1286
rect 127986 -1842 128222 -1606
rect 131586 204818 131822 205054
rect 131586 204498 131822 204734
rect 131586 168818 131822 169054
rect 131586 168498 131822 168734
rect 131586 132818 131822 133054
rect 131586 132498 131822 132734
rect 131586 96818 131822 97054
rect 131586 96498 131822 96734
rect 131586 60818 131822 61054
rect 131586 60498 131822 60734
rect 131586 24818 131822 25054
rect 131586 24498 131822 24734
rect 131586 -3402 131822 -3166
rect 131586 -3722 131822 -3486
rect 135186 208418 135422 208654
rect 135186 208098 135422 208334
rect 135186 172418 135422 172654
rect 135186 172098 135422 172334
rect 135186 136418 135422 136654
rect 135186 136098 135422 136334
rect 135186 100418 135422 100654
rect 135186 100098 135422 100334
rect 135186 64418 135422 64654
rect 135186 64098 135422 64334
rect 135186 28418 135422 28654
rect 135186 28098 135422 28334
rect 135186 -5282 135422 -5046
rect 135186 -5602 135422 -5366
rect 138786 212018 139022 212254
rect 138786 211698 139022 211934
rect 138786 176018 139022 176254
rect 138786 175698 139022 175934
rect 138786 140018 139022 140254
rect 138786 139698 139022 139934
rect 138786 104018 139022 104254
rect 138786 103698 139022 103934
rect 138786 68018 139022 68254
rect 138786 67698 139022 67934
rect 138786 32018 139022 32254
rect 138786 31698 139022 31934
rect 120786 -6222 121022 -5986
rect 120786 -6542 121022 -6306
rect 145986 183218 146222 183454
rect 145986 182898 146222 183134
rect 145986 147218 146222 147454
rect 145986 146898 146222 147134
rect 145986 111218 146222 111454
rect 145986 110898 146222 111134
rect 145986 75218 146222 75454
rect 145986 74898 146222 75134
rect 145986 39218 146222 39454
rect 145986 38898 146222 39134
rect 145986 3218 146222 3454
rect 145986 2898 146222 3134
rect 145986 -582 146222 -346
rect 145986 -902 146222 -666
rect 149586 186818 149822 187054
rect 149586 186498 149822 186734
rect 149586 150818 149822 151054
rect 149586 150498 149822 150734
rect 149586 114818 149822 115054
rect 149586 114498 149822 114734
rect 149586 78818 149822 79054
rect 149586 78498 149822 78734
rect 149586 42818 149822 43054
rect 149586 42498 149822 42734
rect 149586 6818 149822 7054
rect 149586 6498 149822 6734
rect 149586 -2462 149822 -2226
rect 149586 -2782 149822 -2546
rect 153186 190418 153422 190654
rect 153186 190098 153422 190334
rect 153186 154418 153422 154654
rect 153186 154098 153422 154334
rect 153186 118418 153422 118654
rect 153186 118098 153422 118334
rect 153186 82418 153422 82654
rect 153186 82098 153422 82334
rect 153186 46418 153422 46654
rect 153186 46098 153422 46334
rect 153186 10418 153422 10654
rect 153186 10098 153422 10334
rect 153186 -4342 153422 -4106
rect 153186 -4662 153422 -4426
rect 156786 194018 157022 194254
rect 156786 193698 157022 193934
rect 156786 158018 157022 158254
rect 156786 157698 157022 157934
rect 156786 122018 157022 122254
rect 156786 121698 157022 121934
rect 156786 86018 157022 86254
rect 156786 85698 157022 85934
rect 156786 50018 157022 50254
rect 156786 49698 157022 49934
rect 156786 14018 157022 14254
rect 156786 13698 157022 13934
rect 138786 -7162 139022 -6926
rect 138786 -7482 139022 -7246
rect 163986 201218 164222 201454
rect 163986 200898 164222 201134
rect 163986 165218 164222 165454
rect 163986 164898 164222 165134
rect 163986 129218 164222 129454
rect 163986 128898 164222 129134
rect 163986 93218 164222 93454
rect 163986 92898 164222 93134
rect 163986 57218 164222 57454
rect 163986 56898 164222 57134
rect 163986 21218 164222 21454
rect 163986 20898 164222 21134
rect 163986 -1522 164222 -1286
rect 163986 -1842 164222 -1606
rect 167586 204818 167822 205054
rect 167586 204498 167822 204734
rect 167586 168818 167822 169054
rect 167586 168498 167822 168734
rect 167586 132818 167822 133054
rect 167586 132498 167822 132734
rect 167586 96818 167822 97054
rect 167586 96498 167822 96734
rect 167586 60818 167822 61054
rect 167586 60498 167822 60734
rect 167586 24818 167822 25054
rect 167586 24498 167822 24734
rect 167586 -3402 167822 -3166
rect 167586 -3722 167822 -3486
rect 171186 208418 171422 208654
rect 171186 208098 171422 208334
rect 171186 172418 171422 172654
rect 171186 172098 171422 172334
rect 171186 136418 171422 136654
rect 171186 136098 171422 136334
rect 171186 100418 171422 100654
rect 171186 100098 171422 100334
rect 171186 64418 171422 64654
rect 171186 64098 171422 64334
rect 171186 28418 171422 28654
rect 171186 28098 171422 28334
rect 171186 -5282 171422 -5046
rect 171186 -5602 171422 -5366
rect 174786 212018 175022 212254
rect 174786 211698 175022 211934
rect 174786 176018 175022 176254
rect 174786 175698 175022 175934
rect 174786 140018 175022 140254
rect 174786 139698 175022 139934
rect 174786 104018 175022 104254
rect 174786 103698 175022 103934
rect 174786 68018 175022 68254
rect 174786 67698 175022 67934
rect 174786 32018 175022 32254
rect 174786 31698 175022 31934
rect 156786 -6222 157022 -5986
rect 156786 -6542 157022 -6306
rect 181986 183218 182222 183454
rect 181986 182898 182222 183134
rect 181986 147218 182222 147454
rect 181986 146898 182222 147134
rect 181986 111218 182222 111454
rect 181986 110898 182222 111134
rect 181986 75218 182222 75454
rect 181986 74898 182222 75134
rect 181986 39218 182222 39454
rect 181986 38898 182222 39134
rect 181986 3218 182222 3454
rect 181986 2898 182222 3134
rect 181986 -582 182222 -346
rect 181986 -902 182222 -666
rect 185586 186818 185822 187054
rect 185586 186498 185822 186734
rect 185586 150818 185822 151054
rect 185586 150498 185822 150734
rect 185586 114818 185822 115054
rect 185586 114498 185822 114734
rect 185586 78818 185822 79054
rect 185586 78498 185822 78734
rect 185586 42818 185822 43054
rect 185586 42498 185822 42734
rect 185586 6818 185822 7054
rect 185586 6498 185822 6734
rect 185586 -2462 185822 -2226
rect 185586 -2782 185822 -2546
rect 189186 190418 189422 190654
rect 189186 190098 189422 190334
rect 189186 154418 189422 154654
rect 189186 154098 189422 154334
rect 189186 118418 189422 118654
rect 189186 118098 189422 118334
rect 189186 82418 189422 82654
rect 189186 82098 189422 82334
rect 189186 46418 189422 46654
rect 189186 46098 189422 46334
rect 189186 10418 189422 10654
rect 189186 10098 189422 10334
rect 189186 -4342 189422 -4106
rect 189186 -4662 189422 -4426
rect 192786 194018 193022 194254
rect 192786 193698 193022 193934
rect 192786 158018 193022 158254
rect 192786 157698 193022 157934
rect 192786 122018 193022 122254
rect 192786 121698 193022 121934
rect 192786 86018 193022 86254
rect 192786 85698 193022 85934
rect 192786 50018 193022 50254
rect 192786 49698 193022 49934
rect 192786 14018 193022 14254
rect 192786 13698 193022 13934
rect 174786 -7162 175022 -6926
rect 174786 -7482 175022 -7246
rect 199986 201218 200222 201454
rect 199986 200898 200222 201134
rect 199986 165218 200222 165454
rect 199986 164898 200222 165134
rect 199986 129218 200222 129454
rect 199986 128898 200222 129134
rect 199986 93218 200222 93454
rect 199986 92898 200222 93134
rect 199986 57218 200222 57454
rect 199986 56898 200222 57134
rect 199986 21218 200222 21454
rect 199986 20898 200222 21134
rect 199986 -1522 200222 -1286
rect 199986 -1842 200222 -1606
rect 203586 204818 203822 205054
rect 203586 204498 203822 204734
rect 203586 168818 203822 169054
rect 203586 168498 203822 168734
rect 203586 132818 203822 133054
rect 203586 132498 203822 132734
rect 203586 96818 203822 97054
rect 203586 96498 203822 96734
rect 203586 60818 203822 61054
rect 203586 60498 203822 60734
rect 203586 24818 203822 25054
rect 203586 24498 203822 24734
rect 203586 -3402 203822 -3166
rect 203586 -3722 203822 -3486
rect 207186 208418 207422 208654
rect 207186 208098 207422 208334
rect 207186 172418 207422 172654
rect 207186 172098 207422 172334
rect 207186 136418 207422 136654
rect 207186 136098 207422 136334
rect 207186 100418 207422 100654
rect 207186 100098 207422 100334
rect 207186 64418 207422 64654
rect 207186 64098 207422 64334
rect 207186 28418 207422 28654
rect 207186 28098 207422 28334
rect 207186 -5282 207422 -5046
rect 207186 -5602 207422 -5366
rect 210786 212018 211022 212254
rect 210786 211698 211022 211934
rect 210786 176018 211022 176254
rect 210786 175698 211022 175934
rect 210786 140018 211022 140254
rect 210786 139698 211022 139934
rect 210786 104018 211022 104254
rect 210786 103698 211022 103934
rect 210786 68018 211022 68254
rect 210786 67698 211022 67934
rect 210786 32018 211022 32254
rect 210786 31698 211022 31934
rect 192786 -6222 193022 -5986
rect 192786 -6542 193022 -6306
rect 217986 183218 218222 183454
rect 217986 182898 218222 183134
rect 217986 147218 218222 147454
rect 217986 146898 218222 147134
rect 217986 111218 218222 111454
rect 217986 110898 218222 111134
rect 217986 75218 218222 75454
rect 217986 74898 218222 75134
rect 217986 39218 218222 39454
rect 217986 38898 218222 39134
rect 217986 3218 218222 3454
rect 217986 2898 218222 3134
rect 217986 -582 218222 -346
rect 217986 -902 218222 -666
rect 221586 186818 221822 187054
rect 221586 186498 221822 186734
rect 221586 150818 221822 151054
rect 221586 150498 221822 150734
rect 221586 114818 221822 115054
rect 221586 114498 221822 114734
rect 221586 78818 221822 79054
rect 221586 78498 221822 78734
rect 221586 42818 221822 43054
rect 221586 42498 221822 42734
rect 221586 6818 221822 7054
rect 221586 6498 221822 6734
rect 221586 -2462 221822 -2226
rect 221586 -2782 221822 -2546
rect 225186 190418 225422 190654
rect 225186 190098 225422 190334
rect 225186 154418 225422 154654
rect 225186 154098 225422 154334
rect 225186 118418 225422 118654
rect 225186 118098 225422 118334
rect 225186 82418 225422 82654
rect 225186 82098 225422 82334
rect 225186 46418 225422 46654
rect 225186 46098 225422 46334
rect 225186 10418 225422 10654
rect 225186 10098 225422 10334
rect 225186 -4342 225422 -4106
rect 225186 -4662 225422 -4426
rect 228786 194018 229022 194254
rect 228786 193698 229022 193934
rect 228786 158018 229022 158254
rect 228786 157698 229022 157934
rect 228786 122018 229022 122254
rect 228786 121698 229022 121934
rect 228786 86018 229022 86254
rect 228786 85698 229022 85934
rect 228786 50018 229022 50254
rect 228786 49698 229022 49934
rect 228786 14018 229022 14254
rect 228786 13698 229022 13934
rect 210786 -7162 211022 -6926
rect 210786 -7482 211022 -7246
rect 235986 201218 236222 201454
rect 235986 200898 236222 201134
rect 235986 165218 236222 165454
rect 235986 164898 236222 165134
rect 235986 129218 236222 129454
rect 235986 128898 236222 129134
rect 235986 93218 236222 93454
rect 235986 92898 236222 93134
rect 235986 57218 236222 57454
rect 235986 56898 236222 57134
rect 235986 21218 236222 21454
rect 235986 20898 236222 21134
rect 235986 -1522 236222 -1286
rect 235986 -1842 236222 -1606
rect 239586 204818 239822 205054
rect 239586 204498 239822 204734
rect 239586 168818 239822 169054
rect 239586 168498 239822 168734
rect 239586 132818 239822 133054
rect 239586 132498 239822 132734
rect 239586 96818 239822 97054
rect 239586 96498 239822 96734
rect 239586 60818 239822 61054
rect 239586 60498 239822 60734
rect 239586 24818 239822 25054
rect 239586 24498 239822 24734
rect 239586 -3402 239822 -3166
rect 239586 -3722 239822 -3486
rect 243186 208418 243422 208654
rect 243186 208098 243422 208334
rect 243186 172418 243422 172654
rect 243186 172098 243422 172334
rect 243186 136418 243422 136654
rect 243186 136098 243422 136334
rect 243186 100418 243422 100654
rect 243186 100098 243422 100334
rect 243186 64418 243422 64654
rect 243186 64098 243422 64334
rect 243186 28418 243422 28654
rect 243186 28098 243422 28334
rect 243186 -5282 243422 -5046
rect 243186 -5602 243422 -5366
rect 246786 212018 247022 212254
rect 246786 211698 247022 211934
rect 246786 176018 247022 176254
rect 246786 175698 247022 175934
rect 246786 140018 247022 140254
rect 246786 139698 247022 139934
rect 246786 104018 247022 104254
rect 246786 103698 247022 103934
rect 246786 68018 247022 68254
rect 246786 67698 247022 67934
rect 246786 32018 247022 32254
rect 246786 31698 247022 31934
rect 228786 -6222 229022 -5986
rect 228786 -6542 229022 -6306
rect 253986 183218 254222 183454
rect 253986 182898 254222 183134
rect 253986 147218 254222 147454
rect 253986 146898 254222 147134
rect 253986 111218 254222 111454
rect 253986 110898 254222 111134
rect 253986 75218 254222 75454
rect 253986 74898 254222 75134
rect 253986 39218 254222 39454
rect 253986 38898 254222 39134
rect 253986 3218 254222 3454
rect 253986 2898 254222 3134
rect 253986 -582 254222 -346
rect 253986 -902 254222 -666
rect 257586 186818 257822 187054
rect 257586 186498 257822 186734
rect 257586 150818 257822 151054
rect 257586 150498 257822 150734
rect 257586 114818 257822 115054
rect 257586 114498 257822 114734
rect 257586 78818 257822 79054
rect 257586 78498 257822 78734
rect 257586 42818 257822 43054
rect 257586 42498 257822 42734
rect 257586 6818 257822 7054
rect 257586 6498 257822 6734
rect 257586 -2462 257822 -2226
rect 257586 -2782 257822 -2546
rect 261186 190418 261422 190654
rect 261186 190098 261422 190334
rect 261186 154418 261422 154654
rect 261186 154098 261422 154334
rect 261186 118418 261422 118654
rect 261186 118098 261422 118334
rect 261186 82418 261422 82654
rect 261186 82098 261422 82334
rect 261186 46418 261422 46654
rect 261186 46098 261422 46334
rect 261186 10418 261422 10654
rect 261186 10098 261422 10334
rect 261186 -4342 261422 -4106
rect 261186 -4662 261422 -4426
rect 264786 194018 265022 194254
rect 264786 193698 265022 193934
rect 264786 158018 265022 158254
rect 264786 157698 265022 157934
rect 264786 122018 265022 122254
rect 264786 121698 265022 121934
rect 264786 86018 265022 86254
rect 264786 85698 265022 85934
rect 264786 50018 265022 50254
rect 264786 49698 265022 49934
rect 264786 14018 265022 14254
rect 264786 13698 265022 13934
rect 246786 -7162 247022 -6926
rect 246786 -7482 247022 -7246
rect 271986 201218 272222 201454
rect 271986 200898 272222 201134
rect 271986 165218 272222 165454
rect 271986 164898 272222 165134
rect 271986 129218 272222 129454
rect 271986 128898 272222 129134
rect 271986 93218 272222 93454
rect 271986 92898 272222 93134
rect 271986 57218 272222 57454
rect 271986 56898 272222 57134
rect 271986 21218 272222 21454
rect 271986 20898 272222 21134
rect 271986 -1522 272222 -1286
rect 271986 -1842 272222 -1606
rect 275586 204818 275822 205054
rect 275586 204498 275822 204734
rect 275586 168818 275822 169054
rect 275586 168498 275822 168734
rect 275586 132818 275822 133054
rect 275586 132498 275822 132734
rect 275586 96818 275822 97054
rect 275586 96498 275822 96734
rect 275586 60818 275822 61054
rect 275586 60498 275822 60734
rect 275586 24818 275822 25054
rect 275586 24498 275822 24734
rect 275586 -3402 275822 -3166
rect 275586 -3722 275822 -3486
rect 279186 208418 279422 208654
rect 279186 208098 279422 208334
rect 279186 172418 279422 172654
rect 279186 172098 279422 172334
rect 279186 136418 279422 136654
rect 279186 136098 279422 136334
rect 279186 100418 279422 100654
rect 279186 100098 279422 100334
rect 279186 64418 279422 64654
rect 279186 64098 279422 64334
rect 279186 28418 279422 28654
rect 279186 28098 279422 28334
rect 279186 -5282 279422 -5046
rect 279186 -5602 279422 -5366
rect 282786 212018 283022 212254
rect 282786 211698 283022 211934
rect 282786 176018 283022 176254
rect 282786 175698 283022 175934
rect 282786 140018 283022 140254
rect 282786 139698 283022 139934
rect 282786 104018 283022 104254
rect 282786 103698 283022 103934
rect 282786 68018 283022 68254
rect 282786 67698 283022 67934
rect 282786 32018 283022 32254
rect 282786 31698 283022 31934
rect 264786 -6222 265022 -5986
rect 264786 -6542 265022 -6306
rect 289986 183218 290222 183454
rect 289986 182898 290222 183134
rect 289986 147218 290222 147454
rect 289986 146898 290222 147134
rect 289986 111218 290222 111454
rect 289986 110898 290222 111134
rect 289986 75218 290222 75454
rect 289986 74898 290222 75134
rect 289986 39218 290222 39454
rect 289986 38898 290222 39134
rect 289986 3218 290222 3454
rect 289986 2898 290222 3134
rect 289986 -582 290222 -346
rect 289986 -902 290222 -666
rect 293586 186818 293822 187054
rect 293586 186498 293822 186734
rect 293586 150818 293822 151054
rect 293586 150498 293822 150734
rect 293586 114818 293822 115054
rect 293586 114498 293822 114734
rect 293586 78818 293822 79054
rect 293586 78498 293822 78734
rect 293586 42818 293822 43054
rect 293586 42498 293822 42734
rect 293586 6818 293822 7054
rect 293586 6498 293822 6734
rect 293586 -2462 293822 -2226
rect 293586 -2782 293822 -2546
rect 297186 190418 297422 190654
rect 297186 190098 297422 190334
rect 297186 154418 297422 154654
rect 297186 154098 297422 154334
rect 297186 118418 297422 118654
rect 297186 118098 297422 118334
rect 297186 82418 297422 82654
rect 297186 82098 297422 82334
rect 297186 46418 297422 46654
rect 297186 46098 297422 46334
rect 297186 10418 297422 10654
rect 297186 10098 297422 10334
rect 297186 -4342 297422 -4106
rect 297186 -4662 297422 -4426
rect 300786 194018 301022 194254
rect 300786 193698 301022 193934
rect 300786 158018 301022 158254
rect 300786 157698 301022 157934
rect 300786 122018 301022 122254
rect 300786 121698 301022 121934
rect 300786 86018 301022 86254
rect 300786 85698 301022 85934
rect 300786 50018 301022 50254
rect 300786 49698 301022 49934
rect 300786 14018 301022 14254
rect 300786 13698 301022 13934
rect 282786 -7162 283022 -6926
rect 282786 -7482 283022 -7246
rect 307986 201218 308222 201454
rect 307986 200898 308222 201134
rect 307986 165218 308222 165454
rect 307986 164898 308222 165134
rect 307986 129218 308222 129454
rect 307986 128898 308222 129134
rect 307986 93218 308222 93454
rect 307986 92898 308222 93134
rect 307986 57218 308222 57454
rect 307986 56898 308222 57134
rect 307986 21218 308222 21454
rect 307986 20898 308222 21134
rect 307986 -1522 308222 -1286
rect 307986 -1842 308222 -1606
rect 311586 204818 311822 205054
rect 311586 204498 311822 204734
rect 311586 168818 311822 169054
rect 311586 168498 311822 168734
rect 311586 132818 311822 133054
rect 311586 132498 311822 132734
rect 311586 96818 311822 97054
rect 311586 96498 311822 96734
rect 311586 60818 311822 61054
rect 311586 60498 311822 60734
rect 311586 24818 311822 25054
rect 311586 24498 311822 24734
rect 311586 -3402 311822 -3166
rect 311586 -3722 311822 -3486
rect 315186 208418 315422 208654
rect 315186 208098 315422 208334
rect 315186 172418 315422 172654
rect 315186 172098 315422 172334
rect 315186 136418 315422 136654
rect 315186 136098 315422 136334
rect 315186 100418 315422 100654
rect 315186 100098 315422 100334
rect 315186 64418 315422 64654
rect 315186 64098 315422 64334
rect 315186 28418 315422 28654
rect 315186 28098 315422 28334
rect 315186 -5282 315422 -5046
rect 315186 -5602 315422 -5366
rect 318786 212018 319022 212254
rect 318786 211698 319022 211934
rect 318786 176018 319022 176254
rect 318786 175698 319022 175934
rect 318786 140018 319022 140254
rect 318786 139698 319022 139934
rect 318786 104018 319022 104254
rect 318786 103698 319022 103934
rect 318786 68018 319022 68254
rect 318786 67698 319022 67934
rect 318786 32018 319022 32254
rect 318786 31698 319022 31934
rect 300786 -6222 301022 -5986
rect 300786 -6542 301022 -6306
rect 325986 183218 326222 183454
rect 325986 182898 326222 183134
rect 325986 147218 326222 147454
rect 325986 146898 326222 147134
rect 325986 111218 326222 111454
rect 325986 110898 326222 111134
rect 325986 75218 326222 75454
rect 325986 74898 326222 75134
rect 325986 39218 326222 39454
rect 325986 38898 326222 39134
rect 325986 3218 326222 3454
rect 325986 2898 326222 3134
rect 325986 -582 326222 -346
rect 325986 -902 326222 -666
rect 329586 186818 329822 187054
rect 329586 186498 329822 186734
rect 329586 150818 329822 151054
rect 329586 150498 329822 150734
rect 329586 114818 329822 115054
rect 329586 114498 329822 114734
rect 329586 78818 329822 79054
rect 329586 78498 329822 78734
rect 329586 42818 329822 43054
rect 329586 42498 329822 42734
rect 329586 6818 329822 7054
rect 329586 6498 329822 6734
rect 329586 -2462 329822 -2226
rect 329586 -2782 329822 -2546
rect 333186 190418 333422 190654
rect 333186 190098 333422 190334
rect 333186 154418 333422 154654
rect 333186 154098 333422 154334
rect 333186 118418 333422 118654
rect 333186 118098 333422 118334
rect 333186 82418 333422 82654
rect 333186 82098 333422 82334
rect 333186 46418 333422 46654
rect 333186 46098 333422 46334
rect 333186 10418 333422 10654
rect 333186 10098 333422 10334
rect 333186 -4342 333422 -4106
rect 333186 -4662 333422 -4426
rect 336786 194018 337022 194254
rect 336786 193698 337022 193934
rect 336786 158018 337022 158254
rect 336786 157698 337022 157934
rect 336786 122018 337022 122254
rect 336786 121698 337022 121934
rect 336786 86018 337022 86254
rect 336786 85698 337022 85934
rect 336786 50018 337022 50254
rect 336786 49698 337022 49934
rect 336786 14018 337022 14254
rect 336786 13698 337022 13934
rect 318786 -7162 319022 -6926
rect 318786 -7482 319022 -7246
rect 343986 201218 344222 201454
rect 343986 200898 344222 201134
rect 343986 165218 344222 165454
rect 343986 164898 344222 165134
rect 343986 129218 344222 129454
rect 343986 128898 344222 129134
rect 343986 93218 344222 93454
rect 343986 92898 344222 93134
rect 343986 57218 344222 57454
rect 343986 56898 344222 57134
rect 343986 21218 344222 21454
rect 343986 20898 344222 21134
rect 343986 -1522 344222 -1286
rect 343986 -1842 344222 -1606
rect 347586 204818 347822 205054
rect 347586 204498 347822 204734
rect 347586 168818 347822 169054
rect 347586 168498 347822 168734
rect 347586 132818 347822 133054
rect 347586 132498 347822 132734
rect 347586 96818 347822 97054
rect 347586 96498 347822 96734
rect 347586 60818 347822 61054
rect 347586 60498 347822 60734
rect 347586 24818 347822 25054
rect 347586 24498 347822 24734
rect 347586 -3402 347822 -3166
rect 347586 -3722 347822 -3486
rect 351186 208418 351422 208654
rect 351186 208098 351422 208334
rect 351186 172418 351422 172654
rect 351186 172098 351422 172334
rect 351186 136418 351422 136654
rect 351186 136098 351422 136334
rect 351186 100418 351422 100654
rect 351186 100098 351422 100334
rect 351186 64418 351422 64654
rect 351186 64098 351422 64334
rect 351186 28418 351422 28654
rect 351186 28098 351422 28334
rect 351186 -5282 351422 -5046
rect 351186 -5602 351422 -5366
rect 354786 212018 355022 212254
rect 354786 211698 355022 211934
rect 354786 176018 355022 176254
rect 354786 175698 355022 175934
rect 354786 140018 355022 140254
rect 354786 139698 355022 139934
rect 354786 104018 355022 104254
rect 354786 103698 355022 103934
rect 354786 68018 355022 68254
rect 354786 67698 355022 67934
rect 354786 32018 355022 32254
rect 354786 31698 355022 31934
rect 336786 -6222 337022 -5986
rect 336786 -6542 337022 -6306
rect 361986 183218 362222 183454
rect 361986 182898 362222 183134
rect 361986 147218 362222 147454
rect 361986 146898 362222 147134
rect 361986 111218 362222 111454
rect 361986 110898 362222 111134
rect 361986 75218 362222 75454
rect 361986 74898 362222 75134
rect 361986 39218 362222 39454
rect 361986 38898 362222 39134
rect 361986 3218 362222 3454
rect 361986 2898 362222 3134
rect 361986 -582 362222 -346
rect 361986 -902 362222 -666
rect 365586 186818 365822 187054
rect 365586 186498 365822 186734
rect 365586 150818 365822 151054
rect 365586 150498 365822 150734
rect 365586 114818 365822 115054
rect 365586 114498 365822 114734
rect 365586 78818 365822 79054
rect 365586 78498 365822 78734
rect 365586 42818 365822 43054
rect 365586 42498 365822 42734
rect 365586 6818 365822 7054
rect 365586 6498 365822 6734
rect 365586 -2462 365822 -2226
rect 365586 -2782 365822 -2546
rect 369186 190418 369422 190654
rect 369186 190098 369422 190334
rect 369186 154418 369422 154654
rect 369186 154098 369422 154334
rect 369186 118418 369422 118654
rect 369186 118098 369422 118334
rect 369186 82418 369422 82654
rect 369186 82098 369422 82334
rect 369186 46418 369422 46654
rect 369186 46098 369422 46334
rect 369186 10418 369422 10654
rect 369186 10098 369422 10334
rect 369186 -4342 369422 -4106
rect 369186 -4662 369422 -4426
rect 372786 194018 373022 194254
rect 372786 193698 373022 193934
rect 372786 158018 373022 158254
rect 372786 157698 373022 157934
rect 372786 122018 373022 122254
rect 372786 121698 373022 121934
rect 372786 86018 373022 86254
rect 372786 85698 373022 85934
rect 372786 50018 373022 50254
rect 372786 49698 373022 49934
rect 372786 14018 373022 14254
rect 372786 13698 373022 13934
rect 354786 -7162 355022 -6926
rect 354786 -7482 355022 -7246
rect 379986 201218 380222 201454
rect 379986 200898 380222 201134
rect 379986 165218 380222 165454
rect 379986 164898 380222 165134
rect 379986 129218 380222 129454
rect 379986 128898 380222 129134
rect 379986 93218 380222 93454
rect 379986 92898 380222 93134
rect 379986 57218 380222 57454
rect 379986 56898 380222 57134
rect 379986 21218 380222 21454
rect 379986 20898 380222 21134
rect 379986 -1522 380222 -1286
rect 379986 -1842 380222 -1606
rect 383586 204818 383822 205054
rect 383586 204498 383822 204734
rect 383586 168818 383822 169054
rect 383586 168498 383822 168734
rect 383586 132818 383822 133054
rect 383586 132498 383822 132734
rect 383586 96818 383822 97054
rect 383586 96498 383822 96734
rect 383586 60818 383822 61054
rect 383586 60498 383822 60734
rect 383586 24818 383822 25054
rect 383586 24498 383822 24734
rect 383586 -3402 383822 -3166
rect 383586 -3722 383822 -3486
rect 387186 208418 387422 208654
rect 387186 208098 387422 208334
rect 387186 172418 387422 172654
rect 387186 172098 387422 172334
rect 387186 136418 387422 136654
rect 387186 136098 387422 136334
rect 387186 100418 387422 100654
rect 387186 100098 387422 100334
rect 387186 64418 387422 64654
rect 387186 64098 387422 64334
rect 407917 312623 408153 312859
rect 408312 312637 408548 312873
rect 408632 312637 408868 312873
rect 409006 312637 409242 312873
rect 409326 312637 409562 312873
rect 409713 312652 409949 312888
rect 410033 312652 410269 312888
rect 410407 312652 410643 312888
rect 410727 312652 410963 312888
rect 411122 312666 411358 312902
rect 411442 312666 411678 312902
rect 411816 312666 412052 312902
rect 412136 312666 412372 312902
rect 412602 312681 412838 312917
rect 412922 312681 413158 312917
rect 413296 312681 413532 312917
rect 413616 312681 413852 312917
rect 414011 312695 414247 312931
rect 414331 312695 414567 312931
rect 414705 312695 414941 312931
rect 415025 312695 415261 312931
rect 415412 312710 415648 312946
rect 415732 312710 415968 312946
rect 416106 312710 416342 312946
rect 416426 312710 416662 312946
rect 416821 312724 417057 312960
rect 417141 312724 417377 312960
rect 417515 312724 417751 312960
rect 417835 312724 418071 312960
rect 407892 276604 408128 276840
rect 408287 276618 408523 276854
rect 408607 276618 408843 276854
rect 408981 276618 409217 276854
rect 409301 276618 409537 276854
rect 409688 276633 409924 276869
rect 410008 276633 410244 276869
rect 410382 276633 410618 276869
rect 410702 276633 410938 276869
rect 411097 276647 411333 276883
rect 411417 276647 411653 276883
rect 411791 276647 412027 276883
rect 412111 276647 412347 276883
rect 412577 276662 412813 276898
rect 412897 276662 413133 276898
rect 413271 276662 413507 276898
rect 413591 276662 413827 276898
rect 413986 276676 414222 276912
rect 414306 276676 414542 276912
rect 414680 276676 414916 276912
rect 415000 276676 415236 276912
rect 415387 276691 415623 276927
rect 415707 276691 415943 276927
rect 416081 276691 416317 276927
rect 416401 276691 416637 276927
rect 416796 276705 417032 276941
rect 417116 276705 417352 276941
rect 417490 276705 417726 276941
rect 417810 276705 418046 276941
rect 407878 240606 408114 240842
rect 408273 240620 408509 240856
rect 408593 240620 408829 240856
rect 408967 240620 409203 240856
rect 409287 240620 409523 240856
rect 409674 240635 409910 240871
rect 409994 240635 410230 240871
rect 410368 240635 410604 240871
rect 410688 240635 410924 240871
rect 411083 240649 411319 240885
rect 411403 240649 411639 240885
rect 411777 240649 412013 240885
rect 412097 240649 412333 240885
rect 412563 240664 412799 240900
rect 412883 240664 413119 240900
rect 413257 240664 413493 240900
rect 413577 240664 413813 240900
rect 413972 240678 414208 240914
rect 414292 240678 414528 240914
rect 414666 240678 414902 240914
rect 414986 240678 415222 240914
rect 415373 240693 415609 240929
rect 415693 240693 415929 240929
rect 416067 240693 416303 240929
rect 416387 240693 416623 240929
rect 416782 240707 417018 240943
rect 417102 240707 417338 240943
rect 417476 240707 417712 240943
rect 417796 240707 418032 240943
rect 425553 561022 425789 561258
rect 425948 561036 426184 561272
rect 426268 561036 426504 561272
rect 426642 561036 426878 561272
rect 426962 561036 427198 561272
rect 427349 561051 427585 561287
rect 427669 561051 427905 561287
rect 428043 561051 428279 561287
rect 428363 561051 428599 561287
rect 428758 561065 428994 561301
rect 429078 561065 429314 561301
rect 429452 561065 429688 561301
rect 429772 561065 430008 561301
rect 430238 561080 430474 561316
rect 430558 561080 430794 561316
rect 430932 561080 431168 561316
rect 431252 561080 431488 561316
rect 431647 561094 431883 561330
rect 431967 561094 432203 561330
rect 432341 561094 432577 561330
rect 432661 561094 432897 561330
rect 433048 561109 433284 561345
rect 433368 561109 433604 561345
rect 433742 561109 433978 561345
rect 434062 561109 434298 561345
rect 434457 561123 434693 561359
rect 434777 561123 435013 561359
rect 435151 561123 435387 561359
rect 435471 561123 435707 561359
rect 425692 525029 425928 525265
rect 426087 525043 426323 525279
rect 426407 525043 426643 525279
rect 426781 525043 427017 525279
rect 427101 525043 427337 525279
rect 427488 525058 427724 525294
rect 427808 525058 428044 525294
rect 428182 525058 428418 525294
rect 428502 525058 428738 525294
rect 428897 525072 429133 525308
rect 429217 525072 429453 525308
rect 429591 525072 429827 525308
rect 429911 525072 430147 525308
rect 430377 525087 430613 525323
rect 430697 525087 430933 525323
rect 431071 525087 431307 525323
rect 431391 525087 431627 525323
rect 431786 525101 432022 525337
rect 432106 525101 432342 525337
rect 432480 525101 432716 525337
rect 432800 525101 433036 525337
rect 433187 525116 433423 525352
rect 433507 525116 433743 525352
rect 433881 525116 434117 525352
rect 434201 525116 434437 525352
rect 434596 525130 434832 525366
rect 434916 525130 435152 525366
rect 435290 525130 435526 525366
rect 435610 525130 435846 525366
rect 425691 489036 425927 489272
rect 426086 489050 426322 489286
rect 426406 489050 426642 489286
rect 426780 489050 427016 489286
rect 427100 489050 427336 489286
rect 427487 489065 427723 489301
rect 427807 489065 428043 489301
rect 428181 489065 428417 489301
rect 428501 489065 428737 489301
rect 428896 489079 429132 489315
rect 429216 489079 429452 489315
rect 429590 489079 429826 489315
rect 429910 489079 430146 489315
rect 430376 489094 430612 489330
rect 430696 489094 430932 489330
rect 431070 489094 431306 489330
rect 431390 489094 431626 489330
rect 431785 489108 432021 489344
rect 432105 489108 432341 489344
rect 432479 489108 432715 489344
rect 432799 489108 433035 489344
rect 433186 489123 433422 489359
rect 433506 489123 433742 489359
rect 433880 489123 434116 489359
rect 434200 489123 434436 489359
rect 434595 489137 434831 489373
rect 434915 489137 435151 489373
rect 435289 489137 435525 489373
rect 435609 489137 435845 489373
rect 425698 467606 425934 467842
rect 425698 467286 425934 467522
rect 425698 466966 425934 467202
rect 426093 466980 426649 467856
rect 426787 466980 427343 467856
rect 427494 466995 428050 467871
rect 428188 466995 428744 467871
rect 428903 467009 429459 467885
rect 429597 467009 430153 467885
rect 430383 467024 430939 467900
rect 431077 467024 431633 467900
rect 431792 467038 432348 467914
rect 432486 467038 433042 467914
rect 433193 467053 433749 467929
rect 433887 467053 434443 467929
rect 434602 467067 435158 467943
rect 435296 467067 435852 467943
rect 425575 451619 425811 451855
rect 425575 451299 425811 451535
rect 425575 450979 425811 451215
rect 425970 450993 426526 451869
rect 426664 450993 427220 451869
rect 427371 451008 427927 451884
rect 428065 451008 428621 451884
rect 428780 451022 429336 451898
rect 429474 451022 430030 451898
rect 430260 451037 430816 451913
rect 430954 451037 431510 451913
rect 431669 451051 432225 451927
rect 432363 451051 432919 451927
rect 433070 451066 433626 451942
rect 433764 451066 434320 451942
rect 434479 451080 435035 451956
rect 435173 451080 435729 451956
rect 425700 443623 425936 443859
rect 425700 443303 425936 443539
rect 425700 442983 425936 443219
rect 426095 442997 426651 443873
rect 426789 442997 427345 443873
rect 427496 443012 428052 443888
rect 428190 443012 428746 443888
rect 428905 443026 429461 443902
rect 429599 443026 430155 443902
rect 430385 443041 430941 443917
rect 431079 443041 431635 443917
rect 431794 443055 432350 443931
rect 432488 443055 433044 443931
rect 433195 443070 433751 443946
rect 433889 443070 434445 443946
rect 434604 443084 435160 443960
rect 435298 443084 435854 443960
rect 425614 435590 425850 435826
rect 425614 435270 425850 435506
rect 425614 434950 425850 435186
rect 426009 434964 426565 435840
rect 426703 434964 427259 435840
rect 427410 434979 427966 435855
rect 428104 434979 428660 435855
rect 428819 434993 429375 435869
rect 429513 434993 430069 435869
rect 430299 435008 430855 435884
rect 430993 435008 431549 435884
rect 431708 435022 432264 435898
rect 432402 435022 432958 435898
rect 433109 435037 433665 435913
rect 433803 435037 434359 435913
rect 434518 435051 435074 435927
rect 435212 435051 435768 435927
rect 425617 427553 425853 427789
rect 425617 427233 425853 427469
rect 425617 426913 425853 427149
rect 426012 426927 426568 427803
rect 426706 426927 427262 427803
rect 427413 426942 427969 427818
rect 428107 426942 428663 427818
rect 428822 426956 429378 427832
rect 429516 426956 430072 427832
rect 430302 426971 430858 427847
rect 430996 426971 431552 427847
rect 431711 426985 432267 427861
rect 432405 426985 432961 427861
rect 433112 427000 433668 427876
rect 433806 427000 434362 427876
rect 434521 427014 435077 427890
rect 435215 427014 435771 427890
rect 425631 419618 425867 419854
rect 425631 419298 425867 419534
rect 425631 418978 425867 419214
rect 426026 418992 426582 419868
rect 426720 418992 427276 419868
rect 427427 419007 427983 419883
rect 428121 419007 428677 419883
rect 428836 419021 429392 419897
rect 429530 419021 430086 419897
rect 430316 419036 430872 419912
rect 431010 419036 431566 419912
rect 431725 419050 432281 419926
rect 432419 419050 432975 419926
rect 433126 419065 433682 419941
rect 433820 419065 434376 419941
rect 434535 419079 435091 419955
rect 435229 419079 435785 419955
rect 425531 411629 425767 411865
rect 425531 411309 425767 411545
rect 425531 410989 425767 411225
rect 425926 411003 426482 411879
rect 426620 411003 427176 411879
rect 427327 411018 427883 411894
rect 428021 411018 428577 411894
rect 428736 411032 429292 411908
rect 429430 411032 429986 411908
rect 430216 411047 430772 411923
rect 430910 411047 431466 411923
rect 431625 411061 432181 411937
rect 432319 411061 432875 411937
rect 433026 411076 433582 411952
rect 433720 411076 434276 411952
rect 434435 411090 434991 411966
rect 435129 411090 435685 411966
rect 425676 403604 425912 403840
rect 425676 403284 425912 403520
rect 425676 402964 425912 403200
rect 426071 402978 426627 403854
rect 426765 402978 427321 403854
rect 427472 402993 428028 403869
rect 428166 402993 428722 403869
rect 428881 403007 429437 403883
rect 429575 403007 430131 403883
rect 430361 403022 430917 403898
rect 431055 403022 431611 403898
rect 431770 403036 432326 403912
rect 432464 403036 433020 403912
rect 433171 403051 433727 403927
rect 433865 403051 434421 403927
rect 434580 403065 435136 403941
rect 435274 403065 435830 403941
rect 425656 395576 425892 395812
rect 425656 395256 425892 395492
rect 425656 394936 425892 395172
rect 426051 394950 426607 395826
rect 426745 394950 427301 395826
rect 427452 394965 428008 395841
rect 428146 394965 428702 395841
rect 428861 394979 429417 395855
rect 429555 394979 430111 395855
rect 430341 394994 430897 395870
rect 431035 394994 431591 395870
rect 431750 395008 432306 395884
rect 432444 395008 433000 395884
rect 433151 395023 433707 395899
rect 433845 395023 434401 395899
rect 434560 395037 435116 395913
rect 435254 395037 435810 395913
rect 425675 387585 425911 387821
rect 425675 387265 425911 387501
rect 425675 386945 425911 387181
rect 426070 386959 426626 387835
rect 426764 386959 427320 387835
rect 427471 386974 428027 387850
rect 428165 386974 428721 387850
rect 428880 386988 429436 387864
rect 429574 386988 430130 387864
rect 430360 387003 430916 387879
rect 431054 387003 431610 387879
rect 431769 387017 432325 387893
rect 432463 387017 433019 387893
rect 433170 387032 433726 387908
rect 433864 387032 434420 387908
rect 434579 387046 435135 387922
rect 435273 387046 435829 387922
rect 425639 379608 425875 379844
rect 425639 379288 425875 379524
rect 425639 378968 425875 379204
rect 426034 378982 426590 379858
rect 426728 378982 427284 379858
rect 427435 378997 427991 379873
rect 428129 378997 428685 379873
rect 428844 379011 429400 379887
rect 429538 379011 430094 379887
rect 430324 379026 430880 379902
rect 431018 379026 431574 379902
rect 431733 379040 432289 379916
rect 432427 379040 432983 379916
rect 433134 379055 433690 379931
rect 433828 379055 434384 379931
rect 434543 379069 435099 379945
rect 435237 379069 435793 379945
rect 425627 371620 425863 371856
rect 425627 371300 425863 371536
rect 425627 370980 425863 371216
rect 426022 370994 426578 371870
rect 426716 370994 427272 371870
rect 427423 371009 427979 371885
rect 428117 371009 428673 371885
rect 428832 371023 429388 371899
rect 429526 371023 430082 371899
rect 430312 371038 430868 371914
rect 431006 371038 431562 371914
rect 431721 371052 432277 371928
rect 432415 371052 432971 371928
rect 433122 371067 433678 371943
rect 433816 371067 434372 371943
rect 434531 371081 435087 371957
rect 435225 371081 435781 371957
rect 425615 363630 425851 363866
rect 425615 363310 425851 363546
rect 425615 362990 425851 363226
rect 426010 363004 426566 363880
rect 426704 363004 427260 363880
rect 427411 363019 427967 363895
rect 428105 363019 428661 363895
rect 428820 363033 429376 363909
rect 429514 363033 430070 363909
rect 430300 363048 430856 363924
rect 430994 363048 431550 363924
rect 431709 363062 432265 363938
rect 432403 363062 432959 363938
rect 433110 363077 433666 363953
rect 433804 363077 434360 363953
rect 434519 363091 435075 363967
rect 435213 363091 435769 363967
rect 425664 355621 425900 355857
rect 425664 355301 425900 355537
rect 425664 354981 425900 355217
rect 426059 354995 426615 355871
rect 426753 354995 427309 355871
rect 427460 355010 428016 355886
rect 428154 355010 428710 355886
rect 428869 355024 429425 355900
rect 429563 355024 430119 355900
rect 430349 355039 430905 355915
rect 431043 355039 431599 355915
rect 431758 355053 432314 355929
rect 432452 355053 433008 355929
rect 433159 355068 433715 355944
rect 433853 355068 434409 355944
rect 434568 355082 435124 355958
rect 435262 355082 435818 355958
rect 425691 347659 425927 347895
rect 425691 347339 425927 347575
rect 425691 347019 425927 347255
rect 426086 347033 426642 347909
rect 426780 347033 427336 347909
rect 427487 347048 428043 347924
rect 428181 347048 428737 347924
rect 428896 347062 429452 347938
rect 429590 347062 430146 347938
rect 430376 347077 430932 347953
rect 431070 347077 431626 347953
rect 431785 347091 432341 347967
rect 432479 347091 433035 347967
rect 433186 347106 433742 347982
rect 433880 347106 434436 347982
rect 434595 347120 435151 347996
rect 435289 347120 435845 347996
rect 425635 309034 425871 309270
rect 426030 309048 426266 309284
rect 426350 309048 426586 309284
rect 426724 309048 426960 309284
rect 427044 309048 427280 309284
rect 427431 309063 427667 309299
rect 427751 309063 427987 309299
rect 428125 309063 428361 309299
rect 428445 309063 428681 309299
rect 428840 309077 429076 309313
rect 429160 309077 429396 309313
rect 429534 309077 429770 309313
rect 429854 309077 430090 309313
rect 430320 309092 430556 309328
rect 430640 309092 430876 309328
rect 431014 309092 431250 309328
rect 431334 309092 431570 309328
rect 431729 309106 431965 309342
rect 432049 309106 432285 309342
rect 432423 309106 432659 309342
rect 432743 309106 432979 309342
rect 433130 309121 433366 309357
rect 433450 309121 433686 309357
rect 433824 309121 434060 309357
rect 434144 309121 434380 309357
rect 434539 309135 434775 309371
rect 434859 309135 435095 309371
rect 435233 309135 435469 309371
rect 435553 309135 435789 309371
rect 425686 273013 425922 273249
rect 426081 273027 426317 273263
rect 426401 273027 426637 273263
rect 426775 273027 427011 273263
rect 427095 273027 427331 273263
rect 427482 273042 427718 273278
rect 427802 273042 428038 273278
rect 428176 273042 428412 273278
rect 428496 273042 428732 273278
rect 428891 273056 429127 273292
rect 429211 273056 429447 273292
rect 429585 273056 429821 273292
rect 429905 273056 430141 273292
rect 430371 273071 430607 273307
rect 430691 273071 430927 273307
rect 431065 273071 431301 273307
rect 431385 273071 431621 273307
rect 431780 273085 432016 273321
rect 432100 273085 432336 273321
rect 432474 273085 432710 273321
rect 432794 273085 433030 273321
rect 433181 273100 433417 273336
rect 433501 273100 433737 273336
rect 433875 273100 434111 273336
rect 434195 273100 434431 273336
rect 434590 273114 434826 273350
rect 434910 273114 435146 273350
rect 435284 273114 435520 273350
rect 435604 273114 435840 273350
rect 425718 237058 425954 237294
rect 426113 237072 426349 237308
rect 426433 237072 426669 237308
rect 426807 237072 427043 237308
rect 427127 237072 427363 237308
rect 427514 237087 427750 237323
rect 427834 237087 428070 237323
rect 428208 237087 428444 237323
rect 428528 237087 428764 237323
rect 428923 237101 429159 237337
rect 429243 237101 429479 237337
rect 429617 237101 429853 237337
rect 429937 237101 430173 237337
rect 430403 237116 430639 237352
rect 430723 237116 430959 237352
rect 431097 237116 431333 237352
rect 431417 237116 431653 237352
rect 431812 237130 432048 237366
rect 432132 237130 432368 237366
rect 432506 237130 432742 237366
rect 432826 237130 433062 237366
rect 433213 237145 433449 237381
rect 433533 237145 433769 237381
rect 433907 237145 434143 237381
rect 434227 237145 434463 237381
rect 434622 237159 434858 237395
rect 434942 237159 435178 237395
rect 435316 237159 435552 237395
rect 435636 237159 435872 237395
rect 451986 561218 452222 561454
rect 451986 560898 452222 561134
rect 451986 525218 452222 525454
rect 451986 524898 452222 525134
rect 451986 489218 452222 489454
rect 451986 488898 452222 489134
rect 451986 453218 452222 453454
rect 451986 452898 452222 453134
rect 451986 417218 452222 417454
rect 451986 416898 452222 417134
rect 451986 381218 452222 381454
rect 451986 380898 452222 381134
rect 451986 345218 452222 345454
rect 451986 344898 452222 345134
rect 451986 309218 452222 309454
rect 451986 308898 452222 309134
rect 451986 273218 452222 273454
rect 451986 272898 452222 273134
rect 451986 237218 452222 237454
rect 451986 236898 452222 237134
rect 390786 212018 391022 212254
rect 390786 211698 391022 211934
rect 390786 176018 391022 176254
rect 390786 175698 391022 175934
rect 390786 140018 391022 140254
rect 390786 139698 391022 139934
rect 390786 104018 391022 104254
rect 390786 103698 391022 103934
rect 390786 68018 391022 68254
rect 390786 67698 391022 67934
rect 390786 32018 391022 32254
rect 387186 28418 387422 28654
rect 387186 28098 387422 28334
rect 387186 -5282 387422 -5046
rect 387186 -5602 387422 -5366
rect 390786 31698 391022 31934
rect 372786 -6222 373022 -5986
rect 372786 -6542 373022 -6306
rect 397986 183218 398222 183454
rect 397986 182898 398222 183134
rect 397986 147218 398222 147454
rect 397986 146898 398222 147134
rect 397986 111218 398222 111454
rect 397986 110898 398222 111134
rect 397986 75218 398222 75454
rect 397986 74898 398222 75134
rect 397986 39218 398222 39454
rect 397986 38898 398222 39134
rect 397986 3218 398222 3454
rect 397986 2898 398222 3134
rect 397986 -582 398222 -346
rect 397986 -902 398222 -666
rect 401586 186818 401822 187054
rect 401586 186498 401822 186734
rect 401586 150818 401822 151054
rect 401586 150498 401822 150734
rect 401586 114818 401822 115054
rect 401586 114498 401822 114734
rect 401586 78818 401822 79054
rect 401586 78498 401822 78734
rect 401586 42818 401822 43054
rect 401586 42498 401822 42734
rect 401586 6818 401822 7054
rect 401586 6498 401822 6734
rect 401586 -2462 401822 -2226
rect 401586 -2782 401822 -2546
rect 405186 190418 405422 190654
rect 405186 190098 405422 190334
rect 405186 154418 405422 154654
rect 405186 154098 405422 154334
rect 405186 118418 405422 118654
rect 405186 118098 405422 118334
rect 405186 82418 405422 82654
rect 405186 82098 405422 82334
rect 405186 46418 405422 46654
rect 405186 46098 405422 46334
rect 405186 10418 405422 10654
rect 405186 10098 405422 10334
rect 405186 -4342 405422 -4106
rect 405186 -4662 405422 -4426
rect 408786 194018 409022 194254
rect 408786 193698 409022 193934
rect 408786 158018 409022 158254
rect 408786 157698 409022 157934
rect 408786 122018 409022 122254
rect 408786 121698 409022 121934
rect 408786 86018 409022 86254
rect 408786 85698 409022 85934
rect 408786 50018 409022 50254
rect 408786 49698 409022 49934
rect 408786 14018 409022 14254
rect 408786 13698 409022 13934
rect 390786 -7162 391022 -6926
rect 390786 -7482 391022 -7246
rect 415986 201218 416222 201454
rect 415986 200898 416222 201134
rect 415986 165218 416222 165454
rect 415986 164898 416222 165134
rect 415986 129218 416222 129454
rect 415986 128898 416222 129134
rect 415986 93218 416222 93454
rect 415986 92898 416222 93134
rect 415986 57218 416222 57454
rect 415986 56898 416222 57134
rect 415986 21218 416222 21454
rect 415986 20898 416222 21134
rect 415986 -1522 416222 -1286
rect 415986 -1842 416222 -1606
rect 419586 204818 419822 205054
rect 419586 204498 419822 204734
rect 419586 168818 419822 169054
rect 419586 168498 419822 168734
rect 419586 132818 419822 133054
rect 419586 132498 419822 132734
rect 419586 96818 419822 97054
rect 419586 96498 419822 96734
rect 419586 60818 419822 61054
rect 419586 60498 419822 60734
rect 419586 24818 419822 25054
rect 419586 24498 419822 24734
rect 419586 -3402 419822 -3166
rect 419586 -3722 419822 -3486
rect 423186 208418 423422 208654
rect 423186 208098 423422 208334
rect 423186 172418 423422 172654
rect 423186 172098 423422 172334
rect 423186 136418 423422 136654
rect 423186 136098 423422 136334
rect 423186 100418 423422 100654
rect 423186 100098 423422 100334
rect 423186 64418 423422 64654
rect 423186 64098 423422 64334
rect 423186 28418 423422 28654
rect 423186 28098 423422 28334
rect 423186 -5282 423422 -5046
rect 423186 -5602 423422 -5366
rect 426786 212018 427022 212254
rect 426786 211698 427022 211934
rect 426786 176018 427022 176254
rect 426786 175698 427022 175934
rect 426786 140018 427022 140254
rect 426786 139698 427022 139934
rect 426786 104018 427022 104254
rect 426786 103698 427022 103934
rect 426786 68018 427022 68254
rect 426786 67698 427022 67934
rect 426786 32018 427022 32254
rect 426786 31698 427022 31934
rect 408786 -6222 409022 -5986
rect 408786 -6542 409022 -6306
rect 433986 183218 434222 183454
rect 433986 182898 434222 183134
rect 433986 147218 434222 147454
rect 433986 146898 434222 147134
rect 433986 111218 434222 111454
rect 433986 110898 434222 111134
rect 433986 75218 434222 75454
rect 433986 74898 434222 75134
rect 433986 39218 434222 39454
rect 433986 38898 434222 39134
rect 433986 3218 434222 3454
rect 433986 2898 434222 3134
rect 433986 -582 434222 -346
rect 433986 -902 434222 -666
rect 437586 186818 437822 187054
rect 437586 186498 437822 186734
rect 437586 150818 437822 151054
rect 437586 150498 437822 150734
rect 437586 114818 437822 115054
rect 437586 114498 437822 114734
rect 437586 78818 437822 79054
rect 437586 78498 437822 78734
rect 437586 42818 437822 43054
rect 437586 42498 437822 42734
rect 437586 6818 437822 7054
rect 437586 6498 437822 6734
rect 437586 -2462 437822 -2226
rect 437586 -2782 437822 -2546
rect 441186 190418 441422 190654
rect 441186 190098 441422 190334
rect 441186 154418 441422 154654
rect 441186 154098 441422 154334
rect 441186 118418 441422 118654
rect 441186 118098 441422 118334
rect 441186 82418 441422 82654
rect 441186 82098 441422 82334
rect 441186 46418 441422 46654
rect 441186 46098 441422 46334
rect 441186 10418 441422 10654
rect 441186 10098 441422 10334
rect 441186 -4342 441422 -4106
rect 441186 -4662 441422 -4426
rect 444786 194018 445022 194254
rect 444786 193698 445022 193934
rect 444786 158018 445022 158254
rect 444786 157698 445022 157934
rect 444786 122018 445022 122254
rect 444786 121698 445022 121934
rect 444786 86018 445022 86254
rect 444786 85698 445022 85934
rect 444786 50018 445022 50254
rect 444786 49698 445022 49934
rect 444786 14018 445022 14254
rect 444786 13698 445022 13934
rect 426786 -7162 427022 -6926
rect 426786 -7482 427022 -7246
rect 451986 201218 452222 201454
rect 451986 200898 452222 201134
rect 451986 165218 452222 165454
rect 451986 164898 452222 165134
rect 451986 129218 452222 129454
rect 451986 128898 452222 129134
rect 451986 93218 452222 93454
rect 451986 92898 452222 93134
rect 451986 57218 452222 57454
rect 451986 56898 452222 57134
rect 451986 21218 452222 21454
rect 451986 20898 452222 21134
rect 451986 -1522 452222 -1286
rect 451986 -1842 452222 -1606
rect 455586 672818 455822 673054
rect 455586 672498 455822 672734
rect 455586 636818 455822 637054
rect 455586 636498 455822 636734
rect 455586 600818 455822 601054
rect 455586 600498 455822 600734
rect 455586 564818 455822 565054
rect 455586 564498 455822 564734
rect 455586 528818 455822 529054
rect 455586 528498 455822 528734
rect 455586 492818 455822 493054
rect 455586 492498 455822 492734
rect 455586 456818 455822 457054
rect 455586 456498 455822 456734
rect 455586 420818 455822 421054
rect 455586 420498 455822 420734
rect 455586 384818 455822 385054
rect 455586 384498 455822 384734
rect 455586 348818 455822 349054
rect 455586 348498 455822 348734
rect 455586 312818 455822 313054
rect 455586 312498 455822 312734
rect 455586 276818 455822 277054
rect 455586 276498 455822 276734
rect 455586 240818 455822 241054
rect 455586 240498 455822 240734
rect 455586 204818 455822 205054
rect 455586 204498 455822 204734
rect 455586 168818 455822 169054
rect 455586 168498 455822 168734
rect 455586 132818 455822 133054
rect 455586 132498 455822 132734
rect 455586 96818 455822 97054
rect 455586 96498 455822 96734
rect 455586 60818 455822 61054
rect 455586 60498 455822 60734
rect 455586 24818 455822 25054
rect 455586 24498 455822 24734
rect 455586 -3402 455822 -3166
rect 455586 -3722 455822 -3486
rect 459186 676418 459422 676654
rect 459186 676098 459422 676334
rect 459186 640418 459422 640654
rect 459186 640098 459422 640334
rect 459186 604418 459422 604654
rect 459186 604098 459422 604334
rect 459186 568418 459422 568654
rect 459186 568098 459422 568334
rect 459186 532418 459422 532654
rect 459186 532098 459422 532334
rect 459186 496418 459422 496654
rect 459186 496098 459422 496334
rect 459186 460418 459422 460654
rect 459186 460098 459422 460334
rect 459186 424418 459422 424654
rect 459186 424098 459422 424334
rect 459186 388418 459422 388654
rect 459186 388098 459422 388334
rect 459186 352418 459422 352654
rect 459186 352098 459422 352334
rect 459186 316418 459422 316654
rect 459186 316098 459422 316334
rect 459186 280418 459422 280654
rect 459186 280098 459422 280334
rect 459186 244418 459422 244654
rect 459186 244098 459422 244334
rect 459186 208418 459422 208654
rect 459186 208098 459422 208334
rect 459186 172418 459422 172654
rect 459186 172098 459422 172334
rect 459186 136418 459422 136654
rect 459186 136098 459422 136334
rect 459186 100418 459422 100654
rect 459186 100098 459422 100334
rect 459186 64418 459422 64654
rect 459186 64098 459422 64334
rect 459186 28418 459422 28654
rect 459186 28098 459422 28334
rect 459186 -5282 459422 -5046
rect 459186 -5602 459422 -5366
rect 480786 710242 481022 710478
rect 480786 709922 481022 710158
rect 477186 708362 477422 708598
rect 477186 708042 477422 708278
rect 473586 706482 473822 706718
rect 473586 706162 473822 706398
rect 462786 680018 463022 680254
rect 462786 679698 463022 679934
rect 462786 644018 463022 644254
rect 462786 643698 463022 643934
rect 462786 608018 463022 608254
rect 462786 607698 463022 607934
rect 462786 572018 463022 572254
rect 462786 571698 463022 571934
rect 462786 536018 463022 536254
rect 462786 535698 463022 535934
rect 462786 500018 463022 500254
rect 462786 499698 463022 499934
rect 462786 464018 463022 464254
rect 462786 463698 463022 463934
rect 462786 428018 463022 428254
rect 462786 427698 463022 427934
rect 462786 392018 463022 392254
rect 462786 391698 463022 391934
rect 462786 356018 463022 356254
rect 462786 355698 463022 355934
rect 462786 320018 463022 320254
rect 462786 319698 463022 319934
rect 462786 284018 463022 284254
rect 462786 283698 463022 283934
rect 462786 248018 463022 248254
rect 462786 247698 463022 247934
rect 462786 212018 463022 212254
rect 462786 211698 463022 211934
rect 462786 176018 463022 176254
rect 462786 175698 463022 175934
rect 462786 140018 463022 140254
rect 462786 139698 463022 139934
rect 462786 104018 463022 104254
rect 462786 103698 463022 103934
rect 462786 68018 463022 68254
rect 462786 67698 463022 67934
rect 462786 32018 463022 32254
rect 462786 31698 463022 31934
rect 444786 -6222 445022 -5986
rect 444786 -6542 445022 -6306
rect 469986 704602 470222 704838
rect 469986 704282 470222 704518
rect 469986 687218 470222 687454
rect 469986 686898 470222 687134
rect 469986 651218 470222 651454
rect 469986 650898 470222 651134
rect 469986 615218 470222 615454
rect 469986 614898 470222 615134
rect 469986 579218 470222 579454
rect 469986 578898 470222 579134
rect 469986 543218 470222 543454
rect 469986 542898 470222 543134
rect 469986 507218 470222 507454
rect 469986 506898 470222 507134
rect 469986 471218 470222 471454
rect 469986 470898 470222 471134
rect 469986 435218 470222 435454
rect 469986 434898 470222 435134
rect 469986 399218 470222 399454
rect 469986 398898 470222 399134
rect 469986 363218 470222 363454
rect 469986 362898 470222 363134
rect 469986 327218 470222 327454
rect 469986 326898 470222 327134
rect 469986 291218 470222 291454
rect 469986 290898 470222 291134
rect 469986 255218 470222 255454
rect 469986 254898 470222 255134
rect 469986 219218 470222 219454
rect 469986 218898 470222 219134
rect 469986 183218 470222 183454
rect 469986 182898 470222 183134
rect 469986 147218 470222 147454
rect 469986 146898 470222 147134
rect 469986 111218 470222 111454
rect 469986 110898 470222 111134
rect 469986 75218 470222 75454
rect 469986 74898 470222 75134
rect 469986 39218 470222 39454
rect 469986 38898 470222 39134
rect 469986 3218 470222 3454
rect 469986 2898 470222 3134
rect 469986 -582 470222 -346
rect 469986 -902 470222 -666
rect 473586 690818 473822 691054
rect 473586 690498 473822 690734
rect 473586 654818 473822 655054
rect 473586 654498 473822 654734
rect 473586 618818 473822 619054
rect 473586 618498 473822 618734
rect 473586 582818 473822 583054
rect 473586 582498 473822 582734
rect 473586 546818 473822 547054
rect 473586 546498 473822 546734
rect 473586 510818 473822 511054
rect 473586 510498 473822 510734
rect 473586 474818 473822 475054
rect 473586 474498 473822 474734
rect 473586 438818 473822 439054
rect 473586 438498 473822 438734
rect 473586 402818 473822 403054
rect 473586 402498 473822 402734
rect 473586 366818 473822 367054
rect 473586 366498 473822 366734
rect 473586 330818 473822 331054
rect 473586 330498 473822 330734
rect 473586 294818 473822 295054
rect 473586 294498 473822 294734
rect 473586 258818 473822 259054
rect 473586 258498 473822 258734
rect 473586 222818 473822 223054
rect 473586 222498 473822 222734
rect 473586 186818 473822 187054
rect 473586 186498 473822 186734
rect 473586 150818 473822 151054
rect 473586 150498 473822 150734
rect 473586 114818 473822 115054
rect 473586 114498 473822 114734
rect 473586 78818 473822 79054
rect 473586 78498 473822 78734
rect 473586 42818 473822 43054
rect 473586 42498 473822 42734
rect 473586 6818 473822 7054
rect 473586 6498 473822 6734
rect 473586 -2462 473822 -2226
rect 473586 -2782 473822 -2546
rect 477186 694418 477422 694654
rect 477186 694098 477422 694334
rect 477186 658418 477422 658654
rect 477186 658098 477422 658334
rect 477186 622418 477422 622654
rect 477186 622098 477422 622334
rect 477186 586418 477422 586654
rect 477186 586098 477422 586334
rect 477186 550418 477422 550654
rect 477186 550098 477422 550334
rect 477186 514418 477422 514654
rect 477186 514098 477422 514334
rect 477186 478418 477422 478654
rect 477186 478098 477422 478334
rect 477186 442418 477422 442654
rect 477186 442098 477422 442334
rect 477186 406418 477422 406654
rect 477186 406098 477422 406334
rect 477186 370418 477422 370654
rect 477186 370098 477422 370334
rect 477186 334418 477422 334654
rect 477186 334098 477422 334334
rect 477186 298418 477422 298654
rect 477186 298098 477422 298334
rect 477186 262418 477422 262654
rect 477186 262098 477422 262334
rect 477186 226418 477422 226654
rect 477186 226098 477422 226334
rect 477186 190418 477422 190654
rect 477186 190098 477422 190334
rect 477186 154418 477422 154654
rect 477186 154098 477422 154334
rect 477186 118418 477422 118654
rect 477186 118098 477422 118334
rect 477186 82418 477422 82654
rect 477186 82098 477422 82334
rect 477186 46418 477422 46654
rect 477186 46098 477422 46334
rect 477186 10418 477422 10654
rect 477186 10098 477422 10334
rect 477186 -4342 477422 -4106
rect 477186 -4662 477422 -4426
rect 498786 711182 499022 711418
rect 498786 710862 499022 711098
rect 495186 709302 495422 709538
rect 495186 708982 495422 709218
rect 491586 707422 491822 707658
rect 491586 707102 491822 707338
rect 480786 698018 481022 698254
rect 480786 697698 481022 697934
rect 480786 662018 481022 662254
rect 480786 661698 481022 661934
rect 480786 626018 481022 626254
rect 480786 625698 481022 625934
rect 480786 590018 481022 590254
rect 480786 589698 481022 589934
rect 480786 554018 481022 554254
rect 480786 553698 481022 553934
rect 480786 518018 481022 518254
rect 480786 517698 481022 517934
rect 480786 482018 481022 482254
rect 480786 481698 481022 481934
rect 480786 446018 481022 446254
rect 480786 445698 481022 445934
rect 480786 410018 481022 410254
rect 480786 409698 481022 409934
rect 480786 374018 481022 374254
rect 480786 373698 481022 373934
rect 480786 338018 481022 338254
rect 480786 337698 481022 337934
rect 480786 302018 481022 302254
rect 480786 301698 481022 301934
rect 480786 266018 481022 266254
rect 480786 265698 481022 265934
rect 480786 230018 481022 230254
rect 480786 229698 481022 229934
rect 480786 194018 481022 194254
rect 480786 193698 481022 193934
rect 480786 158018 481022 158254
rect 480786 157698 481022 157934
rect 480786 122018 481022 122254
rect 480786 121698 481022 121934
rect 480786 86018 481022 86254
rect 480786 85698 481022 85934
rect 480786 50018 481022 50254
rect 480786 49698 481022 49934
rect 480786 14018 481022 14254
rect 480786 13698 481022 13934
rect 462786 -7162 463022 -6926
rect 462786 -7482 463022 -7246
rect 487986 705542 488222 705778
rect 487986 705222 488222 705458
rect 487986 669218 488222 669454
rect 487986 668898 488222 669134
rect 487986 633218 488222 633454
rect 487986 632898 488222 633134
rect 487986 597218 488222 597454
rect 487986 596898 488222 597134
rect 487986 561218 488222 561454
rect 487986 560898 488222 561134
rect 487986 525218 488222 525454
rect 487986 524898 488222 525134
rect 487986 489218 488222 489454
rect 487986 488898 488222 489134
rect 487986 453218 488222 453454
rect 487986 452898 488222 453134
rect 487986 417218 488222 417454
rect 487986 416898 488222 417134
rect 487986 381218 488222 381454
rect 487986 380898 488222 381134
rect 487986 345218 488222 345454
rect 487986 344898 488222 345134
rect 487986 309218 488222 309454
rect 487986 308898 488222 309134
rect 487986 273218 488222 273454
rect 487986 272898 488222 273134
rect 487986 237218 488222 237454
rect 487986 236898 488222 237134
rect 487986 201218 488222 201454
rect 487986 200898 488222 201134
rect 487986 165218 488222 165454
rect 487986 164898 488222 165134
rect 487986 129218 488222 129454
rect 487986 128898 488222 129134
rect 487986 93218 488222 93454
rect 487986 92898 488222 93134
rect 487986 57218 488222 57454
rect 487986 56898 488222 57134
rect 487986 21218 488222 21454
rect 487986 20898 488222 21134
rect 487986 -1522 488222 -1286
rect 487986 -1842 488222 -1606
rect 491586 672818 491822 673054
rect 491586 672498 491822 672734
rect 491586 636818 491822 637054
rect 491586 636498 491822 636734
rect 491586 600818 491822 601054
rect 491586 600498 491822 600734
rect 491586 564818 491822 565054
rect 491586 564498 491822 564734
rect 491586 528818 491822 529054
rect 491586 528498 491822 528734
rect 491586 492818 491822 493054
rect 491586 492498 491822 492734
rect 491586 456818 491822 457054
rect 491586 456498 491822 456734
rect 491586 420818 491822 421054
rect 491586 420498 491822 420734
rect 491586 384818 491822 385054
rect 491586 384498 491822 384734
rect 491586 348818 491822 349054
rect 491586 348498 491822 348734
rect 491586 312818 491822 313054
rect 491586 312498 491822 312734
rect 491586 276818 491822 277054
rect 491586 276498 491822 276734
rect 491586 240818 491822 241054
rect 491586 240498 491822 240734
rect 491586 204818 491822 205054
rect 491586 204498 491822 204734
rect 491586 168818 491822 169054
rect 491586 168498 491822 168734
rect 491586 132818 491822 133054
rect 491586 132498 491822 132734
rect 491586 96818 491822 97054
rect 491586 96498 491822 96734
rect 491586 60818 491822 61054
rect 491586 60498 491822 60734
rect 491586 24818 491822 25054
rect 491586 24498 491822 24734
rect 491586 -3402 491822 -3166
rect 491586 -3722 491822 -3486
rect 495186 676418 495422 676654
rect 495186 676098 495422 676334
rect 495186 640418 495422 640654
rect 495186 640098 495422 640334
rect 495186 604418 495422 604654
rect 495186 604098 495422 604334
rect 495186 568418 495422 568654
rect 495186 568098 495422 568334
rect 495186 532418 495422 532654
rect 495186 532098 495422 532334
rect 495186 496418 495422 496654
rect 495186 496098 495422 496334
rect 495186 460418 495422 460654
rect 495186 460098 495422 460334
rect 495186 424418 495422 424654
rect 495186 424098 495422 424334
rect 495186 388418 495422 388654
rect 495186 388098 495422 388334
rect 495186 352418 495422 352654
rect 495186 352098 495422 352334
rect 495186 316418 495422 316654
rect 495186 316098 495422 316334
rect 495186 280418 495422 280654
rect 495186 280098 495422 280334
rect 495186 244418 495422 244654
rect 495186 244098 495422 244334
rect 495186 208418 495422 208654
rect 495186 208098 495422 208334
rect 495186 172418 495422 172654
rect 495186 172098 495422 172334
rect 495186 136418 495422 136654
rect 495186 136098 495422 136334
rect 495186 100418 495422 100654
rect 495186 100098 495422 100334
rect 495186 64418 495422 64654
rect 495186 64098 495422 64334
rect 495186 28418 495422 28654
rect 495186 28098 495422 28334
rect 495186 -5282 495422 -5046
rect 495186 -5602 495422 -5366
rect 516786 710242 517022 710478
rect 516786 709922 517022 710158
rect 513186 708362 513422 708598
rect 513186 708042 513422 708278
rect 509586 706482 509822 706718
rect 509586 706162 509822 706398
rect 498786 680018 499022 680254
rect 498786 679698 499022 679934
rect 498786 644018 499022 644254
rect 498786 643698 499022 643934
rect 498786 608018 499022 608254
rect 498786 607698 499022 607934
rect 498786 572018 499022 572254
rect 498786 571698 499022 571934
rect 498786 536018 499022 536254
rect 498786 535698 499022 535934
rect 498786 500018 499022 500254
rect 498786 499698 499022 499934
rect 498786 464018 499022 464254
rect 498786 463698 499022 463934
rect 498786 428018 499022 428254
rect 498786 427698 499022 427934
rect 498786 392018 499022 392254
rect 498786 391698 499022 391934
rect 498786 356018 499022 356254
rect 498786 355698 499022 355934
rect 498786 320018 499022 320254
rect 498786 319698 499022 319934
rect 498786 284018 499022 284254
rect 498786 283698 499022 283934
rect 498786 248018 499022 248254
rect 498786 247698 499022 247934
rect 498786 212018 499022 212254
rect 498786 211698 499022 211934
rect 498786 176018 499022 176254
rect 498786 175698 499022 175934
rect 498786 140018 499022 140254
rect 498786 139698 499022 139934
rect 498786 104018 499022 104254
rect 498786 103698 499022 103934
rect 498786 68018 499022 68254
rect 498786 67698 499022 67934
rect 498786 32018 499022 32254
rect 498786 31698 499022 31934
rect 480786 -6222 481022 -5986
rect 480786 -6542 481022 -6306
rect 505986 704602 506222 704838
rect 505986 704282 506222 704518
rect 505986 687218 506222 687454
rect 505986 686898 506222 687134
rect 505986 651218 506222 651454
rect 505986 650898 506222 651134
rect 505986 615218 506222 615454
rect 505986 614898 506222 615134
rect 505986 579218 506222 579454
rect 505986 578898 506222 579134
rect 505986 543218 506222 543454
rect 505986 542898 506222 543134
rect 505986 507218 506222 507454
rect 505986 506898 506222 507134
rect 505986 471218 506222 471454
rect 505986 470898 506222 471134
rect 505986 435218 506222 435454
rect 505986 434898 506222 435134
rect 505986 399218 506222 399454
rect 505986 398898 506222 399134
rect 505986 363218 506222 363454
rect 505986 362898 506222 363134
rect 505986 327218 506222 327454
rect 505986 326898 506222 327134
rect 505986 291218 506222 291454
rect 505986 290898 506222 291134
rect 505986 255218 506222 255454
rect 505986 254898 506222 255134
rect 505986 219218 506222 219454
rect 505986 218898 506222 219134
rect 505986 183218 506222 183454
rect 505986 182898 506222 183134
rect 505986 147218 506222 147454
rect 505986 146898 506222 147134
rect 505986 111218 506222 111454
rect 505986 110898 506222 111134
rect 505986 75218 506222 75454
rect 505986 74898 506222 75134
rect 505986 39218 506222 39454
rect 505986 38898 506222 39134
rect 505986 3218 506222 3454
rect 505986 2898 506222 3134
rect 505986 -582 506222 -346
rect 505986 -902 506222 -666
rect 509586 690818 509822 691054
rect 509586 690498 509822 690734
rect 509586 654818 509822 655054
rect 509586 654498 509822 654734
rect 509586 618818 509822 619054
rect 509586 618498 509822 618734
rect 509586 582818 509822 583054
rect 509586 582498 509822 582734
rect 509586 546818 509822 547054
rect 509586 546498 509822 546734
rect 509586 510818 509822 511054
rect 509586 510498 509822 510734
rect 509586 474818 509822 475054
rect 509586 474498 509822 474734
rect 509586 438818 509822 439054
rect 509586 438498 509822 438734
rect 509586 402818 509822 403054
rect 509586 402498 509822 402734
rect 509586 366818 509822 367054
rect 509586 366498 509822 366734
rect 509586 330818 509822 331054
rect 509586 330498 509822 330734
rect 509586 294818 509822 295054
rect 509586 294498 509822 294734
rect 509586 258818 509822 259054
rect 509586 258498 509822 258734
rect 509586 222818 509822 223054
rect 509586 222498 509822 222734
rect 509586 186818 509822 187054
rect 509586 186498 509822 186734
rect 509586 150818 509822 151054
rect 509586 150498 509822 150734
rect 509586 114818 509822 115054
rect 509586 114498 509822 114734
rect 509586 78818 509822 79054
rect 509586 78498 509822 78734
rect 509586 42818 509822 43054
rect 509586 42498 509822 42734
rect 509586 6818 509822 7054
rect 509586 6498 509822 6734
rect 509586 -2462 509822 -2226
rect 509586 -2782 509822 -2546
rect 513186 694418 513422 694654
rect 513186 694098 513422 694334
rect 513186 658418 513422 658654
rect 513186 658098 513422 658334
rect 513186 622418 513422 622654
rect 513186 622098 513422 622334
rect 513186 586418 513422 586654
rect 513186 586098 513422 586334
rect 513186 550418 513422 550654
rect 513186 550098 513422 550334
rect 513186 514418 513422 514654
rect 513186 514098 513422 514334
rect 513186 478418 513422 478654
rect 513186 478098 513422 478334
rect 513186 442418 513422 442654
rect 513186 442098 513422 442334
rect 513186 406418 513422 406654
rect 513186 406098 513422 406334
rect 513186 370418 513422 370654
rect 513186 370098 513422 370334
rect 513186 334418 513422 334654
rect 513186 334098 513422 334334
rect 513186 298418 513422 298654
rect 513186 298098 513422 298334
rect 513186 262418 513422 262654
rect 513186 262098 513422 262334
rect 513186 226418 513422 226654
rect 513186 226098 513422 226334
rect 513186 190418 513422 190654
rect 513186 190098 513422 190334
rect 513186 154418 513422 154654
rect 513186 154098 513422 154334
rect 513186 118418 513422 118654
rect 513186 118098 513422 118334
rect 513186 82418 513422 82654
rect 513186 82098 513422 82334
rect 513186 46418 513422 46654
rect 513186 46098 513422 46334
rect 513186 10418 513422 10654
rect 513186 10098 513422 10334
rect 513186 -4342 513422 -4106
rect 513186 -4662 513422 -4426
rect 534786 711182 535022 711418
rect 534786 710862 535022 711098
rect 531186 709302 531422 709538
rect 531186 708982 531422 709218
rect 527586 707422 527822 707658
rect 527586 707102 527822 707338
rect 516786 698018 517022 698254
rect 516786 697698 517022 697934
rect 516786 662018 517022 662254
rect 516786 661698 517022 661934
rect 516786 626018 517022 626254
rect 516786 625698 517022 625934
rect 516786 590018 517022 590254
rect 516786 589698 517022 589934
rect 516786 554018 517022 554254
rect 516786 553698 517022 553934
rect 516786 518018 517022 518254
rect 516786 517698 517022 517934
rect 516786 482018 517022 482254
rect 516786 481698 517022 481934
rect 516786 446018 517022 446254
rect 516786 445698 517022 445934
rect 516786 410018 517022 410254
rect 516786 409698 517022 409934
rect 516786 374018 517022 374254
rect 516786 373698 517022 373934
rect 516786 338018 517022 338254
rect 516786 337698 517022 337934
rect 516786 302018 517022 302254
rect 516786 301698 517022 301934
rect 516786 266018 517022 266254
rect 516786 265698 517022 265934
rect 516786 230018 517022 230254
rect 516786 229698 517022 229934
rect 516786 194018 517022 194254
rect 516786 193698 517022 193934
rect 516786 158018 517022 158254
rect 516786 157698 517022 157934
rect 516786 122018 517022 122254
rect 516786 121698 517022 121934
rect 516786 86018 517022 86254
rect 516786 85698 517022 85934
rect 516786 50018 517022 50254
rect 516786 49698 517022 49934
rect 516786 14018 517022 14254
rect 516786 13698 517022 13934
rect 498786 -7162 499022 -6926
rect 498786 -7482 499022 -7246
rect 523986 705542 524222 705778
rect 523986 705222 524222 705458
rect 523986 669218 524222 669454
rect 523986 668898 524222 669134
rect 523986 633218 524222 633454
rect 523986 632898 524222 633134
rect 523986 597218 524222 597454
rect 523986 596898 524222 597134
rect 523986 561218 524222 561454
rect 523986 560898 524222 561134
rect 523986 525218 524222 525454
rect 523986 524898 524222 525134
rect 523986 489218 524222 489454
rect 523986 488898 524222 489134
rect 523986 453218 524222 453454
rect 523986 452898 524222 453134
rect 523986 417218 524222 417454
rect 523986 416898 524222 417134
rect 523986 381218 524222 381454
rect 523986 380898 524222 381134
rect 523986 345218 524222 345454
rect 523986 344898 524222 345134
rect 523986 309218 524222 309454
rect 523986 308898 524222 309134
rect 523986 273218 524222 273454
rect 523986 272898 524222 273134
rect 523986 237218 524222 237454
rect 523986 236898 524222 237134
rect 523986 201218 524222 201454
rect 523986 200898 524222 201134
rect 523986 165218 524222 165454
rect 523986 164898 524222 165134
rect 523986 129218 524222 129454
rect 523986 128898 524222 129134
rect 523986 93218 524222 93454
rect 523986 92898 524222 93134
rect 523986 57218 524222 57454
rect 523986 56898 524222 57134
rect 523986 21218 524222 21454
rect 523986 20898 524222 21134
rect 523986 -1522 524222 -1286
rect 523986 -1842 524222 -1606
rect 527586 672818 527822 673054
rect 527586 672498 527822 672734
rect 527586 636818 527822 637054
rect 527586 636498 527822 636734
rect 527586 600818 527822 601054
rect 527586 600498 527822 600734
rect 527586 564818 527822 565054
rect 527586 564498 527822 564734
rect 527586 528818 527822 529054
rect 527586 528498 527822 528734
rect 527586 492818 527822 493054
rect 527586 492498 527822 492734
rect 527586 456818 527822 457054
rect 527586 456498 527822 456734
rect 527586 420818 527822 421054
rect 527586 420498 527822 420734
rect 527586 384818 527822 385054
rect 527586 384498 527822 384734
rect 527586 348818 527822 349054
rect 527586 348498 527822 348734
rect 527586 312818 527822 313054
rect 527586 312498 527822 312734
rect 527586 276818 527822 277054
rect 527586 276498 527822 276734
rect 527586 240818 527822 241054
rect 527586 240498 527822 240734
rect 527586 204818 527822 205054
rect 527586 204498 527822 204734
rect 527586 168818 527822 169054
rect 527586 168498 527822 168734
rect 527586 132818 527822 133054
rect 527586 132498 527822 132734
rect 527586 96818 527822 97054
rect 527586 96498 527822 96734
rect 527586 60818 527822 61054
rect 527586 60498 527822 60734
rect 527586 24818 527822 25054
rect 527586 24498 527822 24734
rect 527586 -3402 527822 -3166
rect 527586 -3722 527822 -3486
rect 531186 676418 531422 676654
rect 531186 676098 531422 676334
rect 531186 640418 531422 640654
rect 531186 640098 531422 640334
rect 531186 604418 531422 604654
rect 531186 604098 531422 604334
rect 531186 568418 531422 568654
rect 531186 568098 531422 568334
rect 531186 532418 531422 532654
rect 531186 532098 531422 532334
rect 531186 496418 531422 496654
rect 531186 496098 531422 496334
rect 531186 460418 531422 460654
rect 531186 460098 531422 460334
rect 531186 424418 531422 424654
rect 531186 424098 531422 424334
rect 531186 388418 531422 388654
rect 531186 388098 531422 388334
rect 531186 352418 531422 352654
rect 531186 352098 531422 352334
rect 531186 316418 531422 316654
rect 531186 316098 531422 316334
rect 531186 280418 531422 280654
rect 531186 280098 531422 280334
rect 531186 244418 531422 244654
rect 531186 244098 531422 244334
rect 531186 208418 531422 208654
rect 531186 208098 531422 208334
rect 531186 172418 531422 172654
rect 531186 172098 531422 172334
rect 531186 136418 531422 136654
rect 531186 136098 531422 136334
rect 531186 100418 531422 100654
rect 531186 100098 531422 100334
rect 531186 64418 531422 64654
rect 531186 64098 531422 64334
rect 531186 28418 531422 28654
rect 531186 28098 531422 28334
rect 531186 -5282 531422 -5046
rect 531186 -5602 531422 -5366
rect 552786 710242 553022 710478
rect 552786 709922 553022 710158
rect 549186 708362 549422 708598
rect 549186 708042 549422 708278
rect 545586 706482 545822 706718
rect 545586 706162 545822 706398
rect 534786 680018 535022 680254
rect 534786 679698 535022 679934
rect 534786 644018 535022 644254
rect 534786 643698 535022 643934
rect 534786 608018 535022 608254
rect 534786 607698 535022 607934
rect 534786 572018 535022 572254
rect 534786 571698 535022 571934
rect 534786 536018 535022 536254
rect 534786 535698 535022 535934
rect 534786 500018 535022 500254
rect 534786 499698 535022 499934
rect 534786 464018 535022 464254
rect 534786 463698 535022 463934
rect 534786 428018 535022 428254
rect 534786 427698 535022 427934
rect 534786 392018 535022 392254
rect 534786 391698 535022 391934
rect 534786 356018 535022 356254
rect 534786 355698 535022 355934
rect 534786 320018 535022 320254
rect 534786 319698 535022 319934
rect 534786 284018 535022 284254
rect 534786 283698 535022 283934
rect 534786 248018 535022 248254
rect 534786 247698 535022 247934
rect 534786 212018 535022 212254
rect 534786 211698 535022 211934
rect 534786 176018 535022 176254
rect 534786 175698 535022 175934
rect 534786 140018 535022 140254
rect 534786 139698 535022 139934
rect 534786 104018 535022 104254
rect 534786 103698 535022 103934
rect 534786 68018 535022 68254
rect 534786 67698 535022 67934
rect 534786 32018 535022 32254
rect 534786 31698 535022 31934
rect 516786 -6222 517022 -5986
rect 516786 -6542 517022 -6306
rect 541986 704602 542222 704838
rect 541986 704282 542222 704518
rect 541986 687218 542222 687454
rect 541986 686898 542222 687134
rect 541986 651218 542222 651454
rect 541986 650898 542222 651134
rect 541986 615218 542222 615454
rect 541986 614898 542222 615134
rect 541986 579218 542222 579454
rect 541986 578898 542222 579134
rect 541986 543218 542222 543454
rect 541986 542898 542222 543134
rect 541986 507218 542222 507454
rect 541986 506898 542222 507134
rect 541986 471218 542222 471454
rect 541986 470898 542222 471134
rect 541986 435218 542222 435454
rect 541986 434898 542222 435134
rect 541986 399218 542222 399454
rect 541986 398898 542222 399134
rect 541986 363218 542222 363454
rect 541986 362898 542222 363134
rect 541986 327218 542222 327454
rect 541986 326898 542222 327134
rect 541986 291218 542222 291454
rect 541986 290898 542222 291134
rect 541986 255218 542222 255454
rect 541986 254898 542222 255134
rect 541986 219218 542222 219454
rect 541986 218898 542222 219134
rect 541986 183218 542222 183454
rect 541986 182898 542222 183134
rect 541986 147218 542222 147454
rect 541986 146898 542222 147134
rect 541986 111218 542222 111454
rect 541986 110898 542222 111134
rect 541986 75218 542222 75454
rect 541986 74898 542222 75134
rect 541986 39218 542222 39454
rect 541986 38898 542222 39134
rect 541986 3218 542222 3454
rect 541986 2898 542222 3134
rect 541986 -582 542222 -346
rect 541986 -902 542222 -666
rect 545586 690818 545822 691054
rect 545586 690498 545822 690734
rect 545586 654818 545822 655054
rect 545586 654498 545822 654734
rect 545586 618818 545822 619054
rect 545586 618498 545822 618734
rect 545586 582818 545822 583054
rect 545586 582498 545822 582734
rect 545586 546818 545822 547054
rect 545586 546498 545822 546734
rect 545586 510818 545822 511054
rect 545586 510498 545822 510734
rect 545586 474818 545822 475054
rect 545586 474498 545822 474734
rect 545586 438818 545822 439054
rect 545586 438498 545822 438734
rect 545586 402818 545822 403054
rect 545586 402498 545822 402734
rect 545586 366818 545822 367054
rect 545586 366498 545822 366734
rect 545586 330818 545822 331054
rect 545586 330498 545822 330734
rect 545586 294818 545822 295054
rect 545586 294498 545822 294734
rect 545586 258818 545822 259054
rect 545586 258498 545822 258734
rect 545586 222818 545822 223054
rect 545586 222498 545822 222734
rect 545586 186818 545822 187054
rect 545586 186498 545822 186734
rect 545586 150818 545822 151054
rect 545586 150498 545822 150734
rect 545586 114818 545822 115054
rect 545586 114498 545822 114734
rect 545586 78818 545822 79054
rect 545586 78498 545822 78734
rect 545586 42818 545822 43054
rect 545586 42498 545822 42734
rect 545586 6818 545822 7054
rect 545586 6498 545822 6734
rect 545586 -2462 545822 -2226
rect 545586 -2782 545822 -2546
rect 549186 694418 549422 694654
rect 549186 694098 549422 694334
rect 549186 658418 549422 658654
rect 549186 658098 549422 658334
rect 549186 622418 549422 622654
rect 549186 622098 549422 622334
rect 549186 586418 549422 586654
rect 549186 586098 549422 586334
rect 549186 550418 549422 550654
rect 549186 550098 549422 550334
rect 549186 514418 549422 514654
rect 549186 514098 549422 514334
rect 549186 478418 549422 478654
rect 549186 478098 549422 478334
rect 549186 442418 549422 442654
rect 549186 442098 549422 442334
rect 549186 406418 549422 406654
rect 549186 406098 549422 406334
rect 549186 370418 549422 370654
rect 549186 370098 549422 370334
rect 549186 334418 549422 334654
rect 549186 334098 549422 334334
rect 549186 298418 549422 298654
rect 549186 298098 549422 298334
rect 549186 262418 549422 262654
rect 549186 262098 549422 262334
rect 549186 226418 549422 226654
rect 549186 226098 549422 226334
rect 549186 190418 549422 190654
rect 549186 190098 549422 190334
rect 549186 154418 549422 154654
rect 549186 154098 549422 154334
rect 549186 118418 549422 118654
rect 549186 118098 549422 118334
rect 549186 82418 549422 82654
rect 549186 82098 549422 82334
rect 549186 46418 549422 46654
rect 549186 46098 549422 46334
rect 549186 10418 549422 10654
rect 549186 10098 549422 10334
rect 549186 -4342 549422 -4106
rect 549186 -4662 549422 -4426
rect 570786 711182 571022 711418
rect 570786 710862 571022 711098
rect 567186 709302 567422 709538
rect 567186 708982 567422 709218
rect 563586 707422 563822 707658
rect 563586 707102 563822 707338
rect 552786 698018 553022 698254
rect 552786 697698 553022 697934
rect 552786 662018 553022 662254
rect 552786 661698 553022 661934
rect 552786 626018 553022 626254
rect 552786 625698 553022 625934
rect 552786 590018 553022 590254
rect 552786 589698 553022 589934
rect 552786 554018 553022 554254
rect 552786 553698 553022 553934
rect 552786 518018 553022 518254
rect 552786 517698 553022 517934
rect 552786 482018 553022 482254
rect 552786 481698 553022 481934
rect 552786 446018 553022 446254
rect 552786 445698 553022 445934
rect 552786 410018 553022 410254
rect 552786 409698 553022 409934
rect 552786 374018 553022 374254
rect 552786 373698 553022 373934
rect 552786 338018 553022 338254
rect 552786 337698 553022 337934
rect 552786 302018 553022 302254
rect 552786 301698 553022 301934
rect 552786 266018 553022 266254
rect 552786 265698 553022 265934
rect 552786 230018 553022 230254
rect 552786 229698 553022 229934
rect 552786 194018 553022 194254
rect 552786 193698 553022 193934
rect 552786 158018 553022 158254
rect 552786 157698 553022 157934
rect 552786 122018 553022 122254
rect 552786 121698 553022 121934
rect 552786 86018 553022 86254
rect 552786 85698 553022 85934
rect 552786 50018 553022 50254
rect 552786 49698 553022 49934
rect 552786 14018 553022 14254
rect 552786 13698 553022 13934
rect 534786 -7162 535022 -6926
rect 534786 -7482 535022 -7246
rect 559986 705542 560222 705778
rect 559986 705222 560222 705458
rect 559986 669218 560222 669454
rect 559986 668898 560222 669134
rect 559986 633218 560222 633454
rect 559986 632898 560222 633134
rect 559986 597218 560222 597454
rect 559986 596898 560222 597134
rect 559986 561218 560222 561454
rect 559986 560898 560222 561134
rect 559986 525218 560222 525454
rect 559986 524898 560222 525134
rect 559986 489218 560222 489454
rect 559986 488898 560222 489134
rect 559986 453218 560222 453454
rect 559986 452898 560222 453134
rect 559986 417218 560222 417454
rect 559986 416898 560222 417134
rect 559986 381218 560222 381454
rect 559986 380898 560222 381134
rect 559986 345218 560222 345454
rect 559986 344898 560222 345134
rect 559986 309218 560222 309454
rect 559986 308898 560222 309134
rect 559986 273218 560222 273454
rect 559986 272898 560222 273134
rect 559986 237218 560222 237454
rect 559986 236898 560222 237134
rect 559986 201218 560222 201454
rect 559986 200898 560222 201134
rect 559986 165218 560222 165454
rect 559986 164898 560222 165134
rect 559986 129218 560222 129454
rect 559986 128898 560222 129134
rect 559986 93218 560222 93454
rect 559986 92898 560222 93134
rect 559986 57218 560222 57454
rect 559986 56898 560222 57134
rect 559986 21218 560222 21454
rect 559986 20898 560222 21134
rect 559986 -1522 560222 -1286
rect 559986 -1842 560222 -1606
rect 563586 672818 563822 673054
rect 563586 672498 563822 672734
rect 563586 636818 563822 637054
rect 563586 636498 563822 636734
rect 563586 600818 563822 601054
rect 563586 600498 563822 600734
rect 563586 564818 563822 565054
rect 563586 564498 563822 564734
rect 563586 528818 563822 529054
rect 563586 528498 563822 528734
rect 563586 492818 563822 493054
rect 563586 492498 563822 492734
rect 563586 456818 563822 457054
rect 563586 456498 563822 456734
rect 563586 420818 563822 421054
rect 563586 420498 563822 420734
rect 563586 384818 563822 385054
rect 563586 384498 563822 384734
rect 563586 348818 563822 349054
rect 563586 348498 563822 348734
rect 563586 312818 563822 313054
rect 563586 312498 563822 312734
rect 563586 276818 563822 277054
rect 563586 276498 563822 276734
rect 563586 240818 563822 241054
rect 563586 240498 563822 240734
rect 563586 204818 563822 205054
rect 563586 204498 563822 204734
rect 563586 168818 563822 169054
rect 563586 168498 563822 168734
rect 563586 132818 563822 133054
rect 563586 132498 563822 132734
rect 563586 96818 563822 97054
rect 563586 96498 563822 96734
rect 563586 60818 563822 61054
rect 563586 60498 563822 60734
rect 563586 24818 563822 25054
rect 563586 24498 563822 24734
rect 563586 -3402 563822 -3166
rect 563586 -3722 563822 -3486
rect 567186 676418 567422 676654
rect 567186 676098 567422 676334
rect 567186 640418 567422 640654
rect 567186 640098 567422 640334
rect 567186 604418 567422 604654
rect 567186 604098 567422 604334
rect 567186 568418 567422 568654
rect 567186 568098 567422 568334
rect 567186 532418 567422 532654
rect 567186 532098 567422 532334
rect 567186 496418 567422 496654
rect 567186 496098 567422 496334
rect 567186 460418 567422 460654
rect 567186 460098 567422 460334
rect 567186 424418 567422 424654
rect 567186 424098 567422 424334
rect 567186 388418 567422 388654
rect 567186 388098 567422 388334
rect 567186 352418 567422 352654
rect 567186 352098 567422 352334
rect 567186 316418 567422 316654
rect 567186 316098 567422 316334
rect 567186 280418 567422 280654
rect 567186 280098 567422 280334
rect 567186 244418 567422 244654
rect 567186 244098 567422 244334
rect 567186 208418 567422 208654
rect 567186 208098 567422 208334
rect 567186 172418 567422 172654
rect 567186 172098 567422 172334
rect 567186 136418 567422 136654
rect 567186 136098 567422 136334
rect 567186 100418 567422 100654
rect 567186 100098 567422 100334
rect 567186 64418 567422 64654
rect 567186 64098 567422 64334
rect 567186 28418 567422 28654
rect 567186 28098 567422 28334
rect 567186 -5282 567422 -5046
rect 567186 -5602 567422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 581586 706482 581822 706718
rect 581586 706162 581822 706398
rect 570786 680018 571022 680254
rect 570786 679698 571022 679934
rect 570786 644018 571022 644254
rect 570786 643698 571022 643934
rect 570786 608018 571022 608254
rect 570786 607698 571022 607934
rect 570786 572018 571022 572254
rect 570786 571698 571022 571934
rect 570786 536018 571022 536254
rect 570786 535698 571022 535934
rect 570786 500018 571022 500254
rect 570786 499698 571022 499934
rect 570786 464018 571022 464254
rect 570786 463698 571022 463934
rect 570786 428018 571022 428254
rect 570786 427698 571022 427934
rect 570786 392018 571022 392254
rect 570786 391698 571022 391934
rect 570786 356018 571022 356254
rect 570786 355698 571022 355934
rect 570786 320018 571022 320254
rect 570786 319698 571022 319934
rect 570786 284018 571022 284254
rect 570786 283698 571022 283934
rect 570786 248018 571022 248254
rect 570786 247698 571022 247934
rect 570786 212018 571022 212254
rect 570786 211698 571022 211934
rect 570786 176018 571022 176254
rect 570786 175698 571022 175934
rect 570786 140018 571022 140254
rect 570786 139698 571022 139934
rect 570786 104018 571022 104254
rect 570786 103698 571022 103934
rect 570786 68018 571022 68254
rect 570786 67698 571022 67934
rect 570786 32018 571022 32254
rect 570786 31698 571022 31934
rect 552786 -6222 553022 -5986
rect 552786 -6542 553022 -6306
rect 577986 704602 578222 704838
rect 577986 704282 578222 704518
rect 577986 687218 578222 687454
rect 577986 686898 578222 687134
rect 577986 651218 578222 651454
rect 577986 650898 578222 651134
rect 577986 615218 578222 615454
rect 577986 614898 578222 615134
rect 577986 579218 578222 579454
rect 577986 578898 578222 579134
rect 577986 543218 578222 543454
rect 577986 542898 578222 543134
rect 577986 507218 578222 507454
rect 577986 506898 578222 507134
rect 577986 471218 578222 471454
rect 577986 470898 578222 471134
rect 577986 435218 578222 435454
rect 577986 434898 578222 435134
rect 577986 399218 578222 399454
rect 577986 398898 578222 399134
rect 577986 363218 578222 363454
rect 577986 362898 578222 363134
rect 577986 327218 578222 327454
rect 577986 326898 578222 327134
rect 577986 291218 578222 291454
rect 577986 290898 578222 291134
rect 577986 255218 578222 255454
rect 577986 254898 578222 255134
rect 577986 219218 578222 219454
rect 577986 218898 578222 219134
rect 577986 183218 578222 183454
rect 577986 182898 578222 183134
rect 577986 147218 578222 147454
rect 577986 146898 578222 147134
rect 577986 111218 578222 111454
rect 577986 110898 578222 111134
rect 577986 75218 578222 75454
rect 577986 74898 578222 75134
rect 577986 39218 578222 39454
rect 577986 38898 578222 39134
rect 577986 3218 578222 3454
rect 577986 2898 578222 3134
rect 577986 -582 578222 -346
rect 577986 -902 578222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 581586 690818 581822 691054
rect 581586 690498 581822 690734
rect 581586 654818 581822 655054
rect 581586 654498 581822 654734
rect 581586 618818 581822 619054
rect 581586 618498 581822 618734
rect 581586 582818 581822 583054
rect 581586 582498 581822 582734
rect 581586 546818 581822 547054
rect 581586 546498 581822 546734
rect 581586 510818 581822 511054
rect 581586 510498 581822 510734
rect 581586 474818 581822 475054
rect 581586 474498 581822 474734
rect 581586 438818 581822 439054
rect 581586 438498 581822 438734
rect 581586 402818 581822 403054
rect 581586 402498 581822 402734
rect 581586 366818 581822 367054
rect 581586 366498 581822 366734
rect 581586 330818 581822 331054
rect 581586 330498 581822 330734
rect 581586 294818 581822 295054
rect 581586 294498 581822 294734
rect 581586 258818 581822 259054
rect 581586 258498 581822 258734
rect 581586 222818 581822 223054
rect 581586 222498 581822 222734
rect 581586 186818 581822 187054
rect 581586 186498 581822 186734
rect 581586 150818 581822 151054
rect 581586 150498 581822 150734
rect 581586 114818 581822 115054
rect 581586 114498 581822 114734
rect 581586 78818 581822 79054
rect 581586 78498 581822 78734
rect 581586 42818 581822 43054
rect 581586 42498 581822 42734
rect 581586 6818 581822 7054
rect 581586 6498 581822 6734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 687218 585738 687454
rect 585502 686898 585738 687134
rect 585502 651218 585738 651454
rect 585502 650898 585738 651134
rect 585502 615218 585738 615454
rect 585502 614898 585738 615134
rect 585502 579218 585738 579454
rect 585502 578898 585738 579134
rect 585502 543218 585738 543454
rect 585502 542898 585738 543134
rect 585502 507218 585738 507454
rect 585502 506898 585738 507134
rect 585502 471218 585738 471454
rect 585502 470898 585738 471134
rect 585502 435218 585738 435454
rect 585502 434898 585738 435134
rect 585502 399218 585738 399454
rect 585502 398898 585738 399134
rect 585502 363218 585738 363454
rect 585502 362898 585738 363134
rect 585502 327218 585738 327454
rect 585502 326898 585738 327134
rect 585502 291218 585738 291454
rect 585502 290898 585738 291134
rect 585502 255218 585738 255454
rect 585502 254898 585738 255134
rect 585502 219218 585738 219454
rect 585502 218898 585738 219134
rect 585502 183218 585738 183454
rect 585502 182898 585738 183134
rect 585502 147218 585738 147454
rect 585502 146898 585738 147134
rect 585502 111218 585738 111454
rect 585502 110898 585738 111134
rect 585502 75218 585738 75454
rect 585502 74898 585738 75134
rect 585502 39218 585738 39454
rect 585502 38898 585738 39134
rect 585502 3218 585738 3454
rect 585502 2898 585738 3134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 669218 586678 669454
rect 586442 668898 586678 669134
rect 586442 633218 586678 633454
rect 586442 632898 586678 633134
rect 586442 597218 586678 597454
rect 586442 596898 586678 597134
rect 586442 561218 586678 561454
rect 586442 560898 586678 561134
rect 586442 525218 586678 525454
rect 586442 524898 586678 525134
rect 586442 489218 586678 489454
rect 586442 488898 586678 489134
rect 586442 453218 586678 453454
rect 586442 452898 586678 453134
rect 586442 417218 586678 417454
rect 586442 416898 586678 417134
rect 586442 381218 586678 381454
rect 586442 380898 586678 381134
rect 586442 345218 586678 345454
rect 586442 344898 586678 345134
rect 586442 309218 586678 309454
rect 586442 308898 586678 309134
rect 586442 273218 586678 273454
rect 586442 272898 586678 273134
rect 586442 237218 586678 237454
rect 586442 236898 586678 237134
rect 586442 201218 586678 201454
rect 586442 200898 586678 201134
rect 586442 165218 586678 165454
rect 586442 164898 586678 165134
rect 586442 129218 586678 129454
rect 586442 128898 586678 129134
rect 586442 93218 586678 93454
rect 586442 92898 586678 93134
rect 586442 57218 586678 57454
rect 586442 56898 586678 57134
rect 586442 21218 586678 21454
rect 586442 20898 586678 21134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 690818 587618 691054
rect 587382 690498 587618 690734
rect 587382 654818 587618 655054
rect 587382 654498 587618 654734
rect 587382 618818 587618 619054
rect 587382 618498 587618 618734
rect 587382 582818 587618 583054
rect 587382 582498 587618 582734
rect 587382 546818 587618 547054
rect 587382 546498 587618 546734
rect 587382 510818 587618 511054
rect 587382 510498 587618 510734
rect 587382 474818 587618 475054
rect 587382 474498 587618 474734
rect 587382 438818 587618 439054
rect 587382 438498 587618 438734
rect 587382 402818 587618 403054
rect 587382 402498 587618 402734
rect 587382 366818 587618 367054
rect 587382 366498 587618 366734
rect 587382 330818 587618 331054
rect 587382 330498 587618 330734
rect 587382 294818 587618 295054
rect 587382 294498 587618 294734
rect 587382 258818 587618 259054
rect 587382 258498 587618 258734
rect 587382 222818 587618 223054
rect 587382 222498 587618 222734
rect 587382 186818 587618 187054
rect 587382 186498 587618 186734
rect 587382 150818 587618 151054
rect 587382 150498 587618 150734
rect 587382 114818 587618 115054
rect 587382 114498 587618 114734
rect 587382 78818 587618 79054
rect 587382 78498 587618 78734
rect 587382 42818 587618 43054
rect 587382 42498 587618 42734
rect 587382 6818 587618 7054
rect 587382 6498 587618 6734
rect 581586 -2462 581822 -2226
rect 581586 -2782 581822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 672818 588558 673054
rect 588322 672498 588558 672734
rect 588322 636818 588558 637054
rect 588322 636498 588558 636734
rect 588322 600818 588558 601054
rect 588322 600498 588558 600734
rect 588322 564818 588558 565054
rect 588322 564498 588558 564734
rect 588322 528818 588558 529054
rect 588322 528498 588558 528734
rect 588322 492818 588558 493054
rect 588322 492498 588558 492734
rect 588322 456818 588558 457054
rect 588322 456498 588558 456734
rect 588322 420818 588558 421054
rect 588322 420498 588558 420734
rect 588322 384818 588558 385054
rect 588322 384498 588558 384734
rect 588322 348818 588558 349054
rect 588322 348498 588558 348734
rect 588322 312818 588558 313054
rect 588322 312498 588558 312734
rect 588322 276818 588558 277054
rect 588322 276498 588558 276734
rect 588322 240818 588558 241054
rect 588322 240498 588558 240734
rect 588322 204818 588558 205054
rect 588322 204498 588558 204734
rect 588322 168818 588558 169054
rect 588322 168498 588558 168734
rect 588322 132818 588558 133054
rect 588322 132498 588558 132734
rect 588322 96818 588558 97054
rect 588322 96498 588558 96734
rect 588322 60818 588558 61054
rect 588322 60498 588558 60734
rect 588322 24818 588558 25054
rect 588322 24498 588558 24734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 694418 589498 694654
rect 589262 694098 589498 694334
rect 589262 658418 589498 658654
rect 589262 658098 589498 658334
rect 589262 622418 589498 622654
rect 589262 622098 589498 622334
rect 589262 586418 589498 586654
rect 589262 586098 589498 586334
rect 589262 550418 589498 550654
rect 589262 550098 589498 550334
rect 589262 514418 589498 514654
rect 589262 514098 589498 514334
rect 589262 478418 589498 478654
rect 589262 478098 589498 478334
rect 589262 442418 589498 442654
rect 589262 442098 589498 442334
rect 589262 406418 589498 406654
rect 589262 406098 589498 406334
rect 589262 370418 589498 370654
rect 589262 370098 589498 370334
rect 589262 334418 589498 334654
rect 589262 334098 589498 334334
rect 589262 298418 589498 298654
rect 589262 298098 589498 298334
rect 589262 262418 589498 262654
rect 589262 262098 589498 262334
rect 589262 226418 589498 226654
rect 589262 226098 589498 226334
rect 589262 190418 589498 190654
rect 589262 190098 589498 190334
rect 589262 154418 589498 154654
rect 589262 154098 589498 154334
rect 589262 118418 589498 118654
rect 589262 118098 589498 118334
rect 589262 82418 589498 82654
rect 589262 82098 589498 82334
rect 589262 46418 589498 46654
rect 589262 46098 589498 46334
rect 589262 10418 589498 10654
rect 589262 10098 589498 10334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 676418 590438 676654
rect 590202 676098 590438 676334
rect 590202 640418 590438 640654
rect 590202 640098 590438 640334
rect 590202 604418 590438 604654
rect 590202 604098 590438 604334
rect 590202 568418 590438 568654
rect 590202 568098 590438 568334
rect 590202 532418 590438 532654
rect 590202 532098 590438 532334
rect 590202 496418 590438 496654
rect 590202 496098 590438 496334
rect 590202 460418 590438 460654
rect 590202 460098 590438 460334
rect 590202 424418 590438 424654
rect 590202 424098 590438 424334
rect 590202 388418 590438 388654
rect 590202 388098 590438 388334
rect 590202 352418 590438 352654
rect 590202 352098 590438 352334
rect 590202 316418 590438 316654
rect 590202 316098 590438 316334
rect 590202 280418 590438 280654
rect 590202 280098 590438 280334
rect 590202 244418 590438 244654
rect 590202 244098 590438 244334
rect 590202 208418 590438 208654
rect 590202 208098 590438 208334
rect 590202 172418 590438 172654
rect 590202 172098 590438 172334
rect 590202 136418 590438 136654
rect 590202 136098 590438 136334
rect 590202 100418 590438 100654
rect 590202 100098 590438 100334
rect 590202 64418 590438 64654
rect 590202 64098 590438 64334
rect 590202 28418 590438 28654
rect 590202 28098 590438 28334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 698018 591378 698254
rect 591142 697698 591378 697934
rect 591142 662018 591378 662254
rect 591142 661698 591378 661934
rect 591142 626018 591378 626254
rect 591142 625698 591378 625934
rect 591142 590018 591378 590254
rect 591142 589698 591378 589934
rect 591142 554018 591378 554254
rect 591142 553698 591378 553934
rect 591142 518018 591378 518254
rect 591142 517698 591378 517934
rect 591142 482018 591378 482254
rect 591142 481698 591378 481934
rect 591142 446018 591378 446254
rect 591142 445698 591378 445934
rect 591142 410018 591378 410254
rect 591142 409698 591378 409934
rect 591142 374018 591378 374254
rect 591142 373698 591378 373934
rect 591142 338018 591378 338254
rect 591142 337698 591378 337934
rect 591142 302018 591378 302254
rect 591142 301698 591378 301934
rect 591142 266018 591378 266254
rect 591142 265698 591378 265934
rect 591142 230018 591378 230254
rect 591142 229698 591378 229934
rect 591142 194018 591378 194254
rect 591142 193698 591378 193934
rect 591142 158018 591378 158254
rect 591142 157698 591378 157934
rect 591142 122018 591378 122254
rect 591142 121698 591378 121934
rect 591142 86018 591378 86254
rect 591142 85698 591378 85934
rect 591142 50018 591378 50254
rect 591142 49698 591378 49934
rect 591142 14018 591378 14254
rect 591142 13698 591378 13934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 680018 592318 680254
rect 592082 679698 592318 679934
rect 592082 644018 592318 644254
rect 592082 643698 592318 643934
rect 592082 608018 592318 608254
rect 592082 607698 592318 607934
rect 592082 572018 592318 572254
rect 592082 571698 592318 571934
rect 592082 536018 592318 536254
rect 592082 535698 592318 535934
rect 592082 500018 592318 500254
rect 592082 499698 592318 499934
rect 592082 464018 592318 464254
rect 592082 463698 592318 463934
rect 592082 428018 592318 428254
rect 592082 427698 592318 427934
rect 592082 392018 592318 392254
rect 592082 391698 592318 391934
rect 592082 356018 592318 356254
rect 592082 355698 592318 355934
rect 592082 320018 592318 320254
rect 592082 319698 592318 319934
rect 592082 284018 592318 284254
rect 592082 283698 592318 283934
rect 592082 248018 592318 248254
rect 592082 247698 592318 247934
rect 592082 212018 592318 212254
rect 592082 211698 592318 211934
rect 592082 176018 592318 176254
rect 592082 175698 592318 175934
rect 592082 140018 592318 140254
rect 592082 139698 592318 139934
rect 592082 104018 592318 104254
rect 592082 103698 592318 103934
rect 592082 68018 592318 68254
rect 592082 67698 592318 67934
rect 592082 32018 592318 32254
rect 592082 31698 592318 31934
rect 570786 -7162 571022 -6926
rect 570786 -7482 571022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 30786 711418
rect 31022 711182 66786 711418
rect 67022 711182 102786 711418
rect 103022 711182 138786 711418
rect 139022 711182 174786 711418
rect 175022 711182 210786 711418
rect 211022 711182 246786 711418
rect 247022 711182 282786 711418
rect 283022 711182 318786 711418
rect 319022 711182 354786 711418
rect 355022 711182 390786 711418
rect 391022 711182 426786 711418
rect 427022 711182 462786 711418
rect 463022 711182 498786 711418
rect 499022 711182 534786 711418
rect 535022 711182 570786 711418
rect 571022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 30786 711098
rect 31022 710862 66786 711098
rect 67022 710862 102786 711098
rect 103022 710862 138786 711098
rect 139022 710862 174786 711098
rect 175022 710862 210786 711098
rect 211022 710862 246786 711098
rect 247022 710862 282786 711098
rect 283022 710862 318786 711098
rect 319022 710862 354786 711098
rect 355022 710862 390786 711098
rect 391022 710862 426786 711098
rect 427022 710862 462786 711098
rect 463022 710862 498786 711098
rect 499022 710862 534786 711098
rect 535022 710862 570786 711098
rect 571022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 12786 710478
rect 13022 710242 48786 710478
rect 49022 710242 84786 710478
rect 85022 710242 120786 710478
rect 121022 710242 156786 710478
rect 157022 710242 192786 710478
rect 193022 710242 228786 710478
rect 229022 710242 264786 710478
rect 265022 710242 300786 710478
rect 301022 710242 336786 710478
rect 337022 710242 372786 710478
rect 373022 710242 408786 710478
rect 409022 710242 444786 710478
rect 445022 710242 480786 710478
rect 481022 710242 516786 710478
rect 517022 710242 552786 710478
rect 553022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 12786 710158
rect 13022 709922 48786 710158
rect 49022 709922 84786 710158
rect 85022 709922 120786 710158
rect 121022 709922 156786 710158
rect 157022 709922 192786 710158
rect 193022 709922 228786 710158
rect 229022 709922 264786 710158
rect 265022 709922 300786 710158
rect 301022 709922 336786 710158
rect 337022 709922 372786 710158
rect 373022 709922 408786 710158
rect 409022 709922 444786 710158
rect 445022 709922 480786 710158
rect 481022 709922 516786 710158
rect 517022 709922 552786 710158
rect 553022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 27186 709538
rect 27422 709302 63186 709538
rect 63422 709302 99186 709538
rect 99422 709302 135186 709538
rect 135422 709302 171186 709538
rect 171422 709302 207186 709538
rect 207422 709302 243186 709538
rect 243422 709302 279186 709538
rect 279422 709302 315186 709538
rect 315422 709302 351186 709538
rect 351422 709302 387186 709538
rect 387422 709302 423186 709538
rect 423422 709302 459186 709538
rect 459422 709302 495186 709538
rect 495422 709302 531186 709538
rect 531422 709302 567186 709538
rect 567422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 27186 709218
rect 27422 708982 63186 709218
rect 63422 708982 99186 709218
rect 99422 708982 135186 709218
rect 135422 708982 171186 709218
rect 171422 708982 207186 709218
rect 207422 708982 243186 709218
rect 243422 708982 279186 709218
rect 279422 708982 315186 709218
rect 315422 708982 351186 709218
rect 351422 708982 387186 709218
rect 387422 708982 423186 709218
rect 423422 708982 459186 709218
rect 459422 708982 495186 709218
rect 495422 708982 531186 709218
rect 531422 708982 567186 709218
rect 567422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 9186 708598
rect 9422 708362 45186 708598
rect 45422 708362 81186 708598
rect 81422 708362 117186 708598
rect 117422 708362 153186 708598
rect 153422 708362 189186 708598
rect 189422 708362 225186 708598
rect 225422 708362 261186 708598
rect 261422 708362 297186 708598
rect 297422 708362 333186 708598
rect 333422 708362 369186 708598
rect 369422 708362 405186 708598
rect 405422 708362 441186 708598
rect 441422 708362 477186 708598
rect 477422 708362 513186 708598
rect 513422 708362 549186 708598
rect 549422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 9186 708278
rect 9422 708042 45186 708278
rect 45422 708042 81186 708278
rect 81422 708042 117186 708278
rect 117422 708042 153186 708278
rect 153422 708042 189186 708278
rect 189422 708042 225186 708278
rect 225422 708042 261186 708278
rect 261422 708042 297186 708278
rect 297422 708042 333186 708278
rect 333422 708042 369186 708278
rect 369422 708042 405186 708278
rect 405422 708042 441186 708278
rect 441422 708042 477186 708278
rect 477422 708042 513186 708278
rect 513422 708042 549186 708278
rect 549422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 23586 707658
rect 23822 707422 59586 707658
rect 59822 707422 95586 707658
rect 95822 707422 131586 707658
rect 131822 707422 167586 707658
rect 167822 707422 203586 707658
rect 203822 707422 239586 707658
rect 239822 707422 275586 707658
rect 275822 707422 311586 707658
rect 311822 707422 347586 707658
rect 347822 707422 383586 707658
rect 383822 707422 419586 707658
rect 419822 707422 455586 707658
rect 455822 707422 491586 707658
rect 491822 707422 527586 707658
rect 527822 707422 563586 707658
rect 563822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 23586 707338
rect 23822 707102 59586 707338
rect 59822 707102 95586 707338
rect 95822 707102 131586 707338
rect 131822 707102 167586 707338
rect 167822 707102 203586 707338
rect 203822 707102 239586 707338
rect 239822 707102 275586 707338
rect 275822 707102 311586 707338
rect 311822 707102 347586 707338
rect 347822 707102 383586 707338
rect 383822 707102 419586 707338
rect 419822 707102 455586 707338
rect 455822 707102 491586 707338
rect 491822 707102 527586 707338
rect 527822 707102 563586 707338
rect 563822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 5586 706718
rect 5822 706482 41586 706718
rect 41822 706482 77586 706718
rect 77822 706482 113586 706718
rect 113822 706482 149586 706718
rect 149822 706482 185586 706718
rect 185822 706482 221586 706718
rect 221822 706482 257586 706718
rect 257822 706482 293586 706718
rect 293822 706482 329586 706718
rect 329822 706482 365586 706718
rect 365822 706482 401586 706718
rect 401822 706482 437586 706718
rect 437822 706482 473586 706718
rect 473822 706482 509586 706718
rect 509822 706482 545586 706718
rect 545822 706482 581586 706718
rect 581822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 5586 706398
rect 5822 706162 41586 706398
rect 41822 706162 77586 706398
rect 77822 706162 113586 706398
rect 113822 706162 149586 706398
rect 149822 706162 185586 706398
rect 185822 706162 221586 706398
rect 221822 706162 257586 706398
rect 257822 706162 293586 706398
rect 293822 706162 329586 706398
rect 329822 706162 365586 706398
rect 365822 706162 401586 706398
rect 401822 706162 437586 706398
rect 437822 706162 473586 706398
rect 473822 706162 509586 706398
rect 509822 706162 545586 706398
rect 545822 706162 581586 706398
rect 581822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 19986 705778
rect 20222 705542 55986 705778
rect 56222 705542 91986 705778
rect 92222 705542 127986 705778
rect 128222 705542 163986 705778
rect 164222 705542 199986 705778
rect 200222 705542 235986 705778
rect 236222 705542 271986 705778
rect 272222 705542 307986 705778
rect 308222 705542 343986 705778
rect 344222 705542 379986 705778
rect 380222 705542 415986 705778
rect 416222 705542 451986 705778
rect 452222 705542 487986 705778
rect 488222 705542 523986 705778
rect 524222 705542 559986 705778
rect 560222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 19986 705458
rect 20222 705222 55986 705458
rect 56222 705222 91986 705458
rect 92222 705222 127986 705458
rect 128222 705222 163986 705458
rect 164222 705222 199986 705458
rect 200222 705222 235986 705458
rect 236222 705222 271986 705458
rect 272222 705222 307986 705458
rect 308222 705222 343986 705458
rect 344222 705222 379986 705458
rect 380222 705222 415986 705458
rect 416222 705222 451986 705458
rect 452222 705222 487986 705458
rect 488222 705222 523986 705458
rect 524222 705222 559986 705458
rect 560222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 1986 704838
rect 2222 704602 37986 704838
rect 38222 704602 73986 704838
rect 74222 704602 109986 704838
rect 110222 704602 145986 704838
rect 146222 704602 181986 704838
rect 182222 704602 217986 704838
rect 218222 704602 253986 704838
rect 254222 704602 289986 704838
rect 290222 704602 325986 704838
rect 326222 704602 361986 704838
rect 362222 704602 397986 704838
rect 398222 704602 433986 704838
rect 434222 704602 469986 704838
rect 470222 704602 505986 704838
rect 506222 704602 541986 704838
rect 542222 704602 577986 704838
rect 578222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 1986 704518
rect 2222 704282 37986 704518
rect 38222 704282 73986 704518
rect 74222 704282 109986 704518
rect 110222 704282 145986 704518
rect 146222 704282 181986 704518
rect 182222 704282 217986 704518
rect 218222 704282 253986 704518
rect 254222 704282 289986 704518
rect 290222 704282 325986 704518
rect 326222 704282 361986 704518
rect 362222 704282 397986 704518
rect 398222 704282 433986 704518
rect 434222 704282 469986 704518
rect 470222 704282 505986 704518
rect 506222 704282 541986 704518
rect 542222 704282 577986 704518
rect 578222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect -7636 698276 -7036 698278
rect 12604 698276 13204 698278
rect 48604 698276 49204 698278
rect 84604 698276 85204 698278
rect 120604 698276 121204 698278
rect 156604 698276 157204 698278
rect 192604 698276 193204 698278
rect 228604 698276 229204 698278
rect 264604 698276 265204 698278
rect 300604 698276 301204 698278
rect 336604 698276 337204 698278
rect 372604 698276 373204 698278
rect 408604 698276 409204 698278
rect 444604 698276 445204 698278
rect 480604 698276 481204 698278
rect 516604 698276 517204 698278
rect 552604 698276 553204 698278
rect 590960 698276 591560 698278
rect -8576 698254 592500 698276
rect -8576 698018 -7454 698254
rect -7218 698018 12786 698254
rect 13022 698018 48786 698254
rect 49022 698018 84786 698254
rect 85022 698018 120786 698254
rect 121022 698018 156786 698254
rect 157022 698018 192786 698254
rect 193022 698018 228786 698254
rect 229022 698018 264786 698254
rect 265022 698018 300786 698254
rect 301022 698018 336786 698254
rect 337022 698018 372786 698254
rect 373022 698018 408786 698254
rect 409022 698018 444786 698254
rect 445022 698018 480786 698254
rect 481022 698018 516786 698254
rect 517022 698018 552786 698254
rect 553022 698018 591142 698254
rect 591378 698018 592500 698254
rect -8576 697934 592500 698018
rect -8576 697698 -7454 697934
rect -7218 697698 12786 697934
rect 13022 697698 48786 697934
rect 49022 697698 84786 697934
rect 85022 697698 120786 697934
rect 121022 697698 156786 697934
rect 157022 697698 192786 697934
rect 193022 697698 228786 697934
rect 229022 697698 264786 697934
rect 265022 697698 300786 697934
rect 301022 697698 336786 697934
rect 337022 697698 372786 697934
rect 373022 697698 408786 697934
rect 409022 697698 444786 697934
rect 445022 697698 480786 697934
rect 481022 697698 516786 697934
rect 517022 697698 552786 697934
rect 553022 697698 591142 697934
rect 591378 697698 592500 697934
rect -8576 697676 592500 697698
rect -7636 697674 -7036 697676
rect 12604 697674 13204 697676
rect 48604 697674 49204 697676
rect 84604 697674 85204 697676
rect 120604 697674 121204 697676
rect 156604 697674 157204 697676
rect 192604 697674 193204 697676
rect 228604 697674 229204 697676
rect 264604 697674 265204 697676
rect 300604 697674 301204 697676
rect 336604 697674 337204 697676
rect 372604 697674 373204 697676
rect 408604 697674 409204 697676
rect 444604 697674 445204 697676
rect 480604 697674 481204 697676
rect 516604 697674 517204 697676
rect 552604 697674 553204 697676
rect 590960 697674 591560 697676
rect -5756 694676 -5156 694678
rect 9004 694676 9604 694678
rect 45004 694676 45604 694678
rect 81004 694676 81604 694678
rect 117004 694676 117604 694678
rect 153004 694676 153604 694678
rect 189004 694676 189604 694678
rect 225004 694676 225604 694678
rect 261004 694676 261604 694678
rect 297004 694676 297604 694678
rect 333004 694676 333604 694678
rect 369004 694676 369604 694678
rect 405004 694676 405604 694678
rect 441004 694676 441604 694678
rect 477004 694676 477604 694678
rect 513004 694676 513604 694678
rect 549004 694676 549604 694678
rect 589080 694676 589680 694678
rect -6696 694654 590620 694676
rect -6696 694418 -5574 694654
rect -5338 694418 9186 694654
rect 9422 694418 45186 694654
rect 45422 694418 81186 694654
rect 81422 694418 117186 694654
rect 117422 694418 153186 694654
rect 153422 694418 189186 694654
rect 189422 694418 225186 694654
rect 225422 694418 261186 694654
rect 261422 694418 297186 694654
rect 297422 694418 333186 694654
rect 333422 694418 369186 694654
rect 369422 694418 405186 694654
rect 405422 694418 441186 694654
rect 441422 694418 477186 694654
rect 477422 694418 513186 694654
rect 513422 694418 549186 694654
rect 549422 694418 589262 694654
rect 589498 694418 590620 694654
rect -6696 694334 590620 694418
rect -6696 694098 -5574 694334
rect -5338 694098 9186 694334
rect 9422 694098 45186 694334
rect 45422 694098 81186 694334
rect 81422 694098 117186 694334
rect 117422 694098 153186 694334
rect 153422 694098 189186 694334
rect 189422 694098 225186 694334
rect 225422 694098 261186 694334
rect 261422 694098 297186 694334
rect 297422 694098 333186 694334
rect 333422 694098 369186 694334
rect 369422 694098 405186 694334
rect 405422 694098 441186 694334
rect 441422 694098 477186 694334
rect 477422 694098 513186 694334
rect 513422 694098 549186 694334
rect 549422 694098 589262 694334
rect 589498 694098 590620 694334
rect -6696 694076 590620 694098
rect -5756 694074 -5156 694076
rect 9004 694074 9604 694076
rect 45004 694074 45604 694076
rect 81004 694074 81604 694076
rect 117004 694074 117604 694076
rect 153004 694074 153604 694076
rect 189004 694074 189604 694076
rect 225004 694074 225604 694076
rect 261004 694074 261604 694076
rect 297004 694074 297604 694076
rect 333004 694074 333604 694076
rect 369004 694074 369604 694076
rect 405004 694074 405604 694076
rect 441004 694074 441604 694076
rect 477004 694074 477604 694076
rect 513004 694074 513604 694076
rect 549004 694074 549604 694076
rect 589080 694074 589680 694076
rect -3876 691076 -3276 691078
rect 5404 691076 6004 691078
rect 41404 691076 42004 691078
rect 77404 691076 78004 691078
rect 113404 691076 114004 691078
rect 149404 691076 150004 691078
rect 185404 691076 186004 691078
rect 221404 691076 222004 691078
rect 257404 691076 258004 691078
rect 293404 691076 294004 691078
rect 329404 691076 330004 691078
rect 365404 691076 366004 691078
rect 401404 691076 402004 691078
rect 437404 691076 438004 691078
rect 473404 691076 474004 691078
rect 509404 691076 510004 691078
rect 545404 691076 546004 691078
rect 581404 691076 582004 691078
rect 587200 691076 587800 691078
rect -4816 691054 588740 691076
rect -4816 690818 -3694 691054
rect -3458 690818 5586 691054
rect 5822 690818 41586 691054
rect 41822 690818 77586 691054
rect 77822 690818 113586 691054
rect 113822 690818 149586 691054
rect 149822 690818 185586 691054
rect 185822 690818 221586 691054
rect 221822 690818 257586 691054
rect 257822 690818 293586 691054
rect 293822 690818 329586 691054
rect 329822 690818 365586 691054
rect 365822 690818 401586 691054
rect 401822 690818 437586 691054
rect 437822 690818 473586 691054
rect 473822 690818 509586 691054
rect 509822 690818 545586 691054
rect 545822 690818 581586 691054
rect 581822 690818 587382 691054
rect 587618 690818 588740 691054
rect -4816 690734 588740 690818
rect -4816 690498 -3694 690734
rect -3458 690498 5586 690734
rect 5822 690498 41586 690734
rect 41822 690498 77586 690734
rect 77822 690498 113586 690734
rect 113822 690498 149586 690734
rect 149822 690498 185586 690734
rect 185822 690498 221586 690734
rect 221822 690498 257586 690734
rect 257822 690498 293586 690734
rect 293822 690498 329586 690734
rect 329822 690498 365586 690734
rect 365822 690498 401586 690734
rect 401822 690498 437586 690734
rect 437822 690498 473586 690734
rect 473822 690498 509586 690734
rect 509822 690498 545586 690734
rect 545822 690498 581586 690734
rect 581822 690498 587382 690734
rect 587618 690498 588740 690734
rect -4816 690476 588740 690498
rect -3876 690474 -3276 690476
rect 5404 690474 6004 690476
rect 41404 690474 42004 690476
rect 77404 690474 78004 690476
rect 113404 690474 114004 690476
rect 149404 690474 150004 690476
rect 185404 690474 186004 690476
rect 221404 690474 222004 690476
rect 257404 690474 258004 690476
rect 293404 690474 294004 690476
rect 329404 690474 330004 690476
rect 365404 690474 366004 690476
rect 401404 690474 402004 690476
rect 437404 690474 438004 690476
rect 473404 690474 474004 690476
rect 509404 690474 510004 690476
rect 545404 690474 546004 690476
rect 581404 690474 582004 690476
rect 587200 690474 587800 690476
rect -1996 687476 -1396 687478
rect 1804 687476 2404 687478
rect 37804 687476 38404 687478
rect 73804 687476 74404 687478
rect 109804 687476 110404 687478
rect 145804 687476 146404 687478
rect 181804 687476 182404 687478
rect 217804 687476 218404 687478
rect 253804 687476 254404 687478
rect 289804 687476 290404 687478
rect 325804 687476 326404 687478
rect 361804 687476 362404 687478
rect 397804 687476 398404 687478
rect 433804 687476 434404 687478
rect 469804 687476 470404 687478
rect 505804 687476 506404 687478
rect 541804 687476 542404 687478
rect 577804 687476 578404 687478
rect 585320 687476 585920 687478
rect -2936 687454 586860 687476
rect -2936 687218 -1814 687454
rect -1578 687218 1986 687454
rect 2222 687218 37986 687454
rect 38222 687218 73986 687454
rect 74222 687218 109986 687454
rect 110222 687218 145986 687454
rect 146222 687218 181986 687454
rect 182222 687218 217986 687454
rect 218222 687218 253986 687454
rect 254222 687218 289986 687454
rect 290222 687218 325986 687454
rect 326222 687218 361986 687454
rect 362222 687218 397986 687454
rect 398222 687218 433986 687454
rect 434222 687218 469986 687454
rect 470222 687218 505986 687454
rect 506222 687218 541986 687454
rect 542222 687218 577986 687454
rect 578222 687218 585502 687454
rect 585738 687218 586860 687454
rect -2936 687134 586860 687218
rect -2936 686898 -1814 687134
rect -1578 686898 1986 687134
rect 2222 686898 37986 687134
rect 38222 686898 73986 687134
rect 74222 686898 109986 687134
rect 110222 686898 145986 687134
rect 146222 686898 181986 687134
rect 182222 686898 217986 687134
rect 218222 686898 253986 687134
rect 254222 686898 289986 687134
rect 290222 686898 325986 687134
rect 326222 686898 361986 687134
rect 362222 686898 397986 687134
rect 398222 686898 433986 687134
rect 434222 686898 469986 687134
rect 470222 686898 505986 687134
rect 506222 686898 541986 687134
rect 542222 686898 577986 687134
rect 578222 686898 585502 687134
rect 585738 686898 586860 687134
rect -2936 686876 586860 686898
rect -1996 686874 -1396 686876
rect 1804 686874 2404 686876
rect 37804 686874 38404 686876
rect 73804 686874 74404 686876
rect 109804 686874 110404 686876
rect 145804 686874 146404 686876
rect 181804 686874 182404 686876
rect 217804 686874 218404 686876
rect 253804 686874 254404 686876
rect 289804 686874 290404 686876
rect 325804 686874 326404 686876
rect 361804 686874 362404 686876
rect 397804 686874 398404 686876
rect 433804 686874 434404 686876
rect 469804 686874 470404 686876
rect 505804 686874 506404 686876
rect 541804 686874 542404 686876
rect 577804 686874 578404 686876
rect 585320 686874 585920 686876
rect -8576 680276 -7976 680278
rect 30604 680276 31204 680278
rect 66604 680276 67204 680278
rect 102604 680276 103204 680278
rect 138604 680276 139204 680278
rect 174604 680276 175204 680278
rect 210604 680276 211204 680278
rect 246604 680276 247204 680278
rect 282604 680276 283204 680278
rect 318604 680276 319204 680278
rect 354604 680276 355204 680278
rect 390604 680276 391204 680278
rect 426604 680276 427204 680278
rect 462604 680276 463204 680278
rect 498604 680276 499204 680278
rect 534604 680276 535204 680278
rect 570604 680276 571204 680278
rect 591900 680276 592500 680278
rect -8576 680254 592500 680276
rect -8576 680018 -8394 680254
rect -8158 680018 30786 680254
rect 31022 680018 66786 680254
rect 67022 680018 102786 680254
rect 103022 680018 138786 680254
rect 139022 680018 174786 680254
rect 175022 680018 210786 680254
rect 211022 680018 246786 680254
rect 247022 680018 282786 680254
rect 283022 680018 318786 680254
rect 319022 680018 354786 680254
rect 355022 680018 390786 680254
rect 391022 680018 426786 680254
rect 427022 680018 462786 680254
rect 463022 680018 498786 680254
rect 499022 680018 534786 680254
rect 535022 680018 570786 680254
rect 571022 680018 592082 680254
rect 592318 680018 592500 680254
rect -8576 679934 592500 680018
rect -8576 679698 -8394 679934
rect -8158 679698 30786 679934
rect 31022 679698 66786 679934
rect 67022 679698 102786 679934
rect 103022 679698 138786 679934
rect 139022 679698 174786 679934
rect 175022 679698 210786 679934
rect 211022 679698 246786 679934
rect 247022 679698 282786 679934
rect 283022 679698 318786 679934
rect 319022 679698 354786 679934
rect 355022 679698 390786 679934
rect 391022 679698 426786 679934
rect 427022 679698 462786 679934
rect 463022 679698 498786 679934
rect 499022 679698 534786 679934
rect 535022 679698 570786 679934
rect 571022 679698 592082 679934
rect 592318 679698 592500 679934
rect -8576 679676 592500 679698
rect -8576 679674 -7976 679676
rect 30604 679674 31204 679676
rect 66604 679674 67204 679676
rect 102604 679674 103204 679676
rect 138604 679674 139204 679676
rect 174604 679674 175204 679676
rect 210604 679674 211204 679676
rect 246604 679674 247204 679676
rect 282604 679674 283204 679676
rect 318604 679674 319204 679676
rect 354604 679674 355204 679676
rect 390604 679674 391204 679676
rect 426604 679674 427204 679676
rect 462604 679674 463204 679676
rect 498604 679674 499204 679676
rect 534604 679674 535204 679676
rect 570604 679674 571204 679676
rect 591900 679674 592500 679676
rect -6696 676676 -6096 676678
rect 27004 676676 27604 676678
rect 63004 676676 63604 676678
rect 99004 676676 99604 676678
rect 135004 676676 135604 676678
rect 171004 676676 171604 676678
rect 207004 676676 207604 676678
rect 243004 676676 243604 676678
rect 279004 676676 279604 676678
rect 315004 676676 315604 676678
rect 351004 676676 351604 676678
rect 387004 676676 387604 676678
rect 423004 676676 423604 676678
rect 459004 676676 459604 676678
rect 495004 676676 495604 676678
rect 531004 676676 531604 676678
rect 567004 676676 567604 676678
rect 590020 676676 590620 676678
rect -6696 676654 590620 676676
rect -6696 676418 -6514 676654
rect -6278 676418 27186 676654
rect 27422 676418 63186 676654
rect 63422 676418 99186 676654
rect 99422 676418 135186 676654
rect 135422 676418 171186 676654
rect 171422 676418 207186 676654
rect 207422 676418 243186 676654
rect 243422 676418 279186 676654
rect 279422 676418 315186 676654
rect 315422 676418 351186 676654
rect 351422 676418 387186 676654
rect 387422 676418 423186 676654
rect 423422 676418 459186 676654
rect 459422 676418 495186 676654
rect 495422 676418 531186 676654
rect 531422 676418 567186 676654
rect 567422 676418 590202 676654
rect 590438 676418 590620 676654
rect -6696 676334 590620 676418
rect -6696 676098 -6514 676334
rect -6278 676098 27186 676334
rect 27422 676098 63186 676334
rect 63422 676098 99186 676334
rect 99422 676098 135186 676334
rect 135422 676098 171186 676334
rect 171422 676098 207186 676334
rect 207422 676098 243186 676334
rect 243422 676098 279186 676334
rect 279422 676098 315186 676334
rect 315422 676098 351186 676334
rect 351422 676098 387186 676334
rect 387422 676098 423186 676334
rect 423422 676098 459186 676334
rect 459422 676098 495186 676334
rect 495422 676098 531186 676334
rect 531422 676098 567186 676334
rect 567422 676098 590202 676334
rect 590438 676098 590620 676334
rect -6696 676076 590620 676098
rect -6696 676074 -6096 676076
rect 27004 676074 27604 676076
rect 63004 676074 63604 676076
rect 99004 676074 99604 676076
rect 135004 676074 135604 676076
rect 171004 676074 171604 676076
rect 207004 676074 207604 676076
rect 243004 676074 243604 676076
rect 279004 676074 279604 676076
rect 315004 676074 315604 676076
rect 351004 676074 351604 676076
rect 387004 676074 387604 676076
rect 423004 676074 423604 676076
rect 459004 676074 459604 676076
rect 495004 676074 495604 676076
rect 531004 676074 531604 676076
rect 567004 676074 567604 676076
rect 590020 676074 590620 676076
rect -4816 673076 -4216 673078
rect 23404 673076 24004 673078
rect 59404 673076 60004 673078
rect 95404 673076 96004 673078
rect 131404 673076 132004 673078
rect 167404 673076 168004 673078
rect 203404 673076 204004 673078
rect 239404 673076 240004 673078
rect 275404 673076 276004 673078
rect 311404 673076 312004 673078
rect 347404 673076 348004 673078
rect 383404 673076 384004 673078
rect 419404 673076 420004 673078
rect 455404 673076 456004 673078
rect 491404 673076 492004 673078
rect 527404 673076 528004 673078
rect 563404 673076 564004 673078
rect 588140 673076 588740 673078
rect -4816 673054 588740 673076
rect -4816 672818 -4634 673054
rect -4398 672818 23586 673054
rect 23822 672818 59586 673054
rect 59822 672818 95586 673054
rect 95822 672818 131586 673054
rect 131822 672818 167586 673054
rect 167822 672818 203586 673054
rect 203822 672818 239586 673054
rect 239822 672818 275586 673054
rect 275822 672818 311586 673054
rect 311822 672818 347586 673054
rect 347822 672818 383586 673054
rect 383822 672818 419586 673054
rect 419822 672818 455586 673054
rect 455822 672818 491586 673054
rect 491822 672818 527586 673054
rect 527822 672818 563586 673054
rect 563822 672818 588322 673054
rect 588558 672818 588740 673054
rect -4816 672734 588740 672818
rect -4816 672498 -4634 672734
rect -4398 672498 23586 672734
rect 23822 672498 59586 672734
rect 59822 672498 95586 672734
rect 95822 672498 131586 672734
rect 131822 672498 167586 672734
rect 167822 672498 203586 672734
rect 203822 672498 239586 672734
rect 239822 672498 275586 672734
rect 275822 672498 311586 672734
rect 311822 672498 347586 672734
rect 347822 672498 383586 672734
rect 383822 672498 419586 672734
rect 419822 672498 455586 672734
rect 455822 672498 491586 672734
rect 491822 672498 527586 672734
rect 527822 672498 563586 672734
rect 563822 672498 588322 672734
rect 588558 672498 588740 672734
rect -4816 672476 588740 672498
rect -4816 672474 -4216 672476
rect 23404 672474 24004 672476
rect 59404 672474 60004 672476
rect 95404 672474 96004 672476
rect 131404 672474 132004 672476
rect 167404 672474 168004 672476
rect 203404 672474 204004 672476
rect 239404 672474 240004 672476
rect 275404 672474 276004 672476
rect 311404 672474 312004 672476
rect 347404 672474 348004 672476
rect 383404 672474 384004 672476
rect 419404 672474 420004 672476
rect 455404 672474 456004 672476
rect 491404 672474 492004 672476
rect 527404 672474 528004 672476
rect 563404 672474 564004 672476
rect 588140 672474 588740 672476
rect -2936 669476 -2336 669478
rect 19804 669476 20404 669478
rect 55804 669476 56404 669478
rect 91804 669476 92404 669478
rect 127804 669476 128404 669478
rect 163804 669476 164404 669478
rect 199804 669476 200404 669478
rect 235804 669476 236404 669478
rect 271804 669476 272404 669478
rect 307804 669476 308404 669478
rect 343804 669476 344404 669478
rect 379804 669476 380404 669478
rect 415804 669476 416404 669478
rect 451804 669476 452404 669478
rect 487804 669476 488404 669478
rect 523804 669476 524404 669478
rect 559804 669476 560404 669478
rect 586260 669476 586860 669478
rect -2936 669454 586860 669476
rect -2936 669218 -2754 669454
rect -2518 669218 19986 669454
rect 20222 669218 55986 669454
rect 56222 669218 91986 669454
rect 92222 669218 127986 669454
rect 128222 669218 163986 669454
rect 164222 669218 199986 669454
rect 200222 669218 235986 669454
rect 236222 669218 271986 669454
rect 272222 669218 307986 669454
rect 308222 669218 343986 669454
rect 344222 669218 379986 669454
rect 380222 669218 415986 669454
rect 416222 669218 451986 669454
rect 452222 669218 487986 669454
rect 488222 669218 523986 669454
rect 524222 669218 559986 669454
rect 560222 669218 586442 669454
rect 586678 669218 586860 669454
rect -2936 669134 586860 669218
rect -2936 668898 -2754 669134
rect -2518 668898 19986 669134
rect 20222 668898 55986 669134
rect 56222 668898 91986 669134
rect 92222 668898 127986 669134
rect 128222 668898 163986 669134
rect 164222 668898 199986 669134
rect 200222 668898 235986 669134
rect 236222 668898 271986 669134
rect 272222 668898 307986 669134
rect 308222 668898 343986 669134
rect 344222 668898 379986 669134
rect 380222 668898 415986 669134
rect 416222 668898 451986 669134
rect 452222 668898 487986 669134
rect 488222 668898 523986 669134
rect 524222 668898 559986 669134
rect 560222 668898 586442 669134
rect 586678 668898 586860 669134
rect -2936 668876 586860 668898
rect -2936 668874 -2336 668876
rect 19804 668874 20404 668876
rect 55804 668874 56404 668876
rect 91804 668874 92404 668876
rect 127804 668874 128404 668876
rect 163804 668874 164404 668876
rect 199804 668874 200404 668876
rect 235804 668874 236404 668876
rect 271804 668874 272404 668876
rect 307804 668874 308404 668876
rect 343804 668874 344404 668876
rect 379804 668874 380404 668876
rect 415804 668874 416404 668876
rect 451804 668874 452404 668876
rect 487804 668874 488404 668876
rect 523804 668874 524404 668876
rect 559804 668874 560404 668876
rect 586260 668874 586860 668876
rect -7636 662276 -7036 662278
rect 12604 662276 13204 662278
rect 48604 662276 49204 662278
rect 84604 662276 85204 662278
rect 120604 662276 121204 662278
rect 156604 662276 157204 662278
rect 192604 662276 193204 662278
rect 228604 662276 229204 662278
rect 264604 662276 265204 662278
rect 300604 662276 301204 662278
rect 336604 662276 337204 662278
rect 372604 662276 373204 662278
rect 408604 662276 409204 662278
rect 444604 662276 445204 662278
rect 480604 662276 481204 662278
rect 516604 662276 517204 662278
rect 552604 662276 553204 662278
rect 590960 662276 591560 662278
rect -8576 662254 592500 662276
rect -8576 662018 -7454 662254
rect -7218 662018 12786 662254
rect 13022 662018 48786 662254
rect 49022 662018 84786 662254
rect 85022 662018 120786 662254
rect 121022 662018 156786 662254
rect 157022 662018 192786 662254
rect 193022 662018 228786 662254
rect 229022 662018 264786 662254
rect 265022 662018 300786 662254
rect 301022 662018 336786 662254
rect 337022 662018 372786 662254
rect 373022 662018 408786 662254
rect 409022 662018 444786 662254
rect 445022 662018 480786 662254
rect 481022 662018 516786 662254
rect 517022 662018 552786 662254
rect 553022 662018 591142 662254
rect 591378 662018 592500 662254
rect -8576 661934 592500 662018
rect -8576 661698 -7454 661934
rect -7218 661698 12786 661934
rect 13022 661698 48786 661934
rect 49022 661698 84786 661934
rect 85022 661698 120786 661934
rect 121022 661698 156786 661934
rect 157022 661698 192786 661934
rect 193022 661698 228786 661934
rect 229022 661698 264786 661934
rect 265022 661698 300786 661934
rect 301022 661698 336786 661934
rect 337022 661698 372786 661934
rect 373022 661698 408786 661934
rect 409022 661698 444786 661934
rect 445022 661698 480786 661934
rect 481022 661698 516786 661934
rect 517022 661698 552786 661934
rect 553022 661698 591142 661934
rect 591378 661698 592500 661934
rect -8576 661676 592500 661698
rect -7636 661674 -7036 661676
rect 12604 661674 13204 661676
rect 48604 661674 49204 661676
rect 84604 661674 85204 661676
rect 120604 661674 121204 661676
rect 156604 661674 157204 661676
rect 192604 661674 193204 661676
rect 228604 661674 229204 661676
rect 264604 661674 265204 661676
rect 300604 661674 301204 661676
rect 336604 661674 337204 661676
rect 372604 661674 373204 661676
rect 408604 661674 409204 661676
rect 444604 661674 445204 661676
rect 480604 661674 481204 661676
rect 516604 661674 517204 661676
rect 552604 661674 553204 661676
rect 590960 661674 591560 661676
rect -5756 658676 -5156 658678
rect 9004 658676 9604 658678
rect 45004 658676 45604 658678
rect 81004 658676 81604 658678
rect 117004 658676 117604 658678
rect 153004 658676 153604 658678
rect 189004 658676 189604 658678
rect 225004 658676 225604 658678
rect 261004 658676 261604 658678
rect 297004 658676 297604 658678
rect 333004 658676 333604 658678
rect 369004 658676 369604 658678
rect 405004 658676 405604 658678
rect 441004 658676 441604 658678
rect 477004 658676 477604 658678
rect 513004 658676 513604 658678
rect 549004 658676 549604 658678
rect 589080 658676 589680 658678
rect -6696 658654 590620 658676
rect -6696 658418 -5574 658654
rect -5338 658418 9186 658654
rect 9422 658418 45186 658654
rect 45422 658418 81186 658654
rect 81422 658418 117186 658654
rect 117422 658418 153186 658654
rect 153422 658418 189186 658654
rect 189422 658418 225186 658654
rect 225422 658418 261186 658654
rect 261422 658418 297186 658654
rect 297422 658418 333186 658654
rect 333422 658418 369186 658654
rect 369422 658418 405186 658654
rect 405422 658418 441186 658654
rect 441422 658418 477186 658654
rect 477422 658418 513186 658654
rect 513422 658418 549186 658654
rect 549422 658418 589262 658654
rect 589498 658418 590620 658654
rect -6696 658334 590620 658418
rect -6696 658098 -5574 658334
rect -5338 658098 9186 658334
rect 9422 658098 45186 658334
rect 45422 658098 81186 658334
rect 81422 658098 117186 658334
rect 117422 658098 153186 658334
rect 153422 658098 189186 658334
rect 189422 658098 225186 658334
rect 225422 658098 261186 658334
rect 261422 658098 297186 658334
rect 297422 658098 333186 658334
rect 333422 658098 369186 658334
rect 369422 658098 405186 658334
rect 405422 658098 441186 658334
rect 441422 658098 477186 658334
rect 477422 658098 513186 658334
rect 513422 658098 549186 658334
rect 549422 658098 589262 658334
rect 589498 658098 590620 658334
rect -6696 658076 590620 658098
rect -5756 658074 -5156 658076
rect 9004 658074 9604 658076
rect 45004 658074 45604 658076
rect 81004 658074 81604 658076
rect 117004 658074 117604 658076
rect 153004 658074 153604 658076
rect 189004 658074 189604 658076
rect 225004 658074 225604 658076
rect 261004 658074 261604 658076
rect 297004 658074 297604 658076
rect 333004 658074 333604 658076
rect 369004 658074 369604 658076
rect 405004 658074 405604 658076
rect 441004 658074 441604 658076
rect 477004 658074 477604 658076
rect 513004 658074 513604 658076
rect 549004 658074 549604 658076
rect 589080 658074 589680 658076
rect -3876 655076 -3276 655078
rect 5404 655076 6004 655078
rect 41404 655076 42004 655078
rect 77404 655076 78004 655078
rect 113404 655076 114004 655078
rect 149404 655076 150004 655078
rect 185404 655076 186004 655078
rect 221404 655076 222004 655078
rect 257404 655076 258004 655078
rect 293404 655076 294004 655078
rect 329404 655076 330004 655078
rect 365404 655076 366004 655078
rect 401404 655076 402004 655078
rect 437404 655076 438004 655078
rect 473404 655076 474004 655078
rect 509404 655076 510004 655078
rect 545404 655076 546004 655078
rect 581404 655076 582004 655078
rect 587200 655076 587800 655078
rect -4816 655054 588740 655076
rect -4816 654818 -3694 655054
rect -3458 654818 5586 655054
rect 5822 654818 41586 655054
rect 41822 654818 77586 655054
rect 77822 654818 113586 655054
rect 113822 654818 149586 655054
rect 149822 654818 185586 655054
rect 185822 654818 221586 655054
rect 221822 654818 257586 655054
rect 257822 654818 293586 655054
rect 293822 654818 329586 655054
rect 329822 654818 365586 655054
rect 365822 654818 401586 655054
rect 401822 654818 437586 655054
rect 437822 654818 473586 655054
rect 473822 654818 509586 655054
rect 509822 654818 545586 655054
rect 545822 654818 581586 655054
rect 581822 654818 587382 655054
rect 587618 654818 588740 655054
rect -4816 654734 588740 654818
rect -4816 654498 -3694 654734
rect -3458 654498 5586 654734
rect 5822 654498 41586 654734
rect 41822 654498 77586 654734
rect 77822 654498 113586 654734
rect 113822 654498 149586 654734
rect 149822 654498 185586 654734
rect 185822 654498 221586 654734
rect 221822 654498 257586 654734
rect 257822 654498 293586 654734
rect 293822 654498 329586 654734
rect 329822 654498 365586 654734
rect 365822 654498 401586 654734
rect 401822 654498 437586 654734
rect 437822 654498 473586 654734
rect 473822 654498 509586 654734
rect 509822 654498 545586 654734
rect 545822 654498 581586 654734
rect 581822 654498 587382 654734
rect 587618 654498 588740 654734
rect -4816 654476 588740 654498
rect -3876 654474 -3276 654476
rect 5404 654474 6004 654476
rect 41404 654474 42004 654476
rect 77404 654474 78004 654476
rect 113404 654474 114004 654476
rect 149404 654474 150004 654476
rect 185404 654474 186004 654476
rect 221404 654474 222004 654476
rect 257404 654474 258004 654476
rect 293404 654474 294004 654476
rect 329404 654474 330004 654476
rect 365404 654474 366004 654476
rect 401404 654474 402004 654476
rect 437404 654474 438004 654476
rect 473404 654474 474004 654476
rect 509404 654474 510004 654476
rect 545404 654474 546004 654476
rect 581404 654474 582004 654476
rect 587200 654474 587800 654476
rect -1996 651476 -1396 651478
rect 1804 651476 2404 651478
rect 37804 651476 38404 651478
rect 73804 651476 74404 651478
rect 109804 651476 110404 651478
rect 145804 651476 146404 651478
rect 181804 651476 182404 651478
rect 217804 651476 218404 651478
rect 253804 651476 254404 651478
rect 289804 651476 290404 651478
rect 325804 651476 326404 651478
rect 361804 651476 362404 651478
rect 397804 651476 398404 651478
rect 433804 651476 434404 651478
rect 469804 651476 470404 651478
rect 505804 651476 506404 651478
rect 541804 651476 542404 651478
rect 577804 651476 578404 651478
rect 585320 651476 585920 651478
rect -2936 651454 586860 651476
rect -2936 651218 -1814 651454
rect -1578 651218 1986 651454
rect 2222 651218 37986 651454
rect 38222 651218 73986 651454
rect 74222 651218 109986 651454
rect 110222 651218 145986 651454
rect 146222 651218 181986 651454
rect 182222 651218 217986 651454
rect 218222 651218 253986 651454
rect 254222 651218 289986 651454
rect 290222 651218 325986 651454
rect 326222 651218 361986 651454
rect 362222 651218 397986 651454
rect 398222 651218 433986 651454
rect 434222 651218 469986 651454
rect 470222 651218 505986 651454
rect 506222 651218 541986 651454
rect 542222 651218 577986 651454
rect 578222 651218 585502 651454
rect 585738 651218 586860 651454
rect -2936 651134 586860 651218
rect -2936 650898 -1814 651134
rect -1578 650898 1986 651134
rect 2222 650898 37986 651134
rect 38222 650898 73986 651134
rect 74222 650898 109986 651134
rect 110222 650898 145986 651134
rect 146222 650898 181986 651134
rect 182222 650898 217986 651134
rect 218222 650898 253986 651134
rect 254222 650898 289986 651134
rect 290222 650898 325986 651134
rect 326222 650898 361986 651134
rect 362222 650898 397986 651134
rect 398222 650898 433986 651134
rect 434222 650898 469986 651134
rect 470222 650898 505986 651134
rect 506222 650898 541986 651134
rect 542222 650898 577986 651134
rect 578222 650898 585502 651134
rect 585738 650898 586860 651134
rect -2936 650876 586860 650898
rect -1996 650874 -1396 650876
rect 1804 650874 2404 650876
rect 37804 650874 38404 650876
rect 73804 650874 74404 650876
rect 109804 650874 110404 650876
rect 145804 650874 146404 650876
rect 181804 650874 182404 650876
rect 217804 650874 218404 650876
rect 253804 650874 254404 650876
rect 289804 650874 290404 650876
rect 325804 650874 326404 650876
rect 361804 650874 362404 650876
rect 397804 650874 398404 650876
rect 433804 650874 434404 650876
rect 469804 650874 470404 650876
rect 505804 650874 506404 650876
rect 541804 650874 542404 650876
rect 577804 650874 578404 650876
rect 585320 650874 585920 650876
rect -8576 644276 -7976 644278
rect 30604 644276 31204 644278
rect 66604 644276 67204 644278
rect 102604 644276 103204 644278
rect 138604 644276 139204 644278
rect 174604 644276 175204 644278
rect 210604 644276 211204 644278
rect 246604 644276 247204 644278
rect 282604 644276 283204 644278
rect 318604 644276 319204 644278
rect 354604 644276 355204 644278
rect 390604 644276 391204 644278
rect 426604 644276 427204 644278
rect 462604 644276 463204 644278
rect 498604 644276 499204 644278
rect 534604 644276 535204 644278
rect 570604 644276 571204 644278
rect 591900 644276 592500 644278
rect -8576 644254 592500 644276
rect -8576 644018 -8394 644254
rect -8158 644018 30786 644254
rect 31022 644018 66786 644254
rect 67022 644018 102786 644254
rect 103022 644018 138786 644254
rect 139022 644018 174786 644254
rect 175022 644018 210786 644254
rect 211022 644018 246786 644254
rect 247022 644018 282786 644254
rect 283022 644018 318786 644254
rect 319022 644018 354786 644254
rect 355022 644018 390786 644254
rect 391022 644018 426786 644254
rect 427022 644018 462786 644254
rect 463022 644018 498786 644254
rect 499022 644018 534786 644254
rect 535022 644018 570786 644254
rect 571022 644018 592082 644254
rect 592318 644018 592500 644254
rect -8576 643934 592500 644018
rect -8576 643698 -8394 643934
rect -8158 643698 30786 643934
rect 31022 643698 66786 643934
rect 67022 643698 102786 643934
rect 103022 643698 138786 643934
rect 139022 643698 174786 643934
rect 175022 643698 210786 643934
rect 211022 643698 246786 643934
rect 247022 643698 282786 643934
rect 283022 643698 318786 643934
rect 319022 643698 354786 643934
rect 355022 643698 390786 643934
rect 391022 643698 426786 643934
rect 427022 643698 462786 643934
rect 463022 643698 498786 643934
rect 499022 643698 534786 643934
rect 535022 643698 570786 643934
rect 571022 643698 592082 643934
rect 592318 643698 592500 643934
rect -8576 643676 592500 643698
rect -8576 643674 -7976 643676
rect 30604 643674 31204 643676
rect 66604 643674 67204 643676
rect 102604 643674 103204 643676
rect 138604 643674 139204 643676
rect 174604 643674 175204 643676
rect 210604 643674 211204 643676
rect 246604 643674 247204 643676
rect 282604 643674 283204 643676
rect 318604 643674 319204 643676
rect 354604 643674 355204 643676
rect 390604 643674 391204 643676
rect 426604 643674 427204 643676
rect 462604 643674 463204 643676
rect 498604 643674 499204 643676
rect 534604 643674 535204 643676
rect 570604 643674 571204 643676
rect 591900 643674 592500 643676
rect -6696 640676 -6096 640678
rect 27004 640676 27604 640678
rect 63004 640676 63604 640678
rect 99004 640676 99604 640678
rect 135004 640676 135604 640678
rect 171004 640676 171604 640678
rect 207004 640676 207604 640678
rect 243004 640676 243604 640678
rect 279004 640676 279604 640678
rect 315004 640676 315604 640678
rect 351004 640676 351604 640678
rect 387004 640676 387604 640678
rect 423004 640676 423604 640678
rect 459004 640676 459604 640678
rect 495004 640676 495604 640678
rect 531004 640676 531604 640678
rect 567004 640676 567604 640678
rect 590020 640676 590620 640678
rect -6696 640654 590620 640676
rect -6696 640418 -6514 640654
rect -6278 640418 27186 640654
rect 27422 640418 63186 640654
rect 63422 640418 99186 640654
rect 99422 640418 135186 640654
rect 135422 640418 171186 640654
rect 171422 640418 207186 640654
rect 207422 640418 243186 640654
rect 243422 640418 279186 640654
rect 279422 640418 315186 640654
rect 315422 640418 351186 640654
rect 351422 640418 387186 640654
rect 387422 640418 423186 640654
rect 423422 640418 459186 640654
rect 459422 640418 495186 640654
rect 495422 640418 531186 640654
rect 531422 640418 567186 640654
rect 567422 640418 590202 640654
rect 590438 640418 590620 640654
rect -6696 640334 590620 640418
rect -6696 640098 -6514 640334
rect -6278 640098 27186 640334
rect 27422 640098 63186 640334
rect 63422 640098 99186 640334
rect 99422 640098 135186 640334
rect 135422 640098 171186 640334
rect 171422 640098 207186 640334
rect 207422 640098 243186 640334
rect 243422 640098 279186 640334
rect 279422 640098 315186 640334
rect 315422 640098 351186 640334
rect 351422 640098 387186 640334
rect 387422 640098 423186 640334
rect 423422 640098 459186 640334
rect 459422 640098 495186 640334
rect 495422 640098 531186 640334
rect 531422 640098 567186 640334
rect 567422 640098 590202 640334
rect 590438 640098 590620 640334
rect -6696 640076 590620 640098
rect -6696 640074 -6096 640076
rect 27004 640074 27604 640076
rect 63004 640074 63604 640076
rect 99004 640074 99604 640076
rect 135004 640074 135604 640076
rect 171004 640074 171604 640076
rect 207004 640074 207604 640076
rect 243004 640074 243604 640076
rect 279004 640074 279604 640076
rect 315004 640074 315604 640076
rect 351004 640074 351604 640076
rect 387004 640074 387604 640076
rect 423004 640074 423604 640076
rect 459004 640074 459604 640076
rect 495004 640074 495604 640076
rect 531004 640074 531604 640076
rect 567004 640074 567604 640076
rect 590020 640074 590620 640076
rect -4816 637076 -4216 637078
rect 23404 637076 24004 637078
rect 59404 637076 60004 637078
rect 95404 637076 96004 637078
rect 131404 637076 132004 637078
rect 167404 637076 168004 637078
rect 203404 637076 204004 637078
rect 239404 637076 240004 637078
rect 275404 637076 276004 637078
rect 311404 637076 312004 637078
rect 347404 637076 348004 637078
rect 383404 637076 384004 637078
rect 419404 637076 420004 637078
rect 455404 637076 456004 637078
rect 491404 637076 492004 637078
rect 527404 637076 528004 637078
rect 563404 637076 564004 637078
rect 588140 637076 588740 637078
rect -4816 637054 588740 637076
rect -4816 636818 -4634 637054
rect -4398 636818 23586 637054
rect 23822 636818 59586 637054
rect 59822 636818 95586 637054
rect 95822 636818 131586 637054
rect 131822 636818 167586 637054
rect 167822 636818 203586 637054
rect 203822 636818 239586 637054
rect 239822 636818 275586 637054
rect 275822 636818 311586 637054
rect 311822 636818 347586 637054
rect 347822 636818 383586 637054
rect 383822 636818 419586 637054
rect 419822 636818 455586 637054
rect 455822 636818 491586 637054
rect 491822 636818 527586 637054
rect 527822 636818 563586 637054
rect 563822 636818 588322 637054
rect 588558 636818 588740 637054
rect -4816 636734 588740 636818
rect -4816 636498 -4634 636734
rect -4398 636498 23586 636734
rect 23822 636498 59586 636734
rect 59822 636498 95586 636734
rect 95822 636498 131586 636734
rect 131822 636498 167586 636734
rect 167822 636498 203586 636734
rect 203822 636498 239586 636734
rect 239822 636498 275586 636734
rect 275822 636498 311586 636734
rect 311822 636498 347586 636734
rect 347822 636498 383586 636734
rect 383822 636498 419586 636734
rect 419822 636498 455586 636734
rect 455822 636498 491586 636734
rect 491822 636498 527586 636734
rect 527822 636498 563586 636734
rect 563822 636498 588322 636734
rect 588558 636498 588740 636734
rect -4816 636476 588740 636498
rect -4816 636474 -4216 636476
rect 23404 636474 24004 636476
rect 59404 636474 60004 636476
rect 95404 636474 96004 636476
rect 131404 636474 132004 636476
rect 167404 636474 168004 636476
rect 203404 636474 204004 636476
rect 239404 636474 240004 636476
rect 275404 636474 276004 636476
rect 311404 636474 312004 636476
rect 347404 636474 348004 636476
rect 383404 636474 384004 636476
rect 419404 636474 420004 636476
rect 455404 636474 456004 636476
rect 491404 636474 492004 636476
rect 527404 636474 528004 636476
rect 563404 636474 564004 636476
rect 588140 636474 588740 636476
rect -2936 633476 -2336 633478
rect 19804 633476 20404 633478
rect 55804 633476 56404 633478
rect 91804 633476 92404 633478
rect 127804 633476 128404 633478
rect 163804 633476 164404 633478
rect 199804 633476 200404 633478
rect 235804 633476 236404 633478
rect 271804 633476 272404 633478
rect 307804 633476 308404 633478
rect 343804 633476 344404 633478
rect 379804 633476 380404 633478
rect 415804 633476 416404 633478
rect 451804 633476 452404 633478
rect 487804 633476 488404 633478
rect 523804 633476 524404 633478
rect 559804 633476 560404 633478
rect 586260 633476 586860 633478
rect -2936 633454 586860 633476
rect -2936 633218 -2754 633454
rect -2518 633218 19986 633454
rect 20222 633218 55986 633454
rect 56222 633218 91986 633454
rect 92222 633218 127986 633454
rect 128222 633218 163986 633454
rect 164222 633218 199986 633454
rect 200222 633218 235986 633454
rect 236222 633218 271986 633454
rect 272222 633218 307986 633454
rect 308222 633218 343986 633454
rect 344222 633218 379986 633454
rect 380222 633218 415986 633454
rect 416222 633218 451986 633454
rect 452222 633218 487986 633454
rect 488222 633218 523986 633454
rect 524222 633218 559986 633454
rect 560222 633218 586442 633454
rect 586678 633218 586860 633454
rect -2936 633134 586860 633218
rect -2936 632898 -2754 633134
rect -2518 632898 19986 633134
rect 20222 632898 55986 633134
rect 56222 632898 91986 633134
rect 92222 632898 127986 633134
rect 128222 632898 163986 633134
rect 164222 632898 199986 633134
rect 200222 632898 235986 633134
rect 236222 632898 271986 633134
rect 272222 632898 307986 633134
rect 308222 632898 343986 633134
rect 344222 632898 379986 633134
rect 380222 632898 415986 633134
rect 416222 632898 451986 633134
rect 452222 632898 487986 633134
rect 488222 632898 523986 633134
rect 524222 632898 559986 633134
rect 560222 632898 586442 633134
rect 586678 632898 586860 633134
rect -2936 632876 586860 632898
rect -2936 632874 -2336 632876
rect 19804 632874 20404 632876
rect 55804 632874 56404 632876
rect 91804 632874 92404 632876
rect 127804 632874 128404 632876
rect 163804 632874 164404 632876
rect 199804 632874 200404 632876
rect 235804 632874 236404 632876
rect 271804 632874 272404 632876
rect 307804 632874 308404 632876
rect 343804 632874 344404 632876
rect 379804 632874 380404 632876
rect 415804 632874 416404 632876
rect 451804 632874 452404 632876
rect 487804 632874 488404 632876
rect 523804 632874 524404 632876
rect 559804 632874 560404 632876
rect 586260 632874 586860 632876
rect -7636 626276 -7036 626278
rect 12604 626276 13204 626278
rect 48604 626276 49204 626278
rect 84604 626276 85204 626278
rect 120604 626276 121204 626278
rect 156604 626276 157204 626278
rect 192604 626276 193204 626278
rect 228604 626276 229204 626278
rect 264604 626276 265204 626278
rect 300604 626276 301204 626278
rect 336604 626276 337204 626278
rect 372604 626276 373204 626278
rect 408604 626276 409204 626278
rect 444604 626276 445204 626278
rect 480604 626276 481204 626278
rect 516604 626276 517204 626278
rect 552604 626276 553204 626278
rect 590960 626276 591560 626278
rect -8576 626254 592500 626276
rect -8576 626018 -7454 626254
rect -7218 626018 12786 626254
rect 13022 626018 48786 626254
rect 49022 626018 84786 626254
rect 85022 626018 120786 626254
rect 121022 626018 156786 626254
rect 157022 626018 192786 626254
rect 193022 626018 228786 626254
rect 229022 626018 264786 626254
rect 265022 626018 300786 626254
rect 301022 626018 336786 626254
rect 337022 626018 372786 626254
rect 373022 626018 408786 626254
rect 409022 626018 444786 626254
rect 445022 626018 480786 626254
rect 481022 626018 516786 626254
rect 517022 626018 552786 626254
rect 553022 626018 591142 626254
rect 591378 626018 592500 626254
rect -8576 625934 592500 626018
rect -8576 625698 -7454 625934
rect -7218 625698 12786 625934
rect 13022 625698 48786 625934
rect 49022 625698 84786 625934
rect 85022 625698 120786 625934
rect 121022 625698 156786 625934
rect 157022 625698 192786 625934
rect 193022 625698 228786 625934
rect 229022 625698 264786 625934
rect 265022 625698 300786 625934
rect 301022 625698 336786 625934
rect 337022 625698 372786 625934
rect 373022 625698 408786 625934
rect 409022 625698 444786 625934
rect 445022 625698 480786 625934
rect 481022 625698 516786 625934
rect 517022 625698 552786 625934
rect 553022 625698 591142 625934
rect 591378 625698 592500 625934
rect -8576 625676 592500 625698
rect -7636 625674 -7036 625676
rect 12604 625674 13204 625676
rect 48604 625674 49204 625676
rect 84604 625674 85204 625676
rect 120604 625674 121204 625676
rect 156604 625674 157204 625676
rect 192604 625674 193204 625676
rect 228604 625674 229204 625676
rect 264604 625674 265204 625676
rect 300604 625674 301204 625676
rect 336604 625674 337204 625676
rect 372604 625674 373204 625676
rect 408604 625674 409204 625676
rect 444604 625674 445204 625676
rect 480604 625674 481204 625676
rect 516604 625674 517204 625676
rect 552604 625674 553204 625676
rect 590960 625674 591560 625676
rect -5756 622676 -5156 622678
rect 9004 622676 9604 622678
rect 45004 622676 45604 622678
rect 81004 622676 81604 622678
rect 117004 622676 117604 622678
rect 153004 622676 153604 622678
rect 189004 622676 189604 622678
rect 225004 622676 225604 622678
rect 261004 622676 261604 622678
rect 297004 622676 297604 622678
rect 333004 622676 333604 622678
rect 369004 622676 369604 622678
rect 405004 622676 405604 622678
rect 441004 622676 441604 622678
rect 477004 622676 477604 622678
rect 513004 622676 513604 622678
rect 549004 622676 549604 622678
rect 589080 622676 589680 622678
rect -6696 622654 590620 622676
rect -6696 622418 -5574 622654
rect -5338 622418 9186 622654
rect 9422 622418 45186 622654
rect 45422 622418 81186 622654
rect 81422 622418 117186 622654
rect 117422 622418 153186 622654
rect 153422 622418 189186 622654
rect 189422 622418 225186 622654
rect 225422 622418 261186 622654
rect 261422 622418 297186 622654
rect 297422 622418 333186 622654
rect 333422 622418 369186 622654
rect 369422 622418 405186 622654
rect 405422 622418 441186 622654
rect 441422 622418 477186 622654
rect 477422 622418 513186 622654
rect 513422 622418 549186 622654
rect 549422 622418 589262 622654
rect 589498 622418 590620 622654
rect -6696 622334 590620 622418
rect -6696 622098 -5574 622334
rect -5338 622098 9186 622334
rect 9422 622098 45186 622334
rect 45422 622098 81186 622334
rect 81422 622098 117186 622334
rect 117422 622098 153186 622334
rect 153422 622098 189186 622334
rect 189422 622098 225186 622334
rect 225422 622098 261186 622334
rect 261422 622098 297186 622334
rect 297422 622098 333186 622334
rect 333422 622098 369186 622334
rect 369422 622098 405186 622334
rect 405422 622098 441186 622334
rect 441422 622098 477186 622334
rect 477422 622098 513186 622334
rect 513422 622098 549186 622334
rect 549422 622098 589262 622334
rect 589498 622098 590620 622334
rect -6696 622076 590620 622098
rect -5756 622074 -5156 622076
rect 9004 622074 9604 622076
rect 45004 622074 45604 622076
rect 81004 622074 81604 622076
rect 117004 622074 117604 622076
rect 153004 622074 153604 622076
rect 189004 622074 189604 622076
rect 225004 622074 225604 622076
rect 261004 622074 261604 622076
rect 297004 622074 297604 622076
rect 333004 622074 333604 622076
rect 369004 622074 369604 622076
rect 405004 622074 405604 622076
rect 441004 622074 441604 622076
rect 477004 622074 477604 622076
rect 513004 622074 513604 622076
rect 549004 622074 549604 622076
rect 589080 622074 589680 622076
rect -3876 619076 -3276 619078
rect 5404 619076 6004 619078
rect 41404 619076 42004 619078
rect 77404 619076 78004 619078
rect 113404 619076 114004 619078
rect 149404 619076 150004 619078
rect 185404 619076 186004 619078
rect 221404 619076 222004 619078
rect 257404 619076 258004 619078
rect 293404 619076 294004 619078
rect 329404 619076 330004 619078
rect 365404 619076 366004 619078
rect 401404 619076 402004 619078
rect 437404 619076 438004 619078
rect 473404 619076 474004 619078
rect 509404 619076 510004 619078
rect 545404 619076 546004 619078
rect 581404 619076 582004 619078
rect 587200 619076 587800 619078
rect -4816 619054 588740 619076
rect -4816 618818 -3694 619054
rect -3458 618818 5586 619054
rect 5822 618818 41586 619054
rect 41822 618818 77586 619054
rect 77822 618818 113586 619054
rect 113822 618818 149586 619054
rect 149822 618818 185586 619054
rect 185822 618818 221586 619054
rect 221822 618818 257586 619054
rect 257822 618818 293586 619054
rect 293822 618818 329586 619054
rect 329822 618818 365586 619054
rect 365822 618818 401586 619054
rect 401822 618818 437586 619054
rect 437822 618818 473586 619054
rect 473822 618818 509586 619054
rect 509822 618818 545586 619054
rect 545822 618818 581586 619054
rect 581822 618818 587382 619054
rect 587618 618818 588740 619054
rect -4816 618734 588740 618818
rect -4816 618498 -3694 618734
rect -3458 618498 5586 618734
rect 5822 618498 41586 618734
rect 41822 618498 77586 618734
rect 77822 618498 113586 618734
rect 113822 618498 149586 618734
rect 149822 618498 185586 618734
rect 185822 618498 221586 618734
rect 221822 618498 257586 618734
rect 257822 618498 293586 618734
rect 293822 618498 329586 618734
rect 329822 618498 365586 618734
rect 365822 618498 401586 618734
rect 401822 618498 437586 618734
rect 437822 618498 473586 618734
rect 473822 618498 509586 618734
rect 509822 618498 545586 618734
rect 545822 618498 581586 618734
rect 581822 618498 587382 618734
rect 587618 618498 588740 618734
rect -4816 618476 588740 618498
rect -3876 618474 -3276 618476
rect 5404 618474 6004 618476
rect 41404 618474 42004 618476
rect 77404 618474 78004 618476
rect 113404 618474 114004 618476
rect 149404 618474 150004 618476
rect 185404 618474 186004 618476
rect 221404 618474 222004 618476
rect 257404 618474 258004 618476
rect 293404 618474 294004 618476
rect 329404 618474 330004 618476
rect 365404 618474 366004 618476
rect 401404 618474 402004 618476
rect 437404 618474 438004 618476
rect 473404 618474 474004 618476
rect 509404 618474 510004 618476
rect 545404 618474 546004 618476
rect 581404 618474 582004 618476
rect 587200 618474 587800 618476
rect -1996 615476 -1396 615478
rect 1804 615476 2404 615478
rect 37804 615476 38404 615478
rect 73804 615476 74404 615478
rect 109804 615476 110404 615478
rect 145804 615476 146404 615478
rect 181804 615476 182404 615478
rect 217804 615476 218404 615478
rect 253804 615476 254404 615478
rect 289804 615476 290404 615478
rect 325804 615476 326404 615478
rect 361804 615476 362404 615478
rect 397804 615476 398404 615478
rect 433804 615476 434404 615478
rect 469804 615476 470404 615478
rect 505804 615476 506404 615478
rect 541804 615476 542404 615478
rect 577804 615476 578404 615478
rect 585320 615476 585920 615478
rect -2936 615454 586860 615476
rect -2936 615218 -1814 615454
rect -1578 615218 1986 615454
rect 2222 615218 37986 615454
rect 38222 615218 73986 615454
rect 74222 615218 109986 615454
rect 110222 615218 145986 615454
rect 146222 615218 181986 615454
rect 182222 615218 217986 615454
rect 218222 615218 253986 615454
rect 254222 615218 289986 615454
rect 290222 615218 325986 615454
rect 326222 615218 361986 615454
rect 362222 615218 397986 615454
rect 398222 615218 433986 615454
rect 434222 615218 469986 615454
rect 470222 615218 505986 615454
rect 506222 615218 541986 615454
rect 542222 615218 577986 615454
rect 578222 615218 585502 615454
rect 585738 615218 586860 615454
rect -2936 615134 586860 615218
rect -2936 614898 -1814 615134
rect -1578 614898 1986 615134
rect 2222 614898 37986 615134
rect 38222 614898 73986 615134
rect 74222 614898 109986 615134
rect 110222 614898 145986 615134
rect 146222 614898 181986 615134
rect 182222 614898 217986 615134
rect 218222 614898 253986 615134
rect 254222 614898 289986 615134
rect 290222 614898 325986 615134
rect 326222 614898 361986 615134
rect 362222 614898 397986 615134
rect 398222 614898 433986 615134
rect 434222 614898 469986 615134
rect 470222 614898 505986 615134
rect 506222 614898 541986 615134
rect 542222 614898 577986 615134
rect 578222 614898 585502 615134
rect 585738 614898 586860 615134
rect -2936 614876 586860 614898
rect -1996 614874 -1396 614876
rect 1804 614874 2404 614876
rect 37804 614874 38404 614876
rect 73804 614874 74404 614876
rect 109804 614874 110404 614876
rect 145804 614874 146404 614876
rect 181804 614874 182404 614876
rect 217804 614874 218404 614876
rect 253804 614874 254404 614876
rect 289804 614874 290404 614876
rect 325804 614874 326404 614876
rect 361804 614874 362404 614876
rect 397804 614874 398404 614876
rect 433804 614874 434404 614876
rect 469804 614874 470404 614876
rect 505804 614874 506404 614876
rect 541804 614874 542404 614876
rect 577804 614874 578404 614876
rect 585320 614874 585920 614876
rect -8576 608276 -7976 608278
rect 30604 608276 31204 608278
rect 66604 608276 67204 608278
rect 102604 608276 103204 608278
rect 138604 608276 139204 608278
rect 174604 608276 175204 608278
rect 210604 608276 211204 608278
rect 246604 608276 247204 608278
rect 282604 608276 283204 608278
rect 318604 608276 319204 608278
rect 354604 608276 355204 608278
rect 390604 608276 391204 608278
rect 426604 608276 427204 608278
rect 462604 608276 463204 608278
rect 498604 608276 499204 608278
rect 534604 608276 535204 608278
rect 570604 608276 571204 608278
rect 591900 608276 592500 608278
rect -8576 608254 592500 608276
rect -8576 608018 -8394 608254
rect -8158 608018 30786 608254
rect 31022 608018 66786 608254
rect 67022 608018 102786 608254
rect 103022 608018 138786 608254
rect 139022 608018 174786 608254
rect 175022 608018 210786 608254
rect 211022 608018 246786 608254
rect 247022 608018 282786 608254
rect 283022 608018 318786 608254
rect 319022 608018 354786 608254
rect 355022 608018 390786 608254
rect 391022 608018 426786 608254
rect 427022 608018 462786 608254
rect 463022 608018 498786 608254
rect 499022 608018 534786 608254
rect 535022 608018 570786 608254
rect 571022 608018 592082 608254
rect 592318 608018 592500 608254
rect -8576 607934 592500 608018
rect -8576 607698 -8394 607934
rect -8158 607698 30786 607934
rect 31022 607698 66786 607934
rect 67022 607698 102786 607934
rect 103022 607698 138786 607934
rect 139022 607698 174786 607934
rect 175022 607698 210786 607934
rect 211022 607698 246786 607934
rect 247022 607698 282786 607934
rect 283022 607698 318786 607934
rect 319022 607698 354786 607934
rect 355022 607698 390786 607934
rect 391022 607698 426786 607934
rect 427022 607698 462786 607934
rect 463022 607698 498786 607934
rect 499022 607698 534786 607934
rect 535022 607698 570786 607934
rect 571022 607698 592082 607934
rect 592318 607698 592500 607934
rect -8576 607676 592500 607698
rect -8576 607674 -7976 607676
rect 30604 607674 31204 607676
rect 66604 607674 67204 607676
rect 102604 607674 103204 607676
rect 138604 607674 139204 607676
rect 174604 607674 175204 607676
rect 210604 607674 211204 607676
rect 246604 607674 247204 607676
rect 282604 607674 283204 607676
rect 318604 607674 319204 607676
rect 354604 607674 355204 607676
rect 390604 607674 391204 607676
rect 426604 607674 427204 607676
rect 462604 607674 463204 607676
rect 498604 607674 499204 607676
rect 534604 607674 535204 607676
rect 570604 607674 571204 607676
rect 591900 607674 592500 607676
rect -6696 604676 -6096 604678
rect 27004 604676 27604 604678
rect 63004 604676 63604 604678
rect 99004 604676 99604 604678
rect 135004 604676 135604 604678
rect 171004 604676 171604 604678
rect 207004 604676 207604 604678
rect 243004 604676 243604 604678
rect 279004 604676 279604 604678
rect 315004 604676 315604 604678
rect 351004 604676 351604 604678
rect 387004 604676 387604 604678
rect 423004 604676 423604 604678
rect 459004 604676 459604 604678
rect 495004 604676 495604 604678
rect 531004 604676 531604 604678
rect 567004 604676 567604 604678
rect 590020 604676 590620 604678
rect -6696 604654 590620 604676
rect -6696 604418 -6514 604654
rect -6278 604418 27186 604654
rect 27422 604418 63186 604654
rect 63422 604418 99186 604654
rect 99422 604418 135186 604654
rect 135422 604418 171186 604654
rect 171422 604418 207186 604654
rect 207422 604418 243186 604654
rect 243422 604418 279186 604654
rect 279422 604418 315186 604654
rect 315422 604418 351186 604654
rect 351422 604418 387186 604654
rect 387422 604418 423186 604654
rect 423422 604418 459186 604654
rect 459422 604418 495186 604654
rect 495422 604418 531186 604654
rect 531422 604418 567186 604654
rect 567422 604418 590202 604654
rect 590438 604418 590620 604654
rect -6696 604334 590620 604418
rect -6696 604098 -6514 604334
rect -6278 604098 27186 604334
rect 27422 604098 63186 604334
rect 63422 604098 99186 604334
rect 99422 604098 135186 604334
rect 135422 604098 171186 604334
rect 171422 604098 207186 604334
rect 207422 604098 243186 604334
rect 243422 604098 279186 604334
rect 279422 604098 315186 604334
rect 315422 604098 351186 604334
rect 351422 604098 387186 604334
rect 387422 604098 423186 604334
rect 423422 604098 459186 604334
rect 459422 604098 495186 604334
rect 495422 604098 531186 604334
rect 531422 604098 567186 604334
rect 567422 604098 590202 604334
rect 590438 604098 590620 604334
rect -6696 604076 590620 604098
rect -6696 604074 -6096 604076
rect 27004 604074 27604 604076
rect 63004 604074 63604 604076
rect 99004 604074 99604 604076
rect 135004 604074 135604 604076
rect 171004 604074 171604 604076
rect 207004 604074 207604 604076
rect 243004 604074 243604 604076
rect 279004 604074 279604 604076
rect 315004 604074 315604 604076
rect 351004 604074 351604 604076
rect 387004 604074 387604 604076
rect 423004 604074 423604 604076
rect 459004 604074 459604 604076
rect 495004 604074 495604 604076
rect 531004 604074 531604 604076
rect 567004 604074 567604 604076
rect 590020 604074 590620 604076
rect -4816 601076 -4216 601078
rect 23404 601076 24004 601078
rect 59404 601076 60004 601078
rect 95404 601076 96004 601078
rect 131404 601076 132004 601078
rect 167404 601076 168004 601078
rect 203404 601076 204004 601078
rect 239404 601076 240004 601078
rect 275404 601076 276004 601078
rect 311404 601076 312004 601078
rect 347404 601076 348004 601078
rect 383404 601076 384004 601078
rect 419404 601076 420004 601078
rect 455404 601076 456004 601078
rect 491404 601076 492004 601078
rect 527404 601076 528004 601078
rect 563404 601076 564004 601078
rect 588140 601076 588740 601078
rect -4816 601054 588740 601076
rect -4816 600818 -4634 601054
rect -4398 600818 23586 601054
rect 23822 600818 59586 601054
rect 59822 600818 95586 601054
rect 95822 600818 131586 601054
rect 131822 600818 167586 601054
rect 167822 600818 203586 601054
rect 203822 600818 239586 601054
rect 239822 600818 275586 601054
rect 275822 600818 311586 601054
rect 311822 600818 347586 601054
rect 347822 600818 383586 601054
rect 383822 600818 419586 601054
rect 419822 600818 455586 601054
rect 455822 600818 491586 601054
rect 491822 600818 527586 601054
rect 527822 600818 563586 601054
rect 563822 600818 588322 601054
rect 588558 600818 588740 601054
rect -4816 600734 588740 600818
rect -4816 600498 -4634 600734
rect -4398 600498 23586 600734
rect 23822 600498 59586 600734
rect 59822 600498 95586 600734
rect 95822 600498 131586 600734
rect 131822 600498 167586 600734
rect 167822 600498 203586 600734
rect 203822 600498 239586 600734
rect 239822 600498 275586 600734
rect 275822 600498 311586 600734
rect 311822 600498 347586 600734
rect 347822 600498 383586 600734
rect 383822 600498 419586 600734
rect 419822 600498 455586 600734
rect 455822 600498 491586 600734
rect 491822 600498 527586 600734
rect 527822 600498 563586 600734
rect 563822 600498 588322 600734
rect 588558 600498 588740 600734
rect -4816 600476 588740 600498
rect -4816 600474 -4216 600476
rect 23404 600474 24004 600476
rect 59404 600474 60004 600476
rect 95404 600474 96004 600476
rect 131404 600474 132004 600476
rect 167404 600474 168004 600476
rect 203404 600474 204004 600476
rect 239404 600474 240004 600476
rect 275404 600474 276004 600476
rect 311404 600474 312004 600476
rect 347404 600474 348004 600476
rect 383404 600474 384004 600476
rect 419404 600474 420004 600476
rect 455404 600474 456004 600476
rect 491404 600474 492004 600476
rect 527404 600474 528004 600476
rect 563404 600474 564004 600476
rect 588140 600474 588740 600476
rect -2936 597476 -2336 597478
rect 19804 597476 20404 597478
rect 55804 597476 56404 597478
rect 91804 597476 92404 597478
rect 451804 597476 452404 597478
rect 487804 597476 488404 597478
rect 523804 597476 524404 597478
rect 559804 597476 560404 597478
rect 586260 597476 586860 597478
rect -2936 597454 108000 597476
rect -2936 597218 -2754 597454
rect -2518 597218 19986 597454
rect 20222 597218 55986 597454
rect 56222 597218 91986 597454
rect 92222 597218 108000 597454
rect -2936 597134 108000 597218
rect -2936 596898 -2754 597134
rect -2518 596898 19986 597134
rect 20222 596898 55986 597134
rect 56222 596898 91986 597134
rect 92222 596898 108000 597134
rect -2936 596876 108000 596898
rect 448000 597454 586860 597476
rect 448000 597218 451986 597454
rect 452222 597218 487986 597454
rect 488222 597218 523986 597454
rect 524222 597218 559986 597454
rect 560222 597218 586442 597454
rect 586678 597218 586860 597454
rect 448000 597134 586860 597218
rect 448000 596898 451986 597134
rect 452222 596898 487986 597134
rect 488222 596898 523986 597134
rect 524222 596898 559986 597134
rect 560222 596898 586442 597134
rect 586678 596898 586860 597134
rect 448000 596876 586860 596898
rect -2936 596874 -2336 596876
rect 19804 596874 20404 596876
rect 55804 596874 56404 596876
rect 91804 596874 92404 596876
rect 451804 596874 452404 596876
rect 487804 596874 488404 596876
rect 523804 596874 524404 596876
rect 559804 596874 560404 596876
rect 586260 596874 586860 596876
rect -7636 590276 -7036 590278
rect 12604 590276 13204 590278
rect 48604 590276 49204 590278
rect 84604 590276 85204 590278
rect 480604 590276 481204 590278
rect 516604 590276 517204 590278
rect 552604 590276 553204 590278
rect 590960 590276 591560 590278
rect -8576 590254 108000 590276
rect -8576 590018 -7454 590254
rect -7218 590018 12786 590254
rect 13022 590018 48786 590254
rect 49022 590018 84786 590254
rect 85022 590018 108000 590254
rect -8576 589934 108000 590018
rect -8576 589698 -7454 589934
rect -7218 589698 12786 589934
rect 13022 589698 48786 589934
rect 49022 589698 84786 589934
rect 85022 589698 108000 589934
rect -8576 589676 108000 589698
rect 448000 590254 592500 590276
rect 448000 590018 480786 590254
rect 481022 590018 516786 590254
rect 517022 590018 552786 590254
rect 553022 590018 591142 590254
rect 591378 590018 592500 590254
rect 448000 589934 592500 590018
rect 448000 589698 480786 589934
rect 481022 589698 516786 589934
rect 517022 589698 552786 589934
rect 553022 589698 591142 589934
rect 591378 589698 592500 589934
rect 448000 589676 592500 589698
rect -7636 589674 -7036 589676
rect 12604 589674 13204 589676
rect 48604 589674 49204 589676
rect 84604 589674 85204 589676
rect 480604 589674 481204 589676
rect 516604 589674 517204 589676
rect 552604 589674 553204 589676
rect 590960 589674 591560 589676
rect -5756 586676 -5156 586678
rect 9004 586676 9604 586678
rect 45004 586676 45604 586678
rect 81004 586676 81604 586678
rect 477004 586676 477604 586678
rect 513004 586676 513604 586678
rect 549004 586676 549604 586678
rect 589080 586676 589680 586678
rect -6696 586654 108000 586676
rect -6696 586418 -5574 586654
rect -5338 586418 9186 586654
rect 9422 586418 45186 586654
rect 45422 586418 81186 586654
rect 81422 586418 108000 586654
rect -6696 586334 108000 586418
rect -6696 586098 -5574 586334
rect -5338 586098 9186 586334
rect 9422 586098 45186 586334
rect 45422 586098 81186 586334
rect 81422 586098 108000 586334
rect -6696 586076 108000 586098
rect 448000 586654 590620 586676
rect 448000 586418 477186 586654
rect 477422 586418 513186 586654
rect 513422 586418 549186 586654
rect 549422 586418 589262 586654
rect 589498 586418 590620 586654
rect 448000 586334 590620 586418
rect 448000 586098 477186 586334
rect 477422 586098 513186 586334
rect 513422 586098 549186 586334
rect 549422 586098 589262 586334
rect 589498 586098 590620 586334
rect 448000 586076 590620 586098
rect -5756 586074 -5156 586076
rect 9004 586074 9604 586076
rect 45004 586074 45604 586076
rect 81004 586074 81604 586076
rect 477004 586074 477604 586076
rect 513004 586074 513604 586076
rect 549004 586074 549604 586076
rect 589080 586074 589680 586076
rect -3876 583076 -3276 583078
rect 5404 583076 6004 583078
rect 41404 583076 42004 583078
rect 77404 583076 78004 583078
rect 473404 583076 474004 583078
rect 509404 583076 510004 583078
rect 545404 583076 546004 583078
rect 581404 583076 582004 583078
rect 587200 583076 587800 583078
rect -4816 583054 133883 583076
rect -4816 582818 -3694 583054
rect -3458 582818 5586 583054
rect 5822 582818 41586 583054
rect 41822 582818 77586 583054
rect 77822 583000 133883 583054
rect 77822 582986 132090 583000
rect 77822 582971 130681 582986
rect 77822 582957 129280 582971
rect 77822 582942 127871 582957
rect 77822 582928 126391 582942
rect 77822 582913 124982 582928
rect 77822 582899 123581 582913
rect 77822 582818 123186 582899
rect -4816 582734 123186 582818
rect -4816 582498 -3694 582734
rect -3458 582498 5586 582734
rect 5822 582498 41586 582734
rect 41822 582498 77586 582734
rect 77822 582663 123186 582734
rect 123422 582677 123581 582899
rect 123817 582677 123901 582913
rect 124137 582677 124275 582913
rect 124511 582677 124595 582913
rect 124831 582692 124982 582913
rect 125218 582692 125302 582928
rect 125538 582692 125676 582928
rect 125912 582692 125996 582928
rect 126232 582706 126391 582928
rect 126627 582706 126711 582942
rect 126947 582706 127085 582942
rect 127321 582706 127405 582942
rect 127641 582721 127871 582942
rect 128107 582721 128191 582957
rect 128427 582721 128565 582957
rect 128801 582721 128885 582957
rect 129121 582735 129280 582957
rect 129516 582735 129600 582971
rect 129836 582735 129974 582971
rect 130210 582735 130294 582971
rect 130530 582750 130681 582971
rect 130917 582750 131001 582986
rect 131237 582750 131375 582986
rect 131611 582750 131695 582986
rect 131931 582764 132090 582986
rect 132326 582764 132410 583000
rect 132646 582764 132784 583000
rect 133020 582764 133104 583000
rect 133340 582764 133883 583000
rect 131931 582750 133883 582764
rect 130530 582735 133883 582750
rect 129121 582721 133883 582735
rect 127641 582706 133883 582721
rect 126232 582692 133883 582706
rect 124831 582677 133883 582692
rect 123422 582663 133883 582677
rect 77822 582498 133883 582663
rect -4816 582476 133883 582498
rect 448000 583054 588740 583076
rect 448000 582818 473586 583054
rect 473822 582818 509586 583054
rect 509822 582818 545586 583054
rect 545822 582818 581586 583054
rect 581822 582818 587382 583054
rect 587618 582818 588740 583054
rect 448000 582734 588740 582818
rect 448000 582498 473586 582734
rect 473822 582498 509586 582734
rect 509822 582498 545586 582734
rect 545822 582498 581586 582734
rect 581822 582498 587382 582734
rect 587618 582498 588740 582734
rect 448000 582476 588740 582498
rect -3876 582474 -3276 582476
rect 5404 582474 6004 582476
rect 41404 582474 42004 582476
rect 77404 582474 78004 582476
rect 473404 582474 474004 582476
rect 509404 582474 510004 582476
rect 545404 582474 546004 582476
rect 581404 582474 582004 582476
rect 587200 582474 587800 582476
rect -1996 579476 -1396 579478
rect 1804 579476 2404 579478
rect 37804 579476 38404 579478
rect 73804 579476 74404 579478
rect 469804 579476 470404 579478
rect 505804 579476 506404 579478
rect 541804 579476 542404 579478
rect 577804 579476 578404 579478
rect 585320 579476 585920 579478
rect -2936 579454 151560 579476
rect -2936 579218 -1814 579454
rect -1578 579218 1986 579454
rect 2222 579218 37986 579454
rect 38222 579218 73986 579454
rect 74222 579394 151560 579454
rect 74222 579380 149841 579394
rect 74222 579365 148432 579380
rect 74222 579351 147031 579365
rect 74222 579336 145622 579351
rect 74222 579322 144142 579336
rect 74222 579307 142733 579322
rect 74222 579293 141332 579307
rect 74222 579218 140937 579293
rect -2936 579134 140937 579218
rect -2936 578898 -1814 579134
rect -1578 578898 1986 579134
rect 2222 578898 37986 579134
rect 38222 578898 73986 579134
rect 74222 579057 140937 579134
rect 141173 579071 141332 579293
rect 141568 579071 141652 579307
rect 141888 579071 142026 579307
rect 142262 579071 142346 579307
rect 142582 579086 142733 579307
rect 142969 579086 143053 579322
rect 143289 579086 143427 579322
rect 143663 579086 143747 579322
rect 143983 579100 144142 579322
rect 144378 579100 144462 579336
rect 144698 579100 144836 579336
rect 145072 579100 145156 579336
rect 145392 579115 145622 579336
rect 145858 579115 145942 579351
rect 146178 579115 146316 579351
rect 146552 579115 146636 579351
rect 146872 579129 147031 579351
rect 147267 579129 147351 579365
rect 147587 579129 147725 579365
rect 147961 579129 148045 579365
rect 148281 579144 148432 579365
rect 148668 579144 148752 579380
rect 148988 579144 149126 579380
rect 149362 579144 149446 579380
rect 149682 579158 149841 579380
rect 150077 579158 150161 579394
rect 150397 579158 150535 579394
rect 150771 579158 150855 579394
rect 151091 579158 151560 579394
rect 149682 579144 151560 579158
rect 148281 579129 151560 579144
rect 146872 579115 151560 579129
rect 145392 579100 151560 579115
rect 143983 579086 151560 579100
rect 142582 579071 151560 579086
rect 141173 579057 151560 579071
rect 74222 578898 151560 579057
rect -2936 578876 151560 578898
rect 448000 579454 586860 579476
rect 448000 579218 469986 579454
rect 470222 579218 505986 579454
rect 506222 579218 541986 579454
rect 542222 579218 577986 579454
rect 578222 579218 585502 579454
rect 585738 579218 586860 579454
rect 448000 579134 586860 579218
rect 448000 578898 469986 579134
rect 470222 578898 505986 579134
rect 506222 578898 541986 579134
rect 542222 578898 577986 579134
rect 578222 578898 585502 579134
rect 585738 578898 586860 579134
rect 448000 578876 586860 578898
rect -1996 578874 -1396 578876
rect 1804 578874 2404 578876
rect 37804 578874 38404 578876
rect 73804 578874 74404 578876
rect 469804 578874 470404 578876
rect 505804 578874 506404 578876
rect 541804 578874 542404 578876
rect 577804 578874 578404 578876
rect 585320 578874 585920 578876
rect -8576 572276 -7976 572278
rect 30604 572276 31204 572278
rect 66604 572276 67204 572278
rect 102604 572276 103204 572278
rect 462604 572276 463204 572278
rect 498604 572276 499204 572278
rect 534604 572276 535204 572278
rect 570604 572276 571204 572278
rect 591900 572276 592500 572278
rect -8576 572254 108000 572276
rect -8576 572018 -8394 572254
rect -8158 572018 30786 572254
rect 31022 572018 66786 572254
rect 67022 572018 102786 572254
rect 103022 572018 108000 572254
rect -8576 571934 108000 572018
rect -8576 571698 -8394 571934
rect -8158 571698 30786 571934
rect 31022 571698 66786 571934
rect 67022 571698 102786 571934
rect 103022 571698 108000 571934
rect -8576 571676 108000 571698
rect 448000 572254 592500 572276
rect 448000 572018 462786 572254
rect 463022 572018 498786 572254
rect 499022 572018 534786 572254
rect 535022 572018 570786 572254
rect 571022 572018 592082 572254
rect 592318 572018 592500 572254
rect 448000 571934 592500 572018
rect 448000 571698 462786 571934
rect 463022 571698 498786 571934
rect 499022 571698 534786 571934
rect 535022 571698 570786 571934
rect 571022 571698 592082 571934
rect 592318 571698 592500 571934
rect 448000 571676 592500 571698
rect -8576 571674 -7976 571676
rect 30604 571674 31204 571676
rect 66604 571674 67204 571676
rect 102604 571674 103204 571676
rect 462604 571674 463204 571676
rect 498604 571674 499204 571676
rect 534604 571674 535204 571676
rect 570604 571674 571204 571676
rect 591900 571674 592500 571676
rect -6696 568676 -6096 568678
rect 27004 568676 27604 568678
rect 63004 568676 63604 568678
rect 99004 568676 99604 568678
rect 459004 568676 459604 568678
rect 495004 568676 495604 568678
rect 531004 568676 531604 568678
rect 567004 568676 567604 568678
rect 590020 568676 590620 568678
rect -6696 568654 108000 568676
rect -6696 568418 -6514 568654
rect -6278 568418 27186 568654
rect 27422 568418 63186 568654
rect 63422 568418 99186 568654
rect 99422 568418 108000 568654
rect -6696 568334 108000 568418
rect -6696 568098 -6514 568334
rect -6278 568098 27186 568334
rect 27422 568098 63186 568334
rect 63422 568098 99186 568334
rect 99422 568098 108000 568334
rect -6696 568076 108000 568098
rect 448000 568654 590620 568676
rect 448000 568418 459186 568654
rect 459422 568418 495186 568654
rect 495422 568418 531186 568654
rect 531422 568418 567186 568654
rect 567422 568418 590202 568654
rect 590438 568418 590620 568654
rect 448000 568334 590620 568418
rect 448000 568098 459186 568334
rect 459422 568098 495186 568334
rect 495422 568098 531186 568334
rect 531422 568098 567186 568334
rect 567422 568098 590202 568334
rect 590438 568098 590620 568334
rect 448000 568076 590620 568098
rect -6696 568074 -6096 568076
rect 27004 568074 27604 568076
rect 63004 568074 63604 568076
rect 99004 568074 99604 568076
rect 459004 568074 459604 568076
rect 495004 568074 495604 568076
rect 531004 568074 531604 568076
rect 567004 568074 567604 568076
rect 590020 568074 590620 568076
rect -4816 565076 -4216 565078
rect 23404 565076 24004 565078
rect 59404 565076 60004 565078
rect 95404 565076 96004 565078
rect 455404 565076 456004 565078
rect 491404 565076 492004 565078
rect 527404 565076 528004 565078
rect 563404 565076 564004 565078
rect 588140 565076 588740 565078
rect -4816 565054 108000 565076
rect -4816 564818 -4634 565054
rect -4398 564818 23586 565054
rect 23822 564818 59586 565054
rect 59822 564818 95586 565054
rect 95822 564818 108000 565054
rect -4816 564734 108000 564818
rect -4816 564498 -4634 564734
rect -4398 564498 23586 564734
rect 23822 564498 59586 564734
rect 59822 564498 95586 564734
rect 95822 564498 108000 564734
rect -4816 564476 108000 564498
rect 407589 565054 588740 565076
rect 407589 564959 455586 565054
rect 407589 564945 416812 564959
rect 407589 564930 415403 564945
rect 407589 564916 414002 564930
rect 407589 564901 412593 564916
rect 407589 564887 411113 564901
rect 407589 564872 409704 564887
rect 407589 564858 408303 564872
rect 407589 564622 407908 564858
rect 408144 564636 408303 564858
rect 408539 564636 408623 564872
rect 408859 564636 408997 564872
rect 409233 564636 409317 564872
rect 409553 564651 409704 564872
rect 409940 564651 410024 564887
rect 410260 564651 410398 564887
rect 410634 564651 410718 564887
rect 410954 564665 411113 564887
rect 411349 564665 411433 564901
rect 411669 564665 411807 564901
rect 412043 564665 412127 564901
rect 412363 564680 412593 564901
rect 412829 564680 412913 564916
rect 413149 564680 413287 564916
rect 413523 564680 413607 564916
rect 413843 564694 414002 564916
rect 414238 564694 414322 564930
rect 414558 564694 414696 564930
rect 414932 564694 415016 564930
rect 415252 564709 415403 564930
rect 415639 564709 415723 564945
rect 415959 564709 416097 564945
rect 416333 564709 416417 564945
rect 416653 564723 416812 564945
rect 417048 564723 417132 564959
rect 417368 564723 417506 564959
rect 417742 564723 417826 564959
rect 418062 564818 455586 564959
rect 455822 564818 491586 565054
rect 491822 564818 527586 565054
rect 527822 564818 563586 565054
rect 563822 564818 588322 565054
rect 588558 564818 588740 565054
rect 418062 564734 588740 564818
rect 418062 564723 455586 564734
rect 416653 564709 455586 564723
rect 415252 564694 455586 564709
rect 413843 564680 455586 564694
rect 412363 564665 455586 564680
rect 410954 564651 455586 564665
rect 409553 564636 455586 564651
rect 408144 564622 455586 564636
rect 407589 564498 455586 564622
rect 455822 564498 491586 564734
rect 491822 564498 527586 564734
rect 527822 564498 563586 564734
rect 563822 564498 588322 564734
rect 588558 564498 588740 564734
rect 407589 564476 588740 564498
rect -4816 564474 -4216 564476
rect 23404 564474 24004 564476
rect 59404 564474 60004 564476
rect 95404 564474 96004 564476
rect 455404 564474 456004 564476
rect 491404 564474 492004 564476
rect 527404 564474 528004 564476
rect 563404 564474 564004 564476
rect 588140 564474 588740 564476
rect -2936 561476 -2336 561478
rect 19804 561476 20404 561478
rect 55804 561476 56404 561478
rect 91804 561476 92404 561478
rect 451804 561476 452404 561478
rect 487804 561476 488404 561478
rect 523804 561476 524404 561478
rect 559804 561476 560404 561478
rect 586260 561476 586860 561478
rect -2936 561454 108000 561476
rect -2936 561218 -2754 561454
rect -2518 561218 19986 561454
rect 20222 561218 55986 561454
rect 56222 561218 91986 561454
rect 92222 561218 108000 561454
rect -2936 561134 108000 561218
rect -2936 560898 -2754 561134
rect -2518 560898 19986 561134
rect 20222 560898 55986 561134
rect 56222 560898 91986 561134
rect 92222 560898 108000 561134
rect -2936 560876 108000 560898
rect 425267 561454 586860 561476
rect 425267 561359 451986 561454
rect 425267 561345 434457 561359
rect 425267 561330 433048 561345
rect 425267 561316 431647 561330
rect 425267 561301 430238 561316
rect 425267 561287 428758 561301
rect 425267 561272 427349 561287
rect 425267 561258 425948 561272
rect 425267 561022 425553 561258
rect 425789 561036 425948 561258
rect 426184 561036 426268 561272
rect 426504 561036 426642 561272
rect 426878 561036 426962 561272
rect 427198 561051 427349 561272
rect 427585 561051 427669 561287
rect 427905 561051 428043 561287
rect 428279 561051 428363 561287
rect 428599 561065 428758 561287
rect 428994 561065 429078 561301
rect 429314 561065 429452 561301
rect 429688 561065 429772 561301
rect 430008 561080 430238 561301
rect 430474 561080 430558 561316
rect 430794 561080 430932 561316
rect 431168 561080 431252 561316
rect 431488 561094 431647 561316
rect 431883 561094 431967 561330
rect 432203 561094 432341 561330
rect 432577 561094 432661 561330
rect 432897 561109 433048 561330
rect 433284 561109 433368 561345
rect 433604 561109 433742 561345
rect 433978 561109 434062 561345
rect 434298 561123 434457 561345
rect 434693 561123 434777 561359
rect 435013 561123 435151 561359
rect 435387 561123 435471 561359
rect 435707 561218 451986 561359
rect 452222 561218 487986 561454
rect 488222 561218 523986 561454
rect 524222 561218 559986 561454
rect 560222 561218 586442 561454
rect 586678 561218 586860 561454
rect 435707 561134 586860 561218
rect 435707 561123 451986 561134
rect 434298 561109 451986 561123
rect 432897 561094 451986 561109
rect 431488 561080 451986 561094
rect 430008 561065 451986 561080
rect 428599 561051 451986 561065
rect 427198 561036 451986 561051
rect 425789 561022 451986 561036
rect 425267 560898 451986 561022
rect 452222 560898 487986 561134
rect 488222 560898 523986 561134
rect 524222 560898 559986 561134
rect 560222 560898 586442 561134
rect 586678 560898 586860 561134
rect 425267 560876 586860 560898
rect -2936 560874 -2336 560876
rect 19804 560874 20404 560876
rect 55804 560874 56404 560876
rect 91804 560874 92404 560876
rect 451804 560874 452404 560876
rect 487804 560874 488404 560876
rect 523804 560874 524404 560876
rect 559804 560874 560404 560876
rect 586260 560874 586860 560876
rect -7636 554276 -7036 554278
rect 12604 554276 13204 554278
rect 48604 554276 49204 554278
rect 84604 554276 85204 554278
rect 480604 554276 481204 554278
rect 516604 554276 517204 554278
rect 552604 554276 553204 554278
rect 590960 554276 591560 554278
rect -8576 554254 108000 554276
rect -8576 554018 -7454 554254
rect -7218 554018 12786 554254
rect 13022 554018 48786 554254
rect 49022 554018 84786 554254
rect 85022 554018 108000 554254
rect -8576 553934 108000 554018
rect -8576 553698 -7454 553934
rect -7218 553698 12786 553934
rect 13022 553698 48786 553934
rect 49022 553698 84786 553934
rect 85022 553698 108000 553934
rect -8576 553676 108000 553698
rect 448000 554254 592500 554276
rect 448000 554018 480786 554254
rect 481022 554018 516786 554254
rect 517022 554018 552786 554254
rect 553022 554018 591142 554254
rect 591378 554018 592500 554254
rect 448000 553934 592500 554018
rect 448000 553698 480786 553934
rect 481022 553698 516786 553934
rect 517022 553698 552786 553934
rect 553022 553698 591142 553934
rect 591378 553698 592500 553934
rect 448000 553676 592500 553698
rect -7636 553674 -7036 553676
rect 12604 553674 13204 553676
rect 48604 553674 49204 553676
rect 84604 553674 85204 553676
rect 480604 553674 481204 553676
rect 516604 553674 517204 553676
rect 552604 553674 553204 553676
rect 590960 553674 591560 553676
rect -5756 550676 -5156 550678
rect 9004 550676 9604 550678
rect 45004 550676 45604 550678
rect 81004 550676 81604 550678
rect 477004 550676 477604 550678
rect 513004 550676 513604 550678
rect 549004 550676 549604 550678
rect 589080 550676 589680 550678
rect -6696 550654 108000 550676
rect -6696 550418 -5574 550654
rect -5338 550418 9186 550654
rect 9422 550418 45186 550654
rect 45422 550418 81186 550654
rect 81422 550418 108000 550654
rect -6696 550334 108000 550418
rect -6696 550098 -5574 550334
rect -5338 550098 9186 550334
rect 9422 550098 45186 550334
rect 45422 550098 81186 550334
rect 81422 550098 108000 550334
rect -6696 550076 108000 550098
rect 448000 550654 590620 550676
rect 448000 550418 477186 550654
rect 477422 550418 513186 550654
rect 513422 550418 549186 550654
rect 549422 550418 589262 550654
rect 589498 550418 590620 550654
rect 448000 550334 590620 550418
rect 448000 550098 477186 550334
rect 477422 550098 513186 550334
rect 513422 550098 549186 550334
rect 549422 550098 589262 550334
rect 589498 550098 590620 550334
rect 448000 550076 590620 550098
rect -5756 550074 -5156 550076
rect 9004 550074 9604 550076
rect 45004 550074 45604 550076
rect 81004 550074 81604 550076
rect 477004 550074 477604 550076
rect 513004 550074 513604 550076
rect 549004 550074 549604 550076
rect 589080 550074 589680 550076
rect -3876 547076 -3276 547078
rect 5404 547076 6004 547078
rect 41404 547076 42004 547078
rect 77404 547076 78004 547078
rect 473404 547076 474004 547078
rect 509404 547076 510004 547078
rect 545404 547076 546004 547078
rect 581404 547076 582004 547078
rect 587200 547076 587800 547078
rect -4816 547054 133883 547076
rect -4816 546818 -3694 547054
rect -3458 546818 5586 547054
rect 5822 546818 41586 547054
rect 41822 546818 77586 547054
rect 77822 546976 133883 547054
rect 77822 546962 132177 546976
rect 77822 546947 130768 546962
rect 77822 546933 129367 546947
rect 77822 546918 127958 546933
rect 77822 546904 126478 546918
rect 77822 546889 125069 546904
rect 77822 546875 123668 546889
rect 77822 546818 123273 546875
rect -4816 546734 123273 546818
rect -4816 546498 -3694 546734
rect -3458 546498 5586 546734
rect 5822 546498 41586 546734
rect 41822 546498 77586 546734
rect 77822 546639 123273 546734
rect 123509 546653 123668 546875
rect 123904 546653 123988 546889
rect 124224 546653 124362 546889
rect 124598 546653 124682 546889
rect 124918 546668 125069 546889
rect 125305 546668 125389 546904
rect 125625 546668 125763 546904
rect 125999 546668 126083 546904
rect 126319 546682 126478 546904
rect 126714 546682 126798 546918
rect 127034 546682 127172 546918
rect 127408 546682 127492 546918
rect 127728 546697 127958 546918
rect 128194 546697 128278 546933
rect 128514 546697 128652 546933
rect 128888 546697 128972 546933
rect 129208 546711 129367 546933
rect 129603 546711 129687 546947
rect 129923 546711 130061 546947
rect 130297 546711 130381 546947
rect 130617 546726 130768 546947
rect 131004 546726 131088 546962
rect 131324 546726 131462 546962
rect 131698 546726 131782 546962
rect 132018 546740 132177 546962
rect 132413 546740 132497 546976
rect 132733 546740 132871 546976
rect 133107 546740 133191 546976
rect 133427 546740 133883 546976
rect 132018 546726 133883 546740
rect 130617 546711 133883 546726
rect 129208 546697 133883 546711
rect 127728 546682 133883 546697
rect 126319 546668 133883 546682
rect 124918 546653 133883 546668
rect 123509 546639 133883 546653
rect 77822 546498 133883 546639
rect -4816 546476 133883 546498
rect 448000 547054 588740 547076
rect 448000 546818 473586 547054
rect 473822 546818 509586 547054
rect 509822 546818 545586 547054
rect 545822 546818 581586 547054
rect 581822 546818 587382 547054
rect 587618 546818 588740 547054
rect 448000 546734 588740 546818
rect 448000 546498 473586 546734
rect 473822 546498 509586 546734
rect 509822 546498 545586 546734
rect 545822 546498 581586 546734
rect 581822 546498 587382 546734
rect 587618 546498 588740 546734
rect 448000 546476 588740 546498
rect -3876 546474 -3276 546476
rect 5404 546474 6004 546476
rect 41404 546474 42004 546476
rect 77404 546474 78004 546476
rect 473404 546474 474004 546476
rect 509404 546474 510004 546476
rect 545404 546474 546004 546476
rect 581404 546474 582004 546476
rect 587200 546474 587800 546476
rect -1996 543476 -1396 543478
rect 1804 543476 2404 543478
rect 37804 543476 38404 543478
rect 73804 543476 74404 543478
rect 469804 543476 470404 543478
rect 505804 543476 506404 543478
rect 541804 543476 542404 543478
rect 577804 543476 578404 543478
rect 585320 543476 585920 543478
rect -2936 543454 151560 543476
rect -2936 543218 -1814 543454
rect -1578 543218 1986 543454
rect 2222 543218 37986 543454
rect 38222 543218 73986 543454
rect 74222 543373 151560 543454
rect 74222 543359 149968 543373
rect 74222 543344 148559 543359
rect 74222 543330 147158 543344
rect 74222 543315 145749 543330
rect 74222 543301 144269 543315
rect 74222 543286 142860 543301
rect 74222 543272 141459 543286
rect 74222 543218 141064 543272
rect -2936 543134 141064 543218
rect -2936 542898 -1814 543134
rect -1578 542898 1986 543134
rect 2222 542898 37986 543134
rect 38222 542898 73986 543134
rect 74222 543036 141064 543134
rect 141300 543050 141459 543272
rect 141695 543050 141779 543286
rect 142015 543050 142153 543286
rect 142389 543050 142473 543286
rect 142709 543065 142860 543286
rect 143096 543065 143180 543301
rect 143416 543065 143554 543301
rect 143790 543065 143874 543301
rect 144110 543079 144269 543301
rect 144505 543079 144589 543315
rect 144825 543079 144963 543315
rect 145199 543079 145283 543315
rect 145519 543094 145749 543315
rect 145985 543094 146069 543330
rect 146305 543094 146443 543330
rect 146679 543094 146763 543330
rect 146999 543108 147158 543330
rect 147394 543108 147478 543344
rect 147714 543108 147852 543344
rect 148088 543108 148172 543344
rect 148408 543123 148559 543344
rect 148795 543123 148879 543359
rect 149115 543123 149253 543359
rect 149489 543123 149573 543359
rect 149809 543137 149968 543359
rect 150204 543137 150288 543373
rect 150524 543137 150662 543373
rect 150898 543137 150982 543373
rect 151218 543137 151560 543373
rect 149809 543123 151560 543137
rect 148408 543108 151560 543123
rect 146999 543094 151560 543108
rect 145519 543079 151560 543094
rect 144110 543065 151560 543079
rect 142709 543050 151560 543065
rect 141300 543036 151560 543050
rect 74222 542898 151560 543036
rect -2936 542876 151560 542898
rect 448000 543454 586860 543476
rect 448000 543218 469986 543454
rect 470222 543218 505986 543454
rect 506222 543218 541986 543454
rect 542222 543218 577986 543454
rect 578222 543218 585502 543454
rect 585738 543218 586860 543454
rect 448000 543134 586860 543218
rect 448000 542898 469986 543134
rect 470222 542898 505986 543134
rect 506222 542898 541986 543134
rect 542222 542898 577986 543134
rect 578222 542898 585502 543134
rect 585738 542898 586860 543134
rect 448000 542876 586860 542898
rect -1996 542874 -1396 542876
rect 1804 542874 2404 542876
rect 37804 542874 38404 542876
rect 73804 542874 74404 542876
rect 469804 542874 470404 542876
rect 505804 542874 506404 542876
rect 541804 542874 542404 542876
rect 577804 542874 578404 542876
rect 585320 542874 585920 542876
rect -8576 536276 -7976 536278
rect 30604 536276 31204 536278
rect 66604 536276 67204 536278
rect 102604 536276 103204 536278
rect 462604 536276 463204 536278
rect 498604 536276 499204 536278
rect 534604 536276 535204 536278
rect 570604 536276 571204 536278
rect 591900 536276 592500 536278
rect -8576 536254 108000 536276
rect -8576 536018 -8394 536254
rect -8158 536018 30786 536254
rect 31022 536018 66786 536254
rect 67022 536018 102786 536254
rect 103022 536018 108000 536254
rect -8576 535934 108000 536018
rect -8576 535698 -8394 535934
rect -8158 535698 30786 535934
rect 31022 535698 66786 535934
rect 67022 535698 102786 535934
rect 103022 535698 108000 535934
rect -8576 535676 108000 535698
rect 448000 536254 592500 536276
rect 448000 536018 462786 536254
rect 463022 536018 498786 536254
rect 499022 536018 534786 536254
rect 535022 536018 570786 536254
rect 571022 536018 592082 536254
rect 592318 536018 592500 536254
rect 448000 535934 592500 536018
rect 448000 535698 462786 535934
rect 463022 535698 498786 535934
rect 499022 535698 534786 535934
rect 535022 535698 570786 535934
rect 571022 535698 592082 535934
rect 592318 535698 592500 535934
rect 448000 535676 592500 535698
rect -8576 535674 -7976 535676
rect 30604 535674 31204 535676
rect 66604 535674 67204 535676
rect 102604 535674 103204 535676
rect 462604 535674 463204 535676
rect 498604 535674 499204 535676
rect 534604 535674 535204 535676
rect 570604 535674 571204 535676
rect 591900 535674 592500 535676
rect -6696 532676 -6096 532678
rect 27004 532676 27604 532678
rect 63004 532676 63604 532678
rect 99004 532676 99604 532678
rect 459004 532676 459604 532678
rect 495004 532676 495604 532678
rect 531004 532676 531604 532678
rect 567004 532676 567604 532678
rect 590020 532676 590620 532678
rect -6696 532654 108000 532676
rect -6696 532418 -6514 532654
rect -6278 532418 27186 532654
rect 27422 532418 63186 532654
rect 63422 532418 99186 532654
rect 99422 532418 108000 532654
rect -6696 532334 108000 532418
rect -6696 532098 -6514 532334
rect -6278 532098 27186 532334
rect 27422 532098 63186 532334
rect 63422 532098 99186 532334
rect 99422 532098 108000 532334
rect -6696 532076 108000 532098
rect 448000 532654 590620 532676
rect 448000 532418 459186 532654
rect 459422 532418 495186 532654
rect 495422 532418 531186 532654
rect 531422 532418 567186 532654
rect 567422 532418 590202 532654
rect 590438 532418 590620 532654
rect 448000 532334 590620 532418
rect 448000 532098 459186 532334
rect 459422 532098 495186 532334
rect 495422 532098 531186 532334
rect 531422 532098 567186 532334
rect 567422 532098 590202 532334
rect 590438 532098 590620 532334
rect 448000 532076 590620 532098
rect -6696 532074 -6096 532076
rect 27004 532074 27604 532076
rect 63004 532074 63604 532076
rect 99004 532074 99604 532076
rect 459004 532074 459604 532076
rect 495004 532074 495604 532076
rect 531004 532074 531604 532076
rect 567004 532074 567604 532076
rect 590020 532074 590620 532076
rect -4816 529076 -4216 529078
rect 23404 529076 24004 529078
rect 59404 529076 60004 529078
rect 95404 529076 96004 529078
rect 455404 529076 456004 529078
rect 491404 529076 492004 529078
rect 527404 529076 528004 529078
rect 563404 529076 564004 529078
rect 588140 529076 588740 529078
rect -4816 529054 108000 529076
rect -4816 528818 -4634 529054
rect -4398 528818 23586 529054
rect 23822 528818 59586 529054
rect 59822 528818 95586 529054
rect 95822 528818 108000 529054
rect -4816 528734 108000 528818
rect -4816 528498 -4634 528734
rect -4398 528498 23586 528734
rect 23822 528498 59586 528734
rect 59822 528498 95586 528734
rect 95822 528498 108000 528734
rect -4816 528476 108000 528498
rect 407589 529054 588740 529076
rect 407589 528998 455586 529054
rect 407589 528984 416736 528998
rect 407589 528969 415327 528984
rect 407589 528955 413926 528969
rect 407589 528940 412517 528955
rect 407589 528926 411037 528940
rect 407589 528911 409628 528926
rect 407589 528897 408227 528911
rect 407589 528661 407832 528897
rect 408068 528675 408227 528897
rect 408463 528675 408547 528911
rect 408783 528675 408921 528911
rect 409157 528675 409241 528911
rect 409477 528690 409628 528911
rect 409864 528690 409948 528926
rect 410184 528690 410322 528926
rect 410558 528690 410642 528926
rect 410878 528704 411037 528926
rect 411273 528704 411357 528940
rect 411593 528704 411731 528940
rect 411967 528704 412051 528940
rect 412287 528719 412517 528940
rect 412753 528719 412837 528955
rect 413073 528719 413211 528955
rect 413447 528719 413531 528955
rect 413767 528733 413926 528955
rect 414162 528733 414246 528969
rect 414482 528733 414620 528969
rect 414856 528733 414940 528969
rect 415176 528748 415327 528969
rect 415563 528748 415647 528984
rect 415883 528748 416021 528984
rect 416257 528748 416341 528984
rect 416577 528762 416736 528984
rect 416972 528762 417056 528998
rect 417292 528762 417430 528998
rect 417666 528762 417750 528998
rect 417986 528818 455586 528998
rect 455822 528818 491586 529054
rect 491822 528818 527586 529054
rect 527822 528818 563586 529054
rect 563822 528818 588322 529054
rect 588558 528818 588740 529054
rect 417986 528762 588740 528818
rect 416577 528748 588740 528762
rect 415176 528734 588740 528748
rect 415176 528733 455586 528734
rect 413767 528719 455586 528733
rect 412287 528704 455586 528719
rect 410878 528690 455586 528704
rect 409477 528675 455586 528690
rect 408068 528661 455586 528675
rect 407589 528498 455586 528661
rect 455822 528498 491586 528734
rect 491822 528498 527586 528734
rect 527822 528498 563586 528734
rect 563822 528498 588322 528734
rect 588558 528498 588740 528734
rect 407589 528476 588740 528498
rect -4816 528474 -4216 528476
rect 23404 528474 24004 528476
rect 59404 528474 60004 528476
rect 95404 528474 96004 528476
rect 455404 528474 456004 528476
rect 491404 528474 492004 528476
rect 527404 528474 528004 528476
rect 563404 528474 564004 528476
rect 588140 528474 588740 528476
rect -2936 525476 -2336 525478
rect 19804 525476 20404 525478
rect 55804 525476 56404 525478
rect 91804 525476 92404 525478
rect 451804 525476 452404 525478
rect 487804 525476 488404 525478
rect 523804 525476 524404 525478
rect 559804 525476 560404 525478
rect 586260 525476 586860 525478
rect -2936 525454 108000 525476
rect -2936 525218 -2754 525454
rect -2518 525218 19986 525454
rect 20222 525218 55986 525454
rect 56222 525218 91986 525454
rect 92222 525218 108000 525454
rect -2936 525134 108000 525218
rect -2936 524898 -2754 525134
rect -2518 524898 19986 525134
rect 20222 524898 55986 525134
rect 56222 524898 91986 525134
rect 92222 524898 108000 525134
rect -2936 524876 108000 524898
rect 425267 525454 586860 525476
rect 425267 525366 451986 525454
rect 425267 525352 434596 525366
rect 425267 525337 433187 525352
rect 425267 525323 431786 525337
rect 425267 525308 430377 525323
rect 425267 525294 428897 525308
rect 425267 525279 427488 525294
rect 425267 525265 426087 525279
rect 425267 525029 425692 525265
rect 425928 525043 426087 525265
rect 426323 525043 426407 525279
rect 426643 525043 426781 525279
rect 427017 525043 427101 525279
rect 427337 525058 427488 525279
rect 427724 525058 427808 525294
rect 428044 525058 428182 525294
rect 428418 525058 428502 525294
rect 428738 525072 428897 525294
rect 429133 525072 429217 525308
rect 429453 525072 429591 525308
rect 429827 525072 429911 525308
rect 430147 525087 430377 525308
rect 430613 525087 430697 525323
rect 430933 525087 431071 525323
rect 431307 525087 431391 525323
rect 431627 525101 431786 525323
rect 432022 525101 432106 525337
rect 432342 525101 432480 525337
rect 432716 525101 432800 525337
rect 433036 525116 433187 525337
rect 433423 525116 433507 525352
rect 433743 525116 433881 525352
rect 434117 525116 434201 525352
rect 434437 525130 434596 525352
rect 434832 525130 434916 525366
rect 435152 525130 435290 525366
rect 435526 525130 435610 525366
rect 435846 525218 451986 525366
rect 452222 525218 487986 525454
rect 488222 525218 523986 525454
rect 524222 525218 559986 525454
rect 560222 525218 586442 525454
rect 586678 525218 586860 525454
rect 435846 525134 586860 525218
rect 435846 525130 451986 525134
rect 434437 525116 451986 525130
rect 433036 525101 451986 525116
rect 431627 525087 451986 525101
rect 430147 525072 451986 525087
rect 428738 525058 451986 525072
rect 427337 525043 451986 525058
rect 425928 525029 451986 525043
rect 425267 524898 451986 525029
rect 452222 524898 487986 525134
rect 488222 524898 523986 525134
rect 524222 524898 559986 525134
rect 560222 524898 586442 525134
rect 586678 524898 586860 525134
rect 425267 524876 586860 524898
rect -2936 524874 -2336 524876
rect 19804 524874 20404 524876
rect 55804 524874 56404 524876
rect 91804 524874 92404 524876
rect 451804 524874 452404 524876
rect 487804 524874 488404 524876
rect 523804 524874 524404 524876
rect 559804 524874 560404 524876
rect 586260 524874 586860 524876
rect -7636 518276 -7036 518278
rect 12604 518276 13204 518278
rect 48604 518276 49204 518278
rect 84604 518276 85204 518278
rect 480604 518276 481204 518278
rect 516604 518276 517204 518278
rect 552604 518276 553204 518278
rect 590960 518276 591560 518278
rect -8576 518254 108000 518276
rect -8576 518018 -7454 518254
rect -7218 518018 12786 518254
rect 13022 518018 48786 518254
rect 49022 518018 84786 518254
rect 85022 518018 108000 518254
rect -8576 517934 108000 518018
rect -8576 517698 -7454 517934
rect -7218 517698 12786 517934
rect 13022 517698 48786 517934
rect 49022 517698 84786 517934
rect 85022 517698 108000 517934
rect -8576 517676 108000 517698
rect 448000 518254 592500 518276
rect 448000 518018 480786 518254
rect 481022 518018 516786 518254
rect 517022 518018 552786 518254
rect 553022 518018 591142 518254
rect 591378 518018 592500 518254
rect 448000 517934 592500 518018
rect 448000 517698 480786 517934
rect 481022 517698 516786 517934
rect 517022 517698 552786 517934
rect 553022 517698 591142 517934
rect 591378 517698 592500 517934
rect 448000 517676 592500 517698
rect -7636 517674 -7036 517676
rect 12604 517674 13204 517676
rect 48604 517674 49204 517676
rect 84604 517674 85204 517676
rect 480604 517674 481204 517676
rect 516604 517674 517204 517676
rect 552604 517674 553204 517676
rect 590960 517674 591560 517676
rect -5756 514676 -5156 514678
rect 9004 514676 9604 514678
rect 45004 514676 45604 514678
rect 81004 514676 81604 514678
rect 477004 514676 477604 514678
rect 513004 514676 513604 514678
rect 549004 514676 549604 514678
rect 589080 514676 589680 514678
rect -6696 514654 108000 514676
rect -6696 514418 -5574 514654
rect -5338 514418 9186 514654
rect 9422 514418 45186 514654
rect 45422 514418 81186 514654
rect 81422 514418 108000 514654
rect -6696 514334 108000 514418
rect -6696 514098 -5574 514334
rect -5338 514098 9186 514334
rect 9422 514098 45186 514334
rect 45422 514098 81186 514334
rect 81422 514098 108000 514334
rect -6696 514076 108000 514098
rect 448000 514654 590620 514676
rect 448000 514418 477186 514654
rect 477422 514418 513186 514654
rect 513422 514418 549186 514654
rect 549422 514418 589262 514654
rect 589498 514418 590620 514654
rect 448000 514334 590620 514418
rect 448000 514098 477186 514334
rect 477422 514098 513186 514334
rect 513422 514098 549186 514334
rect 549422 514098 589262 514334
rect 589498 514098 590620 514334
rect 448000 514076 590620 514098
rect -5756 514074 -5156 514076
rect 9004 514074 9604 514076
rect 45004 514074 45604 514076
rect 81004 514074 81604 514076
rect 477004 514074 477604 514076
rect 513004 514074 513604 514076
rect 549004 514074 549604 514076
rect 589080 514074 589680 514076
rect -3876 511076 -3276 511078
rect 5404 511076 6004 511078
rect 41404 511076 42004 511078
rect 77404 511076 78004 511078
rect 473404 511076 474004 511078
rect 509404 511076 510004 511078
rect 545404 511076 546004 511078
rect 581404 511076 582004 511078
rect 587200 511076 587800 511078
rect -4816 511054 133883 511076
rect -4816 510818 -3694 511054
rect -3458 510818 5586 511054
rect 5822 510818 41586 511054
rect 41822 510818 77586 511054
rect 77822 510973 133883 511054
rect 77822 510959 132137 510973
rect 77822 510944 130728 510959
rect 77822 510930 129327 510944
rect 77822 510915 127918 510930
rect 77822 510901 126438 510915
rect 77822 510886 125029 510901
rect 77822 510872 123628 510886
rect 77822 510818 123233 510872
rect -4816 510734 123233 510818
rect -4816 510498 -3694 510734
rect -3458 510498 5586 510734
rect 5822 510498 41586 510734
rect 41822 510498 77586 510734
rect 77822 510636 123233 510734
rect 123469 510650 123628 510872
rect 123864 510650 123948 510886
rect 124184 510650 124322 510886
rect 124558 510650 124642 510886
rect 124878 510665 125029 510886
rect 125265 510665 125349 510901
rect 125585 510665 125723 510901
rect 125959 510665 126043 510901
rect 126279 510679 126438 510901
rect 126674 510679 126758 510915
rect 126994 510679 127132 510915
rect 127368 510679 127452 510915
rect 127688 510694 127918 510915
rect 128154 510694 128238 510930
rect 128474 510694 128612 510930
rect 128848 510694 128932 510930
rect 129168 510708 129327 510930
rect 129563 510708 129647 510944
rect 129883 510708 130021 510944
rect 130257 510708 130341 510944
rect 130577 510723 130728 510944
rect 130964 510723 131048 510959
rect 131284 510723 131422 510959
rect 131658 510723 131742 510959
rect 131978 510737 132137 510959
rect 132373 510737 132457 510973
rect 132693 510737 132831 510973
rect 133067 510737 133151 510973
rect 133387 510737 133883 510973
rect 131978 510723 133883 510737
rect 130577 510708 133883 510723
rect 129168 510694 133883 510708
rect 127688 510679 133883 510694
rect 126279 510665 133883 510679
rect 124878 510650 133883 510665
rect 123469 510636 133883 510650
rect 77822 510498 133883 510636
rect -4816 510476 133883 510498
rect 448000 511054 588740 511076
rect 448000 510818 473586 511054
rect 473822 510818 509586 511054
rect 509822 510818 545586 511054
rect 545822 510818 581586 511054
rect 581822 510818 587382 511054
rect 587618 510818 588740 511054
rect 448000 510734 588740 510818
rect 448000 510498 473586 510734
rect 473822 510498 509586 510734
rect 509822 510498 545586 510734
rect 545822 510498 581586 510734
rect 581822 510498 587382 510734
rect 587618 510498 588740 510734
rect 448000 510476 588740 510498
rect -3876 510474 -3276 510476
rect 5404 510474 6004 510476
rect 41404 510474 42004 510476
rect 77404 510474 78004 510476
rect 473404 510474 474004 510476
rect 509404 510474 510004 510476
rect 545404 510474 546004 510476
rect 581404 510474 582004 510476
rect 587200 510474 587800 510476
rect -1996 507476 -1396 507478
rect 1804 507476 2404 507478
rect 37804 507476 38404 507478
rect 73804 507476 74404 507478
rect 469804 507476 470404 507478
rect 505804 507476 506404 507478
rect 541804 507476 542404 507478
rect 577804 507476 578404 507478
rect 585320 507476 585920 507478
rect -2936 507454 151560 507476
rect -2936 507218 -1814 507454
rect -1578 507218 1986 507454
rect 2222 507218 37986 507454
rect 38222 507218 73986 507454
rect 74222 507406 151560 507454
rect 74222 507392 150152 507406
rect 74222 507377 148743 507392
rect 74222 507363 147342 507377
rect 74222 507348 145933 507363
rect 74222 507334 144453 507348
rect 74222 507319 143044 507334
rect 74222 507305 141643 507319
rect 74222 507218 141248 507305
rect -2936 507134 141248 507218
rect -2936 506898 -1814 507134
rect -1578 506898 1986 507134
rect 2222 506898 37986 507134
rect 38222 506898 73986 507134
rect 74222 507069 141248 507134
rect 141484 507083 141643 507305
rect 141879 507083 141963 507319
rect 142199 507083 142337 507319
rect 142573 507083 142657 507319
rect 142893 507098 143044 507319
rect 143280 507098 143364 507334
rect 143600 507098 143738 507334
rect 143974 507098 144058 507334
rect 144294 507112 144453 507334
rect 144689 507112 144773 507348
rect 145009 507112 145147 507348
rect 145383 507112 145467 507348
rect 145703 507127 145933 507348
rect 146169 507127 146253 507363
rect 146489 507127 146627 507363
rect 146863 507127 146947 507363
rect 147183 507141 147342 507363
rect 147578 507141 147662 507377
rect 147898 507141 148036 507377
rect 148272 507141 148356 507377
rect 148592 507156 148743 507377
rect 148979 507156 149063 507392
rect 149299 507156 149437 507392
rect 149673 507156 149757 507392
rect 149993 507170 150152 507392
rect 150388 507170 150472 507406
rect 150708 507170 150846 507406
rect 151082 507170 151166 507406
rect 151402 507170 151560 507406
rect 149993 507156 151560 507170
rect 148592 507141 151560 507156
rect 147183 507127 151560 507141
rect 145703 507112 151560 507127
rect 144294 507098 151560 507112
rect 142893 507083 151560 507098
rect 141484 507069 151560 507083
rect 74222 506898 151560 507069
rect -2936 506876 151560 506898
rect 448000 507454 586860 507476
rect 448000 507218 469986 507454
rect 470222 507218 505986 507454
rect 506222 507218 541986 507454
rect 542222 507218 577986 507454
rect 578222 507218 585502 507454
rect 585738 507218 586860 507454
rect 448000 507134 586860 507218
rect 448000 506898 469986 507134
rect 470222 506898 505986 507134
rect 506222 506898 541986 507134
rect 542222 506898 577986 507134
rect 578222 506898 585502 507134
rect 585738 506898 586860 507134
rect 448000 506876 586860 506898
rect -1996 506874 -1396 506876
rect 1804 506874 2404 506876
rect 37804 506874 38404 506876
rect 73804 506874 74404 506876
rect 469804 506874 470404 506876
rect 505804 506874 506404 506876
rect 541804 506874 542404 506876
rect 577804 506874 578404 506876
rect 585320 506874 585920 506876
rect -8576 500276 -7976 500278
rect 30604 500276 31204 500278
rect 66604 500276 67204 500278
rect 102604 500276 103204 500278
rect 462604 500276 463204 500278
rect 498604 500276 499204 500278
rect 534604 500276 535204 500278
rect 570604 500276 571204 500278
rect 591900 500276 592500 500278
rect -8576 500254 108000 500276
rect -8576 500018 -8394 500254
rect -8158 500018 30786 500254
rect 31022 500018 66786 500254
rect 67022 500018 102786 500254
rect 103022 500018 108000 500254
rect -8576 499934 108000 500018
rect -8576 499698 -8394 499934
rect -8158 499698 30786 499934
rect 31022 499698 66786 499934
rect 67022 499698 102786 499934
rect 103022 499698 108000 499934
rect -8576 499676 108000 499698
rect 448000 500254 592500 500276
rect 448000 500018 462786 500254
rect 463022 500018 498786 500254
rect 499022 500018 534786 500254
rect 535022 500018 570786 500254
rect 571022 500018 592082 500254
rect 592318 500018 592500 500254
rect 448000 499934 592500 500018
rect 448000 499698 462786 499934
rect 463022 499698 498786 499934
rect 499022 499698 534786 499934
rect 535022 499698 570786 499934
rect 571022 499698 592082 499934
rect 592318 499698 592500 499934
rect 448000 499676 592500 499698
rect -8576 499674 -7976 499676
rect 30604 499674 31204 499676
rect 66604 499674 67204 499676
rect 102604 499674 103204 499676
rect 462604 499674 463204 499676
rect 498604 499674 499204 499676
rect 534604 499674 535204 499676
rect 570604 499674 571204 499676
rect 591900 499674 592500 499676
rect -6696 496676 -6096 496678
rect 27004 496676 27604 496678
rect 63004 496676 63604 496678
rect 99004 496676 99604 496678
rect 459004 496676 459604 496678
rect 495004 496676 495604 496678
rect 531004 496676 531604 496678
rect 567004 496676 567604 496678
rect 590020 496676 590620 496678
rect -6696 496654 108000 496676
rect -6696 496418 -6514 496654
rect -6278 496418 27186 496654
rect 27422 496418 63186 496654
rect 63422 496418 99186 496654
rect 99422 496418 108000 496654
rect -6696 496334 108000 496418
rect -6696 496098 -6514 496334
rect -6278 496098 27186 496334
rect 27422 496098 63186 496334
rect 63422 496098 99186 496334
rect 99422 496098 108000 496334
rect -6696 496076 108000 496098
rect 448000 496654 590620 496676
rect 448000 496418 459186 496654
rect 459422 496418 495186 496654
rect 495422 496418 531186 496654
rect 531422 496418 567186 496654
rect 567422 496418 590202 496654
rect 590438 496418 590620 496654
rect 448000 496334 590620 496418
rect 448000 496098 459186 496334
rect 459422 496098 495186 496334
rect 495422 496098 531186 496334
rect 531422 496098 567186 496334
rect 567422 496098 590202 496334
rect 590438 496098 590620 496334
rect 448000 496076 590620 496098
rect -6696 496074 -6096 496076
rect 27004 496074 27604 496076
rect 63004 496074 63604 496076
rect 99004 496074 99604 496076
rect 459004 496074 459604 496076
rect 495004 496074 495604 496076
rect 531004 496074 531604 496076
rect 567004 496074 567604 496076
rect 590020 496074 590620 496076
rect -4816 493076 -4216 493078
rect 23404 493076 24004 493078
rect 59404 493076 60004 493078
rect 95404 493076 96004 493078
rect 455404 493076 456004 493078
rect 491404 493076 492004 493078
rect 527404 493076 528004 493078
rect 563404 493076 564004 493078
rect 588140 493076 588740 493078
rect -4816 493054 108000 493076
rect -4816 492818 -4634 493054
rect -4398 492818 23586 493054
rect 23822 492818 59586 493054
rect 59822 492818 95586 493054
rect 95822 492818 108000 493054
rect -4816 492734 108000 492818
rect -4816 492498 -4634 492734
rect -4398 492498 23586 492734
rect 23822 492498 59586 492734
rect 59822 492498 95586 492734
rect 95822 492498 108000 492734
rect -4816 492476 108000 492498
rect 407589 493054 588740 493076
rect 407589 492971 455586 493054
rect 407589 492957 416716 492971
rect 407589 492942 415307 492957
rect 407589 492928 413906 492942
rect 407589 492913 412497 492928
rect 407589 492899 411017 492913
rect 407589 492884 409608 492899
rect 407589 492870 408207 492884
rect 407589 492634 407812 492870
rect 408048 492648 408207 492870
rect 408443 492648 408527 492884
rect 408763 492648 408901 492884
rect 409137 492648 409221 492884
rect 409457 492663 409608 492884
rect 409844 492663 409928 492899
rect 410164 492663 410302 492899
rect 410538 492663 410622 492899
rect 410858 492677 411017 492899
rect 411253 492677 411337 492913
rect 411573 492677 411711 492913
rect 411947 492677 412031 492913
rect 412267 492692 412497 492913
rect 412733 492692 412817 492928
rect 413053 492692 413191 492928
rect 413427 492692 413511 492928
rect 413747 492706 413906 492928
rect 414142 492706 414226 492942
rect 414462 492706 414600 492942
rect 414836 492706 414920 492942
rect 415156 492721 415307 492942
rect 415543 492721 415627 492957
rect 415863 492721 416001 492957
rect 416237 492721 416321 492957
rect 416557 492735 416716 492957
rect 416952 492735 417036 492971
rect 417272 492735 417410 492971
rect 417646 492735 417730 492971
rect 417966 492818 455586 492971
rect 455822 492818 491586 493054
rect 491822 492818 527586 493054
rect 527822 492818 563586 493054
rect 563822 492818 588322 493054
rect 588558 492818 588740 493054
rect 417966 492735 588740 492818
rect 416557 492734 588740 492735
rect 416557 492721 455586 492734
rect 415156 492706 455586 492721
rect 413747 492692 455586 492706
rect 412267 492677 455586 492692
rect 410858 492663 455586 492677
rect 409457 492648 455586 492663
rect 408048 492634 455586 492648
rect 407589 492498 455586 492634
rect 455822 492498 491586 492734
rect 491822 492498 527586 492734
rect 527822 492498 563586 492734
rect 563822 492498 588322 492734
rect 588558 492498 588740 492734
rect 407589 492476 588740 492498
rect -4816 492474 -4216 492476
rect 23404 492474 24004 492476
rect 59404 492474 60004 492476
rect 95404 492474 96004 492476
rect 455404 492474 456004 492476
rect 491404 492474 492004 492476
rect 527404 492474 528004 492476
rect 563404 492474 564004 492476
rect 588140 492474 588740 492476
rect -2936 489476 -2336 489478
rect 19804 489476 20404 489478
rect 55804 489476 56404 489478
rect 91804 489476 92404 489478
rect 451804 489476 452404 489478
rect 487804 489476 488404 489478
rect 523804 489476 524404 489478
rect 559804 489476 560404 489478
rect 586260 489476 586860 489478
rect -2936 489454 108000 489476
rect -2936 489218 -2754 489454
rect -2518 489218 19986 489454
rect 20222 489218 55986 489454
rect 56222 489218 91986 489454
rect 92222 489218 108000 489454
rect -2936 489134 108000 489218
rect -2936 488898 -2754 489134
rect -2518 488898 19986 489134
rect 20222 488898 55986 489134
rect 56222 488898 91986 489134
rect 92222 488898 108000 489134
rect -2936 488876 108000 488898
rect 425267 489454 586860 489476
rect 425267 489373 451986 489454
rect 425267 489359 434595 489373
rect 425267 489344 433186 489359
rect 425267 489330 431785 489344
rect 425267 489315 430376 489330
rect 425267 489301 428896 489315
rect 425267 489286 427487 489301
rect 425267 489272 426086 489286
rect 425267 489036 425691 489272
rect 425927 489050 426086 489272
rect 426322 489050 426406 489286
rect 426642 489050 426780 489286
rect 427016 489050 427100 489286
rect 427336 489065 427487 489286
rect 427723 489065 427807 489301
rect 428043 489065 428181 489301
rect 428417 489065 428501 489301
rect 428737 489079 428896 489301
rect 429132 489079 429216 489315
rect 429452 489079 429590 489315
rect 429826 489079 429910 489315
rect 430146 489094 430376 489315
rect 430612 489094 430696 489330
rect 430932 489094 431070 489330
rect 431306 489094 431390 489330
rect 431626 489108 431785 489330
rect 432021 489108 432105 489344
rect 432341 489108 432479 489344
rect 432715 489108 432799 489344
rect 433035 489123 433186 489344
rect 433422 489123 433506 489359
rect 433742 489123 433880 489359
rect 434116 489123 434200 489359
rect 434436 489137 434595 489359
rect 434831 489137 434915 489373
rect 435151 489137 435289 489373
rect 435525 489137 435609 489373
rect 435845 489218 451986 489373
rect 452222 489218 487986 489454
rect 488222 489218 523986 489454
rect 524222 489218 559986 489454
rect 560222 489218 586442 489454
rect 586678 489218 586860 489454
rect 435845 489137 586860 489218
rect 434436 489134 586860 489137
rect 434436 489123 451986 489134
rect 433035 489108 451986 489123
rect 431626 489094 451986 489108
rect 430146 489079 451986 489094
rect 428737 489065 451986 489079
rect 427336 489050 451986 489065
rect 425927 489036 451986 489050
rect 425267 488898 451986 489036
rect 452222 488898 487986 489134
rect 488222 488898 523986 489134
rect 524222 488898 559986 489134
rect 560222 488898 586442 489134
rect 586678 488898 586860 489134
rect 425267 488876 586860 488898
rect -2936 488874 -2336 488876
rect 19804 488874 20404 488876
rect 55804 488874 56404 488876
rect 91804 488874 92404 488876
rect 451804 488874 452404 488876
rect 487804 488874 488404 488876
rect 523804 488874 524404 488876
rect 559804 488874 560404 488876
rect 586260 488874 586860 488876
rect -7636 482276 -7036 482278
rect 12604 482276 13204 482278
rect 48604 482276 49204 482278
rect 84604 482276 85204 482278
rect 480604 482276 481204 482278
rect 516604 482276 517204 482278
rect 552604 482276 553204 482278
rect 590960 482276 591560 482278
rect -8576 482254 108000 482276
rect -8576 482018 -7454 482254
rect -7218 482018 12786 482254
rect 13022 482018 48786 482254
rect 49022 482018 84786 482254
rect 85022 482018 108000 482254
rect -8576 481934 108000 482018
rect -8576 481698 -7454 481934
rect -7218 481698 12786 481934
rect 13022 481698 48786 481934
rect 49022 481698 84786 481934
rect 85022 481698 108000 481934
rect -8576 481676 108000 481698
rect 448000 482254 592500 482276
rect 448000 482018 480786 482254
rect 481022 482018 516786 482254
rect 517022 482018 552786 482254
rect 553022 482018 591142 482254
rect 591378 482018 592500 482254
rect 448000 481934 592500 482018
rect 448000 481698 480786 481934
rect 481022 481698 516786 481934
rect 517022 481698 552786 481934
rect 553022 481698 591142 481934
rect 591378 481698 592500 481934
rect 448000 481676 592500 481698
rect -7636 481674 -7036 481676
rect 12604 481674 13204 481676
rect 48604 481674 49204 481676
rect 84604 481674 85204 481676
rect 480604 481674 481204 481676
rect 516604 481674 517204 481676
rect 552604 481674 553204 481676
rect 590960 481674 591560 481676
rect -5756 478676 -5156 478678
rect 9004 478676 9604 478678
rect 45004 478676 45604 478678
rect 81004 478676 81604 478678
rect 477004 478676 477604 478678
rect 513004 478676 513604 478678
rect 549004 478676 549604 478678
rect 589080 478676 589680 478678
rect -6696 478654 108000 478676
rect -6696 478418 -5574 478654
rect -5338 478418 9186 478654
rect 9422 478418 45186 478654
rect 45422 478418 81186 478654
rect 81422 478418 108000 478654
rect -6696 478334 108000 478418
rect -6696 478098 -5574 478334
rect -5338 478098 9186 478334
rect 9422 478098 45186 478334
rect 45422 478098 81186 478334
rect 81422 478098 108000 478334
rect -6696 478076 108000 478098
rect 448000 478654 590620 478676
rect 448000 478418 477186 478654
rect 477422 478418 513186 478654
rect 513422 478418 549186 478654
rect 549422 478418 589262 478654
rect 589498 478418 590620 478654
rect 448000 478334 590620 478418
rect 448000 478098 477186 478334
rect 477422 478098 513186 478334
rect 513422 478098 549186 478334
rect 549422 478098 589262 478334
rect 589498 478098 590620 478334
rect 448000 478076 590620 478098
rect -5756 478074 -5156 478076
rect 9004 478074 9604 478076
rect 45004 478074 45604 478076
rect 81004 478074 81604 478076
rect 477004 478074 477604 478076
rect 513004 478074 513604 478076
rect 549004 478074 549604 478076
rect 589080 478074 589680 478076
rect -3876 475076 -3276 475078
rect 5404 475076 6004 475078
rect 41404 475076 42004 475078
rect 77404 475076 78004 475078
rect 473404 475076 474004 475078
rect 509404 475076 510004 475078
rect 545404 475076 546004 475078
rect 581404 475076 582004 475078
rect 587200 475076 587800 475078
rect -4816 475054 108000 475076
rect -4816 474818 -3694 475054
rect -3458 474818 5586 475054
rect 5822 474818 41586 475054
rect 41822 474818 77586 475054
rect 77822 474818 108000 475054
rect -4816 474734 108000 474818
rect -4816 474498 -3694 474734
rect -3458 474498 5586 474734
rect 5822 474498 41586 474734
rect 41822 474498 77586 474734
rect 77822 474498 108000 474734
rect -4816 474476 108000 474498
rect 448000 475054 588740 475076
rect 448000 474818 473586 475054
rect 473822 474818 509586 475054
rect 509822 474818 545586 475054
rect 545822 474818 581586 475054
rect 581822 474818 587382 475054
rect 587618 474818 588740 475054
rect 448000 474734 588740 474818
rect 448000 474498 473586 474734
rect 473822 474498 509586 474734
rect 509822 474498 545586 474734
rect 545822 474498 581586 474734
rect 581822 474498 587382 474734
rect 587618 474498 588740 474734
rect 448000 474476 588740 474498
rect -3876 474474 -3276 474476
rect 5404 474474 6004 474476
rect 41404 474474 42004 474476
rect 77404 474474 78004 474476
rect 473404 474474 474004 474476
rect 509404 474474 510004 474476
rect 545404 474474 546004 474476
rect 581404 474474 582004 474476
rect 587200 474474 587800 474476
rect -1996 471476 -1396 471478
rect 1804 471476 2404 471478
rect 37804 471476 38404 471478
rect 73804 471476 74404 471478
rect -2936 471454 108000 471476
rect -2936 471218 -1814 471454
rect -1578 471218 1986 471454
rect 2222 471218 37986 471454
rect 38222 471218 73986 471454
rect 74222 471218 108000 471454
rect -2936 471134 108000 471218
rect -2936 470898 -1814 471134
rect -1578 470898 1986 471134
rect 2222 470898 37986 471134
rect 38222 470898 73986 471134
rect 74222 470898 108000 471134
rect 469804 471476 470404 471478
rect 505804 471476 506404 471478
rect 541804 471476 542404 471478
rect 577804 471476 578404 471478
rect 585320 471476 585920 471478
rect 448000 471454 586860 471476
rect 448000 471218 469986 471454
rect 470222 471218 505986 471454
rect 506222 471218 541986 471454
rect 542222 471218 577986 471454
rect 578222 471218 585502 471454
rect 585738 471218 586860 471454
rect 448000 471134 586860 471218
rect -2936 470876 108000 470898
rect 448000 470898 469986 471134
rect 470222 470898 505986 471134
rect 506222 470898 541986 471134
rect 542222 470898 577986 471134
rect 578222 470898 585502 471134
rect 585738 470898 586860 471134
rect 448000 470876 586860 470898
rect -1996 470874 -1396 470876
rect 1804 470874 2404 470876
rect 37804 470874 38404 470876
rect 73804 470874 74404 470876
rect 469804 470874 470404 470876
rect 505804 470874 506404 470876
rect 541804 470874 542404 470876
rect 577804 470874 578404 470876
rect 585320 470874 585920 470876
rect -8576 464276 -7976 464278
rect 30604 464276 31204 464278
rect 66604 464276 67204 464278
rect 102604 464276 103204 464278
rect 462604 464276 463204 464278
rect 498604 464276 499204 464278
rect 534604 464276 535204 464278
rect 570604 464276 571204 464278
rect 591900 464276 592500 464278
rect -8576 464254 108000 464276
rect -8576 464018 -8394 464254
rect -8158 464018 30786 464254
rect 31022 464018 66786 464254
rect 67022 464018 102786 464254
rect 103022 464018 108000 464254
rect -8576 463934 108000 464018
rect 448000 464254 592500 464276
rect 448000 464018 462786 464254
rect 463022 464018 498786 464254
rect 499022 464018 534786 464254
rect 535022 464018 570786 464254
rect 571022 464018 592082 464254
rect 592318 464018 592500 464254
rect -8576 463698 -8394 463934
rect -8158 463698 30786 463934
rect 31022 463698 66786 463934
rect 67022 463698 102786 463934
rect 103022 463698 108000 463934
rect -8576 463676 108000 463698
rect -8576 463674 -7976 463676
rect 30604 463674 31204 463676
rect 66604 463674 67204 463676
rect 102604 463674 103204 463676
rect 448000 463934 592500 464018
rect 448000 463698 462786 463934
rect 463022 463698 498786 463934
rect 499022 463698 534786 463934
rect 535022 463698 570786 463934
rect 571022 463698 592082 463934
rect 592318 463698 592500 463934
rect 448000 463676 592500 463698
rect 462604 463674 463204 463676
rect 498604 463674 499204 463676
rect 534604 463674 535204 463676
rect 570604 463674 571204 463676
rect 591900 463674 592500 463676
rect -6696 460676 -6096 460678
rect 27004 460676 27604 460678
rect 63004 460676 63604 460678
rect 99004 460676 99604 460678
rect -6696 460654 108000 460676
rect -6696 460418 -6514 460654
rect -6278 460418 27186 460654
rect 27422 460418 63186 460654
rect 63422 460418 99186 460654
rect 99422 460418 108000 460654
rect 459004 460676 459604 460678
rect 495004 460676 495604 460678
rect 531004 460676 531604 460678
rect 567004 460676 567604 460678
rect 590020 460676 590620 460678
rect 448000 460654 590620 460676
rect -6696 460334 108000 460418
rect -6696 460098 -6514 460334
rect -6278 460098 27186 460334
rect 27422 460098 63186 460334
rect 63422 460098 99186 460334
rect 99422 460098 108000 460334
rect -6696 460076 108000 460098
rect 448000 460418 459186 460654
rect 459422 460418 495186 460654
rect 495422 460418 531186 460654
rect 531422 460418 567186 460654
rect 567422 460418 590202 460654
rect 590438 460418 590620 460654
rect 448000 460334 590620 460418
rect 448000 460098 459186 460334
rect 459422 460098 495186 460334
rect 495422 460098 531186 460334
rect 531422 460098 567186 460334
rect 567422 460098 590202 460334
rect 590438 460098 590620 460334
rect 448000 460076 590620 460098
rect -6696 460074 -6096 460076
rect 27004 460074 27604 460076
rect 63004 460074 63604 460076
rect 99004 460074 99604 460076
rect 459004 460074 459604 460076
rect 495004 460074 495604 460076
rect 531004 460074 531604 460076
rect 567004 460074 567604 460076
rect 590020 460074 590620 460076
rect -4816 457076 -4216 457078
rect 23404 457076 24004 457078
rect 59404 457076 60004 457078
rect 95404 457076 96004 457078
rect -4816 457054 108000 457076
rect -4816 456818 -4634 457054
rect -4398 456818 23586 457054
rect 23822 456818 59586 457054
rect 59822 456818 95586 457054
rect 95822 456818 108000 457054
rect -4816 456734 108000 456818
rect -4816 456498 -4634 456734
rect -4398 456498 23586 456734
rect 23822 456498 59586 456734
rect 59822 456498 95586 456734
rect 95822 456498 108000 456734
rect 455404 457076 456004 457078
rect 491404 457076 492004 457078
rect 527404 457076 528004 457078
rect 563404 457076 564004 457078
rect 588140 457076 588740 457078
rect 448000 457054 588740 457076
rect 448000 456818 455586 457054
rect 455822 456818 491586 457054
rect 491822 456818 527586 457054
rect 527822 456818 563586 457054
rect 563822 456818 588322 457054
rect 588558 456818 588740 457054
rect 448000 456734 588740 456818
rect -4816 456476 108000 456498
rect 448000 456498 455586 456734
rect 455822 456498 491586 456734
rect 491822 456498 527586 456734
rect 527822 456498 563586 456734
rect 563822 456498 588322 456734
rect 588558 456498 588740 456734
rect 448000 456476 588740 456498
rect -4816 456474 -4216 456476
rect 23404 456474 24004 456476
rect 59404 456474 60004 456476
rect 95404 456474 96004 456476
rect 455404 456474 456004 456476
rect 491404 456474 492004 456476
rect 527404 456474 528004 456476
rect 563404 456474 564004 456476
rect 588140 456474 588740 456476
rect -2936 453476 -2336 453478
rect 19804 453476 20404 453478
rect 55804 453476 56404 453478
rect 91804 453476 92404 453478
rect -2936 453454 108000 453476
rect -2936 453218 -2754 453454
rect -2518 453218 19986 453454
rect 20222 453218 55986 453454
rect 56222 453218 91986 453454
rect 92222 453218 108000 453454
rect -2936 453134 108000 453218
rect -2936 452898 -2754 453134
rect -2518 452898 19986 453134
rect 20222 452898 55986 453134
rect 56222 452898 91986 453134
rect 92222 452898 108000 453134
rect -2936 452876 108000 452898
rect -2936 452874 -2336 452876
rect 19804 452874 20404 452876
rect 55804 452874 56404 452876
rect 91804 452874 92404 452876
rect 451804 453476 452404 453478
rect 487804 453476 488404 453478
rect 523804 453476 524404 453478
rect 559804 453476 560404 453478
rect 586260 453476 586860 453478
rect 448000 453454 586860 453476
rect 448000 453218 451986 453454
rect 452222 453218 487986 453454
rect 488222 453218 523986 453454
rect 524222 453218 559986 453454
rect 560222 453218 586442 453454
rect 586678 453218 586860 453454
rect 448000 453134 586860 453218
rect 448000 452898 451986 453134
rect 452222 452898 487986 453134
rect 488222 452898 523986 453134
rect 524222 452898 559986 453134
rect 560222 452898 586442 453134
rect 586678 452898 586860 453134
rect 448000 452876 586860 452898
rect 451804 452874 452404 452876
rect 487804 452874 488404 452876
rect 523804 452874 524404 452876
rect 559804 452874 560404 452876
rect 586260 452874 586860 452876
rect -7636 446276 -7036 446278
rect 12604 446276 13204 446278
rect 48604 446276 49204 446278
rect 84604 446276 85204 446278
rect 480604 446276 481204 446278
rect 516604 446276 517204 446278
rect 552604 446276 553204 446278
rect 590960 446276 591560 446278
rect -8576 446254 108000 446276
rect -8576 446018 -7454 446254
rect -7218 446018 12786 446254
rect 13022 446018 48786 446254
rect 49022 446018 84786 446254
rect 85022 446018 108000 446254
rect -8576 445934 108000 446018
rect -8576 445698 -7454 445934
rect -7218 445698 12786 445934
rect 13022 445698 48786 445934
rect 49022 445698 84786 445934
rect 85022 445698 108000 445934
rect -8576 445676 108000 445698
rect 448000 446254 592500 446276
rect 448000 446018 480786 446254
rect 481022 446018 516786 446254
rect 517022 446018 552786 446254
rect 553022 446018 591142 446254
rect 591378 446018 592500 446254
rect 448000 445934 592500 446018
rect 448000 445698 480786 445934
rect 481022 445698 516786 445934
rect 517022 445698 552786 445934
rect 553022 445698 591142 445934
rect 591378 445698 592500 445934
rect 448000 445676 592500 445698
rect -7636 445674 -7036 445676
rect 12604 445674 13204 445676
rect 48604 445674 49204 445676
rect 84604 445674 85204 445676
rect 480604 445674 481204 445676
rect 516604 445674 517204 445676
rect 552604 445674 553204 445676
rect 590960 445674 591560 445676
rect -5756 442676 -5156 442678
rect 9004 442676 9604 442678
rect 45004 442676 45604 442678
rect 81004 442676 81604 442678
rect 477004 442676 477604 442678
rect 513004 442676 513604 442678
rect 549004 442676 549604 442678
rect 589080 442676 589680 442678
rect -6696 442654 108000 442676
rect -6696 442418 -5574 442654
rect -5338 442418 9186 442654
rect 9422 442418 45186 442654
rect 45422 442418 81186 442654
rect 81422 442418 108000 442654
rect -6696 442334 108000 442418
rect -6696 442098 -5574 442334
rect -5338 442098 9186 442334
rect 9422 442098 45186 442334
rect 45422 442098 81186 442334
rect 81422 442098 108000 442334
rect -6696 442076 108000 442098
rect 448000 442654 590620 442676
rect 448000 442418 477186 442654
rect 477422 442418 513186 442654
rect 513422 442418 549186 442654
rect 549422 442418 589262 442654
rect 589498 442418 590620 442654
rect 448000 442334 590620 442418
rect 448000 442098 477186 442334
rect 477422 442098 513186 442334
rect 513422 442098 549186 442334
rect 549422 442098 589262 442334
rect 589498 442098 590620 442334
rect 448000 442076 590620 442098
rect -5756 442074 -5156 442076
rect 9004 442074 9604 442076
rect 45004 442074 45604 442076
rect 81004 442074 81604 442076
rect 477004 442074 477604 442076
rect 513004 442074 513604 442076
rect 549004 442074 549604 442076
rect 589080 442074 589680 442076
rect -3876 439076 -3276 439078
rect 5404 439076 6004 439078
rect 41404 439076 42004 439078
rect 77404 439076 78004 439078
rect -4816 439054 108000 439076
rect -4816 438818 -3694 439054
rect -3458 438818 5586 439054
rect 5822 438818 41586 439054
rect 41822 438818 77586 439054
rect 77822 438818 108000 439054
rect 473404 439076 474004 439078
rect 509404 439076 510004 439078
rect 545404 439076 546004 439078
rect 581404 439076 582004 439078
rect 587200 439076 587800 439078
rect 448000 439054 588740 439076
rect -4816 438734 108000 438818
rect -4816 438498 -3694 438734
rect -3458 438498 5586 438734
rect 5822 438498 41586 438734
rect 41822 438498 77586 438734
rect 77822 438498 108000 438734
rect -4816 438476 108000 438498
rect 448000 438818 473586 439054
rect 473822 438818 509586 439054
rect 509822 438818 545586 439054
rect 545822 438818 581586 439054
rect 581822 438818 587382 439054
rect 587618 438818 588740 439054
rect 448000 438734 588740 438818
rect 448000 438498 473586 438734
rect 473822 438498 509586 438734
rect 509822 438498 545586 438734
rect 545822 438498 581586 438734
rect 581822 438498 587382 438734
rect 587618 438498 588740 438734
rect 448000 438476 588740 438498
rect -3876 438474 -3276 438476
rect 5404 438474 6004 438476
rect 41404 438474 42004 438476
rect 77404 438474 78004 438476
rect 473404 438474 474004 438476
rect 509404 438474 510004 438476
rect 545404 438474 546004 438476
rect 581404 438474 582004 438476
rect 587200 438474 587800 438476
rect -1996 435476 -1396 435478
rect 1804 435476 2404 435478
rect 37804 435476 38404 435478
rect 73804 435476 74404 435478
rect -2936 435454 108000 435476
rect -2936 435218 -1814 435454
rect -1578 435218 1986 435454
rect 2222 435218 37986 435454
rect 38222 435218 73986 435454
rect 74222 435218 108000 435454
rect -2936 435134 108000 435218
rect -2936 434898 -1814 435134
rect -1578 434898 1986 435134
rect 2222 434898 37986 435134
rect 38222 434898 73986 435134
rect 74222 434898 108000 435134
rect 469804 435476 470404 435478
rect 505804 435476 506404 435478
rect 541804 435476 542404 435478
rect 577804 435476 578404 435478
rect 585320 435476 585920 435478
rect 448000 435454 586860 435476
rect 448000 435218 469986 435454
rect 470222 435218 505986 435454
rect 506222 435218 541986 435454
rect 542222 435218 577986 435454
rect 578222 435218 585502 435454
rect 585738 435218 586860 435454
rect 448000 435134 586860 435218
rect -2936 434876 108000 434898
rect 448000 434898 469986 435134
rect 470222 434898 505986 435134
rect 506222 434898 541986 435134
rect 542222 434898 577986 435134
rect 578222 434898 585502 435134
rect 585738 434898 586860 435134
rect 448000 434876 586860 434898
rect -1996 434874 -1396 434876
rect 1804 434874 2404 434876
rect 37804 434874 38404 434876
rect 73804 434874 74404 434876
rect 469804 434874 470404 434876
rect 505804 434874 506404 434876
rect 541804 434874 542404 434876
rect 577804 434874 578404 434876
rect 585320 434874 585920 434876
rect -8576 428276 -7976 428278
rect 30604 428276 31204 428278
rect 66604 428276 67204 428278
rect 102604 428276 103204 428278
rect 462604 428276 463204 428278
rect 498604 428276 499204 428278
rect 534604 428276 535204 428278
rect 570604 428276 571204 428278
rect 591900 428276 592500 428278
rect -8576 428254 108000 428276
rect -8576 428018 -8394 428254
rect -8158 428018 30786 428254
rect 31022 428018 66786 428254
rect 67022 428018 102786 428254
rect 103022 428018 108000 428254
rect -8576 427934 108000 428018
rect -8576 427698 -8394 427934
rect -8158 427698 30786 427934
rect 31022 427698 66786 427934
rect 67022 427698 102786 427934
rect 103022 427698 108000 427934
rect 448000 428254 592500 428276
rect 448000 428018 462786 428254
rect 463022 428018 498786 428254
rect 499022 428018 534786 428254
rect 535022 428018 570786 428254
rect 571022 428018 592082 428254
rect 592318 428018 592500 428254
rect 448000 427934 592500 428018
rect -8576 427676 108000 427698
rect -8576 427674 -7976 427676
rect 30604 427674 31204 427676
rect 66604 427674 67204 427676
rect 102604 427674 103204 427676
rect 448000 427698 462786 427934
rect 463022 427698 498786 427934
rect 499022 427698 534786 427934
rect 535022 427698 570786 427934
rect 571022 427698 592082 427934
rect 592318 427698 592500 427934
rect 448000 427676 592500 427698
rect 462604 427674 463204 427676
rect 498604 427674 499204 427676
rect 534604 427674 535204 427676
rect 570604 427674 571204 427676
rect 591900 427674 592500 427676
rect -6696 424676 -6096 424678
rect 27004 424676 27604 424678
rect 63004 424676 63604 424678
rect 99004 424676 99604 424678
rect 459004 424676 459604 424678
rect 495004 424676 495604 424678
rect 531004 424676 531604 424678
rect 567004 424676 567604 424678
rect 590020 424676 590620 424678
rect -6696 424654 108000 424676
rect -6696 424418 -6514 424654
rect -6278 424418 27186 424654
rect 27422 424418 63186 424654
rect 63422 424418 99186 424654
rect 99422 424418 108000 424654
rect -6696 424334 108000 424418
rect -6696 424098 -6514 424334
rect -6278 424098 27186 424334
rect 27422 424098 63186 424334
rect 63422 424098 99186 424334
rect 99422 424098 108000 424334
rect -6696 424076 108000 424098
rect 448000 424654 590620 424676
rect 448000 424418 459186 424654
rect 459422 424418 495186 424654
rect 495422 424418 531186 424654
rect 531422 424418 567186 424654
rect 567422 424418 590202 424654
rect 590438 424418 590620 424654
rect 448000 424334 590620 424418
rect 448000 424098 459186 424334
rect 459422 424098 495186 424334
rect 495422 424098 531186 424334
rect 531422 424098 567186 424334
rect 567422 424098 590202 424334
rect 590438 424098 590620 424334
rect 448000 424076 590620 424098
rect -6696 424074 -6096 424076
rect 27004 424074 27604 424076
rect 63004 424074 63604 424076
rect 99004 424074 99604 424076
rect 459004 424074 459604 424076
rect 495004 424074 495604 424076
rect 531004 424074 531604 424076
rect 567004 424074 567604 424076
rect 590020 424074 590620 424076
rect -4816 421076 -4216 421078
rect 23404 421076 24004 421078
rect 59404 421076 60004 421078
rect 95404 421076 96004 421078
rect -4816 421054 108000 421076
rect -4816 420818 -4634 421054
rect -4398 420818 23586 421054
rect 23822 420818 59586 421054
rect 59822 420818 95586 421054
rect 95822 420818 108000 421054
rect -4816 420734 108000 420818
rect -4816 420498 -4634 420734
rect -4398 420498 23586 420734
rect 23822 420498 59586 420734
rect 59822 420498 95586 420734
rect 95822 420498 108000 420734
rect 455404 421076 456004 421078
rect 491404 421076 492004 421078
rect 527404 421076 528004 421078
rect 563404 421076 564004 421078
rect 588140 421076 588740 421078
rect 448000 421054 588740 421076
rect 448000 420818 455586 421054
rect 455822 420818 491586 421054
rect 491822 420818 527586 421054
rect 527822 420818 563586 421054
rect 563822 420818 588322 421054
rect 588558 420818 588740 421054
rect 448000 420734 588740 420818
rect -4816 420476 108000 420498
rect 448000 420498 455586 420734
rect 455822 420498 491586 420734
rect 491822 420498 527586 420734
rect 527822 420498 563586 420734
rect 563822 420498 588322 420734
rect 588558 420498 588740 420734
rect 448000 420476 588740 420498
rect -4816 420474 -4216 420476
rect 23404 420474 24004 420476
rect 59404 420474 60004 420476
rect 95404 420474 96004 420476
rect 455404 420474 456004 420476
rect 491404 420474 492004 420476
rect 527404 420474 528004 420476
rect 563404 420474 564004 420476
rect 588140 420474 588740 420476
rect -2936 417476 -2336 417478
rect 19804 417476 20404 417478
rect 55804 417476 56404 417478
rect 91804 417476 92404 417478
rect -2936 417454 108000 417476
rect -2936 417218 -2754 417454
rect -2518 417218 19986 417454
rect 20222 417218 55986 417454
rect 56222 417218 91986 417454
rect 92222 417218 108000 417454
rect -2936 417134 108000 417218
rect -2936 416898 -2754 417134
rect -2518 416898 19986 417134
rect 20222 416898 55986 417134
rect 56222 416898 91986 417134
rect 92222 416898 108000 417134
rect -2936 416876 108000 416898
rect -2936 416874 -2336 416876
rect 19804 416874 20404 416876
rect 55804 416874 56404 416876
rect 91804 416874 92404 416876
rect 451804 417476 452404 417478
rect 487804 417476 488404 417478
rect 523804 417476 524404 417478
rect 559804 417476 560404 417478
rect 586260 417476 586860 417478
rect 448000 417454 586860 417476
rect 448000 417218 451986 417454
rect 452222 417218 487986 417454
rect 488222 417218 523986 417454
rect 524222 417218 559986 417454
rect 560222 417218 586442 417454
rect 586678 417218 586860 417454
rect 448000 417134 586860 417218
rect 448000 416898 451986 417134
rect 452222 416898 487986 417134
rect 488222 416898 523986 417134
rect 524222 416898 559986 417134
rect 560222 416898 586442 417134
rect 586678 416898 586860 417134
rect 448000 416876 586860 416898
rect 451804 416874 452404 416876
rect 487804 416874 488404 416876
rect 523804 416874 524404 416876
rect 559804 416874 560404 416876
rect 586260 416874 586860 416876
rect -7636 410276 -7036 410278
rect 12604 410276 13204 410278
rect 48604 410276 49204 410278
rect 84604 410276 85204 410278
rect 480604 410276 481204 410278
rect 516604 410276 517204 410278
rect 552604 410276 553204 410278
rect 590960 410276 591560 410278
rect -8576 410254 108000 410276
rect -8576 410018 -7454 410254
rect -7218 410018 12786 410254
rect 13022 410018 48786 410254
rect 49022 410018 84786 410254
rect 85022 410018 108000 410254
rect -8576 409934 108000 410018
rect -8576 409698 -7454 409934
rect -7218 409698 12786 409934
rect 13022 409698 48786 409934
rect 49022 409698 84786 409934
rect 85022 409698 108000 409934
rect -8576 409676 108000 409698
rect 448000 410254 592500 410276
rect 448000 410018 480786 410254
rect 481022 410018 516786 410254
rect 517022 410018 552786 410254
rect 553022 410018 591142 410254
rect 591378 410018 592500 410254
rect 448000 409934 592500 410018
rect 448000 409698 480786 409934
rect 481022 409698 516786 409934
rect 517022 409698 552786 409934
rect 553022 409698 591142 409934
rect 591378 409698 592500 409934
rect 448000 409676 592500 409698
rect -7636 409674 -7036 409676
rect 12604 409674 13204 409676
rect 48604 409674 49204 409676
rect 84604 409674 85204 409676
rect 480604 409674 481204 409676
rect 516604 409674 517204 409676
rect 552604 409674 553204 409676
rect 590960 409674 591560 409676
rect -5756 406676 -5156 406678
rect 9004 406676 9604 406678
rect 45004 406676 45604 406678
rect 81004 406676 81604 406678
rect 477004 406676 477604 406678
rect 513004 406676 513604 406678
rect 549004 406676 549604 406678
rect 589080 406676 589680 406678
rect -6696 406654 108000 406676
rect -6696 406418 -5574 406654
rect -5338 406418 9186 406654
rect 9422 406418 45186 406654
rect 45422 406418 81186 406654
rect 81422 406418 108000 406654
rect -6696 406334 108000 406418
rect -6696 406098 -5574 406334
rect -5338 406098 9186 406334
rect 9422 406098 45186 406334
rect 45422 406098 81186 406334
rect 81422 406098 108000 406334
rect -6696 406076 108000 406098
rect 448000 406654 590620 406676
rect 448000 406418 477186 406654
rect 477422 406418 513186 406654
rect 513422 406418 549186 406654
rect 549422 406418 589262 406654
rect 589498 406418 590620 406654
rect 448000 406334 590620 406418
rect 448000 406098 477186 406334
rect 477422 406098 513186 406334
rect 513422 406098 549186 406334
rect 549422 406098 589262 406334
rect 589498 406098 590620 406334
rect 448000 406076 590620 406098
rect -5756 406074 -5156 406076
rect 9004 406074 9604 406076
rect 45004 406074 45604 406076
rect 81004 406074 81604 406076
rect 477004 406074 477604 406076
rect 513004 406074 513604 406076
rect 549004 406074 549604 406076
rect 589080 406074 589680 406076
rect -3876 403076 -3276 403078
rect 5404 403076 6004 403078
rect 41404 403076 42004 403078
rect 77404 403076 78004 403078
rect -4816 403054 108000 403076
rect -4816 402818 -3694 403054
rect -3458 402818 5586 403054
rect 5822 402818 41586 403054
rect 41822 402818 77586 403054
rect 77822 402818 108000 403054
rect 473404 403076 474004 403078
rect 509404 403076 510004 403078
rect 545404 403076 546004 403078
rect 581404 403076 582004 403078
rect 587200 403076 587800 403078
rect 448000 403054 588740 403076
rect -4816 402734 108000 402818
rect -4816 402498 -3694 402734
rect -3458 402498 5586 402734
rect 5822 402498 41586 402734
rect 41822 402498 77586 402734
rect 77822 402498 108000 402734
rect -4816 402476 108000 402498
rect 448000 402818 473586 403054
rect 473822 402818 509586 403054
rect 509822 402818 545586 403054
rect 545822 402818 581586 403054
rect 581822 402818 587382 403054
rect 587618 402818 588740 403054
rect 448000 402734 588740 402818
rect 448000 402498 473586 402734
rect 473822 402498 509586 402734
rect 509822 402498 545586 402734
rect 545822 402498 581586 402734
rect 581822 402498 587382 402734
rect 587618 402498 588740 402734
rect 448000 402476 588740 402498
rect -3876 402474 -3276 402476
rect 5404 402474 6004 402476
rect 41404 402474 42004 402476
rect 77404 402474 78004 402476
rect 473404 402474 474004 402476
rect 509404 402474 510004 402476
rect 545404 402474 546004 402476
rect 581404 402474 582004 402476
rect 587200 402474 587800 402476
rect -1996 399476 -1396 399478
rect 1804 399476 2404 399478
rect 37804 399476 38404 399478
rect 73804 399476 74404 399478
rect -2936 399454 108000 399476
rect -2936 399218 -1814 399454
rect -1578 399218 1986 399454
rect 2222 399218 37986 399454
rect 38222 399218 73986 399454
rect 74222 399218 108000 399454
rect -2936 399134 108000 399218
rect -2936 398898 -1814 399134
rect -1578 398898 1986 399134
rect 2222 398898 37986 399134
rect 38222 398898 73986 399134
rect 74222 398898 108000 399134
rect 469804 399476 470404 399478
rect 505804 399476 506404 399478
rect 541804 399476 542404 399478
rect 577804 399476 578404 399478
rect 585320 399476 585920 399478
rect 448000 399454 586860 399476
rect 448000 399218 469986 399454
rect 470222 399218 505986 399454
rect 506222 399218 541986 399454
rect 542222 399218 577986 399454
rect 578222 399218 585502 399454
rect 585738 399218 586860 399454
rect 448000 399134 586860 399218
rect -2936 398876 108000 398898
rect 448000 398898 469986 399134
rect 470222 398898 505986 399134
rect 506222 398898 541986 399134
rect 542222 398898 577986 399134
rect 578222 398898 585502 399134
rect 585738 398898 586860 399134
rect 448000 398876 586860 398898
rect -1996 398874 -1396 398876
rect 1804 398874 2404 398876
rect 37804 398874 38404 398876
rect 73804 398874 74404 398876
rect 469804 398874 470404 398876
rect 505804 398874 506404 398876
rect 541804 398874 542404 398876
rect 577804 398874 578404 398876
rect 585320 398874 585920 398876
rect -8576 392276 -7976 392278
rect 30604 392276 31204 392278
rect 66604 392276 67204 392278
rect 102604 392276 103204 392278
rect 462604 392276 463204 392278
rect 498604 392276 499204 392278
rect 534604 392276 535204 392278
rect 570604 392276 571204 392278
rect 591900 392276 592500 392278
rect -8576 392254 108000 392276
rect -8576 392018 -8394 392254
rect -8158 392018 30786 392254
rect 31022 392018 66786 392254
rect 67022 392018 102786 392254
rect 103022 392018 108000 392254
rect -8576 391934 108000 392018
rect 448000 392254 592500 392276
rect 448000 392018 462786 392254
rect 463022 392018 498786 392254
rect 499022 392018 534786 392254
rect 535022 392018 570786 392254
rect 571022 392018 592082 392254
rect 592318 392018 592500 392254
rect -8576 391698 -8394 391934
rect -8158 391698 30786 391934
rect 31022 391698 66786 391934
rect 67022 391698 102786 391934
rect 103022 391698 108000 391934
rect -8576 391676 108000 391698
rect -8576 391674 -7976 391676
rect 30604 391674 31204 391676
rect 66604 391674 67204 391676
rect 102604 391674 103204 391676
rect 448000 391934 592500 392018
rect 448000 391698 462786 391934
rect 463022 391698 498786 391934
rect 499022 391698 534786 391934
rect 535022 391698 570786 391934
rect 571022 391698 592082 391934
rect 592318 391698 592500 391934
rect 448000 391676 592500 391698
rect 462604 391674 463204 391676
rect 498604 391674 499204 391676
rect 534604 391674 535204 391676
rect 570604 391674 571204 391676
rect 591900 391674 592500 391676
rect -6696 388676 -6096 388678
rect 27004 388676 27604 388678
rect 63004 388676 63604 388678
rect 99004 388676 99604 388678
rect -6696 388654 108000 388676
rect -6696 388418 -6514 388654
rect -6278 388418 27186 388654
rect 27422 388418 63186 388654
rect 63422 388418 99186 388654
rect 99422 388418 108000 388654
rect 459004 388676 459604 388678
rect 495004 388676 495604 388678
rect 531004 388676 531604 388678
rect 567004 388676 567604 388678
rect 590020 388676 590620 388678
rect 448000 388654 590620 388676
rect -6696 388334 108000 388418
rect -6696 388098 -6514 388334
rect -6278 388098 27186 388334
rect 27422 388098 63186 388334
rect 63422 388098 99186 388334
rect 99422 388098 108000 388334
rect -6696 388076 108000 388098
rect 448000 388418 459186 388654
rect 459422 388418 495186 388654
rect 495422 388418 531186 388654
rect 531422 388418 567186 388654
rect 567422 388418 590202 388654
rect 590438 388418 590620 388654
rect 448000 388334 590620 388418
rect 448000 388098 459186 388334
rect 459422 388098 495186 388334
rect 495422 388098 531186 388334
rect 531422 388098 567186 388334
rect 567422 388098 590202 388334
rect 590438 388098 590620 388334
rect 448000 388076 590620 388098
rect -6696 388074 -6096 388076
rect 27004 388074 27604 388076
rect 63004 388074 63604 388076
rect 99004 388074 99604 388076
rect 459004 388074 459604 388076
rect 495004 388074 495604 388076
rect 531004 388074 531604 388076
rect 567004 388074 567604 388076
rect 590020 388074 590620 388076
rect -4816 385076 -4216 385078
rect 23404 385076 24004 385078
rect 59404 385076 60004 385078
rect 95404 385076 96004 385078
rect -4816 385054 108000 385076
rect -4816 384818 -4634 385054
rect -4398 384818 23586 385054
rect 23822 384818 59586 385054
rect 59822 384818 95586 385054
rect 95822 384818 108000 385054
rect -4816 384734 108000 384818
rect -4816 384498 -4634 384734
rect -4398 384498 23586 384734
rect 23822 384498 59586 384734
rect 59822 384498 95586 384734
rect 95822 384498 108000 384734
rect 455404 385076 456004 385078
rect 491404 385076 492004 385078
rect 527404 385076 528004 385078
rect 563404 385076 564004 385078
rect 588140 385076 588740 385078
rect 448000 385054 588740 385076
rect 448000 384818 455586 385054
rect 455822 384818 491586 385054
rect 491822 384818 527586 385054
rect 527822 384818 563586 385054
rect 563822 384818 588322 385054
rect 588558 384818 588740 385054
rect 448000 384734 588740 384818
rect -4816 384476 108000 384498
rect 448000 384498 455586 384734
rect 455822 384498 491586 384734
rect 491822 384498 527586 384734
rect 527822 384498 563586 384734
rect 563822 384498 588322 384734
rect 588558 384498 588740 384734
rect 448000 384476 588740 384498
rect -4816 384474 -4216 384476
rect 23404 384474 24004 384476
rect 59404 384474 60004 384476
rect 95404 384474 96004 384476
rect 455404 384474 456004 384476
rect 491404 384474 492004 384476
rect 527404 384474 528004 384476
rect 563404 384474 564004 384476
rect 588140 384474 588740 384476
rect -2936 381476 -2336 381478
rect 19804 381476 20404 381478
rect 55804 381476 56404 381478
rect 91804 381476 92404 381478
rect -2936 381454 108000 381476
rect -2936 381218 -2754 381454
rect -2518 381218 19986 381454
rect 20222 381218 55986 381454
rect 56222 381218 91986 381454
rect 92222 381218 108000 381454
rect -2936 381134 108000 381218
rect -2936 380898 -2754 381134
rect -2518 380898 19986 381134
rect 20222 380898 55986 381134
rect 56222 380898 91986 381134
rect 92222 380898 108000 381134
rect -2936 380876 108000 380898
rect -2936 380874 -2336 380876
rect 19804 380874 20404 380876
rect 55804 380874 56404 380876
rect 91804 380874 92404 380876
rect 451804 381476 452404 381478
rect 487804 381476 488404 381478
rect 523804 381476 524404 381478
rect 559804 381476 560404 381478
rect 586260 381476 586860 381478
rect 448000 381454 586860 381476
rect 448000 381218 451986 381454
rect 452222 381218 487986 381454
rect 488222 381218 523986 381454
rect 524222 381218 559986 381454
rect 560222 381218 586442 381454
rect 586678 381218 586860 381454
rect 448000 381134 586860 381218
rect 448000 380898 451986 381134
rect 452222 380898 487986 381134
rect 488222 380898 523986 381134
rect 524222 380898 559986 381134
rect 560222 380898 586442 381134
rect 586678 380898 586860 381134
rect 448000 380876 586860 380898
rect 451804 380874 452404 380876
rect 487804 380874 488404 380876
rect 523804 380874 524404 380876
rect 559804 380874 560404 380876
rect 586260 380874 586860 380876
rect -7636 374276 -7036 374278
rect 12604 374276 13204 374278
rect 48604 374276 49204 374278
rect 84604 374276 85204 374278
rect 480604 374276 481204 374278
rect 516604 374276 517204 374278
rect 552604 374276 553204 374278
rect 590960 374276 591560 374278
rect -8576 374254 108000 374276
rect -8576 374018 -7454 374254
rect -7218 374018 12786 374254
rect 13022 374018 48786 374254
rect 49022 374018 84786 374254
rect 85022 374018 108000 374254
rect -8576 373934 108000 374018
rect -8576 373698 -7454 373934
rect -7218 373698 12786 373934
rect 13022 373698 48786 373934
rect 49022 373698 84786 373934
rect 85022 373698 108000 373934
rect -8576 373676 108000 373698
rect 448000 374254 592500 374276
rect 448000 374018 480786 374254
rect 481022 374018 516786 374254
rect 517022 374018 552786 374254
rect 553022 374018 591142 374254
rect 591378 374018 592500 374254
rect 448000 373934 592500 374018
rect 448000 373698 480786 373934
rect 481022 373698 516786 373934
rect 517022 373698 552786 373934
rect 553022 373698 591142 373934
rect 591378 373698 592500 373934
rect 448000 373676 592500 373698
rect -7636 373674 -7036 373676
rect 12604 373674 13204 373676
rect 48604 373674 49204 373676
rect 84604 373674 85204 373676
rect 480604 373674 481204 373676
rect 516604 373674 517204 373676
rect 552604 373674 553204 373676
rect 590960 373674 591560 373676
rect -5756 370676 -5156 370678
rect 9004 370676 9604 370678
rect 45004 370676 45604 370678
rect 81004 370676 81604 370678
rect 477004 370676 477604 370678
rect 513004 370676 513604 370678
rect 549004 370676 549604 370678
rect 589080 370676 589680 370678
rect -6696 370654 108000 370676
rect -6696 370418 -5574 370654
rect -5338 370418 9186 370654
rect 9422 370418 45186 370654
rect 45422 370418 81186 370654
rect 81422 370418 108000 370654
rect -6696 370334 108000 370418
rect -6696 370098 -5574 370334
rect -5338 370098 9186 370334
rect 9422 370098 45186 370334
rect 45422 370098 81186 370334
rect 81422 370098 108000 370334
rect -6696 370076 108000 370098
rect 448000 370654 590620 370676
rect 448000 370418 477186 370654
rect 477422 370418 513186 370654
rect 513422 370418 549186 370654
rect 549422 370418 589262 370654
rect 589498 370418 590620 370654
rect 448000 370334 590620 370418
rect 448000 370098 477186 370334
rect 477422 370098 513186 370334
rect 513422 370098 549186 370334
rect 549422 370098 589262 370334
rect 589498 370098 590620 370334
rect 448000 370076 590620 370098
rect -5756 370074 -5156 370076
rect 9004 370074 9604 370076
rect 45004 370074 45604 370076
rect 81004 370074 81604 370076
rect 477004 370074 477604 370076
rect 513004 370074 513604 370076
rect 549004 370074 549604 370076
rect 589080 370074 589680 370076
rect -3876 367076 -3276 367078
rect 5404 367076 6004 367078
rect 41404 367076 42004 367078
rect 77404 367076 78004 367078
rect -4816 367054 108000 367076
rect -4816 366818 -3694 367054
rect -3458 366818 5586 367054
rect 5822 366818 41586 367054
rect 41822 366818 77586 367054
rect 77822 366818 108000 367054
rect 473404 367076 474004 367078
rect 509404 367076 510004 367078
rect 545404 367076 546004 367078
rect 581404 367076 582004 367078
rect 587200 367076 587800 367078
rect 448000 367054 588740 367076
rect -4816 366734 108000 366818
rect -4816 366498 -3694 366734
rect -3458 366498 5586 366734
rect 5822 366498 41586 366734
rect 41822 366498 77586 366734
rect 77822 366498 108000 366734
rect -4816 366476 108000 366498
rect 448000 366818 473586 367054
rect 473822 366818 509586 367054
rect 509822 366818 545586 367054
rect 545822 366818 581586 367054
rect 581822 366818 587382 367054
rect 587618 366818 588740 367054
rect 448000 366734 588740 366818
rect 448000 366498 473586 366734
rect 473822 366498 509586 366734
rect 509822 366498 545586 366734
rect 545822 366498 581586 366734
rect 581822 366498 587382 366734
rect 587618 366498 588740 366734
rect 448000 366476 588740 366498
rect -3876 366474 -3276 366476
rect 5404 366474 6004 366476
rect 41404 366474 42004 366476
rect 77404 366474 78004 366476
rect 473404 366474 474004 366476
rect 509404 366474 510004 366476
rect 545404 366474 546004 366476
rect 581404 366474 582004 366476
rect 587200 366474 587800 366476
rect -1996 363476 -1396 363478
rect 1804 363476 2404 363478
rect 37804 363476 38404 363478
rect 73804 363476 74404 363478
rect -2936 363454 108000 363476
rect -2936 363218 -1814 363454
rect -1578 363218 1986 363454
rect 2222 363218 37986 363454
rect 38222 363218 73986 363454
rect 74222 363218 108000 363454
rect -2936 363134 108000 363218
rect -2936 362898 -1814 363134
rect -1578 362898 1986 363134
rect 2222 362898 37986 363134
rect 38222 362898 73986 363134
rect 74222 362898 108000 363134
rect 469804 363476 470404 363478
rect 505804 363476 506404 363478
rect 541804 363476 542404 363478
rect 577804 363476 578404 363478
rect 585320 363476 585920 363478
rect 448000 363454 586860 363476
rect 448000 363218 469986 363454
rect 470222 363218 505986 363454
rect 506222 363218 541986 363454
rect 542222 363218 577986 363454
rect 578222 363218 585502 363454
rect 585738 363218 586860 363454
rect 448000 363134 586860 363218
rect -2936 362876 108000 362898
rect 448000 362898 469986 363134
rect 470222 362898 505986 363134
rect 506222 362898 541986 363134
rect 542222 362898 577986 363134
rect 578222 362898 585502 363134
rect 585738 362898 586860 363134
rect 448000 362876 586860 362898
rect -1996 362874 -1396 362876
rect 1804 362874 2404 362876
rect 37804 362874 38404 362876
rect 73804 362874 74404 362876
rect 469804 362874 470404 362876
rect 505804 362874 506404 362876
rect 541804 362874 542404 362876
rect 577804 362874 578404 362876
rect 585320 362874 585920 362876
rect -8576 356276 -7976 356278
rect 30604 356276 31204 356278
rect 66604 356276 67204 356278
rect 102604 356276 103204 356278
rect 462604 356276 463204 356278
rect 498604 356276 499204 356278
rect 534604 356276 535204 356278
rect 570604 356276 571204 356278
rect 591900 356276 592500 356278
rect -8576 356254 108000 356276
rect -8576 356018 -8394 356254
rect -8158 356018 30786 356254
rect 31022 356018 66786 356254
rect 67022 356018 102786 356254
rect 103022 356018 108000 356254
rect -8576 355934 108000 356018
rect 448000 356254 592500 356276
rect 448000 356018 462786 356254
rect 463022 356018 498786 356254
rect 499022 356018 534786 356254
rect 535022 356018 570786 356254
rect 571022 356018 592082 356254
rect 592318 356018 592500 356254
rect -8576 355698 -8394 355934
rect -8158 355698 30786 355934
rect 31022 355698 66786 355934
rect 67022 355698 102786 355934
rect 103022 355698 108000 355934
rect -8576 355676 108000 355698
rect -8576 355674 -7976 355676
rect 30604 355674 31204 355676
rect 66604 355674 67204 355676
rect 102604 355674 103204 355676
rect 448000 355934 592500 356018
rect 448000 355698 462786 355934
rect 463022 355698 498786 355934
rect 499022 355698 534786 355934
rect 535022 355698 570786 355934
rect 571022 355698 592082 355934
rect 592318 355698 592500 355934
rect 448000 355676 592500 355698
rect 462604 355674 463204 355676
rect 498604 355674 499204 355676
rect 534604 355674 535204 355676
rect 570604 355674 571204 355676
rect 591900 355674 592500 355676
rect -6696 352676 -6096 352678
rect 27004 352676 27604 352678
rect 63004 352676 63604 352678
rect 99004 352676 99604 352678
rect -6696 352654 108000 352676
rect -6696 352418 -6514 352654
rect -6278 352418 27186 352654
rect 27422 352418 63186 352654
rect 63422 352418 99186 352654
rect 99422 352418 108000 352654
rect 459004 352676 459604 352678
rect 495004 352676 495604 352678
rect 531004 352676 531604 352678
rect 567004 352676 567604 352678
rect 590020 352676 590620 352678
rect 448000 352654 590620 352676
rect -6696 352334 108000 352418
rect -6696 352098 -6514 352334
rect -6278 352098 27186 352334
rect 27422 352098 63186 352334
rect 63422 352098 99186 352334
rect 99422 352098 108000 352334
rect -6696 352076 108000 352098
rect 448000 352418 459186 352654
rect 459422 352418 495186 352654
rect 495422 352418 531186 352654
rect 531422 352418 567186 352654
rect 567422 352418 590202 352654
rect 590438 352418 590620 352654
rect 448000 352334 590620 352418
rect 448000 352098 459186 352334
rect 459422 352098 495186 352334
rect 495422 352098 531186 352334
rect 531422 352098 567186 352334
rect 567422 352098 590202 352334
rect 590438 352098 590620 352334
rect 448000 352076 590620 352098
rect -6696 352074 -6096 352076
rect 27004 352074 27604 352076
rect 63004 352074 63604 352076
rect 99004 352074 99604 352076
rect 459004 352074 459604 352076
rect 495004 352074 495604 352076
rect 531004 352074 531604 352076
rect 567004 352074 567604 352076
rect 590020 352074 590620 352076
rect -4816 349076 -4216 349078
rect 23404 349076 24004 349078
rect 59404 349076 60004 349078
rect 95404 349076 96004 349078
rect -4816 349054 108000 349076
rect -4816 348818 -4634 349054
rect -4398 348818 23586 349054
rect 23822 348818 59586 349054
rect 59822 348818 95586 349054
rect 95822 348818 108000 349054
rect -4816 348734 108000 348818
rect -4816 348498 -4634 348734
rect -4398 348498 23586 348734
rect 23822 348498 59586 348734
rect 59822 348498 95586 348734
rect 95822 348498 108000 348734
rect 455404 349076 456004 349078
rect 491404 349076 492004 349078
rect 527404 349076 528004 349078
rect 563404 349076 564004 349078
rect 588140 349076 588740 349078
rect 448000 349054 588740 349076
rect 448000 348818 455586 349054
rect 455822 348818 491586 349054
rect 491822 348818 527586 349054
rect 527822 348818 563586 349054
rect 563822 348818 588322 349054
rect 588558 348818 588740 349054
rect 448000 348734 588740 348818
rect -4816 348476 108000 348498
rect 448000 348498 455586 348734
rect 455822 348498 491586 348734
rect 491822 348498 527586 348734
rect 527822 348498 563586 348734
rect 563822 348498 588322 348734
rect 588558 348498 588740 348734
rect 448000 348476 588740 348498
rect -4816 348474 -4216 348476
rect 23404 348474 24004 348476
rect 59404 348474 60004 348476
rect 95404 348474 96004 348476
rect 455404 348474 456004 348476
rect 491404 348474 492004 348476
rect 527404 348474 528004 348476
rect 563404 348474 564004 348476
rect 588140 348474 588740 348476
rect -2936 345476 -2336 345478
rect 19804 345476 20404 345478
rect 55804 345476 56404 345478
rect 91804 345476 92404 345478
rect -2936 345454 108000 345476
rect -2936 345218 -2754 345454
rect -2518 345218 19986 345454
rect 20222 345218 55986 345454
rect 56222 345218 91986 345454
rect 92222 345218 108000 345454
rect -2936 345134 108000 345218
rect -2936 344898 -2754 345134
rect -2518 344898 19986 345134
rect 20222 344898 55986 345134
rect 56222 344898 91986 345134
rect 92222 344898 108000 345134
rect -2936 344876 108000 344898
rect -2936 344874 -2336 344876
rect 19804 344874 20404 344876
rect 55804 344874 56404 344876
rect 91804 344874 92404 344876
rect 451804 345476 452404 345478
rect 487804 345476 488404 345478
rect 523804 345476 524404 345478
rect 559804 345476 560404 345478
rect 586260 345476 586860 345478
rect 448000 345454 586860 345476
rect 448000 345218 451986 345454
rect 452222 345218 487986 345454
rect 488222 345218 523986 345454
rect 524222 345218 559986 345454
rect 560222 345218 586442 345454
rect 586678 345218 586860 345454
rect 448000 345134 586860 345218
rect 448000 344898 451986 345134
rect 452222 344898 487986 345134
rect 488222 344898 523986 345134
rect 524222 344898 559986 345134
rect 560222 344898 586442 345134
rect 586678 344898 586860 345134
rect 448000 344876 586860 344898
rect 451804 344874 452404 344876
rect 487804 344874 488404 344876
rect 523804 344874 524404 344876
rect 559804 344874 560404 344876
rect 586260 344874 586860 344876
rect -7636 338276 -7036 338278
rect 12604 338276 13204 338278
rect 48604 338276 49204 338278
rect 84604 338276 85204 338278
rect 480604 338276 481204 338278
rect 516604 338276 517204 338278
rect 552604 338276 553204 338278
rect 590960 338276 591560 338278
rect -8576 338254 108000 338276
rect -8576 338018 -7454 338254
rect -7218 338018 12786 338254
rect 13022 338018 48786 338254
rect 49022 338018 84786 338254
rect 85022 338018 108000 338254
rect -8576 337934 108000 338018
rect -8576 337698 -7454 337934
rect -7218 337698 12786 337934
rect 13022 337698 48786 337934
rect 49022 337698 84786 337934
rect 85022 337698 108000 337934
rect -8576 337676 108000 337698
rect 448000 338254 592500 338276
rect 448000 338018 480786 338254
rect 481022 338018 516786 338254
rect 517022 338018 552786 338254
rect 553022 338018 591142 338254
rect 591378 338018 592500 338254
rect 448000 337934 592500 338018
rect 448000 337698 480786 337934
rect 481022 337698 516786 337934
rect 517022 337698 552786 337934
rect 553022 337698 591142 337934
rect 591378 337698 592500 337934
rect 448000 337676 592500 337698
rect -7636 337674 -7036 337676
rect 12604 337674 13204 337676
rect 48604 337674 49204 337676
rect 84604 337674 85204 337676
rect 480604 337674 481204 337676
rect 516604 337674 517204 337676
rect 552604 337674 553204 337676
rect 590960 337674 591560 337676
rect -5756 334676 -5156 334678
rect 9004 334676 9604 334678
rect 45004 334676 45604 334678
rect 81004 334676 81604 334678
rect 477004 334676 477604 334678
rect 513004 334676 513604 334678
rect 549004 334676 549604 334678
rect 589080 334676 589680 334678
rect -6696 334654 108000 334676
rect -6696 334418 -5574 334654
rect -5338 334418 9186 334654
rect 9422 334418 45186 334654
rect 45422 334418 81186 334654
rect 81422 334418 108000 334654
rect -6696 334334 108000 334418
rect -6696 334098 -5574 334334
rect -5338 334098 9186 334334
rect 9422 334098 45186 334334
rect 45422 334098 81186 334334
rect 81422 334098 108000 334334
rect -6696 334076 108000 334098
rect 448000 334654 590620 334676
rect 448000 334418 477186 334654
rect 477422 334418 513186 334654
rect 513422 334418 549186 334654
rect 549422 334418 589262 334654
rect 589498 334418 590620 334654
rect 448000 334334 590620 334418
rect 448000 334098 477186 334334
rect 477422 334098 513186 334334
rect 513422 334098 549186 334334
rect 549422 334098 589262 334334
rect 589498 334098 590620 334334
rect 448000 334076 590620 334098
rect -5756 334074 -5156 334076
rect 9004 334074 9604 334076
rect 45004 334074 45604 334076
rect 81004 334074 81604 334076
rect 477004 334074 477604 334076
rect 513004 334074 513604 334076
rect 549004 334074 549604 334076
rect 589080 334074 589680 334076
rect -3876 331076 -3276 331078
rect 5404 331076 6004 331078
rect 41404 331076 42004 331078
rect 77404 331076 78004 331078
rect 473404 331076 474004 331078
rect 509404 331076 510004 331078
rect 545404 331076 546004 331078
rect 581404 331076 582004 331078
rect 587200 331076 587800 331078
rect -4816 331054 133883 331076
rect -4816 330818 -3694 331054
rect -3458 330818 5586 331054
rect 5822 330818 41586 331054
rect 41822 330818 77586 331054
rect 77822 330947 133883 331054
rect 77822 330933 132359 330947
rect 77822 330918 130950 330933
rect 77822 330904 129549 330918
rect 77822 330889 128140 330904
rect 77822 330875 126660 330889
rect 77822 330860 125251 330875
rect 77822 330846 123850 330860
rect 77822 330818 123455 330846
rect -4816 330734 123455 330818
rect -4816 330498 -3694 330734
rect -3458 330498 5586 330734
rect 5822 330498 41586 330734
rect 41822 330498 77586 330734
rect 77822 330610 123455 330734
rect 123691 330624 123850 330846
rect 124086 330624 124170 330860
rect 124406 330624 124544 330860
rect 124780 330624 124864 330860
rect 125100 330639 125251 330860
rect 125487 330639 125571 330875
rect 125807 330639 125945 330875
rect 126181 330639 126265 330875
rect 126501 330653 126660 330875
rect 126896 330653 126980 330889
rect 127216 330653 127354 330889
rect 127590 330653 127674 330889
rect 127910 330668 128140 330889
rect 128376 330668 128460 330904
rect 128696 330668 128834 330904
rect 129070 330668 129154 330904
rect 129390 330682 129549 330904
rect 129785 330682 129869 330918
rect 130105 330682 130243 330918
rect 130479 330682 130563 330918
rect 130799 330697 130950 330918
rect 131186 330697 131270 330933
rect 131506 330697 131644 330933
rect 131880 330697 131964 330933
rect 132200 330711 132359 330933
rect 132595 330711 132679 330947
rect 132915 330711 133053 330947
rect 133289 330711 133373 330947
rect 133609 330711 133883 330947
rect 132200 330697 133883 330711
rect 130799 330682 133883 330697
rect 129390 330668 133883 330682
rect 127910 330653 133883 330668
rect 126501 330639 133883 330653
rect 125100 330624 133883 330639
rect 123691 330610 133883 330624
rect 77822 330498 133883 330610
rect -4816 330476 133883 330498
rect 448000 331054 588740 331076
rect 448000 330818 473586 331054
rect 473822 330818 509586 331054
rect 509822 330818 545586 331054
rect 545822 330818 581586 331054
rect 581822 330818 587382 331054
rect 587618 330818 588740 331054
rect 448000 330734 588740 330818
rect 448000 330498 473586 330734
rect 473822 330498 509586 330734
rect 509822 330498 545586 330734
rect 545822 330498 581586 330734
rect 581822 330498 587382 330734
rect 587618 330498 588740 330734
rect 448000 330476 588740 330498
rect -3876 330474 -3276 330476
rect 5404 330474 6004 330476
rect 41404 330474 42004 330476
rect 77404 330474 78004 330476
rect 473404 330474 474004 330476
rect 509404 330474 510004 330476
rect 545404 330474 546004 330476
rect 581404 330474 582004 330476
rect 587200 330474 587800 330476
rect -1996 327476 -1396 327478
rect 1804 327476 2404 327478
rect 37804 327476 38404 327478
rect 73804 327476 74404 327478
rect 469804 327476 470404 327478
rect 505804 327476 506404 327478
rect 541804 327476 542404 327478
rect 577804 327476 578404 327478
rect 585320 327476 585920 327478
rect -2936 327454 151560 327476
rect -2936 327218 -1814 327454
rect -1578 327218 1986 327454
rect 2222 327218 37986 327454
rect 38222 327218 73986 327454
rect 74222 327368 151560 327454
rect 74222 327354 150048 327368
rect 74222 327339 148639 327354
rect 74222 327325 147238 327339
rect 74222 327310 145829 327325
rect 74222 327296 144349 327310
rect 74222 327281 142940 327296
rect 74222 327267 141539 327281
rect 74222 327218 141144 327267
rect -2936 327134 141144 327218
rect -2936 326898 -1814 327134
rect -1578 326898 1986 327134
rect 2222 326898 37986 327134
rect 38222 326898 73986 327134
rect 74222 327031 141144 327134
rect 141380 327045 141539 327267
rect 141775 327045 141859 327281
rect 142095 327045 142233 327281
rect 142469 327045 142553 327281
rect 142789 327060 142940 327281
rect 143176 327060 143260 327296
rect 143496 327060 143634 327296
rect 143870 327060 143954 327296
rect 144190 327074 144349 327296
rect 144585 327074 144669 327310
rect 144905 327074 145043 327310
rect 145279 327074 145363 327310
rect 145599 327089 145829 327310
rect 146065 327089 146149 327325
rect 146385 327089 146523 327325
rect 146759 327089 146843 327325
rect 147079 327103 147238 327325
rect 147474 327103 147558 327339
rect 147794 327103 147932 327339
rect 148168 327103 148252 327339
rect 148488 327118 148639 327339
rect 148875 327118 148959 327354
rect 149195 327118 149333 327354
rect 149569 327118 149653 327354
rect 149889 327132 150048 327354
rect 150284 327132 150368 327368
rect 150604 327132 150742 327368
rect 150978 327132 151062 327368
rect 151298 327132 151560 327368
rect 149889 327118 151560 327132
rect 148488 327103 151560 327118
rect 147079 327089 151560 327103
rect 145599 327074 151560 327089
rect 144190 327060 151560 327074
rect 142789 327045 151560 327060
rect 141380 327031 151560 327045
rect 74222 326898 151560 327031
rect -2936 326876 151560 326898
rect 448000 327454 586860 327476
rect 448000 327218 469986 327454
rect 470222 327218 505986 327454
rect 506222 327218 541986 327454
rect 542222 327218 577986 327454
rect 578222 327218 585502 327454
rect 585738 327218 586860 327454
rect 448000 327134 586860 327218
rect 448000 326898 469986 327134
rect 470222 326898 505986 327134
rect 506222 326898 541986 327134
rect 542222 326898 577986 327134
rect 578222 326898 585502 327134
rect 585738 326898 586860 327134
rect 448000 326876 586860 326898
rect -1996 326874 -1396 326876
rect 1804 326874 2404 326876
rect 37804 326874 38404 326876
rect 73804 326874 74404 326876
rect 469804 326874 470404 326876
rect 505804 326874 506404 326876
rect 541804 326874 542404 326876
rect 577804 326874 578404 326876
rect 585320 326874 585920 326876
rect -8576 320276 -7976 320278
rect 30604 320276 31204 320278
rect 66604 320276 67204 320278
rect 102604 320276 103204 320278
rect 462604 320276 463204 320278
rect 498604 320276 499204 320278
rect 534604 320276 535204 320278
rect 570604 320276 571204 320278
rect 591900 320276 592500 320278
rect -8576 320254 108000 320276
rect -8576 320018 -8394 320254
rect -8158 320018 30786 320254
rect 31022 320018 66786 320254
rect 67022 320018 102786 320254
rect 103022 320018 108000 320254
rect -8576 319934 108000 320018
rect -8576 319698 -8394 319934
rect -8158 319698 30786 319934
rect 31022 319698 66786 319934
rect 67022 319698 102786 319934
rect 103022 319698 108000 319934
rect -8576 319676 108000 319698
rect 448000 320254 592500 320276
rect 448000 320018 462786 320254
rect 463022 320018 498786 320254
rect 499022 320018 534786 320254
rect 535022 320018 570786 320254
rect 571022 320018 592082 320254
rect 592318 320018 592500 320254
rect 448000 319934 592500 320018
rect 448000 319698 462786 319934
rect 463022 319698 498786 319934
rect 499022 319698 534786 319934
rect 535022 319698 570786 319934
rect 571022 319698 592082 319934
rect 592318 319698 592500 319934
rect 448000 319676 592500 319698
rect -8576 319674 -7976 319676
rect 30604 319674 31204 319676
rect 66604 319674 67204 319676
rect 102604 319674 103204 319676
rect 462604 319674 463204 319676
rect 498604 319674 499204 319676
rect 534604 319674 535204 319676
rect 570604 319674 571204 319676
rect 591900 319674 592500 319676
rect -6696 316676 -6096 316678
rect 27004 316676 27604 316678
rect 63004 316676 63604 316678
rect 99004 316676 99604 316678
rect 459004 316676 459604 316678
rect 495004 316676 495604 316678
rect 531004 316676 531604 316678
rect 567004 316676 567604 316678
rect 590020 316676 590620 316678
rect -6696 316654 108000 316676
rect -6696 316418 -6514 316654
rect -6278 316418 27186 316654
rect 27422 316418 63186 316654
rect 63422 316418 99186 316654
rect 99422 316418 108000 316654
rect -6696 316334 108000 316418
rect -6696 316098 -6514 316334
rect -6278 316098 27186 316334
rect 27422 316098 63186 316334
rect 63422 316098 99186 316334
rect 99422 316098 108000 316334
rect -6696 316076 108000 316098
rect 448000 316654 590620 316676
rect 448000 316418 459186 316654
rect 459422 316418 495186 316654
rect 495422 316418 531186 316654
rect 531422 316418 567186 316654
rect 567422 316418 590202 316654
rect 590438 316418 590620 316654
rect 448000 316334 590620 316418
rect 448000 316098 459186 316334
rect 459422 316098 495186 316334
rect 495422 316098 531186 316334
rect 531422 316098 567186 316334
rect 567422 316098 590202 316334
rect 590438 316098 590620 316334
rect 448000 316076 590620 316098
rect -6696 316074 -6096 316076
rect 27004 316074 27604 316076
rect 63004 316074 63604 316076
rect 99004 316074 99604 316076
rect 459004 316074 459604 316076
rect 495004 316074 495604 316076
rect 531004 316074 531604 316076
rect 567004 316074 567604 316076
rect 590020 316074 590620 316076
rect -4816 313076 -4216 313078
rect 23404 313076 24004 313078
rect 59404 313076 60004 313078
rect 95404 313076 96004 313078
rect 455404 313076 456004 313078
rect 491404 313076 492004 313078
rect 527404 313076 528004 313078
rect 563404 313076 564004 313078
rect 588140 313076 588740 313078
rect -4816 313054 108000 313076
rect -4816 312818 -4634 313054
rect -4398 312818 23586 313054
rect 23822 312818 59586 313054
rect 59822 312818 95586 313054
rect 95822 312818 108000 313054
rect -4816 312734 108000 312818
rect -4816 312498 -4634 312734
rect -4398 312498 23586 312734
rect 23822 312498 59586 312734
rect 59822 312498 95586 312734
rect 95822 312498 108000 312734
rect -4816 312476 108000 312498
rect 407589 313054 588740 313076
rect 407589 312960 455586 313054
rect 407589 312946 416821 312960
rect 407589 312931 415412 312946
rect 407589 312917 414011 312931
rect 407589 312902 412602 312917
rect 407589 312888 411122 312902
rect 407589 312873 409713 312888
rect 407589 312859 408312 312873
rect 407589 312623 407917 312859
rect 408153 312637 408312 312859
rect 408548 312637 408632 312873
rect 408868 312637 409006 312873
rect 409242 312637 409326 312873
rect 409562 312652 409713 312873
rect 409949 312652 410033 312888
rect 410269 312652 410407 312888
rect 410643 312652 410727 312888
rect 410963 312666 411122 312888
rect 411358 312666 411442 312902
rect 411678 312666 411816 312902
rect 412052 312666 412136 312902
rect 412372 312681 412602 312902
rect 412838 312681 412922 312917
rect 413158 312681 413296 312917
rect 413532 312681 413616 312917
rect 413852 312695 414011 312917
rect 414247 312695 414331 312931
rect 414567 312695 414705 312931
rect 414941 312695 415025 312931
rect 415261 312710 415412 312931
rect 415648 312710 415732 312946
rect 415968 312710 416106 312946
rect 416342 312710 416426 312946
rect 416662 312724 416821 312946
rect 417057 312724 417141 312960
rect 417377 312724 417515 312960
rect 417751 312724 417835 312960
rect 418071 312818 455586 312960
rect 455822 312818 491586 313054
rect 491822 312818 527586 313054
rect 527822 312818 563586 313054
rect 563822 312818 588322 313054
rect 588558 312818 588740 313054
rect 418071 312734 588740 312818
rect 418071 312724 455586 312734
rect 416662 312710 455586 312724
rect 415261 312695 455586 312710
rect 413852 312681 455586 312695
rect 412372 312666 455586 312681
rect 410963 312652 455586 312666
rect 409562 312637 455586 312652
rect 408153 312623 455586 312637
rect 407589 312498 455586 312623
rect 455822 312498 491586 312734
rect 491822 312498 527586 312734
rect 527822 312498 563586 312734
rect 563822 312498 588322 312734
rect 588558 312498 588740 312734
rect 407589 312476 588740 312498
rect -4816 312474 -4216 312476
rect 23404 312474 24004 312476
rect 59404 312474 60004 312476
rect 95404 312474 96004 312476
rect 455404 312474 456004 312476
rect 491404 312474 492004 312476
rect 527404 312474 528004 312476
rect 563404 312474 564004 312476
rect 588140 312474 588740 312476
rect -2936 309476 -2336 309478
rect 19804 309476 20404 309478
rect 55804 309476 56404 309478
rect 91804 309476 92404 309478
rect 451804 309476 452404 309478
rect 487804 309476 488404 309478
rect 523804 309476 524404 309478
rect 559804 309476 560404 309478
rect 586260 309476 586860 309478
rect -2936 309454 108000 309476
rect -2936 309218 -2754 309454
rect -2518 309218 19986 309454
rect 20222 309218 55986 309454
rect 56222 309218 91986 309454
rect 92222 309218 108000 309454
rect -2936 309134 108000 309218
rect -2936 308898 -2754 309134
rect -2518 308898 19986 309134
rect 20222 308898 55986 309134
rect 56222 308898 91986 309134
rect 92222 308898 108000 309134
rect -2936 308876 108000 308898
rect 425267 309454 586860 309476
rect 425267 309371 451986 309454
rect 425267 309357 434539 309371
rect 425267 309342 433130 309357
rect 425267 309328 431729 309342
rect 425267 309313 430320 309328
rect 425267 309299 428840 309313
rect 425267 309284 427431 309299
rect 425267 309270 426030 309284
rect 425267 309034 425635 309270
rect 425871 309048 426030 309270
rect 426266 309048 426350 309284
rect 426586 309048 426724 309284
rect 426960 309048 427044 309284
rect 427280 309063 427431 309284
rect 427667 309063 427751 309299
rect 427987 309063 428125 309299
rect 428361 309063 428445 309299
rect 428681 309077 428840 309299
rect 429076 309077 429160 309313
rect 429396 309077 429534 309313
rect 429770 309077 429854 309313
rect 430090 309092 430320 309313
rect 430556 309092 430640 309328
rect 430876 309092 431014 309328
rect 431250 309092 431334 309328
rect 431570 309106 431729 309328
rect 431965 309106 432049 309342
rect 432285 309106 432423 309342
rect 432659 309106 432743 309342
rect 432979 309121 433130 309342
rect 433366 309121 433450 309357
rect 433686 309121 433824 309357
rect 434060 309121 434144 309357
rect 434380 309135 434539 309357
rect 434775 309135 434859 309371
rect 435095 309135 435233 309371
rect 435469 309135 435553 309371
rect 435789 309218 451986 309371
rect 452222 309218 487986 309454
rect 488222 309218 523986 309454
rect 524222 309218 559986 309454
rect 560222 309218 586442 309454
rect 586678 309218 586860 309454
rect 435789 309135 586860 309218
rect 434380 309134 586860 309135
rect 434380 309121 451986 309134
rect 432979 309106 451986 309121
rect 431570 309092 451986 309106
rect 430090 309077 451986 309092
rect 428681 309063 451986 309077
rect 427280 309048 451986 309063
rect 425871 309034 451986 309048
rect 425267 308898 451986 309034
rect 452222 308898 487986 309134
rect 488222 308898 523986 309134
rect 524222 308898 559986 309134
rect 560222 308898 586442 309134
rect 586678 308898 586860 309134
rect 425267 308876 586860 308898
rect -2936 308874 -2336 308876
rect 19804 308874 20404 308876
rect 55804 308874 56404 308876
rect 91804 308874 92404 308876
rect 451804 308874 452404 308876
rect 487804 308874 488404 308876
rect 523804 308874 524404 308876
rect 559804 308874 560404 308876
rect 586260 308874 586860 308876
rect -7636 302276 -7036 302278
rect 12604 302276 13204 302278
rect 48604 302276 49204 302278
rect 84604 302276 85204 302278
rect 480604 302276 481204 302278
rect 516604 302276 517204 302278
rect 552604 302276 553204 302278
rect 590960 302276 591560 302278
rect -8576 302254 108000 302276
rect -8576 302018 -7454 302254
rect -7218 302018 12786 302254
rect 13022 302018 48786 302254
rect 49022 302018 84786 302254
rect 85022 302018 108000 302254
rect -8576 301934 108000 302018
rect -8576 301698 -7454 301934
rect -7218 301698 12786 301934
rect 13022 301698 48786 301934
rect 49022 301698 84786 301934
rect 85022 301698 108000 301934
rect -8576 301676 108000 301698
rect 448000 302254 592500 302276
rect 448000 302018 480786 302254
rect 481022 302018 516786 302254
rect 517022 302018 552786 302254
rect 553022 302018 591142 302254
rect 591378 302018 592500 302254
rect 448000 301934 592500 302018
rect 448000 301698 480786 301934
rect 481022 301698 516786 301934
rect 517022 301698 552786 301934
rect 553022 301698 591142 301934
rect 591378 301698 592500 301934
rect 448000 301676 592500 301698
rect -7636 301674 -7036 301676
rect 12604 301674 13204 301676
rect 48604 301674 49204 301676
rect 84604 301674 85204 301676
rect 480604 301674 481204 301676
rect 516604 301674 517204 301676
rect 552604 301674 553204 301676
rect 590960 301674 591560 301676
rect -5756 298676 -5156 298678
rect 9004 298676 9604 298678
rect 45004 298676 45604 298678
rect 81004 298676 81604 298678
rect 477004 298676 477604 298678
rect 513004 298676 513604 298678
rect 549004 298676 549604 298678
rect 589080 298676 589680 298678
rect -6696 298654 108000 298676
rect -6696 298418 -5574 298654
rect -5338 298418 9186 298654
rect 9422 298418 45186 298654
rect 45422 298418 81186 298654
rect 81422 298418 108000 298654
rect -6696 298334 108000 298418
rect -6696 298098 -5574 298334
rect -5338 298098 9186 298334
rect 9422 298098 45186 298334
rect 45422 298098 81186 298334
rect 81422 298098 108000 298334
rect -6696 298076 108000 298098
rect 448000 298654 590620 298676
rect 448000 298418 477186 298654
rect 477422 298418 513186 298654
rect 513422 298418 549186 298654
rect 549422 298418 589262 298654
rect 589498 298418 590620 298654
rect 448000 298334 590620 298418
rect 448000 298098 477186 298334
rect 477422 298098 513186 298334
rect 513422 298098 549186 298334
rect 549422 298098 589262 298334
rect 589498 298098 590620 298334
rect 448000 298076 590620 298098
rect -5756 298074 -5156 298076
rect 9004 298074 9604 298076
rect 45004 298074 45604 298076
rect 81004 298074 81604 298076
rect 477004 298074 477604 298076
rect 513004 298074 513604 298076
rect 549004 298074 549604 298076
rect 589080 298074 589680 298076
rect -3876 295076 -3276 295078
rect 5404 295076 6004 295078
rect 41404 295076 42004 295078
rect 77404 295076 78004 295078
rect 473404 295076 474004 295078
rect 509404 295076 510004 295078
rect 545404 295076 546004 295078
rect 581404 295076 582004 295078
rect 587200 295076 587800 295078
rect -4816 295054 133883 295076
rect -4816 294818 -3694 295054
rect -3458 294818 5586 295054
rect 5822 294818 41586 295054
rect 41822 294818 77586 295054
rect 77822 294944 133883 295054
rect 77822 294930 132376 294944
rect 77822 294915 130967 294930
rect 77822 294901 129566 294915
rect 77822 294886 128157 294901
rect 77822 294872 126677 294886
rect 77822 294857 125268 294872
rect 77822 294843 123867 294857
rect 77822 294818 123472 294843
rect -4816 294734 123472 294818
rect -4816 294498 -3694 294734
rect -3458 294498 5586 294734
rect 5822 294498 41586 294734
rect 41822 294498 77586 294734
rect 77822 294607 123472 294734
rect 123708 294621 123867 294843
rect 124103 294621 124187 294857
rect 124423 294621 124561 294857
rect 124797 294621 124881 294857
rect 125117 294636 125268 294857
rect 125504 294636 125588 294872
rect 125824 294636 125962 294872
rect 126198 294636 126282 294872
rect 126518 294650 126677 294872
rect 126913 294650 126997 294886
rect 127233 294650 127371 294886
rect 127607 294650 127691 294886
rect 127927 294665 128157 294886
rect 128393 294665 128477 294901
rect 128713 294665 128851 294901
rect 129087 294665 129171 294901
rect 129407 294679 129566 294901
rect 129802 294679 129886 294915
rect 130122 294679 130260 294915
rect 130496 294679 130580 294915
rect 130816 294694 130967 294915
rect 131203 294694 131287 294930
rect 131523 294694 131661 294930
rect 131897 294694 131981 294930
rect 132217 294708 132376 294930
rect 132612 294708 132696 294944
rect 132932 294708 133070 294944
rect 133306 294708 133390 294944
rect 133626 294708 133883 294944
rect 132217 294694 133883 294708
rect 130816 294679 133883 294694
rect 129407 294665 133883 294679
rect 127927 294650 133883 294665
rect 126518 294636 133883 294650
rect 125117 294621 133883 294636
rect 123708 294607 133883 294621
rect 77822 294498 133883 294607
rect -4816 294476 133883 294498
rect 448000 295054 588740 295076
rect 448000 294818 473586 295054
rect 473822 294818 509586 295054
rect 509822 294818 545586 295054
rect 545822 294818 581586 295054
rect 581822 294818 587382 295054
rect 587618 294818 588740 295054
rect 448000 294734 588740 294818
rect 448000 294498 473586 294734
rect 473822 294498 509586 294734
rect 509822 294498 545586 294734
rect 545822 294498 581586 294734
rect 581822 294498 587382 294734
rect 587618 294498 588740 294734
rect 448000 294476 588740 294498
rect -3876 294474 -3276 294476
rect 5404 294474 6004 294476
rect 41404 294474 42004 294476
rect 77404 294474 78004 294476
rect 473404 294474 474004 294476
rect 509404 294474 510004 294476
rect 545404 294474 546004 294476
rect 581404 294474 582004 294476
rect 587200 294474 587800 294476
rect -1996 291476 -1396 291478
rect 1804 291476 2404 291478
rect 37804 291476 38404 291478
rect 73804 291476 74404 291478
rect 469804 291476 470404 291478
rect 505804 291476 506404 291478
rect 541804 291476 542404 291478
rect 577804 291476 578404 291478
rect 585320 291476 585920 291478
rect -2936 291454 151560 291476
rect -2936 291218 -1814 291454
rect -1578 291218 1986 291454
rect 2222 291218 37986 291454
rect 38222 291218 73986 291454
rect 74222 291335 151560 291454
rect 74222 291321 149921 291335
rect 74222 291306 148512 291321
rect 74222 291292 147111 291306
rect 74222 291277 145702 291292
rect 74222 291263 144222 291277
rect 74222 291248 142813 291263
rect 74222 291234 141412 291248
rect 74222 291218 141017 291234
rect -2936 291134 141017 291218
rect -2936 290898 -1814 291134
rect -1578 290898 1986 291134
rect 2222 290898 37986 291134
rect 38222 290898 73986 291134
rect 74222 290998 141017 291134
rect 141253 291012 141412 291234
rect 141648 291012 141732 291248
rect 141968 291012 142106 291248
rect 142342 291012 142426 291248
rect 142662 291027 142813 291248
rect 143049 291027 143133 291263
rect 143369 291027 143507 291263
rect 143743 291027 143827 291263
rect 144063 291041 144222 291263
rect 144458 291041 144542 291277
rect 144778 291041 144916 291277
rect 145152 291041 145236 291277
rect 145472 291056 145702 291277
rect 145938 291056 146022 291292
rect 146258 291056 146396 291292
rect 146632 291056 146716 291292
rect 146952 291070 147111 291292
rect 147347 291070 147431 291306
rect 147667 291070 147805 291306
rect 148041 291070 148125 291306
rect 148361 291085 148512 291306
rect 148748 291085 148832 291321
rect 149068 291085 149206 291321
rect 149442 291085 149526 291321
rect 149762 291099 149921 291321
rect 150157 291099 150241 291335
rect 150477 291099 150615 291335
rect 150851 291099 150935 291335
rect 151171 291099 151560 291335
rect 149762 291085 151560 291099
rect 148361 291070 151560 291085
rect 146952 291056 151560 291070
rect 145472 291041 151560 291056
rect 144063 291027 151560 291041
rect 142662 291012 151560 291027
rect 141253 290998 151560 291012
rect 74222 290898 151560 290998
rect -2936 290876 151560 290898
rect 448000 291454 586860 291476
rect 448000 291218 469986 291454
rect 470222 291218 505986 291454
rect 506222 291218 541986 291454
rect 542222 291218 577986 291454
rect 578222 291218 585502 291454
rect 585738 291218 586860 291454
rect 448000 291134 586860 291218
rect 448000 290898 469986 291134
rect 470222 290898 505986 291134
rect 506222 290898 541986 291134
rect 542222 290898 577986 291134
rect 578222 290898 585502 291134
rect 585738 290898 586860 291134
rect 448000 290876 586860 290898
rect -1996 290874 -1396 290876
rect 1804 290874 2404 290876
rect 37804 290874 38404 290876
rect 73804 290874 74404 290876
rect 469804 290874 470404 290876
rect 505804 290874 506404 290876
rect 541804 290874 542404 290876
rect 577804 290874 578404 290876
rect 585320 290874 585920 290876
rect -8576 284276 -7976 284278
rect 30604 284276 31204 284278
rect 66604 284276 67204 284278
rect 102604 284276 103204 284278
rect 462604 284276 463204 284278
rect 498604 284276 499204 284278
rect 534604 284276 535204 284278
rect 570604 284276 571204 284278
rect 591900 284276 592500 284278
rect -8576 284254 108000 284276
rect -8576 284018 -8394 284254
rect -8158 284018 30786 284254
rect 31022 284018 66786 284254
rect 67022 284018 102786 284254
rect 103022 284018 108000 284254
rect -8576 283934 108000 284018
rect -8576 283698 -8394 283934
rect -8158 283698 30786 283934
rect 31022 283698 66786 283934
rect 67022 283698 102786 283934
rect 103022 283698 108000 283934
rect -8576 283676 108000 283698
rect 448000 284254 592500 284276
rect 448000 284018 462786 284254
rect 463022 284018 498786 284254
rect 499022 284018 534786 284254
rect 535022 284018 570786 284254
rect 571022 284018 592082 284254
rect 592318 284018 592500 284254
rect 448000 283934 592500 284018
rect 448000 283698 462786 283934
rect 463022 283698 498786 283934
rect 499022 283698 534786 283934
rect 535022 283698 570786 283934
rect 571022 283698 592082 283934
rect 592318 283698 592500 283934
rect 448000 283676 592500 283698
rect -8576 283674 -7976 283676
rect 30604 283674 31204 283676
rect 66604 283674 67204 283676
rect 102604 283674 103204 283676
rect 462604 283674 463204 283676
rect 498604 283674 499204 283676
rect 534604 283674 535204 283676
rect 570604 283674 571204 283676
rect 591900 283674 592500 283676
rect -6696 280676 -6096 280678
rect 27004 280676 27604 280678
rect 63004 280676 63604 280678
rect 99004 280676 99604 280678
rect 459004 280676 459604 280678
rect 495004 280676 495604 280678
rect 531004 280676 531604 280678
rect 567004 280676 567604 280678
rect 590020 280676 590620 280678
rect -6696 280654 108000 280676
rect -6696 280418 -6514 280654
rect -6278 280418 27186 280654
rect 27422 280418 63186 280654
rect 63422 280418 99186 280654
rect 99422 280418 108000 280654
rect -6696 280334 108000 280418
rect -6696 280098 -6514 280334
rect -6278 280098 27186 280334
rect 27422 280098 63186 280334
rect 63422 280098 99186 280334
rect 99422 280098 108000 280334
rect -6696 280076 108000 280098
rect 448000 280654 590620 280676
rect 448000 280418 459186 280654
rect 459422 280418 495186 280654
rect 495422 280418 531186 280654
rect 531422 280418 567186 280654
rect 567422 280418 590202 280654
rect 590438 280418 590620 280654
rect 448000 280334 590620 280418
rect 448000 280098 459186 280334
rect 459422 280098 495186 280334
rect 495422 280098 531186 280334
rect 531422 280098 567186 280334
rect 567422 280098 590202 280334
rect 590438 280098 590620 280334
rect 448000 280076 590620 280098
rect -6696 280074 -6096 280076
rect 27004 280074 27604 280076
rect 63004 280074 63604 280076
rect 99004 280074 99604 280076
rect 459004 280074 459604 280076
rect 495004 280074 495604 280076
rect 531004 280074 531604 280076
rect 567004 280074 567604 280076
rect 590020 280074 590620 280076
rect -4816 277076 -4216 277078
rect 23404 277076 24004 277078
rect 59404 277076 60004 277078
rect 95404 277076 96004 277078
rect 455404 277076 456004 277078
rect 491404 277076 492004 277078
rect 527404 277076 528004 277078
rect 563404 277076 564004 277078
rect 588140 277076 588740 277078
rect -4816 277054 108000 277076
rect -4816 276818 -4634 277054
rect -4398 276818 23586 277054
rect 23822 276818 59586 277054
rect 59822 276818 95586 277054
rect 95822 276818 108000 277054
rect -4816 276734 108000 276818
rect -4816 276498 -4634 276734
rect -4398 276498 23586 276734
rect 23822 276498 59586 276734
rect 59822 276498 95586 276734
rect 95822 276498 108000 276734
rect -4816 276476 108000 276498
rect 407589 277054 588740 277076
rect 407589 276941 455586 277054
rect 407589 276927 416796 276941
rect 407589 276912 415387 276927
rect 407589 276898 413986 276912
rect 407589 276883 412577 276898
rect 407589 276869 411097 276883
rect 407589 276854 409688 276869
rect 407589 276840 408287 276854
rect 407589 276604 407892 276840
rect 408128 276618 408287 276840
rect 408523 276618 408607 276854
rect 408843 276618 408981 276854
rect 409217 276618 409301 276854
rect 409537 276633 409688 276854
rect 409924 276633 410008 276869
rect 410244 276633 410382 276869
rect 410618 276633 410702 276869
rect 410938 276647 411097 276869
rect 411333 276647 411417 276883
rect 411653 276647 411791 276883
rect 412027 276647 412111 276883
rect 412347 276662 412577 276883
rect 412813 276662 412897 276898
rect 413133 276662 413271 276898
rect 413507 276662 413591 276898
rect 413827 276676 413986 276898
rect 414222 276676 414306 276912
rect 414542 276676 414680 276912
rect 414916 276676 415000 276912
rect 415236 276691 415387 276912
rect 415623 276691 415707 276927
rect 415943 276691 416081 276927
rect 416317 276691 416401 276927
rect 416637 276705 416796 276927
rect 417032 276705 417116 276941
rect 417352 276705 417490 276941
rect 417726 276705 417810 276941
rect 418046 276818 455586 276941
rect 455822 276818 491586 277054
rect 491822 276818 527586 277054
rect 527822 276818 563586 277054
rect 563822 276818 588322 277054
rect 588558 276818 588740 277054
rect 418046 276734 588740 276818
rect 418046 276705 455586 276734
rect 416637 276691 455586 276705
rect 415236 276676 455586 276691
rect 413827 276662 455586 276676
rect 412347 276647 455586 276662
rect 410938 276633 455586 276647
rect 409537 276618 455586 276633
rect 408128 276604 455586 276618
rect 407589 276498 455586 276604
rect 455822 276498 491586 276734
rect 491822 276498 527586 276734
rect 527822 276498 563586 276734
rect 563822 276498 588322 276734
rect 588558 276498 588740 276734
rect 407589 276476 588740 276498
rect -4816 276474 -4216 276476
rect 23404 276474 24004 276476
rect 59404 276474 60004 276476
rect 95404 276474 96004 276476
rect 455404 276474 456004 276476
rect 491404 276474 492004 276476
rect 527404 276474 528004 276476
rect 563404 276474 564004 276476
rect 588140 276474 588740 276476
rect -2936 273476 -2336 273478
rect 19804 273476 20404 273478
rect 55804 273476 56404 273478
rect 91804 273476 92404 273478
rect 451804 273476 452404 273478
rect 487804 273476 488404 273478
rect 523804 273476 524404 273478
rect 559804 273476 560404 273478
rect 586260 273476 586860 273478
rect -2936 273454 108000 273476
rect -2936 273218 -2754 273454
rect -2518 273218 19986 273454
rect 20222 273218 55986 273454
rect 56222 273218 91986 273454
rect 92222 273218 108000 273454
rect -2936 273134 108000 273218
rect -2936 272898 -2754 273134
rect -2518 272898 19986 273134
rect 20222 272898 55986 273134
rect 56222 272898 91986 273134
rect 92222 272898 108000 273134
rect -2936 272876 108000 272898
rect 425267 273454 586860 273476
rect 425267 273350 451986 273454
rect 425267 273336 434590 273350
rect 425267 273321 433181 273336
rect 425267 273307 431780 273321
rect 425267 273292 430371 273307
rect 425267 273278 428891 273292
rect 425267 273263 427482 273278
rect 425267 273249 426081 273263
rect 425267 273013 425686 273249
rect 425922 273027 426081 273249
rect 426317 273027 426401 273263
rect 426637 273027 426775 273263
rect 427011 273027 427095 273263
rect 427331 273042 427482 273263
rect 427718 273042 427802 273278
rect 428038 273042 428176 273278
rect 428412 273042 428496 273278
rect 428732 273056 428891 273278
rect 429127 273056 429211 273292
rect 429447 273056 429585 273292
rect 429821 273056 429905 273292
rect 430141 273071 430371 273292
rect 430607 273071 430691 273307
rect 430927 273071 431065 273307
rect 431301 273071 431385 273307
rect 431621 273085 431780 273307
rect 432016 273085 432100 273321
rect 432336 273085 432474 273321
rect 432710 273085 432794 273321
rect 433030 273100 433181 273321
rect 433417 273100 433501 273336
rect 433737 273100 433875 273336
rect 434111 273100 434195 273336
rect 434431 273114 434590 273336
rect 434826 273114 434910 273350
rect 435146 273114 435284 273350
rect 435520 273114 435604 273350
rect 435840 273218 451986 273350
rect 452222 273218 487986 273454
rect 488222 273218 523986 273454
rect 524222 273218 559986 273454
rect 560222 273218 586442 273454
rect 586678 273218 586860 273454
rect 435840 273134 586860 273218
rect 435840 273114 451986 273134
rect 434431 273100 451986 273114
rect 433030 273085 451986 273100
rect 431621 273071 451986 273085
rect 430141 273056 451986 273071
rect 428732 273042 451986 273056
rect 427331 273027 451986 273042
rect 425922 273013 451986 273027
rect 425267 272898 451986 273013
rect 452222 272898 487986 273134
rect 488222 272898 523986 273134
rect 524222 272898 559986 273134
rect 560222 272898 586442 273134
rect 586678 272898 586860 273134
rect 425267 272876 586860 272898
rect -2936 272874 -2336 272876
rect 19804 272874 20404 272876
rect 55804 272874 56404 272876
rect 91804 272874 92404 272876
rect 451804 272874 452404 272876
rect 487804 272874 488404 272876
rect 523804 272874 524404 272876
rect 559804 272874 560404 272876
rect 586260 272874 586860 272876
rect -7636 266276 -7036 266278
rect 12604 266276 13204 266278
rect 48604 266276 49204 266278
rect 84604 266276 85204 266278
rect 480604 266276 481204 266278
rect 516604 266276 517204 266278
rect 552604 266276 553204 266278
rect 590960 266276 591560 266278
rect -8576 266254 108000 266276
rect -8576 266018 -7454 266254
rect -7218 266018 12786 266254
rect 13022 266018 48786 266254
rect 49022 266018 84786 266254
rect 85022 266018 108000 266254
rect -8576 265934 108000 266018
rect -8576 265698 -7454 265934
rect -7218 265698 12786 265934
rect 13022 265698 48786 265934
rect 49022 265698 84786 265934
rect 85022 265698 108000 265934
rect -8576 265676 108000 265698
rect 448000 266254 592500 266276
rect 448000 266018 480786 266254
rect 481022 266018 516786 266254
rect 517022 266018 552786 266254
rect 553022 266018 591142 266254
rect 591378 266018 592500 266254
rect 448000 265934 592500 266018
rect 448000 265698 480786 265934
rect 481022 265698 516786 265934
rect 517022 265698 552786 265934
rect 553022 265698 591142 265934
rect 591378 265698 592500 265934
rect 448000 265676 592500 265698
rect -7636 265674 -7036 265676
rect 12604 265674 13204 265676
rect 48604 265674 49204 265676
rect 84604 265674 85204 265676
rect 480604 265674 481204 265676
rect 516604 265674 517204 265676
rect 552604 265674 553204 265676
rect 590960 265674 591560 265676
rect -5756 262676 -5156 262678
rect 9004 262676 9604 262678
rect 45004 262676 45604 262678
rect 81004 262676 81604 262678
rect 477004 262676 477604 262678
rect 513004 262676 513604 262678
rect 549004 262676 549604 262678
rect 589080 262676 589680 262678
rect -6696 262654 108000 262676
rect -6696 262418 -5574 262654
rect -5338 262418 9186 262654
rect 9422 262418 45186 262654
rect 45422 262418 81186 262654
rect 81422 262418 108000 262654
rect -6696 262334 108000 262418
rect -6696 262098 -5574 262334
rect -5338 262098 9186 262334
rect 9422 262098 45186 262334
rect 45422 262098 81186 262334
rect 81422 262098 108000 262334
rect -6696 262076 108000 262098
rect 448000 262654 590620 262676
rect 448000 262418 477186 262654
rect 477422 262418 513186 262654
rect 513422 262418 549186 262654
rect 549422 262418 589262 262654
rect 589498 262418 590620 262654
rect 448000 262334 590620 262418
rect 448000 262098 477186 262334
rect 477422 262098 513186 262334
rect 513422 262098 549186 262334
rect 549422 262098 589262 262334
rect 589498 262098 590620 262334
rect 448000 262076 590620 262098
rect -5756 262074 -5156 262076
rect 9004 262074 9604 262076
rect 45004 262074 45604 262076
rect 81004 262074 81604 262076
rect 477004 262074 477604 262076
rect 513004 262074 513604 262076
rect 549004 262074 549604 262076
rect 589080 262074 589680 262076
rect -3876 259076 -3276 259078
rect 5404 259076 6004 259078
rect 41404 259076 42004 259078
rect 77404 259076 78004 259078
rect 473404 259076 474004 259078
rect 509404 259076 510004 259078
rect 545404 259076 546004 259078
rect 581404 259076 582004 259078
rect 587200 259076 587800 259078
rect -4816 259054 133883 259076
rect -4816 258818 -3694 259054
rect -3458 258818 5586 259054
rect 5822 258818 41586 259054
rect 41822 258818 77586 259054
rect 77822 258944 133883 259054
rect 77822 258930 132142 258944
rect 77822 258915 130733 258930
rect 77822 258901 129332 258915
rect 77822 258886 127923 258901
rect 77822 258872 126443 258886
rect 77822 258857 125034 258872
rect 77822 258843 123633 258857
rect 77822 258818 123238 258843
rect -4816 258734 123238 258818
rect -4816 258498 -3694 258734
rect -3458 258498 5586 258734
rect 5822 258498 41586 258734
rect 41822 258498 77586 258734
rect 77822 258607 123238 258734
rect 123474 258621 123633 258843
rect 123869 258621 123953 258857
rect 124189 258621 124327 258857
rect 124563 258621 124647 258857
rect 124883 258636 125034 258857
rect 125270 258636 125354 258872
rect 125590 258636 125728 258872
rect 125964 258636 126048 258872
rect 126284 258650 126443 258872
rect 126679 258650 126763 258886
rect 126999 258650 127137 258886
rect 127373 258650 127457 258886
rect 127693 258665 127923 258886
rect 128159 258665 128243 258901
rect 128479 258665 128617 258901
rect 128853 258665 128937 258901
rect 129173 258679 129332 258901
rect 129568 258679 129652 258915
rect 129888 258679 130026 258915
rect 130262 258679 130346 258915
rect 130582 258694 130733 258915
rect 130969 258694 131053 258930
rect 131289 258694 131427 258930
rect 131663 258694 131747 258930
rect 131983 258708 132142 258930
rect 132378 258708 132462 258944
rect 132698 258708 132836 258944
rect 133072 258708 133156 258944
rect 133392 258708 133883 258944
rect 131983 258694 133883 258708
rect 130582 258679 133883 258694
rect 129173 258665 133883 258679
rect 127693 258650 133883 258665
rect 126284 258636 133883 258650
rect 124883 258621 133883 258636
rect 123474 258607 133883 258621
rect 77822 258498 133883 258607
rect -4816 258476 133883 258498
rect 448000 259054 588740 259076
rect 448000 258818 473586 259054
rect 473822 258818 509586 259054
rect 509822 258818 545586 259054
rect 545822 258818 581586 259054
rect 581822 258818 587382 259054
rect 587618 258818 588740 259054
rect 448000 258734 588740 258818
rect 448000 258498 473586 258734
rect 473822 258498 509586 258734
rect 509822 258498 545586 258734
rect 545822 258498 581586 258734
rect 581822 258498 587382 258734
rect 587618 258498 588740 258734
rect 448000 258476 588740 258498
rect -3876 258474 -3276 258476
rect 5404 258474 6004 258476
rect 41404 258474 42004 258476
rect 77404 258474 78004 258476
rect 473404 258474 474004 258476
rect 509404 258474 510004 258476
rect 545404 258474 546004 258476
rect 581404 258474 582004 258476
rect 587200 258474 587800 258476
rect -1996 255476 -1396 255478
rect 1804 255476 2404 255478
rect 37804 255476 38404 255478
rect 73804 255476 74404 255478
rect 469804 255476 470404 255478
rect 505804 255476 506404 255478
rect 541804 255476 542404 255478
rect 577804 255476 578404 255478
rect 585320 255476 585920 255478
rect -2936 255454 151560 255476
rect -2936 255218 -1814 255454
rect -1578 255218 1986 255454
rect 2222 255218 37986 255454
rect 38222 255218 73986 255454
rect 74222 255325 151560 255454
rect 74222 255311 149949 255325
rect 74222 255296 148540 255311
rect 74222 255282 147139 255296
rect 74222 255267 145730 255282
rect 74222 255253 144250 255267
rect 74222 255238 142841 255253
rect 74222 255224 141440 255238
rect 74222 255218 141045 255224
rect -2936 255134 141045 255218
rect -2936 254898 -1814 255134
rect -1578 254898 1986 255134
rect 2222 254898 37986 255134
rect 38222 254898 73986 255134
rect 74222 254988 141045 255134
rect 141281 255002 141440 255224
rect 141676 255002 141760 255238
rect 141996 255002 142134 255238
rect 142370 255002 142454 255238
rect 142690 255017 142841 255238
rect 143077 255017 143161 255253
rect 143397 255017 143535 255253
rect 143771 255017 143855 255253
rect 144091 255031 144250 255253
rect 144486 255031 144570 255267
rect 144806 255031 144944 255267
rect 145180 255031 145264 255267
rect 145500 255046 145730 255267
rect 145966 255046 146050 255282
rect 146286 255046 146424 255282
rect 146660 255046 146744 255282
rect 146980 255060 147139 255282
rect 147375 255060 147459 255296
rect 147695 255060 147833 255296
rect 148069 255060 148153 255296
rect 148389 255075 148540 255296
rect 148776 255075 148860 255311
rect 149096 255075 149234 255311
rect 149470 255075 149554 255311
rect 149790 255089 149949 255311
rect 150185 255089 150269 255325
rect 150505 255089 150643 255325
rect 150879 255089 150963 255325
rect 151199 255089 151560 255325
rect 149790 255075 151560 255089
rect 148389 255060 151560 255075
rect 146980 255046 151560 255060
rect 145500 255031 151560 255046
rect 144091 255017 151560 255031
rect 142690 255002 151560 255017
rect 141281 254988 151560 255002
rect 74222 254898 151560 254988
rect -2936 254876 151560 254898
rect 448000 255454 586860 255476
rect 448000 255218 469986 255454
rect 470222 255218 505986 255454
rect 506222 255218 541986 255454
rect 542222 255218 577986 255454
rect 578222 255218 585502 255454
rect 585738 255218 586860 255454
rect 448000 255134 586860 255218
rect 448000 254898 469986 255134
rect 470222 254898 505986 255134
rect 506222 254898 541986 255134
rect 542222 254898 577986 255134
rect 578222 254898 585502 255134
rect 585738 254898 586860 255134
rect 448000 254876 586860 254898
rect -1996 254874 -1396 254876
rect 1804 254874 2404 254876
rect 37804 254874 38404 254876
rect 73804 254874 74404 254876
rect 469804 254874 470404 254876
rect 505804 254874 506404 254876
rect 541804 254874 542404 254876
rect 577804 254874 578404 254876
rect 585320 254874 585920 254876
rect -8576 248276 -7976 248278
rect 30604 248276 31204 248278
rect 66604 248276 67204 248278
rect 102604 248276 103204 248278
rect 462604 248276 463204 248278
rect 498604 248276 499204 248278
rect 534604 248276 535204 248278
rect 570604 248276 571204 248278
rect 591900 248276 592500 248278
rect -8576 248254 108000 248276
rect -8576 248018 -8394 248254
rect -8158 248018 30786 248254
rect 31022 248018 66786 248254
rect 67022 248018 102786 248254
rect 103022 248018 108000 248254
rect -8576 247934 108000 248018
rect -8576 247698 -8394 247934
rect -8158 247698 30786 247934
rect 31022 247698 66786 247934
rect 67022 247698 102786 247934
rect 103022 247698 108000 247934
rect -8576 247676 108000 247698
rect 448000 248254 592500 248276
rect 448000 248018 462786 248254
rect 463022 248018 498786 248254
rect 499022 248018 534786 248254
rect 535022 248018 570786 248254
rect 571022 248018 592082 248254
rect 592318 248018 592500 248254
rect 448000 247934 592500 248018
rect 448000 247698 462786 247934
rect 463022 247698 498786 247934
rect 499022 247698 534786 247934
rect 535022 247698 570786 247934
rect 571022 247698 592082 247934
rect 592318 247698 592500 247934
rect 448000 247676 592500 247698
rect -8576 247674 -7976 247676
rect 30604 247674 31204 247676
rect 66604 247674 67204 247676
rect 102604 247674 103204 247676
rect 462604 247674 463204 247676
rect 498604 247674 499204 247676
rect 534604 247674 535204 247676
rect 570604 247674 571204 247676
rect 591900 247674 592500 247676
rect -6696 244676 -6096 244678
rect 27004 244676 27604 244678
rect 63004 244676 63604 244678
rect 99004 244676 99604 244678
rect 459004 244676 459604 244678
rect 495004 244676 495604 244678
rect 531004 244676 531604 244678
rect 567004 244676 567604 244678
rect 590020 244676 590620 244678
rect -6696 244654 108000 244676
rect -6696 244418 -6514 244654
rect -6278 244418 27186 244654
rect 27422 244418 63186 244654
rect 63422 244418 99186 244654
rect 99422 244418 108000 244654
rect -6696 244334 108000 244418
rect -6696 244098 -6514 244334
rect -6278 244098 27186 244334
rect 27422 244098 63186 244334
rect 63422 244098 99186 244334
rect 99422 244098 108000 244334
rect -6696 244076 108000 244098
rect 448000 244654 590620 244676
rect 448000 244418 459186 244654
rect 459422 244418 495186 244654
rect 495422 244418 531186 244654
rect 531422 244418 567186 244654
rect 567422 244418 590202 244654
rect 590438 244418 590620 244654
rect 448000 244334 590620 244418
rect 448000 244098 459186 244334
rect 459422 244098 495186 244334
rect 495422 244098 531186 244334
rect 531422 244098 567186 244334
rect 567422 244098 590202 244334
rect 590438 244098 590620 244334
rect 448000 244076 590620 244098
rect -6696 244074 -6096 244076
rect 27004 244074 27604 244076
rect 63004 244074 63604 244076
rect 99004 244074 99604 244076
rect 459004 244074 459604 244076
rect 495004 244074 495604 244076
rect 531004 244074 531604 244076
rect 567004 244074 567604 244076
rect 590020 244074 590620 244076
rect -4816 241076 -4216 241078
rect 23404 241076 24004 241078
rect 59404 241076 60004 241078
rect 95404 241076 96004 241078
rect 455404 241076 456004 241078
rect 491404 241076 492004 241078
rect 527404 241076 528004 241078
rect 563404 241076 564004 241078
rect 588140 241076 588740 241078
rect -4816 241054 108000 241076
rect -4816 240818 -4634 241054
rect -4398 240818 23586 241054
rect 23822 240818 59586 241054
rect 59822 240818 95586 241054
rect 95822 240818 108000 241054
rect -4816 240734 108000 240818
rect -4816 240498 -4634 240734
rect -4398 240498 23586 240734
rect 23822 240498 59586 240734
rect 59822 240498 95586 240734
rect 95822 240498 108000 240734
rect -4816 240476 108000 240498
rect 407589 241054 588740 241076
rect 407589 240943 455586 241054
rect 407589 240929 416782 240943
rect 407589 240914 415373 240929
rect 407589 240900 413972 240914
rect 407589 240885 412563 240900
rect 407589 240871 411083 240885
rect 407589 240856 409674 240871
rect 407589 240842 408273 240856
rect 407589 240606 407878 240842
rect 408114 240620 408273 240842
rect 408509 240620 408593 240856
rect 408829 240620 408967 240856
rect 409203 240620 409287 240856
rect 409523 240635 409674 240856
rect 409910 240635 409994 240871
rect 410230 240635 410368 240871
rect 410604 240635 410688 240871
rect 410924 240649 411083 240871
rect 411319 240649 411403 240885
rect 411639 240649 411777 240885
rect 412013 240649 412097 240885
rect 412333 240664 412563 240885
rect 412799 240664 412883 240900
rect 413119 240664 413257 240900
rect 413493 240664 413577 240900
rect 413813 240678 413972 240900
rect 414208 240678 414292 240914
rect 414528 240678 414666 240914
rect 414902 240678 414986 240914
rect 415222 240693 415373 240914
rect 415609 240693 415693 240929
rect 415929 240693 416067 240929
rect 416303 240693 416387 240929
rect 416623 240707 416782 240929
rect 417018 240707 417102 240943
rect 417338 240707 417476 240943
rect 417712 240707 417796 240943
rect 418032 240818 455586 240943
rect 455822 240818 491586 241054
rect 491822 240818 527586 241054
rect 527822 240818 563586 241054
rect 563822 240818 588322 241054
rect 588558 240818 588740 241054
rect 418032 240734 588740 240818
rect 418032 240707 455586 240734
rect 416623 240693 455586 240707
rect 415222 240678 455586 240693
rect 413813 240664 455586 240678
rect 412333 240649 455586 240664
rect 410924 240635 455586 240649
rect 409523 240620 455586 240635
rect 408114 240606 455586 240620
rect 407589 240498 455586 240606
rect 455822 240498 491586 240734
rect 491822 240498 527586 240734
rect 527822 240498 563586 240734
rect 563822 240498 588322 240734
rect 588558 240498 588740 240734
rect 407589 240476 588740 240498
rect -4816 240474 -4216 240476
rect 23404 240474 24004 240476
rect 59404 240474 60004 240476
rect 95404 240474 96004 240476
rect 455404 240474 456004 240476
rect 491404 240474 492004 240476
rect 527404 240474 528004 240476
rect 563404 240474 564004 240476
rect 588140 240474 588740 240476
rect -2936 237476 -2336 237478
rect 19804 237476 20404 237478
rect 55804 237476 56404 237478
rect 91804 237476 92404 237478
rect 451804 237476 452404 237478
rect 487804 237476 488404 237478
rect 523804 237476 524404 237478
rect 559804 237476 560404 237478
rect 586260 237476 586860 237478
rect -2936 237454 108000 237476
rect -2936 237218 -2754 237454
rect -2518 237218 19986 237454
rect 20222 237218 55986 237454
rect 56222 237218 91986 237454
rect 92222 237218 108000 237454
rect -2936 237134 108000 237218
rect -2936 236898 -2754 237134
rect -2518 236898 19986 237134
rect 20222 236898 55986 237134
rect 56222 236898 91986 237134
rect 92222 236898 108000 237134
rect -2936 236876 108000 236898
rect 425267 237454 586860 237476
rect 425267 237395 451986 237454
rect 425267 237381 434622 237395
rect 425267 237366 433213 237381
rect 425267 237352 431812 237366
rect 425267 237337 430403 237352
rect 425267 237323 428923 237337
rect 425267 237308 427514 237323
rect 425267 237294 426113 237308
rect 425267 237058 425718 237294
rect 425954 237072 426113 237294
rect 426349 237072 426433 237308
rect 426669 237072 426807 237308
rect 427043 237072 427127 237308
rect 427363 237087 427514 237308
rect 427750 237087 427834 237323
rect 428070 237087 428208 237323
rect 428444 237087 428528 237323
rect 428764 237101 428923 237323
rect 429159 237101 429243 237337
rect 429479 237101 429617 237337
rect 429853 237101 429937 237337
rect 430173 237116 430403 237337
rect 430639 237116 430723 237352
rect 430959 237116 431097 237352
rect 431333 237116 431417 237352
rect 431653 237130 431812 237352
rect 432048 237130 432132 237366
rect 432368 237130 432506 237366
rect 432742 237130 432826 237366
rect 433062 237145 433213 237366
rect 433449 237145 433533 237381
rect 433769 237145 433907 237381
rect 434143 237145 434227 237381
rect 434463 237159 434622 237381
rect 434858 237159 434942 237395
rect 435178 237159 435316 237395
rect 435552 237159 435636 237395
rect 435872 237218 451986 237395
rect 452222 237218 487986 237454
rect 488222 237218 523986 237454
rect 524222 237218 559986 237454
rect 560222 237218 586442 237454
rect 586678 237218 586860 237454
rect 435872 237159 586860 237218
rect 434463 237145 586860 237159
rect 433062 237134 586860 237145
rect 433062 237130 451986 237134
rect 431653 237116 451986 237130
rect 430173 237101 451986 237116
rect 428764 237087 451986 237101
rect 427363 237072 451986 237087
rect 425954 237058 451986 237072
rect 425267 236898 451986 237058
rect 452222 236898 487986 237134
rect 488222 236898 523986 237134
rect 524222 236898 559986 237134
rect 560222 236898 586442 237134
rect 586678 236898 586860 237134
rect 425267 236876 586860 236898
rect -2936 236874 -2336 236876
rect 19804 236874 20404 236876
rect 55804 236874 56404 236876
rect 91804 236874 92404 236876
rect 451804 236874 452404 236876
rect 487804 236874 488404 236876
rect 523804 236874 524404 236876
rect 559804 236874 560404 236876
rect 586260 236874 586860 236876
rect -7636 230276 -7036 230278
rect 12604 230276 13204 230278
rect 48604 230276 49204 230278
rect 84604 230276 85204 230278
rect 480604 230276 481204 230278
rect 516604 230276 517204 230278
rect 552604 230276 553204 230278
rect 590960 230276 591560 230278
rect -8576 230254 108000 230276
rect -8576 230018 -7454 230254
rect -7218 230018 12786 230254
rect 13022 230018 48786 230254
rect 49022 230018 84786 230254
rect 85022 230018 108000 230254
rect -8576 229934 108000 230018
rect -8576 229698 -7454 229934
rect -7218 229698 12786 229934
rect 13022 229698 48786 229934
rect 49022 229698 84786 229934
rect 85022 229698 108000 229934
rect -8576 229676 108000 229698
rect 448000 230254 592500 230276
rect 448000 230018 480786 230254
rect 481022 230018 516786 230254
rect 517022 230018 552786 230254
rect 553022 230018 591142 230254
rect 591378 230018 592500 230254
rect 448000 229934 592500 230018
rect 448000 229698 480786 229934
rect 481022 229698 516786 229934
rect 517022 229698 552786 229934
rect 553022 229698 591142 229934
rect 591378 229698 592500 229934
rect 448000 229676 592500 229698
rect -7636 229674 -7036 229676
rect 12604 229674 13204 229676
rect 48604 229674 49204 229676
rect 84604 229674 85204 229676
rect 480604 229674 481204 229676
rect 516604 229674 517204 229676
rect 552604 229674 553204 229676
rect 590960 229674 591560 229676
rect -5756 226676 -5156 226678
rect 9004 226676 9604 226678
rect 45004 226676 45604 226678
rect 81004 226676 81604 226678
rect 477004 226676 477604 226678
rect 513004 226676 513604 226678
rect 549004 226676 549604 226678
rect 589080 226676 589680 226678
rect -6696 226654 108000 226676
rect -6696 226418 -5574 226654
rect -5338 226418 9186 226654
rect 9422 226418 45186 226654
rect 45422 226418 81186 226654
rect 81422 226418 108000 226654
rect -6696 226334 108000 226418
rect -6696 226098 -5574 226334
rect -5338 226098 9186 226334
rect 9422 226098 45186 226334
rect 45422 226098 81186 226334
rect 81422 226098 108000 226334
rect -6696 226076 108000 226098
rect 448000 226654 590620 226676
rect 448000 226418 477186 226654
rect 477422 226418 513186 226654
rect 513422 226418 549186 226654
rect 549422 226418 589262 226654
rect 589498 226418 590620 226654
rect 448000 226334 590620 226418
rect 448000 226098 477186 226334
rect 477422 226098 513186 226334
rect 513422 226098 549186 226334
rect 549422 226098 589262 226334
rect 589498 226098 590620 226334
rect 448000 226076 590620 226098
rect -5756 226074 -5156 226076
rect 9004 226074 9604 226076
rect 45004 226074 45604 226076
rect 81004 226074 81604 226076
rect 477004 226074 477604 226076
rect 513004 226074 513604 226076
rect 549004 226074 549604 226076
rect 589080 226074 589680 226076
rect -3876 223076 -3276 223078
rect 5404 223076 6004 223078
rect 41404 223076 42004 223078
rect 77404 223076 78004 223078
rect 473404 223076 474004 223078
rect 509404 223076 510004 223078
rect 545404 223076 546004 223078
rect 581404 223076 582004 223078
rect 587200 223076 587800 223078
rect -4816 223054 108000 223076
rect -4816 222818 -3694 223054
rect -3458 222818 5586 223054
rect 5822 222818 41586 223054
rect 41822 222818 77586 223054
rect 77822 222818 108000 223054
rect -4816 222734 108000 222818
rect -4816 222498 -3694 222734
rect -3458 222498 5586 222734
rect 5822 222498 41586 222734
rect 41822 222498 77586 222734
rect 77822 222498 108000 222734
rect -4816 222476 108000 222498
rect 448000 223054 588740 223076
rect 448000 222818 473586 223054
rect 473822 222818 509586 223054
rect 509822 222818 545586 223054
rect 545822 222818 581586 223054
rect 581822 222818 587382 223054
rect 587618 222818 588740 223054
rect 448000 222734 588740 222818
rect 448000 222498 473586 222734
rect 473822 222498 509586 222734
rect 509822 222498 545586 222734
rect 545822 222498 581586 222734
rect 581822 222498 587382 222734
rect 587618 222498 588740 222734
rect 448000 222476 588740 222498
rect -3876 222474 -3276 222476
rect 5404 222474 6004 222476
rect 41404 222474 42004 222476
rect 77404 222474 78004 222476
rect 473404 222474 474004 222476
rect 509404 222474 510004 222476
rect 545404 222474 546004 222476
rect 581404 222474 582004 222476
rect 587200 222474 587800 222476
rect -1996 219476 -1396 219478
rect 1804 219476 2404 219478
rect 37804 219476 38404 219478
rect 73804 219476 74404 219478
rect 469804 219476 470404 219478
rect 505804 219476 506404 219478
rect 541804 219476 542404 219478
rect 577804 219476 578404 219478
rect 585320 219476 585920 219478
rect -2936 219454 108000 219476
rect -2936 219218 -1814 219454
rect -1578 219218 1986 219454
rect 2222 219218 37986 219454
rect 38222 219218 73986 219454
rect 74222 219218 108000 219454
rect -2936 219134 108000 219218
rect -2936 218898 -1814 219134
rect -1578 218898 1986 219134
rect 2222 218898 37986 219134
rect 38222 218898 73986 219134
rect 74222 218898 108000 219134
rect -2936 218876 108000 218898
rect 448000 219454 586860 219476
rect 448000 219218 469986 219454
rect 470222 219218 505986 219454
rect 506222 219218 541986 219454
rect 542222 219218 577986 219454
rect 578222 219218 585502 219454
rect 585738 219218 586860 219454
rect 448000 219134 586860 219218
rect 448000 218898 469986 219134
rect 470222 218898 505986 219134
rect 506222 218898 541986 219134
rect 542222 218898 577986 219134
rect 578222 218898 585502 219134
rect 585738 218898 586860 219134
rect 448000 218876 586860 218898
rect -1996 218874 -1396 218876
rect 1804 218874 2404 218876
rect 37804 218874 38404 218876
rect 73804 218874 74404 218876
rect 469804 218874 470404 218876
rect 505804 218874 506404 218876
rect 541804 218874 542404 218876
rect 577804 218874 578404 218876
rect 585320 218874 585920 218876
rect -8576 212276 -7976 212278
rect 30604 212276 31204 212278
rect 66604 212276 67204 212278
rect 102604 212276 103204 212278
rect 138604 212276 139204 212278
rect 174604 212276 175204 212278
rect 210604 212276 211204 212278
rect 246604 212276 247204 212278
rect 282604 212276 283204 212278
rect 318604 212276 319204 212278
rect 354604 212276 355204 212278
rect 390604 212276 391204 212278
rect 426604 212276 427204 212278
rect 462604 212276 463204 212278
rect 498604 212276 499204 212278
rect 534604 212276 535204 212278
rect 570604 212276 571204 212278
rect 591900 212276 592500 212278
rect -8576 212254 592500 212276
rect -8576 212018 -8394 212254
rect -8158 212018 30786 212254
rect 31022 212018 66786 212254
rect 67022 212018 102786 212254
rect 103022 212018 138786 212254
rect 139022 212018 174786 212254
rect 175022 212018 210786 212254
rect 211022 212018 246786 212254
rect 247022 212018 282786 212254
rect 283022 212018 318786 212254
rect 319022 212018 354786 212254
rect 355022 212018 390786 212254
rect 391022 212018 426786 212254
rect 427022 212018 462786 212254
rect 463022 212018 498786 212254
rect 499022 212018 534786 212254
rect 535022 212018 570786 212254
rect 571022 212018 592082 212254
rect 592318 212018 592500 212254
rect -8576 211934 592500 212018
rect -8576 211698 -8394 211934
rect -8158 211698 30786 211934
rect 31022 211698 66786 211934
rect 67022 211698 102786 211934
rect 103022 211698 138786 211934
rect 139022 211698 174786 211934
rect 175022 211698 210786 211934
rect 211022 211698 246786 211934
rect 247022 211698 282786 211934
rect 283022 211698 318786 211934
rect 319022 211698 354786 211934
rect 355022 211698 390786 211934
rect 391022 211698 426786 211934
rect 427022 211698 462786 211934
rect 463022 211698 498786 211934
rect 499022 211698 534786 211934
rect 535022 211698 570786 211934
rect 571022 211698 592082 211934
rect 592318 211698 592500 211934
rect -8576 211676 592500 211698
rect -8576 211674 -7976 211676
rect 30604 211674 31204 211676
rect 66604 211674 67204 211676
rect 102604 211674 103204 211676
rect 138604 211674 139204 211676
rect 174604 211674 175204 211676
rect 210604 211674 211204 211676
rect 246604 211674 247204 211676
rect 282604 211674 283204 211676
rect 318604 211674 319204 211676
rect 354604 211674 355204 211676
rect 390604 211674 391204 211676
rect 426604 211674 427204 211676
rect 462604 211674 463204 211676
rect 498604 211674 499204 211676
rect 534604 211674 535204 211676
rect 570604 211674 571204 211676
rect 591900 211674 592500 211676
rect -6696 208676 -6096 208678
rect 27004 208676 27604 208678
rect 63004 208676 63604 208678
rect 99004 208676 99604 208678
rect 135004 208676 135604 208678
rect 171004 208676 171604 208678
rect 207004 208676 207604 208678
rect 243004 208676 243604 208678
rect 279004 208676 279604 208678
rect 315004 208676 315604 208678
rect 351004 208676 351604 208678
rect 387004 208676 387604 208678
rect 423004 208676 423604 208678
rect 459004 208676 459604 208678
rect 495004 208676 495604 208678
rect 531004 208676 531604 208678
rect 567004 208676 567604 208678
rect 590020 208676 590620 208678
rect -6696 208654 590620 208676
rect -6696 208418 -6514 208654
rect -6278 208418 27186 208654
rect 27422 208418 63186 208654
rect 63422 208418 99186 208654
rect 99422 208418 135186 208654
rect 135422 208418 171186 208654
rect 171422 208418 207186 208654
rect 207422 208418 243186 208654
rect 243422 208418 279186 208654
rect 279422 208418 315186 208654
rect 315422 208418 351186 208654
rect 351422 208418 387186 208654
rect 387422 208418 423186 208654
rect 423422 208418 459186 208654
rect 459422 208418 495186 208654
rect 495422 208418 531186 208654
rect 531422 208418 567186 208654
rect 567422 208418 590202 208654
rect 590438 208418 590620 208654
rect -6696 208334 590620 208418
rect -6696 208098 -6514 208334
rect -6278 208098 27186 208334
rect 27422 208098 63186 208334
rect 63422 208098 99186 208334
rect 99422 208098 135186 208334
rect 135422 208098 171186 208334
rect 171422 208098 207186 208334
rect 207422 208098 243186 208334
rect 243422 208098 279186 208334
rect 279422 208098 315186 208334
rect 315422 208098 351186 208334
rect 351422 208098 387186 208334
rect 387422 208098 423186 208334
rect 423422 208098 459186 208334
rect 459422 208098 495186 208334
rect 495422 208098 531186 208334
rect 531422 208098 567186 208334
rect 567422 208098 590202 208334
rect 590438 208098 590620 208334
rect -6696 208076 590620 208098
rect -6696 208074 -6096 208076
rect 27004 208074 27604 208076
rect 63004 208074 63604 208076
rect 99004 208074 99604 208076
rect 135004 208074 135604 208076
rect 171004 208074 171604 208076
rect 207004 208074 207604 208076
rect 243004 208074 243604 208076
rect 279004 208074 279604 208076
rect 315004 208074 315604 208076
rect 351004 208074 351604 208076
rect 387004 208074 387604 208076
rect 423004 208074 423604 208076
rect 459004 208074 459604 208076
rect 495004 208074 495604 208076
rect 531004 208074 531604 208076
rect 567004 208074 567604 208076
rect 590020 208074 590620 208076
rect -4816 205076 -4216 205078
rect 23404 205076 24004 205078
rect 59404 205076 60004 205078
rect 95404 205076 96004 205078
rect 131404 205076 132004 205078
rect 167404 205076 168004 205078
rect 203404 205076 204004 205078
rect 239404 205076 240004 205078
rect 275404 205076 276004 205078
rect 311404 205076 312004 205078
rect 347404 205076 348004 205078
rect 383404 205076 384004 205078
rect 419404 205076 420004 205078
rect 455404 205076 456004 205078
rect 491404 205076 492004 205078
rect 527404 205076 528004 205078
rect 563404 205076 564004 205078
rect 588140 205076 588740 205078
rect -4816 205054 588740 205076
rect -4816 204818 -4634 205054
rect -4398 204818 23586 205054
rect 23822 204818 59586 205054
rect 59822 204818 95586 205054
rect 95822 204818 131586 205054
rect 131822 204818 167586 205054
rect 167822 204818 203586 205054
rect 203822 204818 239586 205054
rect 239822 204818 275586 205054
rect 275822 204818 311586 205054
rect 311822 204818 347586 205054
rect 347822 204818 383586 205054
rect 383822 204818 419586 205054
rect 419822 204818 455586 205054
rect 455822 204818 491586 205054
rect 491822 204818 527586 205054
rect 527822 204818 563586 205054
rect 563822 204818 588322 205054
rect 588558 204818 588740 205054
rect -4816 204734 588740 204818
rect -4816 204498 -4634 204734
rect -4398 204498 23586 204734
rect 23822 204498 59586 204734
rect 59822 204498 95586 204734
rect 95822 204498 131586 204734
rect 131822 204498 167586 204734
rect 167822 204498 203586 204734
rect 203822 204498 239586 204734
rect 239822 204498 275586 204734
rect 275822 204498 311586 204734
rect 311822 204498 347586 204734
rect 347822 204498 383586 204734
rect 383822 204498 419586 204734
rect 419822 204498 455586 204734
rect 455822 204498 491586 204734
rect 491822 204498 527586 204734
rect 527822 204498 563586 204734
rect 563822 204498 588322 204734
rect 588558 204498 588740 204734
rect -4816 204476 588740 204498
rect -4816 204474 -4216 204476
rect 23404 204474 24004 204476
rect 59404 204474 60004 204476
rect 95404 204474 96004 204476
rect 131404 204474 132004 204476
rect 167404 204474 168004 204476
rect 203404 204474 204004 204476
rect 239404 204474 240004 204476
rect 275404 204474 276004 204476
rect 311404 204474 312004 204476
rect 347404 204474 348004 204476
rect 383404 204474 384004 204476
rect 419404 204474 420004 204476
rect 455404 204474 456004 204476
rect 491404 204474 492004 204476
rect 527404 204474 528004 204476
rect 563404 204474 564004 204476
rect 588140 204474 588740 204476
rect -2936 201476 -2336 201478
rect 19804 201476 20404 201478
rect 55804 201476 56404 201478
rect 91804 201476 92404 201478
rect 127804 201476 128404 201478
rect 163804 201476 164404 201478
rect 199804 201476 200404 201478
rect 235804 201476 236404 201478
rect 271804 201476 272404 201478
rect 307804 201476 308404 201478
rect 343804 201476 344404 201478
rect 379804 201476 380404 201478
rect 415804 201476 416404 201478
rect 451804 201476 452404 201478
rect 487804 201476 488404 201478
rect 523804 201476 524404 201478
rect 559804 201476 560404 201478
rect 586260 201476 586860 201478
rect -2936 201454 586860 201476
rect -2936 201218 -2754 201454
rect -2518 201218 19986 201454
rect 20222 201218 55986 201454
rect 56222 201218 91986 201454
rect 92222 201218 127986 201454
rect 128222 201218 163986 201454
rect 164222 201218 199986 201454
rect 200222 201218 235986 201454
rect 236222 201218 271986 201454
rect 272222 201218 307986 201454
rect 308222 201218 343986 201454
rect 344222 201218 379986 201454
rect 380222 201218 415986 201454
rect 416222 201218 451986 201454
rect 452222 201218 487986 201454
rect 488222 201218 523986 201454
rect 524222 201218 559986 201454
rect 560222 201218 586442 201454
rect 586678 201218 586860 201454
rect -2936 201134 586860 201218
rect -2936 200898 -2754 201134
rect -2518 200898 19986 201134
rect 20222 200898 55986 201134
rect 56222 200898 91986 201134
rect 92222 200898 127986 201134
rect 128222 200898 163986 201134
rect 164222 200898 199986 201134
rect 200222 200898 235986 201134
rect 236222 200898 271986 201134
rect 272222 200898 307986 201134
rect 308222 200898 343986 201134
rect 344222 200898 379986 201134
rect 380222 200898 415986 201134
rect 416222 200898 451986 201134
rect 452222 200898 487986 201134
rect 488222 200898 523986 201134
rect 524222 200898 559986 201134
rect 560222 200898 586442 201134
rect 586678 200898 586860 201134
rect -2936 200876 586860 200898
rect -2936 200874 -2336 200876
rect 19804 200874 20404 200876
rect 55804 200874 56404 200876
rect 91804 200874 92404 200876
rect 127804 200874 128404 200876
rect 163804 200874 164404 200876
rect 199804 200874 200404 200876
rect 235804 200874 236404 200876
rect 271804 200874 272404 200876
rect 307804 200874 308404 200876
rect 343804 200874 344404 200876
rect 379804 200874 380404 200876
rect 415804 200874 416404 200876
rect 451804 200874 452404 200876
rect 487804 200874 488404 200876
rect 523804 200874 524404 200876
rect 559804 200874 560404 200876
rect 586260 200874 586860 200876
rect -7636 194276 -7036 194278
rect 12604 194276 13204 194278
rect 48604 194276 49204 194278
rect 84604 194276 85204 194278
rect 120604 194276 121204 194278
rect 156604 194276 157204 194278
rect 192604 194276 193204 194278
rect 228604 194276 229204 194278
rect 264604 194276 265204 194278
rect 300604 194276 301204 194278
rect 336604 194276 337204 194278
rect 372604 194276 373204 194278
rect 408604 194276 409204 194278
rect 444604 194276 445204 194278
rect 480604 194276 481204 194278
rect 516604 194276 517204 194278
rect 552604 194276 553204 194278
rect 590960 194276 591560 194278
rect -8576 194254 592500 194276
rect -8576 194018 -7454 194254
rect -7218 194018 12786 194254
rect 13022 194018 48786 194254
rect 49022 194018 84786 194254
rect 85022 194018 120786 194254
rect 121022 194018 156786 194254
rect 157022 194018 192786 194254
rect 193022 194018 228786 194254
rect 229022 194018 264786 194254
rect 265022 194018 300786 194254
rect 301022 194018 336786 194254
rect 337022 194018 372786 194254
rect 373022 194018 408786 194254
rect 409022 194018 444786 194254
rect 445022 194018 480786 194254
rect 481022 194018 516786 194254
rect 517022 194018 552786 194254
rect 553022 194018 591142 194254
rect 591378 194018 592500 194254
rect -8576 193934 592500 194018
rect -8576 193698 -7454 193934
rect -7218 193698 12786 193934
rect 13022 193698 48786 193934
rect 49022 193698 84786 193934
rect 85022 193698 120786 193934
rect 121022 193698 156786 193934
rect 157022 193698 192786 193934
rect 193022 193698 228786 193934
rect 229022 193698 264786 193934
rect 265022 193698 300786 193934
rect 301022 193698 336786 193934
rect 337022 193698 372786 193934
rect 373022 193698 408786 193934
rect 409022 193698 444786 193934
rect 445022 193698 480786 193934
rect 481022 193698 516786 193934
rect 517022 193698 552786 193934
rect 553022 193698 591142 193934
rect 591378 193698 592500 193934
rect -8576 193676 592500 193698
rect -7636 193674 -7036 193676
rect 12604 193674 13204 193676
rect 48604 193674 49204 193676
rect 84604 193674 85204 193676
rect 120604 193674 121204 193676
rect 156604 193674 157204 193676
rect 192604 193674 193204 193676
rect 228604 193674 229204 193676
rect 264604 193674 265204 193676
rect 300604 193674 301204 193676
rect 336604 193674 337204 193676
rect 372604 193674 373204 193676
rect 408604 193674 409204 193676
rect 444604 193674 445204 193676
rect 480604 193674 481204 193676
rect 516604 193674 517204 193676
rect 552604 193674 553204 193676
rect 590960 193674 591560 193676
rect -5756 190676 -5156 190678
rect 9004 190676 9604 190678
rect 45004 190676 45604 190678
rect 81004 190676 81604 190678
rect 117004 190676 117604 190678
rect 153004 190676 153604 190678
rect 189004 190676 189604 190678
rect 225004 190676 225604 190678
rect 261004 190676 261604 190678
rect 297004 190676 297604 190678
rect 333004 190676 333604 190678
rect 369004 190676 369604 190678
rect 405004 190676 405604 190678
rect 441004 190676 441604 190678
rect 477004 190676 477604 190678
rect 513004 190676 513604 190678
rect 549004 190676 549604 190678
rect 589080 190676 589680 190678
rect -6696 190654 590620 190676
rect -6696 190418 -5574 190654
rect -5338 190418 9186 190654
rect 9422 190418 45186 190654
rect 45422 190418 81186 190654
rect 81422 190418 117186 190654
rect 117422 190418 153186 190654
rect 153422 190418 189186 190654
rect 189422 190418 225186 190654
rect 225422 190418 261186 190654
rect 261422 190418 297186 190654
rect 297422 190418 333186 190654
rect 333422 190418 369186 190654
rect 369422 190418 405186 190654
rect 405422 190418 441186 190654
rect 441422 190418 477186 190654
rect 477422 190418 513186 190654
rect 513422 190418 549186 190654
rect 549422 190418 589262 190654
rect 589498 190418 590620 190654
rect -6696 190334 590620 190418
rect -6696 190098 -5574 190334
rect -5338 190098 9186 190334
rect 9422 190098 45186 190334
rect 45422 190098 81186 190334
rect 81422 190098 117186 190334
rect 117422 190098 153186 190334
rect 153422 190098 189186 190334
rect 189422 190098 225186 190334
rect 225422 190098 261186 190334
rect 261422 190098 297186 190334
rect 297422 190098 333186 190334
rect 333422 190098 369186 190334
rect 369422 190098 405186 190334
rect 405422 190098 441186 190334
rect 441422 190098 477186 190334
rect 477422 190098 513186 190334
rect 513422 190098 549186 190334
rect 549422 190098 589262 190334
rect 589498 190098 590620 190334
rect -6696 190076 590620 190098
rect -5756 190074 -5156 190076
rect 9004 190074 9604 190076
rect 45004 190074 45604 190076
rect 81004 190074 81604 190076
rect 117004 190074 117604 190076
rect 153004 190074 153604 190076
rect 189004 190074 189604 190076
rect 225004 190074 225604 190076
rect 261004 190074 261604 190076
rect 297004 190074 297604 190076
rect 333004 190074 333604 190076
rect 369004 190074 369604 190076
rect 405004 190074 405604 190076
rect 441004 190074 441604 190076
rect 477004 190074 477604 190076
rect 513004 190074 513604 190076
rect 549004 190074 549604 190076
rect 589080 190074 589680 190076
rect -3876 187076 -3276 187078
rect 5404 187076 6004 187078
rect 41404 187076 42004 187078
rect 77404 187076 78004 187078
rect 113404 187076 114004 187078
rect 149404 187076 150004 187078
rect 185404 187076 186004 187078
rect 221404 187076 222004 187078
rect 257404 187076 258004 187078
rect 293404 187076 294004 187078
rect 329404 187076 330004 187078
rect 365404 187076 366004 187078
rect 401404 187076 402004 187078
rect 437404 187076 438004 187078
rect 473404 187076 474004 187078
rect 509404 187076 510004 187078
rect 545404 187076 546004 187078
rect 581404 187076 582004 187078
rect 587200 187076 587800 187078
rect -4816 187054 588740 187076
rect -4816 186818 -3694 187054
rect -3458 186818 5586 187054
rect 5822 186818 41586 187054
rect 41822 186818 77586 187054
rect 77822 186818 113586 187054
rect 113822 186818 149586 187054
rect 149822 186818 185586 187054
rect 185822 186818 221586 187054
rect 221822 186818 257586 187054
rect 257822 186818 293586 187054
rect 293822 186818 329586 187054
rect 329822 186818 365586 187054
rect 365822 186818 401586 187054
rect 401822 186818 437586 187054
rect 437822 186818 473586 187054
rect 473822 186818 509586 187054
rect 509822 186818 545586 187054
rect 545822 186818 581586 187054
rect 581822 186818 587382 187054
rect 587618 186818 588740 187054
rect -4816 186734 588740 186818
rect -4816 186498 -3694 186734
rect -3458 186498 5586 186734
rect 5822 186498 41586 186734
rect 41822 186498 77586 186734
rect 77822 186498 113586 186734
rect 113822 186498 149586 186734
rect 149822 186498 185586 186734
rect 185822 186498 221586 186734
rect 221822 186498 257586 186734
rect 257822 186498 293586 186734
rect 293822 186498 329586 186734
rect 329822 186498 365586 186734
rect 365822 186498 401586 186734
rect 401822 186498 437586 186734
rect 437822 186498 473586 186734
rect 473822 186498 509586 186734
rect 509822 186498 545586 186734
rect 545822 186498 581586 186734
rect 581822 186498 587382 186734
rect 587618 186498 588740 186734
rect -4816 186476 588740 186498
rect -3876 186474 -3276 186476
rect 5404 186474 6004 186476
rect 41404 186474 42004 186476
rect 77404 186474 78004 186476
rect 113404 186474 114004 186476
rect 149404 186474 150004 186476
rect 185404 186474 186004 186476
rect 221404 186474 222004 186476
rect 257404 186474 258004 186476
rect 293404 186474 294004 186476
rect 329404 186474 330004 186476
rect 365404 186474 366004 186476
rect 401404 186474 402004 186476
rect 437404 186474 438004 186476
rect 473404 186474 474004 186476
rect 509404 186474 510004 186476
rect 545404 186474 546004 186476
rect 581404 186474 582004 186476
rect 587200 186474 587800 186476
rect -1996 183476 -1396 183478
rect 1804 183476 2404 183478
rect 37804 183476 38404 183478
rect 73804 183476 74404 183478
rect 109804 183476 110404 183478
rect 145804 183476 146404 183478
rect 181804 183476 182404 183478
rect 217804 183476 218404 183478
rect 253804 183476 254404 183478
rect 289804 183476 290404 183478
rect 325804 183476 326404 183478
rect 361804 183476 362404 183478
rect 397804 183476 398404 183478
rect 433804 183476 434404 183478
rect 469804 183476 470404 183478
rect 505804 183476 506404 183478
rect 541804 183476 542404 183478
rect 577804 183476 578404 183478
rect 585320 183476 585920 183478
rect -2936 183454 586860 183476
rect -2936 183218 -1814 183454
rect -1578 183218 1986 183454
rect 2222 183218 37986 183454
rect 38222 183218 73986 183454
rect 74222 183218 109986 183454
rect 110222 183218 145986 183454
rect 146222 183218 181986 183454
rect 182222 183218 217986 183454
rect 218222 183218 253986 183454
rect 254222 183218 289986 183454
rect 290222 183218 325986 183454
rect 326222 183218 361986 183454
rect 362222 183218 397986 183454
rect 398222 183218 433986 183454
rect 434222 183218 469986 183454
rect 470222 183218 505986 183454
rect 506222 183218 541986 183454
rect 542222 183218 577986 183454
rect 578222 183218 585502 183454
rect 585738 183218 586860 183454
rect -2936 183134 586860 183218
rect -2936 182898 -1814 183134
rect -1578 182898 1986 183134
rect 2222 182898 37986 183134
rect 38222 182898 73986 183134
rect 74222 182898 109986 183134
rect 110222 182898 145986 183134
rect 146222 182898 181986 183134
rect 182222 182898 217986 183134
rect 218222 182898 253986 183134
rect 254222 182898 289986 183134
rect 290222 182898 325986 183134
rect 326222 182898 361986 183134
rect 362222 182898 397986 183134
rect 398222 182898 433986 183134
rect 434222 182898 469986 183134
rect 470222 182898 505986 183134
rect 506222 182898 541986 183134
rect 542222 182898 577986 183134
rect 578222 182898 585502 183134
rect 585738 182898 586860 183134
rect -2936 182876 586860 182898
rect -1996 182874 -1396 182876
rect 1804 182874 2404 182876
rect 37804 182874 38404 182876
rect 73804 182874 74404 182876
rect 109804 182874 110404 182876
rect 145804 182874 146404 182876
rect 181804 182874 182404 182876
rect 217804 182874 218404 182876
rect 253804 182874 254404 182876
rect 289804 182874 290404 182876
rect 325804 182874 326404 182876
rect 361804 182874 362404 182876
rect 397804 182874 398404 182876
rect 433804 182874 434404 182876
rect 469804 182874 470404 182876
rect 505804 182874 506404 182876
rect 541804 182874 542404 182876
rect 577804 182874 578404 182876
rect 585320 182874 585920 182876
rect -8576 176276 -7976 176278
rect 30604 176276 31204 176278
rect 66604 176276 67204 176278
rect 102604 176276 103204 176278
rect 138604 176276 139204 176278
rect 174604 176276 175204 176278
rect 210604 176276 211204 176278
rect 246604 176276 247204 176278
rect 282604 176276 283204 176278
rect 318604 176276 319204 176278
rect 354604 176276 355204 176278
rect 390604 176276 391204 176278
rect 426604 176276 427204 176278
rect 462604 176276 463204 176278
rect 498604 176276 499204 176278
rect 534604 176276 535204 176278
rect 570604 176276 571204 176278
rect 591900 176276 592500 176278
rect -8576 176254 592500 176276
rect -8576 176018 -8394 176254
rect -8158 176018 30786 176254
rect 31022 176018 66786 176254
rect 67022 176018 102786 176254
rect 103022 176018 138786 176254
rect 139022 176018 174786 176254
rect 175022 176018 210786 176254
rect 211022 176018 246786 176254
rect 247022 176018 282786 176254
rect 283022 176018 318786 176254
rect 319022 176018 354786 176254
rect 355022 176018 390786 176254
rect 391022 176018 426786 176254
rect 427022 176018 462786 176254
rect 463022 176018 498786 176254
rect 499022 176018 534786 176254
rect 535022 176018 570786 176254
rect 571022 176018 592082 176254
rect 592318 176018 592500 176254
rect -8576 175934 592500 176018
rect -8576 175698 -8394 175934
rect -8158 175698 30786 175934
rect 31022 175698 66786 175934
rect 67022 175698 102786 175934
rect 103022 175698 138786 175934
rect 139022 175698 174786 175934
rect 175022 175698 210786 175934
rect 211022 175698 246786 175934
rect 247022 175698 282786 175934
rect 283022 175698 318786 175934
rect 319022 175698 354786 175934
rect 355022 175698 390786 175934
rect 391022 175698 426786 175934
rect 427022 175698 462786 175934
rect 463022 175698 498786 175934
rect 499022 175698 534786 175934
rect 535022 175698 570786 175934
rect 571022 175698 592082 175934
rect 592318 175698 592500 175934
rect -8576 175676 592500 175698
rect -8576 175674 -7976 175676
rect 30604 175674 31204 175676
rect 66604 175674 67204 175676
rect 102604 175674 103204 175676
rect 138604 175674 139204 175676
rect 174604 175674 175204 175676
rect 210604 175674 211204 175676
rect 246604 175674 247204 175676
rect 282604 175674 283204 175676
rect 318604 175674 319204 175676
rect 354604 175674 355204 175676
rect 390604 175674 391204 175676
rect 426604 175674 427204 175676
rect 462604 175674 463204 175676
rect 498604 175674 499204 175676
rect 534604 175674 535204 175676
rect 570604 175674 571204 175676
rect 591900 175674 592500 175676
rect -6696 172676 -6096 172678
rect 27004 172676 27604 172678
rect 63004 172676 63604 172678
rect 99004 172676 99604 172678
rect 135004 172676 135604 172678
rect 171004 172676 171604 172678
rect 207004 172676 207604 172678
rect 243004 172676 243604 172678
rect 279004 172676 279604 172678
rect 315004 172676 315604 172678
rect 351004 172676 351604 172678
rect 387004 172676 387604 172678
rect 423004 172676 423604 172678
rect 459004 172676 459604 172678
rect 495004 172676 495604 172678
rect 531004 172676 531604 172678
rect 567004 172676 567604 172678
rect 590020 172676 590620 172678
rect -6696 172654 590620 172676
rect -6696 172418 -6514 172654
rect -6278 172418 27186 172654
rect 27422 172418 63186 172654
rect 63422 172418 99186 172654
rect 99422 172418 135186 172654
rect 135422 172418 171186 172654
rect 171422 172418 207186 172654
rect 207422 172418 243186 172654
rect 243422 172418 279186 172654
rect 279422 172418 315186 172654
rect 315422 172418 351186 172654
rect 351422 172418 387186 172654
rect 387422 172418 423186 172654
rect 423422 172418 459186 172654
rect 459422 172418 495186 172654
rect 495422 172418 531186 172654
rect 531422 172418 567186 172654
rect 567422 172418 590202 172654
rect 590438 172418 590620 172654
rect -6696 172334 590620 172418
rect -6696 172098 -6514 172334
rect -6278 172098 27186 172334
rect 27422 172098 63186 172334
rect 63422 172098 99186 172334
rect 99422 172098 135186 172334
rect 135422 172098 171186 172334
rect 171422 172098 207186 172334
rect 207422 172098 243186 172334
rect 243422 172098 279186 172334
rect 279422 172098 315186 172334
rect 315422 172098 351186 172334
rect 351422 172098 387186 172334
rect 387422 172098 423186 172334
rect 423422 172098 459186 172334
rect 459422 172098 495186 172334
rect 495422 172098 531186 172334
rect 531422 172098 567186 172334
rect 567422 172098 590202 172334
rect 590438 172098 590620 172334
rect -6696 172076 590620 172098
rect -6696 172074 -6096 172076
rect 27004 172074 27604 172076
rect 63004 172074 63604 172076
rect 99004 172074 99604 172076
rect 135004 172074 135604 172076
rect 171004 172074 171604 172076
rect 207004 172074 207604 172076
rect 243004 172074 243604 172076
rect 279004 172074 279604 172076
rect 315004 172074 315604 172076
rect 351004 172074 351604 172076
rect 387004 172074 387604 172076
rect 423004 172074 423604 172076
rect 459004 172074 459604 172076
rect 495004 172074 495604 172076
rect 531004 172074 531604 172076
rect 567004 172074 567604 172076
rect 590020 172074 590620 172076
rect -4816 169076 -4216 169078
rect 23404 169076 24004 169078
rect 59404 169076 60004 169078
rect 95404 169076 96004 169078
rect 131404 169076 132004 169078
rect 167404 169076 168004 169078
rect 203404 169076 204004 169078
rect 239404 169076 240004 169078
rect 275404 169076 276004 169078
rect 311404 169076 312004 169078
rect 347404 169076 348004 169078
rect 383404 169076 384004 169078
rect 419404 169076 420004 169078
rect 455404 169076 456004 169078
rect 491404 169076 492004 169078
rect 527404 169076 528004 169078
rect 563404 169076 564004 169078
rect 588140 169076 588740 169078
rect -4816 169054 588740 169076
rect -4816 168818 -4634 169054
rect -4398 168818 23586 169054
rect 23822 168818 59586 169054
rect 59822 168818 95586 169054
rect 95822 168818 131586 169054
rect 131822 168818 167586 169054
rect 167822 168818 203586 169054
rect 203822 168818 239586 169054
rect 239822 168818 275586 169054
rect 275822 168818 311586 169054
rect 311822 168818 347586 169054
rect 347822 168818 383586 169054
rect 383822 168818 419586 169054
rect 419822 168818 455586 169054
rect 455822 168818 491586 169054
rect 491822 168818 527586 169054
rect 527822 168818 563586 169054
rect 563822 168818 588322 169054
rect 588558 168818 588740 169054
rect -4816 168734 588740 168818
rect -4816 168498 -4634 168734
rect -4398 168498 23586 168734
rect 23822 168498 59586 168734
rect 59822 168498 95586 168734
rect 95822 168498 131586 168734
rect 131822 168498 167586 168734
rect 167822 168498 203586 168734
rect 203822 168498 239586 168734
rect 239822 168498 275586 168734
rect 275822 168498 311586 168734
rect 311822 168498 347586 168734
rect 347822 168498 383586 168734
rect 383822 168498 419586 168734
rect 419822 168498 455586 168734
rect 455822 168498 491586 168734
rect 491822 168498 527586 168734
rect 527822 168498 563586 168734
rect 563822 168498 588322 168734
rect 588558 168498 588740 168734
rect -4816 168476 588740 168498
rect -4816 168474 -4216 168476
rect 23404 168474 24004 168476
rect 59404 168474 60004 168476
rect 95404 168474 96004 168476
rect 131404 168474 132004 168476
rect 167404 168474 168004 168476
rect 203404 168474 204004 168476
rect 239404 168474 240004 168476
rect 275404 168474 276004 168476
rect 311404 168474 312004 168476
rect 347404 168474 348004 168476
rect 383404 168474 384004 168476
rect 419404 168474 420004 168476
rect 455404 168474 456004 168476
rect 491404 168474 492004 168476
rect 527404 168474 528004 168476
rect 563404 168474 564004 168476
rect 588140 168474 588740 168476
rect -2936 165476 -2336 165478
rect 19804 165476 20404 165478
rect 55804 165476 56404 165478
rect 91804 165476 92404 165478
rect 127804 165476 128404 165478
rect 163804 165476 164404 165478
rect 199804 165476 200404 165478
rect 235804 165476 236404 165478
rect 271804 165476 272404 165478
rect 307804 165476 308404 165478
rect 343804 165476 344404 165478
rect 379804 165476 380404 165478
rect 415804 165476 416404 165478
rect 451804 165476 452404 165478
rect 487804 165476 488404 165478
rect 523804 165476 524404 165478
rect 559804 165476 560404 165478
rect 586260 165476 586860 165478
rect -2936 165454 586860 165476
rect -2936 165218 -2754 165454
rect -2518 165218 19986 165454
rect 20222 165218 55986 165454
rect 56222 165218 91986 165454
rect 92222 165218 127986 165454
rect 128222 165218 163986 165454
rect 164222 165218 199986 165454
rect 200222 165218 235986 165454
rect 236222 165218 271986 165454
rect 272222 165218 307986 165454
rect 308222 165218 343986 165454
rect 344222 165218 379986 165454
rect 380222 165218 415986 165454
rect 416222 165218 451986 165454
rect 452222 165218 487986 165454
rect 488222 165218 523986 165454
rect 524222 165218 559986 165454
rect 560222 165218 586442 165454
rect 586678 165218 586860 165454
rect -2936 165134 586860 165218
rect -2936 164898 -2754 165134
rect -2518 164898 19986 165134
rect 20222 164898 55986 165134
rect 56222 164898 91986 165134
rect 92222 164898 127986 165134
rect 128222 164898 163986 165134
rect 164222 164898 199986 165134
rect 200222 164898 235986 165134
rect 236222 164898 271986 165134
rect 272222 164898 307986 165134
rect 308222 164898 343986 165134
rect 344222 164898 379986 165134
rect 380222 164898 415986 165134
rect 416222 164898 451986 165134
rect 452222 164898 487986 165134
rect 488222 164898 523986 165134
rect 524222 164898 559986 165134
rect 560222 164898 586442 165134
rect 586678 164898 586860 165134
rect -2936 164876 586860 164898
rect -2936 164874 -2336 164876
rect 19804 164874 20404 164876
rect 55804 164874 56404 164876
rect 91804 164874 92404 164876
rect 127804 164874 128404 164876
rect 163804 164874 164404 164876
rect 199804 164874 200404 164876
rect 235804 164874 236404 164876
rect 271804 164874 272404 164876
rect 307804 164874 308404 164876
rect 343804 164874 344404 164876
rect 379804 164874 380404 164876
rect 415804 164874 416404 164876
rect 451804 164874 452404 164876
rect 487804 164874 488404 164876
rect 523804 164874 524404 164876
rect 559804 164874 560404 164876
rect 586260 164874 586860 164876
rect -7636 158276 -7036 158278
rect 12604 158276 13204 158278
rect 48604 158276 49204 158278
rect 84604 158276 85204 158278
rect 120604 158276 121204 158278
rect 156604 158276 157204 158278
rect 192604 158276 193204 158278
rect 228604 158276 229204 158278
rect 264604 158276 265204 158278
rect 300604 158276 301204 158278
rect 336604 158276 337204 158278
rect 372604 158276 373204 158278
rect 408604 158276 409204 158278
rect 444604 158276 445204 158278
rect 480604 158276 481204 158278
rect 516604 158276 517204 158278
rect 552604 158276 553204 158278
rect 590960 158276 591560 158278
rect -8576 158254 592500 158276
rect -8576 158018 -7454 158254
rect -7218 158018 12786 158254
rect 13022 158018 48786 158254
rect 49022 158018 84786 158254
rect 85022 158018 120786 158254
rect 121022 158018 156786 158254
rect 157022 158018 192786 158254
rect 193022 158018 228786 158254
rect 229022 158018 264786 158254
rect 265022 158018 300786 158254
rect 301022 158018 336786 158254
rect 337022 158018 372786 158254
rect 373022 158018 408786 158254
rect 409022 158018 444786 158254
rect 445022 158018 480786 158254
rect 481022 158018 516786 158254
rect 517022 158018 552786 158254
rect 553022 158018 591142 158254
rect 591378 158018 592500 158254
rect -8576 157934 592500 158018
rect -8576 157698 -7454 157934
rect -7218 157698 12786 157934
rect 13022 157698 48786 157934
rect 49022 157698 84786 157934
rect 85022 157698 120786 157934
rect 121022 157698 156786 157934
rect 157022 157698 192786 157934
rect 193022 157698 228786 157934
rect 229022 157698 264786 157934
rect 265022 157698 300786 157934
rect 301022 157698 336786 157934
rect 337022 157698 372786 157934
rect 373022 157698 408786 157934
rect 409022 157698 444786 157934
rect 445022 157698 480786 157934
rect 481022 157698 516786 157934
rect 517022 157698 552786 157934
rect 553022 157698 591142 157934
rect 591378 157698 592500 157934
rect -8576 157676 592500 157698
rect -7636 157674 -7036 157676
rect 12604 157674 13204 157676
rect 48604 157674 49204 157676
rect 84604 157674 85204 157676
rect 120604 157674 121204 157676
rect 156604 157674 157204 157676
rect 192604 157674 193204 157676
rect 228604 157674 229204 157676
rect 264604 157674 265204 157676
rect 300604 157674 301204 157676
rect 336604 157674 337204 157676
rect 372604 157674 373204 157676
rect 408604 157674 409204 157676
rect 444604 157674 445204 157676
rect 480604 157674 481204 157676
rect 516604 157674 517204 157676
rect 552604 157674 553204 157676
rect 590960 157674 591560 157676
rect -5756 154676 -5156 154678
rect 9004 154676 9604 154678
rect 45004 154676 45604 154678
rect 81004 154676 81604 154678
rect 117004 154676 117604 154678
rect 153004 154676 153604 154678
rect 189004 154676 189604 154678
rect 225004 154676 225604 154678
rect 261004 154676 261604 154678
rect 297004 154676 297604 154678
rect 333004 154676 333604 154678
rect 369004 154676 369604 154678
rect 405004 154676 405604 154678
rect 441004 154676 441604 154678
rect 477004 154676 477604 154678
rect 513004 154676 513604 154678
rect 549004 154676 549604 154678
rect 589080 154676 589680 154678
rect -6696 154654 590620 154676
rect -6696 154418 -5574 154654
rect -5338 154418 9186 154654
rect 9422 154418 45186 154654
rect 45422 154418 81186 154654
rect 81422 154418 117186 154654
rect 117422 154418 153186 154654
rect 153422 154418 189186 154654
rect 189422 154418 225186 154654
rect 225422 154418 261186 154654
rect 261422 154418 297186 154654
rect 297422 154418 333186 154654
rect 333422 154418 369186 154654
rect 369422 154418 405186 154654
rect 405422 154418 441186 154654
rect 441422 154418 477186 154654
rect 477422 154418 513186 154654
rect 513422 154418 549186 154654
rect 549422 154418 589262 154654
rect 589498 154418 590620 154654
rect -6696 154334 590620 154418
rect -6696 154098 -5574 154334
rect -5338 154098 9186 154334
rect 9422 154098 45186 154334
rect 45422 154098 81186 154334
rect 81422 154098 117186 154334
rect 117422 154098 153186 154334
rect 153422 154098 189186 154334
rect 189422 154098 225186 154334
rect 225422 154098 261186 154334
rect 261422 154098 297186 154334
rect 297422 154098 333186 154334
rect 333422 154098 369186 154334
rect 369422 154098 405186 154334
rect 405422 154098 441186 154334
rect 441422 154098 477186 154334
rect 477422 154098 513186 154334
rect 513422 154098 549186 154334
rect 549422 154098 589262 154334
rect 589498 154098 590620 154334
rect -6696 154076 590620 154098
rect -5756 154074 -5156 154076
rect 9004 154074 9604 154076
rect 45004 154074 45604 154076
rect 81004 154074 81604 154076
rect 117004 154074 117604 154076
rect 153004 154074 153604 154076
rect 189004 154074 189604 154076
rect 225004 154074 225604 154076
rect 261004 154074 261604 154076
rect 297004 154074 297604 154076
rect 333004 154074 333604 154076
rect 369004 154074 369604 154076
rect 405004 154074 405604 154076
rect 441004 154074 441604 154076
rect 477004 154074 477604 154076
rect 513004 154074 513604 154076
rect 549004 154074 549604 154076
rect 589080 154074 589680 154076
rect -3876 151076 -3276 151078
rect 5404 151076 6004 151078
rect 41404 151076 42004 151078
rect 77404 151076 78004 151078
rect 113404 151076 114004 151078
rect 149404 151076 150004 151078
rect 185404 151076 186004 151078
rect 221404 151076 222004 151078
rect 257404 151076 258004 151078
rect 293404 151076 294004 151078
rect 329404 151076 330004 151078
rect 365404 151076 366004 151078
rect 401404 151076 402004 151078
rect 437404 151076 438004 151078
rect 473404 151076 474004 151078
rect 509404 151076 510004 151078
rect 545404 151076 546004 151078
rect 581404 151076 582004 151078
rect 587200 151076 587800 151078
rect -4816 151054 588740 151076
rect -4816 150818 -3694 151054
rect -3458 150818 5586 151054
rect 5822 150818 41586 151054
rect 41822 150818 77586 151054
rect 77822 150818 113586 151054
rect 113822 150818 149586 151054
rect 149822 150818 185586 151054
rect 185822 150818 221586 151054
rect 221822 150818 257586 151054
rect 257822 150818 293586 151054
rect 293822 150818 329586 151054
rect 329822 150818 365586 151054
rect 365822 150818 401586 151054
rect 401822 150818 437586 151054
rect 437822 150818 473586 151054
rect 473822 150818 509586 151054
rect 509822 150818 545586 151054
rect 545822 150818 581586 151054
rect 581822 150818 587382 151054
rect 587618 150818 588740 151054
rect -4816 150734 588740 150818
rect -4816 150498 -3694 150734
rect -3458 150498 5586 150734
rect 5822 150498 41586 150734
rect 41822 150498 77586 150734
rect 77822 150498 113586 150734
rect 113822 150498 149586 150734
rect 149822 150498 185586 150734
rect 185822 150498 221586 150734
rect 221822 150498 257586 150734
rect 257822 150498 293586 150734
rect 293822 150498 329586 150734
rect 329822 150498 365586 150734
rect 365822 150498 401586 150734
rect 401822 150498 437586 150734
rect 437822 150498 473586 150734
rect 473822 150498 509586 150734
rect 509822 150498 545586 150734
rect 545822 150498 581586 150734
rect 581822 150498 587382 150734
rect 587618 150498 588740 150734
rect -4816 150476 588740 150498
rect -3876 150474 -3276 150476
rect 5404 150474 6004 150476
rect 41404 150474 42004 150476
rect 77404 150474 78004 150476
rect 113404 150474 114004 150476
rect 149404 150474 150004 150476
rect 185404 150474 186004 150476
rect 221404 150474 222004 150476
rect 257404 150474 258004 150476
rect 293404 150474 294004 150476
rect 329404 150474 330004 150476
rect 365404 150474 366004 150476
rect 401404 150474 402004 150476
rect 437404 150474 438004 150476
rect 473404 150474 474004 150476
rect 509404 150474 510004 150476
rect 545404 150474 546004 150476
rect 581404 150474 582004 150476
rect 587200 150474 587800 150476
rect -1996 147476 -1396 147478
rect 1804 147476 2404 147478
rect 37804 147476 38404 147478
rect 73804 147476 74404 147478
rect 109804 147476 110404 147478
rect 145804 147476 146404 147478
rect 181804 147476 182404 147478
rect 217804 147476 218404 147478
rect 253804 147476 254404 147478
rect 289804 147476 290404 147478
rect 325804 147476 326404 147478
rect 361804 147476 362404 147478
rect 397804 147476 398404 147478
rect 433804 147476 434404 147478
rect 469804 147476 470404 147478
rect 505804 147476 506404 147478
rect 541804 147476 542404 147478
rect 577804 147476 578404 147478
rect 585320 147476 585920 147478
rect -2936 147454 586860 147476
rect -2936 147218 -1814 147454
rect -1578 147218 1986 147454
rect 2222 147218 37986 147454
rect 38222 147218 73986 147454
rect 74222 147218 109986 147454
rect 110222 147218 145986 147454
rect 146222 147218 181986 147454
rect 182222 147218 217986 147454
rect 218222 147218 253986 147454
rect 254222 147218 289986 147454
rect 290222 147218 325986 147454
rect 326222 147218 361986 147454
rect 362222 147218 397986 147454
rect 398222 147218 433986 147454
rect 434222 147218 469986 147454
rect 470222 147218 505986 147454
rect 506222 147218 541986 147454
rect 542222 147218 577986 147454
rect 578222 147218 585502 147454
rect 585738 147218 586860 147454
rect -2936 147134 586860 147218
rect -2936 146898 -1814 147134
rect -1578 146898 1986 147134
rect 2222 146898 37986 147134
rect 38222 146898 73986 147134
rect 74222 146898 109986 147134
rect 110222 146898 145986 147134
rect 146222 146898 181986 147134
rect 182222 146898 217986 147134
rect 218222 146898 253986 147134
rect 254222 146898 289986 147134
rect 290222 146898 325986 147134
rect 326222 146898 361986 147134
rect 362222 146898 397986 147134
rect 398222 146898 433986 147134
rect 434222 146898 469986 147134
rect 470222 146898 505986 147134
rect 506222 146898 541986 147134
rect 542222 146898 577986 147134
rect 578222 146898 585502 147134
rect 585738 146898 586860 147134
rect -2936 146876 586860 146898
rect -1996 146874 -1396 146876
rect 1804 146874 2404 146876
rect 37804 146874 38404 146876
rect 73804 146874 74404 146876
rect 109804 146874 110404 146876
rect 145804 146874 146404 146876
rect 181804 146874 182404 146876
rect 217804 146874 218404 146876
rect 253804 146874 254404 146876
rect 289804 146874 290404 146876
rect 325804 146874 326404 146876
rect 361804 146874 362404 146876
rect 397804 146874 398404 146876
rect 433804 146874 434404 146876
rect 469804 146874 470404 146876
rect 505804 146874 506404 146876
rect 541804 146874 542404 146876
rect 577804 146874 578404 146876
rect 585320 146874 585920 146876
rect -8576 140276 -7976 140278
rect 30604 140276 31204 140278
rect 66604 140276 67204 140278
rect 102604 140276 103204 140278
rect 138604 140276 139204 140278
rect 174604 140276 175204 140278
rect 210604 140276 211204 140278
rect 246604 140276 247204 140278
rect 282604 140276 283204 140278
rect 318604 140276 319204 140278
rect 354604 140276 355204 140278
rect 390604 140276 391204 140278
rect 426604 140276 427204 140278
rect 462604 140276 463204 140278
rect 498604 140276 499204 140278
rect 534604 140276 535204 140278
rect 570604 140276 571204 140278
rect 591900 140276 592500 140278
rect -8576 140254 592500 140276
rect -8576 140018 -8394 140254
rect -8158 140018 30786 140254
rect 31022 140018 66786 140254
rect 67022 140018 102786 140254
rect 103022 140018 138786 140254
rect 139022 140018 174786 140254
rect 175022 140018 210786 140254
rect 211022 140018 246786 140254
rect 247022 140018 282786 140254
rect 283022 140018 318786 140254
rect 319022 140018 354786 140254
rect 355022 140018 390786 140254
rect 391022 140018 426786 140254
rect 427022 140018 462786 140254
rect 463022 140018 498786 140254
rect 499022 140018 534786 140254
rect 535022 140018 570786 140254
rect 571022 140018 592082 140254
rect 592318 140018 592500 140254
rect -8576 139934 592500 140018
rect -8576 139698 -8394 139934
rect -8158 139698 30786 139934
rect 31022 139698 66786 139934
rect 67022 139698 102786 139934
rect 103022 139698 138786 139934
rect 139022 139698 174786 139934
rect 175022 139698 210786 139934
rect 211022 139698 246786 139934
rect 247022 139698 282786 139934
rect 283022 139698 318786 139934
rect 319022 139698 354786 139934
rect 355022 139698 390786 139934
rect 391022 139698 426786 139934
rect 427022 139698 462786 139934
rect 463022 139698 498786 139934
rect 499022 139698 534786 139934
rect 535022 139698 570786 139934
rect 571022 139698 592082 139934
rect 592318 139698 592500 139934
rect -8576 139676 592500 139698
rect -8576 139674 -7976 139676
rect 30604 139674 31204 139676
rect 66604 139674 67204 139676
rect 102604 139674 103204 139676
rect 138604 139674 139204 139676
rect 174604 139674 175204 139676
rect 210604 139674 211204 139676
rect 246604 139674 247204 139676
rect 282604 139674 283204 139676
rect 318604 139674 319204 139676
rect 354604 139674 355204 139676
rect 390604 139674 391204 139676
rect 426604 139674 427204 139676
rect 462604 139674 463204 139676
rect 498604 139674 499204 139676
rect 534604 139674 535204 139676
rect 570604 139674 571204 139676
rect 591900 139674 592500 139676
rect -6696 136676 -6096 136678
rect 27004 136676 27604 136678
rect 63004 136676 63604 136678
rect 99004 136676 99604 136678
rect 135004 136676 135604 136678
rect 171004 136676 171604 136678
rect 207004 136676 207604 136678
rect 243004 136676 243604 136678
rect 279004 136676 279604 136678
rect 315004 136676 315604 136678
rect 351004 136676 351604 136678
rect 387004 136676 387604 136678
rect 423004 136676 423604 136678
rect 459004 136676 459604 136678
rect 495004 136676 495604 136678
rect 531004 136676 531604 136678
rect 567004 136676 567604 136678
rect 590020 136676 590620 136678
rect -6696 136654 590620 136676
rect -6696 136418 -6514 136654
rect -6278 136418 27186 136654
rect 27422 136418 63186 136654
rect 63422 136418 99186 136654
rect 99422 136418 135186 136654
rect 135422 136418 171186 136654
rect 171422 136418 207186 136654
rect 207422 136418 243186 136654
rect 243422 136418 279186 136654
rect 279422 136418 315186 136654
rect 315422 136418 351186 136654
rect 351422 136418 387186 136654
rect 387422 136418 423186 136654
rect 423422 136418 459186 136654
rect 459422 136418 495186 136654
rect 495422 136418 531186 136654
rect 531422 136418 567186 136654
rect 567422 136418 590202 136654
rect 590438 136418 590620 136654
rect -6696 136334 590620 136418
rect -6696 136098 -6514 136334
rect -6278 136098 27186 136334
rect 27422 136098 63186 136334
rect 63422 136098 99186 136334
rect 99422 136098 135186 136334
rect 135422 136098 171186 136334
rect 171422 136098 207186 136334
rect 207422 136098 243186 136334
rect 243422 136098 279186 136334
rect 279422 136098 315186 136334
rect 315422 136098 351186 136334
rect 351422 136098 387186 136334
rect 387422 136098 423186 136334
rect 423422 136098 459186 136334
rect 459422 136098 495186 136334
rect 495422 136098 531186 136334
rect 531422 136098 567186 136334
rect 567422 136098 590202 136334
rect 590438 136098 590620 136334
rect -6696 136076 590620 136098
rect -6696 136074 -6096 136076
rect 27004 136074 27604 136076
rect 63004 136074 63604 136076
rect 99004 136074 99604 136076
rect 135004 136074 135604 136076
rect 171004 136074 171604 136076
rect 207004 136074 207604 136076
rect 243004 136074 243604 136076
rect 279004 136074 279604 136076
rect 315004 136074 315604 136076
rect 351004 136074 351604 136076
rect 387004 136074 387604 136076
rect 423004 136074 423604 136076
rect 459004 136074 459604 136076
rect 495004 136074 495604 136076
rect 531004 136074 531604 136076
rect 567004 136074 567604 136076
rect 590020 136074 590620 136076
rect -4816 133076 -4216 133078
rect 23404 133076 24004 133078
rect 59404 133076 60004 133078
rect 95404 133076 96004 133078
rect 131404 133076 132004 133078
rect 167404 133076 168004 133078
rect 203404 133076 204004 133078
rect 239404 133076 240004 133078
rect 275404 133076 276004 133078
rect 311404 133076 312004 133078
rect 347404 133076 348004 133078
rect 383404 133076 384004 133078
rect 419404 133076 420004 133078
rect 455404 133076 456004 133078
rect 491404 133076 492004 133078
rect 527404 133076 528004 133078
rect 563404 133076 564004 133078
rect 588140 133076 588740 133078
rect -4816 133054 588740 133076
rect -4816 132818 -4634 133054
rect -4398 132818 23586 133054
rect 23822 132818 59586 133054
rect 59822 132818 95586 133054
rect 95822 132818 131586 133054
rect 131822 132818 167586 133054
rect 167822 132818 203586 133054
rect 203822 132818 239586 133054
rect 239822 132818 275586 133054
rect 275822 132818 311586 133054
rect 311822 132818 347586 133054
rect 347822 132818 383586 133054
rect 383822 132818 419586 133054
rect 419822 132818 455586 133054
rect 455822 132818 491586 133054
rect 491822 132818 527586 133054
rect 527822 132818 563586 133054
rect 563822 132818 588322 133054
rect 588558 132818 588740 133054
rect -4816 132734 588740 132818
rect -4816 132498 -4634 132734
rect -4398 132498 23586 132734
rect 23822 132498 59586 132734
rect 59822 132498 95586 132734
rect 95822 132498 131586 132734
rect 131822 132498 167586 132734
rect 167822 132498 203586 132734
rect 203822 132498 239586 132734
rect 239822 132498 275586 132734
rect 275822 132498 311586 132734
rect 311822 132498 347586 132734
rect 347822 132498 383586 132734
rect 383822 132498 419586 132734
rect 419822 132498 455586 132734
rect 455822 132498 491586 132734
rect 491822 132498 527586 132734
rect 527822 132498 563586 132734
rect 563822 132498 588322 132734
rect 588558 132498 588740 132734
rect -4816 132476 588740 132498
rect -4816 132474 -4216 132476
rect 23404 132474 24004 132476
rect 59404 132474 60004 132476
rect 95404 132474 96004 132476
rect 131404 132474 132004 132476
rect 167404 132474 168004 132476
rect 203404 132474 204004 132476
rect 239404 132474 240004 132476
rect 275404 132474 276004 132476
rect 311404 132474 312004 132476
rect 347404 132474 348004 132476
rect 383404 132474 384004 132476
rect 419404 132474 420004 132476
rect 455404 132474 456004 132476
rect 491404 132474 492004 132476
rect 527404 132474 528004 132476
rect 563404 132474 564004 132476
rect 588140 132474 588740 132476
rect -2936 129476 -2336 129478
rect 19804 129476 20404 129478
rect 55804 129476 56404 129478
rect 91804 129476 92404 129478
rect 127804 129476 128404 129478
rect 163804 129476 164404 129478
rect 199804 129476 200404 129478
rect 235804 129476 236404 129478
rect 271804 129476 272404 129478
rect 307804 129476 308404 129478
rect 343804 129476 344404 129478
rect 379804 129476 380404 129478
rect 415804 129476 416404 129478
rect 451804 129476 452404 129478
rect 487804 129476 488404 129478
rect 523804 129476 524404 129478
rect 559804 129476 560404 129478
rect 586260 129476 586860 129478
rect -2936 129454 586860 129476
rect -2936 129218 -2754 129454
rect -2518 129218 19986 129454
rect 20222 129218 55986 129454
rect 56222 129218 91986 129454
rect 92222 129218 127986 129454
rect 128222 129218 163986 129454
rect 164222 129218 199986 129454
rect 200222 129218 235986 129454
rect 236222 129218 271986 129454
rect 272222 129218 307986 129454
rect 308222 129218 343986 129454
rect 344222 129218 379986 129454
rect 380222 129218 415986 129454
rect 416222 129218 451986 129454
rect 452222 129218 487986 129454
rect 488222 129218 523986 129454
rect 524222 129218 559986 129454
rect 560222 129218 586442 129454
rect 586678 129218 586860 129454
rect -2936 129134 586860 129218
rect -2936 128898 -2754 129134
rect -2518 128898 19986 129134
rect 20222 128898 55986 129134
rect 56222 128898 91986 129134
rect 92222 128898 127986 129134
rect 128222 128898 163986 129134
rect 164222 128898 199986 129134
rect 200222 128898 235986 129134
rect 236222 128898 271986 129134
rect 272222 128898 307986 129134
rect 308222 128898 343986 129134
rect 344222 128898 379986 129134
rect 380222 128898 415986 129134
rect 416222 128898 451986 129134
rect 452222 128898 487986 129134
rect 488222 128898 523986 129134
rect 524222 128898 559986 129134
rect 560222 128898 586442 129134
rect 586678 128898 586860 129134
rect -2936 128876 586860 128898
rect -2936 128874 -2336 128876
rect 19804 128874 20404 128876
rect 55804 128874 56404 128876
rect 91804 128874 92404 128876
rect 127804 128874 128404 128876
rect 163804 128874 164404 128876
rect 199804 128874 200404 128876
rect 235804 128874 236404 128876
rect 271804 128874 272404 128876
rect 307804 128874 308404 128876
rect 343804 128874 344404 128876
rect 379804 128874 380404 128876
rect 415804 128874 416404 128876
rect 451804 128874 452404 128876
rect 487804 128874 488404 128876
rect 523804 128874 524404 128876
rect 559804 128874 560404 128876
rect 586260 128874 586860 128876
rect -7636 122276 -7036 122278
rect 12604 122276 13204 122278
rect 48604 122276 49204 122278
rect 84604 122276 85204 122278
rect 120604 122276 121204 122278
rect 156604 122276 157204 122278
rect 192604 122276 193204 122278
rect 228604 122276 229204 122278
rect 264604 122276 265204 122278
rect 300604 122276 301204 122278
rect 336604 122276 337204 122278
rect 372604 122276 373204 122278
rect 408604 122276 409204 122278
rect 444604 122276 445204 122278
rect 480604 122276 481204 122278
rect 516604 122276 517204 122278
rect 552604 122276 553204 122278
rect 590960 122276 591560 122278
rect -8576 122254 592500 122276
rect -8576 122018 -7454 122254
rect -7218 122018 12786 122254
rect 13022 122018 48786 122254
rect 49022 122018 84786 122254
rect 85022 122018 120786 122254
rect 121022 122018 156786 122254
rect 157022 122018 192786 122254
rect 193022 122018 228786 122254
rect 229022 122018 264786 122254
rect 265022 122018 300786 122254
rect 301022 122018 336786 122254
rect 337022 122018 372786 122254
rect 373022 122018 408786 122254
rect 409022 122018 444786 122254
rect 445022 122018 480786 122254
rect 481022 122018 516786 122254
rect 517022 122018 552786 122254
rect 553022 122018 591142 122254
rect 591378 122018 592500 122254
rect -8576 121934 592500 122018
rect -8576 121698 -7454 121934
rect -7218 121698 12786 121934
rect 13022 121698 48786 121934
rect 49022 121698 84786 121934
rect 85022 121698 120786 121934
rect 121022 121698 156786 121934
rect 157022 121698 192786 121934
rect 193022 121698 228786 121934
rect 229022 121698 264786 121934
rect 265022 121698 300786 121934
rect 301022 121698 336786 121934
rect 337022 121698 372786 121934
rect 373022 121698 408786 121934
rect 409022 121698 444786 121934
rect 445022 121698 480786 121934
rect 481022 121698 516786 121934
rect 517022 121698 552786 121934
rect 553022 121698 591142 121934
rect 591378 121698 592500 121934
rect -8576 121676 592500 121698
rect -7636 121674 -7036 121676
rect 12604 121674 13204 121676
rect 48604 121674 49204 121676
rect 84604 121674 85204 121676
rect 120604 121674 121204 121676
rect 156604 121674 157204 121676
rect 192604 121674 193204 121676
rect 228604 121674 229204 121676
rect 264604 121674 265204 121676
rect 300604 121674 301204 121676
rect 336604 121674 337204 121676
rect 372604 121674 373204 121676
rect 408604 121674 409204 121676
rect 444604 121674 445204 121676
rect 480604 121674 481204 121676
rect 516604 121674 517204 121676
rect 552604 121674 553204 121676
rect 590960 121674 591560 121676
rect -5756 118676 -5156 118678
rect 9004 118676 9604 118678
rect 45004 118676 45604 118678
rect 81004 118676 81604 118678
rect 117004 118676 117604 118678
rect 153004 118676 153604 118678
rect 189004 118676 189604 118678
rect 225004 118676 225604 118678
rect 261004 118676 261604 118678
rect 297004 118676 297604 118678
rect 333004 118676 333604 118678
rect 369004 118676 369604 118678
rect 405004 118676 405604 118678
rect 441004 118676 441604 118678
rect 477004 118676 477604 118678
rect 513004 118676 513604 118678
rect 549004 118676 549604 118678
rect 589080 118676 589680 118678
rect -6696 118654 590620 118676
rect -6696 118418 -5574 118654
rect -5338 118418 9186 118654
rect 9422 118418 45186 118654
rect 45422 118418 81186 118654
rect 81422 118418 117186 118654
rect 117422 118418 153186 118654
rect 153422 118418 189186 118654
rect 189422 118418 225186 118654
rect 225422 118418 261186 118654
rect 261422 118418 297186 118654
rect 297422 118418 333186 118654
rect 333422 118418 369186 118654
rect 369422 118418 405186 118654
rect 405422 118418 441186 118654
rect 441422 118418 477186 118654
rect 477422 118418 513186 118654
rect 513422 118418 549186 118654
rect 549422 118418 589262 118654
rect 589498 118418 590620 118654
rect -6696 118334 590620 118418
rect -6696 118098 -5574 118334
rect -5338 118098 9186 118334
rect 9422 118098 45186 118334
rect 45422 118098 81186 118334
rect 81422 118098 117186 118334
rect 117422 118098 153186 118334
rect 153422 118098 189186 118334
rect 189422 118098 225186 118334
rect 225422 118098 261186 118334
rect 261422 118098 297186 118334
rect 297422 118098 333186 118334
rect 333422 118098 369186 118334
rect 369422 118098 405186 118334
rect 405422 118098 441186 118334
rect 441422 118098 477186 118334
rect 477422 118098 513186 118334
rect 513422 118098 549186 118334
rect 549422 118098 589262 118334
rect 589498 118098 590620 118334
rect -6696 118076 590620 118098
rect -5756 118074 -5156 118076
rect 9004 118074 9604 118076
rect 45004 118074 45604 118076
rect 81004 118074 81604 118076
rect 117004 118074 117604 118076
rect 153004 118074 153604 118076
rect 189004 118074 189604 118076
rect 225004 118074 225604 118076
rect 261004 118074 261604 118076
rect 297004 118074 297604 118076
rect 333004 118074 333604 118076
rect 369004 118074 369604 118076
rect 405004 118074 405604 118076
rect 441004 118074 441604 118076
rect 477004 118074 477604 118076
rect 513004 118074 513604 118076
rect 549004 118074 549604 118076
rect 589080 118074 589680 118076
rect -3876 115076 -3276 115078
rect 5404 115076 6004 115078
rect 41404 115076 42004 115078
rect 77404 115076 78004 115078
rect 113404 115076 114004 115078
rect 149404 115076 150004 115078
rect 185404 115076 186004 115078
rect 221404 115076 222004 115078
rect 257404 115076 258004 115078
rect 293404 115076 294004 115078
rect 329404 115076 330004 115078
rect 365404 115076 366004 115078
rect 401404 115076 402004 115078
rect 437404 115076 438004 115078
rect 473404 115076 474004 115078
rect 509404 115076 510004 115078
rect 545404 115076 546004 115078
rect 581404 115076 582004 115078
rect 587200 115076 587800 115078
rect -4816 115054 588740 115076
rect -4816 114818 -3694 115054
rect -3458 114818 5586 115054
rect 5822 114818 41586 115054
rect 41822 114818 77586 115054
rect 77822 114818 113586 115054
rect 113822 114818 149586 115054
rect 149822 114818 185586 115054
rect 185822 114818 221586 115054
rect 221822 114818 257586 115054
rect 257822 114818 293586 115054
rect 293822 114818 329586 115054
rect 329822 114818 365586 115054
rect 365822 114818 401586 115054
rect 401822 114818 437586 115054
rect 437822 114818 473586 115054
rect 473822 114818 509586 115054
rect 509822 114818 545586 115054
rect 545822 114818 581586 115054
rect 581822 114818 587382 115054
rect 587618 114818 588740 115054
rect -4816 114734 588740 114818
rect -4816 114498 -3694 114734
rect -3458 114498 5586 114734
rect 5822 114498 41586 114734
rect 41822 114498 77586 114734
rect 77822 114498 113586 114734
rect 113822 114498 149586 114734
rect 149822 114498 185586 114734
rect 185822 114498 221586 114734
rect 221822 114498 257586 114734
rect 257822 114498 293586 114734
rect 293822 114498 329586 114734
rect 329822 114498 365586 114734
rect 365822 114498 401586 114734
rect 401822 114498 437586 114734
rect 437822 114498 473586 114734
rect 473822 114498 509586 114734
rect 509822 114498 545586 114734
rect 545822 114498 581586 114734
rect 581822 114498 587382 114734
rect 587618 114498 588740 114734
rect -4816 114476 588740 114498
rect -3876 114474 -3276 114476
rect 5404 114474 6004 114476
rect 41404 114474 42004 114476
rect 77404 114474 78004 114476
rect 113404 114474 114004 114476
rect 149404 114474 150004 114476
rect 185404 114474 186004 114476
rect 221404 114474 222004 114476
rect 257404 114474 258004 114476
rect 293404 114474 294004 114476
rect 329404 114474 330004 114476
rect 365404 114474 366004 114476
rect 401404 114474 402004 114476
rect 437404 114474 438004 114476
rect 473404 114474 474004 114476
rect 509404 114474 510004 114476
rect 545404 114474 546004 114476
rect 581404 114474 582004 114476
rect 587200 114474 587800 114476
rect -1996 111476 -1396 111478
rect 1804 111476 2404 111478
rect 37804 111476 38404 111478
rect 73804 111476 74404 111478
rect 109804 111476 110404 111478
rect 145804 111476 146404 111478
rect 181804 111476 182404 111478
rect 217804 111476 218404 111478
rect 253804 111476 254404 111478
rect 289804 111476 290404 111478
rect 325804 111476 326404 111478
rect 361804 111476 362404 111478
rect 397804 111476 398404 111478
rect 433804 111476 434404 111478
rect 469804 111476 470404 111478
rect 505804 111476 506404 111478
rect 541804 111476 542404 111478
rect 577804 111476 578404 111478
rect 585320 111476 585920 111478
rect -2936 111454 586860 111476
rect -2936 111218 -1814 111454
rect -1578 111218 1986 111454
rect 2222 111218 37986 111454
rect 38222 111218 73986 111454
rect 74222 111218 109986 111454
rect 110222 111218 145986 111454
rect 146222 111218 181986 111454
rect 182222 111218 217986 111454
rect 218222 111218 253986 111454
rect 254222 111218 289986 111454
rect 290222 111218 325986 111454
rect 326222 111218 361986 111454
rect 362222 111218 397986 111454
rect 398222 111218 433986 111454
rect 434222 111218 469986 111454
rect 470222 111218 505986 111454
rect 506222 111218 541986 111454
rect 542222 111218 577986 111454
rect 578222 111218 585502 111454
rect 585738 111218 586860 111454
rect -2936 111134 586860 111218
rect -2936 110898 -1814 111134
rect -1578 110898 1986 111134
rect 2222 110898 37986 111134
rect 38222 110898 73986 111134
rect 74222 110898 109986 111134
rect 110222 110898 145986 111134
rect 146222 110898 181986 111134
rect 182222 110898 217986 111134
rect 218222 110898 253986 111134
rect 254222 110898 289986 111134
rect 290222 110898 325986 111134
rect 326222 110898 361986 111134
rect 362222 110898 397986 111134
rect 398222 110898 433986 111134
rect 434222 110898 469986 111134
rect 470222 110898 505986 111134
rect 506222 110898 541986 111134
rect 542222 110898 577986 111134
rect 578222 110898 585502 111134
rect 585738 110898 586860 111134
rect -2936 110876 586860 110898
rect -1996 110874 -1396 110876
rect 1804 110874 2404 110876
rect 37804 110874 38404 110876
rect 73804 110874 74404 110876
rect 109804 110874 110404 110876
rect 145804 110874 146404 110876
rect 181804 110874 182404 110876
rect 217804 110874 218404 110876
rect 253804 110874 254404 110876
rect 289804 110874 290404 110876
rect 325804 110874 326404 110876
rect 361804 110874 362404 110876
rect 397804 110874 398404 110876
rect 433804 110874 434404 110876
rect 469804 110874 470404 110876
rect 505804 110874 506404 110876
rect 541804 110874 542404 110876
rect 577804 110874 578404 110876
rect 585320 110874 585920 110876
rect -8576 104276 -7976 104278
rect 30604 104276 31204 104278
rect 66604 104276 67204 104278
rect 102604 104276 103204 104278
rect 138604 104276 139204 104278
rect 174604 104276 175204 104278
rect 210604 104276 211204 104278
rect 246604 104276 247204 104278
rect 282604 104276 283204 104278
rect 318604 104276 319204 104278
rect 354604 104276 355204 104278
rect 390604 104276 391204 104278
rect 426604 104276 427204 104278
rect 462604 104276 463204 104278
rect 498604 104276 499204 104278
rect 534604 104276 535204 104278
rect 570604 104276 571204 104278
rect 591900 104276 592500 104278
rect -8576 104254 592500 104276
rect -8576 104018 -8394 104254
rect -8158 104018 30786 104254
rect 31022 104018 66786 104254
rect 67022 104018 102786 104254
rect 103022 104018 138786 104254
rect 139022 104018 174786 104254
rect 175022 104018 210786 104254
rect 211022 104018 246786 104254
rect 247022 104018 282786 104254
rect 283022 104018 318786 104254
rect 319022 104018 354786 104254
rect 355022 104018 390786 104254
rect 391022 104018 426786 104254
rect 427022 104018 462786 104254
rect 463022 104018 498786 104254
rect 499022 104018 534786 104254
rect 535022 104018 570786 104254
rect 571022 104018 592082 104254
rect 592318 104018 592500 104254
rect -8576 103934 592500 104018
rect -8576 103698 -8394 103934
rect -8158 103698 30786 103934
rect 31022 103698 66786 103934
rect 67022 103698 102786 103934
rect 103022 103698 138786 103934
rect 139022 103698 174786 103934
rect 175022 103698 210786 103934
rect 211022 103698 246786 103934
rect 247022 103698 282786 103934
rect 283022 103698 318786 103934
rect 319022 103698 354786 103934
rect 355022 103698 390786 103934
rect 391022 103698 426786 103934
rect 427022 103698 462786 103934
rect 463022 103698 498786 103934
rect 499022 103698 534786 103934
rect 535022 103698 570786 103934
rect 571022 103698 592082 103934
rect 592318 103698 592500 103934
rect -8576 103676 592500 103698
rect -8576 103674 -7976 103676
rect 30604 103674 31204 103676
rect 66604 103674 67204 103676
rect 102604 103674 103204 103676
rect 138604 103674 139204 103676
rect 174604 103674 175204 103676
rect 210604 103674 211204 103676
rect 246604 103674 247204 103676
rect 282604 103674 283204 103676
rect 318604 103674 319204 103676
rect 354604 103674 355204 103676
rect 390604 103674 391204 103676
rect 426604 103674 427204 103676
rect 462604 103674 463204 103676
rect 498604 103674 499204 103676
rect 534604 103674 535204 103676
rect 570604 103674 571204 103676
rect 591900 103674 592500 103676
rect -6696 100676 -6096 100678
rect 27004 100676 27604 100678
rect 63004 100676 63604 100678
rect 99004 100676 99604 100678
rect 135004 100676 135604 100678
rect 171004 100676 171604 100678
rect 207004 100676 207604 100678
rect 243004 100676 243604 100678
rect 279004 100676 279604 100678
rect 315004 100676 315604 100678
rect 351004 100676 351604 100678
rect 387004 100676 387604 100678
rect 423004 100676 423604 100678
rect 459004 100676 459604 100678
rect 495004 100676 495604 100678
rect 531004 100676 531604 100678
rect 567004 100676 567604 100678
rect 590020 100676 590620 100678
rect -6696 100654 590620 100676
rect -6696 100418 -6514 100654
rect -6278 100418 27186 100654
rect 27422 100418 63186 100654
rect 63422 100418 99186 100654
rect 99422 100418 135186 100654
rect 135422 100418 171186 100654
rect 171422 100418 207186 100654
rect 207422 100418 243186 100654
rect 243422 100418 279186 100654
rect 279422 100418 315186 100654
rect 315422 100418 351186 100654
rect 351422 100418 387186 100654
rect 387422 100418 423186 100654
rect 423422 100418 459186 100654
rect 459422 100418 495186 100654
rect 495422 100418 531186 100654
rect 531422 100418 567186 100654
rect 567422 100418 590202 100654
rect 590438 100418 590620 100654
rect -6696 100334 590620 100418
rect -6696 100098 -6514 100334
rect -6278 100098 27186 100334
rect 27422 100098 63186 100334
rect 63422 100098 99186 100334
rect 99422 100098 135186 100334
rect 135422 100098 171186 100334
rect 171422 100098 207186 100334
rect 207422 100098 243186 100334
rect 243422 100098 279186 100334
rect 279422 100098 315186 100334
rect 315422 100098 351186 100334
rect 351422 100098 387186 100334
rect 387422 100098 423186 100334
rect 423422 100098 459186 100334
rect 459422 100098 495186 100334
rect 495422 100098 531186 100334
rect 531422 100098 567186 100334
rect 567422 100098 590202 100334
rect 590438 100098 590620 100334
rect -6696 100076 590620 100098
rect -6696 100074 -6096 100076
rect 27004 100074 27604 100076
rect 63004 100074 63604 100076
rect 99004 100074 99604 100076
rect 135004 100074 135604 100076
rect 171004 100074 171604 100076
rect 207004 100074 207604 100076
rect 243004 100074 243604 100076
rect 279004 100074 279604 100076
rect 315004 100074 315604 100076
rect 351004 100074 351604 100076
rect 387004 100074 387604 100076
rect 423004 100074 423604 100076
rect 459004 100074 459604 100076
rect 495004 100074 495604 100076
rect 531004 100074 531604 100076
rect 567004 100074 567604 100076
rect 590020 100074 590620 100076
rect -4816 97076 -4216 97078
rect 23404 97076 24004 97078
rect 59404 97076 60004 97078
rect 95404 97076 96004 97078
rect 131404 97076 132004 97078
rect 167404 97076 168004 97078
rect 203404 97076 204004 97078
rect 239404 97076 240004 97078
rect 275404 97076 276004 97078
rect 311404 97076 312004 97078
rect 347404 97076 348004 97078
rect 383404 97076 384004 97078
rect 419404 97076 420004 97078
rect 455404 97076 456004 97078
rect 491404 97076 492004 97078
rect 527404 97076 528004 97078
rect 563404 97076 564004 97078
rect 588140 97076 588740 97078
rect -4816 97054 588740 97076
rect -4816 96818 -4634 97054
rect -4398 96818 23586 97054
rect 23822 96818 59586 97054
rect 59822 96818 95586 97054
rect 95822 96818 131586 97054
rect 131822 96818 167586 97054
rect 167822 96818 203586 97054
rect 203822 96818 239586 97054
rect 239822 96818 275586 97054
rect 275822 96818 311586 97054
rect 311822 96818 347586 97054
rect 347822 96818 383586 97054
rect 383822 96818 419586 97054
rect 419822 96818 455586 97054
rect 455822 96818 491586 97054
rect 491822 96818 527586 97054
rect 527822 96818 563586 97054
rect 563822 96818 588322 97054
rect 588558 96818 588740 97054
rect -4816 96734 588740 96818
rect -4816 96498 -4634 96734
rect -4398 96498 23586 96734
rect 23822 96498 59586 96734
rect 59822 96498 95586 96734
rect 95822 96498 131586 96734
rect 131822 96498 167586 96734
rect 167822 96498 203586 96734
rect 203822 96498 239586 96734
rect 239822 96498 275586 96734
rect 275822 96498 311586 96734
rect 311822 96498 347586 96734
rect 347822 96498 383586 96734
rect 383822 96498 419586 96734
rect 419822 96498 455586 96734
rect 455822 96498 491586 96734
rect 491822 96498 527586 96734
rect 527822 96498 563586 96734
rect 563822 96498 588322 96734
rect 588558 96498 588740 96734
rect -4816 96476 588740 96498
rect -4816 96474 -4216 96476
rect 23404 96474 24004 96476
rect 59404 96474 60004 96476
rect 95404 96474 96004 96476
rect 131404 96474 132004 96476
rect 167404 96474 168004 96476
rect 203404 96474 204004 96476
rect 239404 96474 240004 96476
rect 275404 96474 276004 96476
rect 311404 96474 312004 96476
rect 347404 96474 348004 96476
rect 383404 96474 384004 96476
rect 419404 96474 420004 96476
rect 455404 96474 456004 96476
rect 491404 96474 492004 96476
rect 527404 96474 528004 96476
rect 563404 96474 564004 96476
rect 588140 96474 588740 96476
rect -2936 93476 -2336 93478
rect 19804 93476 20404 93478
rect 55804 93476 56404 93478
rect 91804 93476 92404 93478
rect 127804 93476 128404 93478
rect 163804 93476 164404 93478
rect 199804 93476 200404 93478
rect 235804 93476 236404 93478
rect 271804 93476 272404 93478
rect 307804 93476 308404 93478
rect 343804 93476 344404 93478
rect 379804 93476 380404 93478
rect 415804 93476 416404 93478
rect 451804 93476 452404 93478
rect 487804 93476 488404 93478
rect 523804 93476 524404 93478
rect 559804 93476 560404 93478
rect 586260 93476 586860 93478
rect -2936 93454 586860 93476
rect -2936 93218 -2754 93454
rect -2518 93218 19986 93454
rect 20222 93218 55986 93454
rect 56222 93218 91986 93454
rect 92222 93218 127986 93454
rect 128222 93218 163986 93454
rect 164222 93218 199986 93454
rect 200222 93218 235986 93454
rect 236222 93218 271986 93454
rect 272222 93218 307986 93454
rect 308222 93218 343986 93454
rect 344222 93218 379986 93454
rect 380222 93218 415986 93454
rect 416222 93218 451986 93454
rect 452222 93218 487986 93454
rect 488222 93218 523986 93454
rect 524222 93218 559986 93454
rect 560222 93218 586442 93454
rect 586678 93218 586860 93454
rect -2936 93134 586860 93218
rect -2936 92898 -2754 93134
rect -2518 92898 19986 93134
rect 20222 92898 55986 93134
rect 56222 92898 91986 93134
rect 92222 92898 127986 93134
rect 128222 92898 163986 93134
rect 164222 92898 199986 93134
rect 200222 92898 235986 93134
rect 236222 92898 271986 93134
rect 272222 92898 307986 93134
rect 308222 92898 343986 93134
rect 344222 92898 379986 93134
rect 380222 92898 415986 93134
rect 416222 92898 451986 93134
rect 452222 92898 487986 93134
rect 488222 92898 523986 93134
rect 524222 92898 559986 93134
rect 560222 92898 586442 93134
rect 586678 92898 586860 93134
rect -2936 92876 586860 92898
rect -2936 92874 -2336 92876
rect 19804 92874 20404 92876
rect 55804 92874 56404 92876
rect 91804 92874 92404 92876
rect 127804 92874 128404 92876
rect 163804 92874 164404 92876
rect 199804 92874 200404 92876
rect 235804 92874 236404 92876
rect 271804 92874 272404 92876
rect 307804 92874 308404 92876
rect 343804 92874 344404 92876
rect 379804 92874 380404 92876
rect 415804 92874 416404 92876
rect 451804 92874 452404 92876
rect 487804 92874 488404 92876
rect 523804 92874 524404 92876
rect 559804 92874 560404 92876
rect 586260 92874 586860 92876
rect -7636 86276 -7036 86278
rect 12604 86276 13204 86278
rect 48604 86276 49204 86278
rect 84604 86276 85204 86278
rect 120604 86276 121204 86278
rect 156604 86276 157204 86278
rect 192604 86276 193204 86278
rect 228604 86276 229204 86278
rect 264604 86276 265204 86278
rect 300604 86276 301204 86278
rect 336604 86276 337204 86278
rect 372604 86276 373204 86278
rect 408604 86276 409204 86278
rect 444604 86276 445204 86278
rect 480604 86276 481204 86278
rect 516604 86276 517204 86278
rect 552604 86276 553204 86278
rect 590960 86276 591560 86278
rect -8576 86254 592500 86276
rect -8576 86018 -7454 86254
rect -7218 86018 12786 86254
rect 13022 86018 48786 86254
rect 49022 86018 84786 86254
rect 85022 86018 120786 86254
rect 121022 86018 156786 86254
rect 157022 86018 192786 86254
rect 193022 86018 228786 86254
rect 229022 86018 264786 86254
rect 265022 86018 300786 86254
rect 301022 86018 336786 86254
rect 337022 86018 372786 86254
rect 373022 86018 408786 86254
rect 409022 86018 444786 86254
rect 445022 86018 480786 86254
rect 481022 86018 516786 86254
rect 517022 86018 552786 86254
rect 553022 86018 591142 86254
rect 591378 86018 592500 86254
rect -8576 85934 592500 86018
rect -8576 85698 -7454 85934
rect -7218 85698 12786 85934
rect 13022 85698 48786 85934
rect 49022 85698 84786 85934
rect 85022 85698 120786 85934
rect 121022 85698 156786 85934
rect 157022 85698 192786 85934
rect 193022 85698 228786 85934
rect 229022 85698 264786 85934
rect 265022 85698 300786 85934
rect 301022 85698 336786 85934
rect 337022 85698 372786 85934
rect 373022 85698 408786 85934
rect 409022 85698 444786 85934
rect 445022 85698 480786 85934
rect 481022 85698 516786 85934
rect 517022 85698 552786 85934
rect 553022 85698 591142 85934
rect 591378 85698 592500 85934
rect -8576 85676 592500 85698
rect -7636 85674 -7036 85676
rect 12604 85674 13204 85676
rect 48604 85674 49204 85676
rect 84604 85674 85204 85676
rect 120604 85674 121204 85676
rect 156604 85674 157204 85676
rect 192604 85674 193204 85676
rect 228604 85674 229204 85676
rect 264604 85674 265204 85676
rect 300604 85674 301204 85676
rect 336604 85674 337204 85676
rect 372604 85674 373204 85676
rect 408604 85674 409204 85676
rect 444604 85674 445204 85676
rect 480604 85674 481204 85676
rect 516604 85674 517204 85676
rect 552604 85674 553204 85676
rect 590960 85674 591560 85676
rect -5756 82676 -5156 82678
rect 9004 82676 9604 82678
rect 45004 82676 45604 82678
rect 81004 82676 81604 82678
rect 117004 82676 117604 82678
rect 153004 82676 153604 82678
rect 189004 82676 189604 82678
rect 225004 82676 225604 82678
rect 261004 82676 261604 82678
rect 297004 82676 297604 82678
rect 333004 82676 333604 82678
rect 369004 82676 369604 82678
rect 405004 82676 405604 82678
rect 441004 82676 441604 82678
rect 477004 82676 477604 82678
rect 513004 82676 513604 82678
rect 549004 82676 549604 82678
rect 589080 82676 589680 82678
rect -6696 82654 590620 82676
rect -6696 82418 -5574 82654
rect -5338 82418 9186 82654
rect 9422 82418 45186 82654
rect 45422 82418 81186 82654
rect 81422 82418 117186 82654
rect 117422 82418 153186 82654
rect 153422 82418 189186 82654
rect 189422 82418 225186 82654
rect 225422 82418 261186 82654
rect 261422 82418 297186 82654
rect 297422 82418 333186 82654
rect 333422 82418 369186 82654
rect 369422 82418 405186 82654
rect 405422 82418 441186 82654
rect 441422 82418 477186 82654
rect 477422 82418 513186 82654
rect 513422 82418 549186 82654
rect 549422 82418 589262 82654
rect 589498 82418 590620 82654
rect -6696 82334 590620 82418
rect -6696 82098 -5574 82334
rect -5338 82098 9186 82334
rect 9422 82098 45186 82334
rect 45422 82098 81186 82334
rect 81422 82098 117186 82334
rect 117422 82098 153186 82334
rect 153422 82098 189186 82334
rect 189422 82098 225186 82334
rect 225422 82098 261186 82334
rect 261422 82098 297186 82334
rect 297422 82098 333186 82334
rect 333422 82098 369186 82334
rect 369422 82098 405186 82334
rect 405422 82098 441186 82334
rect 441422 82098 477186 82334
rect 477422 82098 513186 82334
rect 513422 82098 549186 82334
rect 549422 82098 589262 82334
rect 589498 82098 590620 82334
rect -6696 82076 590620 82098
rect -5756 82074 -5156 82076
rect 9004 82074 9604 82076
rect 45004 82074 45604 82076
rect 81004 82074 81604 82076
rect 117004 82074 117604 82076
rect 153004 82074 153604 82076
rect 189004 82074 189604 82076
rect 225004 82074 225604 82076
rect 261004 82074 261604 82076
rect 297004 82074 297604 82076
rect 333004 82074 333604 82076
rect 369004 82074 369604 82076
rect 405004 82074 405604 82076
rect 441004 82074 441604 82076
rect 477004 82074 477604 82076
rect 513004 82074 513604 82076
rect 549004 82074 549604 82076
rect 589080 82074 589680 82076
rect -3876 79076 -3276 79078
rect 5404 79076 6004 79078
rect 41404 79076 42004 79078
rect 77404 79076 78004 79078
rect 113404 79076 114004 79078
rect 149404 79076 150004 79078
rect 185404 79076 186004 79078
rect 221404 79076 222004 79078
rect 257404 79076 258004 79078
rect 293404 79076 294004 79078
rect 329404 79076 330004 79078
rect 365404 79076 366004 79078
rect 401404 79076 402004 79078
rect 437404 79076 438004 79078
rect 473404 79076 474004 79078
rect 509404 79076 510004 79078
rect 545404 79076 546004 79078
rect 581404 79076 582004 79078
rect 587200 79076 587800 79078
rect -4816 79054 588740 79076
rect -4816 78818 -3694 79054
rect -3458 78818 5586 79054
rect 5822 78818 41586 79054
rect 41822 78818 77586 79054
rect 77822 78818 113586 79054
rect 113822 78818 149586 79054
rect 149822 78818 185586 79054
rect 185822 78818 221586 79054
rect 221822 78818 257586 79054
rect 257822 78818 293586 79054
rect 293822 78818 329586 79054
rect 329822 78818 365586 79054
rect 365822 78818 401586 79054
rect 401822 78818 437586 79054
rect 437822 78818 473586 79054
rect 473822 78818 509586 79054
rect 509822 78818 545586 79054
rect 545822 78818 581586 79054
rect 581822 78818 587382 79054
rect 587618 78818 588740 79054
rect -4816 78734 588740 78818
rect -4816 78498 -3694 78734
rect -3458 78498 5586 78734
rect 5822 78498 41586 78734
rect 41822 78498 77586 78734
rect 77822 78498 113586 78734
rect 113822 78498 149586 78734
rect 149822 78498 185586 78734
rect 185822 78498 221586 78734
rect 221822 78498 257586 78734
rect 257822 78498 293586 78734
rect 293822 78498 329586 78734
rect 329822 78498 365586 78734
rect 365822 78498 401586 78734
rect 401822 78498 437586 78734
rect 437822 78498 473586 78734
rect 473822 78498 509586 78734
rect 509822 78498 545586 78734
rect 545822 78498 581586 78734
rect 581822 78498 587382 78734
rect 587618 78498 588740 78734
rect -4816 78476 588740 78498
rect -3876 78474 -3276 78476
rect 5404 78474 6004 78476
rect 41404 78474 42004 78476
rect 77404 78474 78004 78476
rect 113404 78474 114004 78476
rect 149404 78474 150004 78476
rect 185404 78474 186004 78476
rect 221404 78474 222004 78476
rect 257404 78474 258004 78476
rect 293404 78474 294004 78476
rect 329404 78474 330004 78476
rect 365404 78474 366004 78476
rect 401404 78474 402004 78476
rect 437404 78474 438004 78476
rect 473404 78474 474004 78476
rect 509404 78474 510004 78476
rect 545404 78474 546004 78476
rect 581404 78474 582004 78476
rect 587200 78474 587800 78476
rect -1996 75476 -1396 75478
rect 1804 75476 2404 75478
rect 37804 75476 38404 75478
rect 73804 75476 74404 75478
rect 109804 75476 110404 75478
rect 145804 75476 146404 75478
rect 181804 75476 182404 75478
rect 217804 75476 218404 75478
rect 253804 75476 254404 75478
rect 289804 75476 290404 75478
rect 325804 75476 326404 75478
rect 361804 75476 362404 75478
rect 397804 75476 398404 75478
rect 433804 75476 434404 75478
rect 469804 75476 470404 75478
rect 505804 75476 506404 75478
rect 541804 75476 542404 75478
rect 577804 75476 578404 75478
rect 585320 75476 585920 75478
rect -2936 75454 586860 75476
rect -2936 75218 -1814 75454
rect -1578 75218 1986 75454
rect 2222 75218 37986 75454
rect 38222 75218 73986 75454
rect 74222 75218 109986 75454
rect 110222 75218 145986 75454
rect 146222 75218 181986 75454
rect 182222 75218 217986 75454
rect 218222 75218 253986 75454
rect 254222 75218 289986 75454
rect 290222 75218 325986 75454
rect 326222 75218 361986 75454
rect 362222 75218 397986 75454
rect 398222 75218 433986 75454
rect 434222 75218 469986 75454
rect 470222 75218 505986 75454
rect 506222 75218 541986 75454
rect 542222 75218 577986 75454
rect 578222 75218 585502 75454
rect 585738 75218 586860 75454
rect -2936 75134 586860 75218
rect -2936 74898 -1814 75134
rect -1578 74898 1986 75134
rect 2222 74898 37986 75134
rect 38222 74898 73986 75134
rect 74222 74898 109986 75134
rect 110222 74898 145986 75134
rect 146222 74898 181986 75134
rect 182222 74898 217986 75134
rect 218222 74898 253986 75134
rect 254222 74898 289986 75134
rect 290222 74898 325986 75134
rect 326222 74898 361986 75134
rect 362222 74898 397986 75134
rect 398222 74898 433986 75134
rect 434222 74898 469986 75134
rect 470222 74898 505986 75134
rect 506222 74898 541986 75134
rect 542222 74898 577986 75134
rect 578222 74898 585502 75134
rect 585738 74898 586860 75134
rect -2936 74876 586860 74898
rect -1996 74874 -1396 74876
rect 1804 74874 2404 74876
rect 37804 74874 38404 74876
rect 73804 74874 74404 74876
rect 109804 74874 110404 74876
rect 145804 74874 146404 74876
rect 181804 74874 182404 74876
rect 217804 74874 218404 74876
rect 253804 74874 254404 74876
rect 289804 74874 290404 74876
rect 325804 74874 326404 74876
rect 361804 74874 362404 74876
rect 397804 74874 398404 74876
rect 433804 74874 434404 74876
rect 469804 74874 470404 74876
rect 505804 74874 506404 74876
rect 541804 74874 542404 74876
rect 577804 74874 578404 74876
rect 585320 74874 585920 74876
rect -8576 68276 -7976 68278
rect 30604 68276 31204 68278
rect 66604 68276 67204 68278
rect 102604 68276 103204 68278
rect 138604 68276 139204 68278
rect 174604 68276 175204 68278
rect 210604 68276 211204 68278
rect 246604 68276 247204 68278
rect 282604 68276 283204 68278
rect 318604 68276 319204 68278
rect 354604 68276 355204 68278
rect 390604 68276 391204 68278
rect 426604 68276 427204 68278
rect 462604 68276 463204 68278
rect 498604 68276 499204 68278
rect 534604 68276 535204 68278
rect 570604 68276 571204 68278
rect 591900 68276 592500 68278
rect -8576 68254 592500 68276
rect -8576 68018 -8394 68254
rect -8158 68018 30786 68254
rect 31022 68018 66786 68254
rect 67022 68018 102786 68254
rect 103022 68018 138786 68254
rect 139022 68018 174786 68254
rect 175022 68018 210786 68254
rect 211022 68018 246786 68254
rect 247022 68018 282786 68254
rect 283022 68018 318786 68254
rect 319022 68018 354786 68254
rect 355022 68018 390786 68254
rect 391022 68018 426786 68254
rect 427022 68018 462786 68254
rect 463022 68018 498786 68254
rect 499022 68018 534786 68254
rect 535022 68018 570786 68254
rect 571022 68018 592082 68254
rect 592318 68018 592500 68254
rect -8576 67934 592500 68018
rect -8576 67698 -8394 67934
rect -8158 67698 30786 67934
rect 31022 67698 66786 67934
rect 67022 67698 102786 67934
rect 103022 67698 138786 67934
rect 139022 67698 174786 67934
rect 175022 67698 210786 67934
rect 211022 67698 246786 67934
rect 247022 67698 282786 67934
rect 283022 67698 318786 67934
rect 319022 67698 354786 67934
rect 355022 67698 390786 67934
rect 391022 67698 426786 67934
rect 427022 67698 462786 67934
rect 463022 67698 498786 67934
rect 499022 67698 534786 67934
rect 535022 67698 570786 67934
rect 571022 67698 592082 67934
rect 592318 67698 592500 67934
rect -8576 67676 592500 67698
rect -8576 67674 -7976 67676
rect 30604 67674 31204 67676
rect 66604 67674 67204 67676
rect 102604 67674 103204 67676
rect 138604 67674 139204 67676
rect 174604 67674 175204 67676
rect 210604 67674 211204 67676
rect 246604 67674 247204 67676
rect 282604 67674 283204 67676
rect 318604 67674 319204 67676
rect 354604 67674 355204 67676
rect 390604 67674 391204 67676
rect 426604 67674 427204 67676
rect 462604 67674 463204 67676
rect 498604 67674 499204 67676
rect 534604 67674 535204 67676
rect 570604 67674 571204 67676
rect 591900 67674 592500 67676
rect -6696 64676 -6096 64678
rect 27004 64676 27604 64678
rect 63004 64676 63604 64678
rect 99004 64676 99604 64678
rect 135004 64676 135604 64678
rect 171004 64676 171604 64678
rect 207004 64676 207604 64678
rect 243004 64676 243604 64678
rect 279004 64676 279604 64678
rect 315004 64676 315604 64678
rect 351004 64676 351604 64678
rect 387004 64676 387604 64678
rect 423004 64676 423604 64678
rect 459004 64676 459604 64678
rect 495004 64676 495604 64678
rect 531004 64676 531604 64678
rect 567004 64676 567604 64678
rect 590020 64676 590620 64678
rect -6696 64654 590620 64676
rect -6696 64418 -6514 64654
rect -6278 64418 27186 64654
rect 27422 64418 63186 64654
rect 63422 64418 99186 64654
rect 99422 64418 135186 64654
rect 135422 64418 171186 64654
rect 171422 64418 207186 64654
rect 207422 64418 243186 64654
rect 243422 64418 279186 64654
rect 279422 64418 315186 64654
rect 315422 64418 351186 64654
rect 351422 64418 387186 64654
rect 387422 64418 423186 64654
rect 423422 64418 459186 64654
rect 459422 64418 495186 64654
rect 495422 64418 531186 64654
rect 531422 64418 567186 64654
rect 567422 64418 590202 64654
rect 590438 64418 590620 64654
rect -6696 64334 590620 64418
rect -6696 64098 -6514 64334
rect -6278 64098 27186 64334
rect 27422 64098 63186 64334
rect 63422 64098 99186 64334
rect 99422 64098 135186 64334
rect 135422 64098 171186 64334
rect 171422 64098 207186 64334
rect 207422 64098 243186 64334
rect 243422 64098 279186 64334
rect 279422 64098 315186 64334
rect 315422 64098 351186 64334
rect 351422 64098 387186 64334
rect 387422 64098 423186 64334
rect 423422 64098 459186 64334
rect 459422 64098 495186 64334
rect 495422 64098 531186 64334
rect 531422 64098 567186 64334
rect 567422 64098 590202 64334
rect 590438 64098 590620 64334
rect -6696 64076 590620 64098
rect -6696 64074 -6096 64076
rect 27004 64074 27604 64076
rect 63004 64074 63604 64076
rect 99004 64074 99604 64076
rect 135004 64074 135604 64076
rect 171004 64074 171604 64076
rect 207004 64074 207604 64076
rect 243004 64074 243604 64076
rect 279004 64074 279604 64076
rect 315004 64074 315604 64076
rect 351004 64074 351604 64076
rect 387004 64074 387604 64076
rect 423004 64074 423604 64076
rect 459004 64074 459604 64076
rect 495004 64074 495604 64076
rect 531004 64074 531604 64076
rect 567004 64074 567604 64076
rect 590020 64074 590620 64076
rect -4816 61076 -4216 61078
rect 23404 61076 24004 61078
rect 59404 61076 60004 61078
rect 95404 61076 96004 61078
rect 131404 61076 132004 61078
rect 167404 61076 168004 61078
rect 203404 61076 204004 61078
rect 239404 61076 240004 61078
rect 275404 61076 276004 61078
rect 311404 61076 312004 61078
rect 347404 61076 348004 61078
rect 383404 61076 384004 61078
rect 419404 61076 420004 61078
rect 455404 61076 456004 61078
rect 491404 61076 492004 61078
rect 527404 61076 528004 61078
rect 563404 61076 564004 61078
rect 588140 61076 588740 61078
rect -4816 61054 588740 61076
rect -4816 60818 -4634 61054
rect -4398 60818 23586 61054
rect 23822 60818 59586 61054
rect 59822 60818 95586 61054
rect 95822 60818 131586 61054
rect 131822 60818 167586 61054
rect 167822 60818 203586 61054
rect 203822 60818 239586 61054
rect 239822 60818 275586 61054
rect 275822 60818 311586 61054
rect 311822 60818 347586 61054
rect 347822 60818 383586 61054
rect 383822 60818 419586 61054
rect 419822 60818 455586 61054
rect 455822 60818 491586 61054
rect 491822 60818 527586 61054
rect 527822 60818 563586 61054
rect 563822 60818 588322 61054
rect 588558 60818 588740 61054
rect -4816 60734 588740 60818
rect -4816 60498 -4634 60734
rect -4398 60498 23586 60734
rect 23822 60498 59586 60734
rect 59822 60498 95586 60734
rect 95822 60498 131586 60734
rect 131822 60498 167586 60734
rect 167822 60498 203586 60734
rect 203822 60498 239586 60734
rect 239822 60498 275586 60734
rect 275822 60498 311586 60734
rect 311822 60498 347586 60734
rect 347822 60498 383586 60734
rect 383822 60498 419586 60734
rect 419822 60498 455586 60734
rect 455822 60498 491586 60734
rect 491822 60498 527586 60734
rect 527822 60498 563586 60734
rect 563822 60498 588322 60734
rect 588558 60498 588740 60734
rect -4816 60476 588740 60498
rect -4816 60474 -4216 60476
rect 23404 60474 24004 60476
rect 59404 60474 60004 60476
rect 95404 60474 96004 60476
rect 131404 60474 132004 60476
rect 167404 60474 168004 60476
rect 203404 60474 204004 60476
rect 239404 60474 240004 60476
rect 275404 60474 276004 60476
rect 311404 60474 312004 60476
rect 347404 60474 348004 60476
rect 383404 60474 384004 60476
rect 419404 60474 420004 60476
rect 455404 60474 456004 60476
rect 491404 60474 492004 60476
rect 527404 60474 528004 60476
rect 563404 60474 564004 60476
rect 588140 60474 588740 60476
rect -2936 57476 -2336 57478
rect 19804 57476 20404 57478
rect 55804 57476 56404 57478
rect 91804 57476 92404 57478
rect 127804 57476 128404 57478
rect 163804 57476 164404 57478
rect 199804 57476 200404 57478
rect 235804 57476 236404 57478
rect 271804 57476 272404 57478
rect 307804 57476 308404 57478
rect 343804 57476 344404 57478
rect 379804 57476 380404 57478
rect 415804 57476 416404 57478
rect 451804 57476 452404 57478
rect 487804 57476 488404 57478
rect 523804 57476 524404 57478
rect 559804 57476 560404 57478
rect 586260 57476 586860 57478
rect -2936 57454 586860 57476
rect -2936 57218 -2754 57454
rect -2518 57218 19986 57454
rect 20222 57218 55986 57454
rect 56222 57218 91986 57454
rect 92222 57218 127986 57454
rect 128222 57218 163986 57454
rect 164222 57218 199986 57454
rect 200222 57218 235986 57454
rect 236222 57218 271986 57454
rect 272222 57218 307986 57454
rect 308222 57218 343986 57454
rect 344222 57218 379986 57454
rect 380222 57218 415986 57454
rect 416222 57218 451986 57454
rect 452222 57218 487986 57454
rect 488222 57218 523986 57454
rect 524222 57218 559986 57454
rect 560222 57218 586442 57454
rect 586678 57218 586860 57454
rect -2936 57134 586860 57218
rect -2936 56898 -2754 57134
rect -2518 56898 19986 57134
rect 20222 56898 55986 57134
rect 56222 56898 91986 57134
rect 92222 56898 127986 57134
rect 128222 56898 163986 57134
rect 164222 56898 199986 57134
rect 200222 56898 235986 57134
rect 236222 56898 271986 57134
rect 272222 56898 307986 57134
rect 308222 56898 343986 57134
rect 344222 56898 379986 57134
rect 380222 56898 415986 57134
rect 416222 56898 451986 57134
rect 452222 56898 487986 57134
rect 488222 56898 523986 57134
rect 524222 56898 559986 57134
rect 560222 56898 586442 57134
rect 586678 56898 586860 57134
rect -2936 56876 586860 56898
rect -2936 56874 -2336 56876
rect 19804 56874 20404 56876
rect 55804 56874 56404 56876
rect 91804 56874 92404 56876
rect 127804 56874 128404 56876
rect 163804 56874 164404 56876
rect 199804 56874 200404 56876
rect 235804 56874 236404 56876
rect 271804 56874 272404 56876
rect 307804 56874 308404 56876
rect 343804 56874 344404 56876
rect 379804 56874 380404 56876
rect 415804 56874 416404 56876
rect 451804 56874 452404 56876
rect 487804 56874 488404 56876
rect 523804 56874 524404 56876
rect 559804 56874 560404 56876
rect 586260 56874 586860 56876
rect -7636 50276 -7036 50278
rect 12604 50276 13204 50278
rect 48604 50276 49204 50278
rect 84604 50276 85204 50278
rect 120604 50276 121204 50278
rect 156604 50276 157204 50278
rect 192604 50276 193204 50278
rect 228604 50276 229204 50278
rect 264604 50276 265204 50278
rect 300604 50276 301204 50278
rect 336604 50276 337204 50278
rect 372604 50276 373204 50278
rect 408604 50276 409204 50278
rect 444604 50276 445204 50278
rect 480604 50276 481204 50278
rect 516604 50276 517204 50278
rect 552604 50276 553204 50278
rect 590960 50276 591560 50278
rect -8576 50254 592500 50276
rect -8576 50018 -7454 50254
rect -7218 50018 12786 50254
rect 13022 50018 48786 50254
rect 49022 50018 84786 50254
rect 85022 50018 120786 50254
rect 121022 50018 156786 50254
rect 157022 50018 192786 50254
rect 193022 50018 228786 50254
rect 229022 50018 264786 50254
rect 265022 50018 300786 50254
rect 301022 50018 336786 50254
rect 337022 50018 372786 50254
rect 373022 50018 408786 50254
rect 409022 50018 444786 50254
rect 445022 50018 480786 50254
rect 481022 50018 516786 50254
rect 517022 50018 552786 50254
rect 553022 50018 591142 50254
rect 591378 50018 592500 50254
rect -8576 49934 592500 50018
rect -8576 49698 -7454 49934
rect -7218 49698 12786 49934
rect 13022 49698 48786 49934
rect 49022 49698 84786 49934
rect 85022 49698 120786 49934
rect 121022 49698 156786 49934
rect 157022 49698 192786 49934
rect 193022 49698 228786 49934
rect 229022 49698 264786 49934
rect 265022 49698 300786 49934
rect 301022 49698 336786 49934
rect 337022 49698 372786 49934
rect 373022 49698 408786 49934
rect 409022 49698 444786 49934
rect 445022 49698 480786 49934
rect 481022 49698 516786 49934
rect 517022 49698 552786 49934
rect 553022 49698 591142 49934
rect 591378 49698 592500 49934
rect -8576 49676 592500 49698
rect -7636 49674 -7036 49676
rect 12604 49674 13204 49676
rect 48604 49674 49204 49676
rect 84604 49674 85204 49676
rect 120604 49674 121204 49676
rect 156604 49674 157204 49676
rect 192604 49674 193204 49676
rect 228604 49674 229204 49676
rect 264604 49674 265204 49676
rect 300604 49674 301204 49676
rect 336604 49674 337204 49676
rect 372604 49674 373204 49676
rect 408604 49674 409204 49676
rect 444604 49674 445204 49676
rect 480604 49674 481204 49676
rect 516604 49674 517204 49676
rect 552604 49674 553204 49676
rect 590960 49674 591560 49676
rect -5756 46676 -5156 46678
rect 9004 46676 9604 46678
rect 45004 46676 45604 46678
rect 81004 46676 81604 46678
rect 117004 46676 117604 46678
rect 153004 46676 153604 46678
rect 189004 46676 189604 46678
rect 225004 46676 225604 46678
rect 261004 46676 261604 46678
rect 297004 46676 297604 46678
rect 333004 46676 333604 46678
rect 369004 46676 369604 46678
rect 405004 46676 405604 46678
rect 441004 46676 441604 46678
rect 477004 46676 477604 46678
rect 513004 46676 513604 46678
rect 549004 46676 549604 46678
rect 589080 46676 589680 46678
rect -6696 46654 590620 46676
rect -6696 46418 -5574 46654
rect -5338 46418 9186 46654
rect 9422 46418 45186 46654
rect 45422 46418 81186 46654
rect 81422 46418 117186 46654
rect 117422 46418 153186 46654
rect 153422 46418 189186 46654
rect 189422 46418 225186 46654
rect 225422 46418 261186 46654
rect 261422 46418 297186 46654
rect 297422 46418 333186 46654
rect 333422 46418 369186 46654
rect 369422 46418 405186 46654
rect 405422 46418 441186 46654
rect 441422 46418 477186 46654
rect 477422 46418 513186 46654
rect 513422 46418 549186 46654
rect 549422 46418 589262 46654
rect 589498 46418 590620 46654
rect -6696 46334 590620 46418
rect -6696 46098 -5574 46334
rect -5338 46098 9186 46334
rect 9422 46098 45186 46334
rect 45422 46098 81186 46334
rect 81422 46098 117186 46334
rect 117422 46098 153186 46334
rect 153422 46098 189186 46334
rect 189422 46098 225186 46334
rect 225422 46098 261186 46334
rect 261422 46098 297186 46334
rect 297422 46098 333186 46334
rect 333422 46098 369186 46334
rect 369422 46098 405186 46334
rect 405422 46098 441186 46334
rect 441422 46098 477186 46334
rect 477422 46098 513186 46334
rect 513422 46098 549186 46334
rect 549422 46098 589262 46334
rect 589498 46098 590620 46334
rect -6696 46076 590620 46098
rect -5756 46074 -5156 46076
rect 9004 46074 9604 46076
rect 45004 46074 45604 46076
rect 81004 46074 81604 46076
rect 117004 46074 117604 46076
rect 153004 46074 153604 46076
rect 189004 46074 189604 46076
rect 225004 46074 225604 46076
rect 261004 46074 261604 46076
rect 297004 46074 297604 46076
rect 333004 46074 333604 46076
rect 369004 46074 369604 46076
rect 405004 46074 405604 46076
rect 441004 46074 441604 46076
rect 477004 46074 477604 46076
rect 513004 46074 513604 46076
rect 549004 46074 549604 46076
rect 589080 46074 589680 46076
rect -3876 43076 -3276 43078
rect 5404 43076 6004 43078
rect 41404 43076 42004 43078
rect 77404 43076 78004 43078
rect 113404 43076 114004 43078
rect 149404 43076 150004 43078
rect 185404 43076 186004 43078
rect 221404 43076 222004 43078
rect 257404 43076 258004 43078
rect 293404 43076 294004 43078
rect 329404 43076 330004 43078
rect 365404 43076 366004 43078
rect 401404 43076 402004 43078
rect 437404 43076 438004 43078
rect 473404 43076 474004 43078
rect 509404 43076 510004 43078
rect 545404 43076 546004 43078
rect 581404 43076 582004 43078
rect 587200 43076 587800 43078
rect -4816 43054 588740 43076
rect -4816 42818 -3694 43054
rect -3458 42818 5586 43054
rect 5822 42818 41586 43054
rect 41822 42818 77586 43054
rect 77822 42818 113586 43054
rect 113822 42818 149586 43054
rect 149822 42818 185586 43054
rect 185822 42818 221586 43054
rect 221822 42818 257586 43054
rect 257822 42818 293586 43054
rect 293822 42818 329586 43054
rect 329822 42818 365586 43054
rect 365822 42818 401586 43054
rect 401822 42818 437586 43054
rect 437822 42818 473586 43054
rect 473822 42818 509586 43054
rect 509822 42818 545586 43054
rect 545822 42818 581586 43054
rect 581822 42818 587382 43054
rect 587618 42818 588740 43054
rect -4816 42734 588740 42818
rect -4816 42498 -3694 42734
rect -3458 42498 5586 42734
rect 5822 42498 41586 42734
rect 41822 42498 77586 42734
rect 77822 42498 113586 42734
rect 113822 42498 149586 42734
rect 149822 42498 185586 42734
rect 185822 42498 221586 42734
rect 221822 42498 257586 42734
rect 257822 42498 293586 42734
rect 293822 42498 329586 42734
rect 329822 42498 365586 42734
rect 365822 42498 401586 42734
rect 401822 42498 437586 42734
rect 437822 42498 473586 42734
rect 473822 42498 509586 42734
rect 509822 42498 545586 42734
rect 545822 42498 581586 42734
rect 581822 42498 587382 42734
rect 587618 42498 588740 42734
rect -4816 42476 588740 42498
rect -3876 42474 -3276 42476
rect 5404 42474 6004 42476
rect 41404 42474 42004 42476
rect 77404 42474 78004 42476
rect 113404 42474 114004 42476
rect 149404 42474 150004 42476
rect 185404 42474 186004 42476
rect 221404 42474 222004 42476
rect 257404 42474 258004 42476
rect 293404 42474 294004 42476
rect 329404 42474 330004 42476
rect 365404 42474 366004 42476
rect 401404 42474 402004 42476
rect 437404 42474 438004 42476
rect 473404 42474 474004 42476
rect 509404 42474 510004 42476
rect 545404 42474 546004 42476
rect 581404 42474 582004 42476
rect 587200 42474 587800 42476
rect -1996 39476 -1396 39478
rect 1804 39476 2404 39478
rect 37804 39476 38404 39478
rect 73804 39476 74404 39478
rect 109804 39476 110404 39478
rect 145804 39476 146404 39478
rect 181804 39476 182404 39478
rect 217804 39476 218404 39478
rect 253804 39476 254404 39478
rect 289804 39476 290404 39478
rect 325804 39476 326404 39478
rect 361804 39476 362404 39478
rect 397804 39476 398404 39478
rect 433804 39476 434404 39478
rect 469804 39476 470404 39478
rect 505804 39476 506404 39478
rect 541804 39476 542404 39478
rect 577804 39476 578404 39478
rect 585320 39476 585920 39478
rect -2936 39454 586860 39476
rect -2936 39218 -1814 39454
rect -1578 39218 1986 39454
rect 2222 39218 37986 39454
rect 38222 39218 73986 39454
rect 74222 39218 109986 39454
rect 110222 39218 145986 39454
rect 146222 39218 181986 39454
rect 182222 39218 217986 39454
rect 218222 39218 253986 39454
rect 254222 39218 289986 39454
rect 290222 39218 325986 39454
rect 326222 39218 361986 39454
rect 362222 39218 397986 39454
rect 398222 39218 433986 39454
rect 434222 39218 469986 39454
rect 470222 39218 505986 39454
rect 506222 39218 541986 39454
rect 542222 39218 577986 39454
rect 578222 39218 585502 39454
rect 585738 39218 586860 39454
rect -2936 39134 586860 39218
rect -2936 38898 -1814 39134
rect -1578 38898 1986 39134
rect 2222 38898 37986 39134
rect 38222 38898 73986 39134
rect 74222 38898 109986 39134
rect 110222 38898 145986 39134
rect 146222 38898 181986 39134
rect 182222 38898 217986 39134
rect 218222 38898 253986 39134
rect 254222 38898 289986 39134
rect 290222 38898 325986 39134
rect 326222 38898 361986 39134
rect 362222 38898 397986 39134
rect 398222 38898 433986 39134
rect 434222 38898 469986 39134
rect 470222 38898 505986 39134
rect 506222 38898 541986 39134
rect 542222 38898 577986 39134
rect 578222 38898 585502 39134
rect 585738 38898 586860 39134
rect -2936 38876 586860 38898
rect -1996 38874 -1396 38876
rect 1804 38874 2404 38876
rect 37804 38874 38404 38876
rect 73804 38874 74404 38876
rect 109804 38874 110404 38876
rect 145804 38874 146404 38876
rect 181804 38874 182404 38876
rect 217804 38874 218404 38876
rect 253804 38874 254404 38876
rect 289804 38874 290404 38876
rect 325804 38874 326404 38876
rect 361804 38874 362404 38876
rect 397804 38874 398404 38876
rect 433804 38874 434404 38876
rect 469804 38874 470404 38876
rect 505804 38874 506404 38876
rect 541804 38874 542404 38876
rect 577804 38874 578404 38876
rect 585320 38874 585920 38876
rect -8576 32276 -7976 32278
rect 30604 32276 31204 32278
rect 66604 32276 67204 32278
rect 102604 32276 103204 32278
rect 138604 32276 139204 32278
rect 174604 32276 175204 32278
rect 210604 32276 211204 32278
rect 246604 32276 247204 32278
rect 282604 32276 283204 32278
rect 318604 32276 319204 32278
rect 354604 32276 355204 32278
rect 390604 32276 391204 32278
rect 426604 32276 427204 32278
rect 462604 32276 463204 32278
rect 498604 32276 499204 32278
rect 534604 32276 535204 32278
rect 570604 32276 571204 32278
rect 591900 32276 592500 32278
rect -8576 32254 592500 32276
rect -8576 32018 -8394 32254
rect -8158 32018 30786 32254
rect 31022 32018 66786 32254
rect 67022 32018 102786 32254
rect 103022 32018 138786 32254
rect 139022 32018 174786 32254
rect 175022 32018 210786 32254
rect 211022 32018 246786 32254
rect 247022 32018 282786 32254
rect 283022 32018 318786 32254
rect 319022 32018 354786 32254
rect 355022 32018 390786 32254
rect 391022 32018 426786 32254
rect 427022 32018 462786 32254
rect 463022 32018 498786 32254
rect 499022 32018 534786 32254
rect 535022 32018 570786 32254
rect 571022 32018 592082 32254
rect 592318 32018 592500 32254
rect -8576 31934 592500 32018
rect -8576 31698 -8394 31934
rect -8158 31698 30786 31934
rect 31022 31698 66786 31934
rect 67022 31698 102786 31934
rect 103022 31698 138786 31934
rect 139022 31698 174786 31934
rect 175022 31698 210786 31934
rect 211022 31698 246786 31934
rect 247022 31698 282786 31934
rect 283022 31698 318786 31934
rect 319022 31698 354786 31934
rect 355022 31698 390786 31934
rect 391022 31698 426786 31934
rect 427022 31698 462786 31934
rect 463022 31698 498786 31934
rect 499022 31698 534786 31934
rect 535022 31698 570786 31934
rect 571022 31698 592082 31934
rect 592318 31698 592500 31934
rect -8576 31676 592500 31698
rect -8576 31674 -7976 31676
rect 30604 31674 31204 31676
rect 66604 31674 67204 31676
rect 102604 31674 103204 31676
rect 138604 31674 139204 31676
rect 174604 31674 175204 31676
rect 210604 31674 211204 31676
rect 246604 31674 247204 31676
rect 282604 31674 283204 31676
rect 318604 31674 319204 31676
rect 354604 31674 355204 31676
rect 390604 31674 391204 31676
rect 426604 31674 427204 31676
rect 462604 31674 463204 31676
rect 498604 31674 499204 31676
rect 534604 31674 535204 31676
rect 570604 31674 571204 31676
rect 591900 31674 592500 31676
rect -6696 28676 -6096 28678
rect 27004 28676 27604 28678
rect 63004 28676 63604 28678
rect 99004 28676 99604 28678
rect 135004 28676 135604 28678
rect 171004 28676 171604 28678
rect 207004 28676 207604 28678
rect 243004 28676 243604 28678
rect 279004 28676 279604 28678
rect 315004 28676 315604 28678
rect 351004 28676 351604 28678
rect 387004 28676 387604 28678
rect 423004 28676 423604 28678
rect 459004 28676 459604 28678
rect 495004 28676 495604 28678
rect 531004 28676 531604 28678
rect 567004 28676 567604 28678
rect 590020 28676 590620 28678
rect -6696 28654 590620 28676
rect -6696 28418 -6514 28654
rect -6278 28418 27186 28654
rect 27422 28418 63186 28654
rect 63422 28418 99186 28654
rect 99422 28418 135186 28654
rect 135422 28418 171186 28654
rect 171422 28418 207186 28654
rect 207422 28418 243186 28654
rect 243422 28418 279186 28654
rect 279422 28418 315186 28654
rect 315422 28418 351186 28654
rect 351422 28418 387186 28654
rect 387422 28418 423186 28654
rect 423422 28418 459186 28654
rect 459422 28418 495186 28654
rect 495422 28418 531186 28654
rect 531422 28418 567186 28654
rect 567422 28418 590202 28654
rect 590438 28418 590620 28654
rect -6696 28334 590620 28418
rect -6696 28098 -6514 28334
rect -6278 28098 27186 28334
rect 27422 28098 63186 28334
rect 63422 28098 99186 28334
rect 99422 28098 135186 28334
rect 135422 28098 171186 28334
rect 171422 28098 207186 28334
rect 207422 28098 243186 28334
rect 243422 28098 279186 28334
rect 279422 28098 315186 28334
rect 315422 28098 351186 28334
rect 351422 28098 387186 28334
rect 387422 28098 423186 28334
rect 423422 28098 459186 28334
rect 459422 28098 495186 28334
rect 495422 28098 531186 28334
rect 531422 28098 567186 28334
rect 567422 28098 590202 28334
rect 590438 28098 590620 28334
rect -6696 28076 590620 28098
rect -6696 28074 -6096 28076
rect 27004 28074 27604 28076
rect 63004 28074 63604 28076
rect 99004 28074 99604 28076
rect 135004 28074 135604 28076
rect 171004 28074 171604 28076
rect 207004 28074 207604 28076
rect 243004 28074 243604 28076
rect 279004 28074 279604 28076
rect 315004 28074 315604 28076
rect 351004 28074 351604 28076
rect 387004 28074 387604 28076
rect 423004 28074 423604 28076
rect 459004 28074 459604 28076
rect 495004 28074 495604 28076
rect 531004 28074 531604 28076
rect 567004 28074 567604 28076
rect 590020 28074 590620 28076
rect -4816 25076 -4216 25078
rect 23404 25076 24004 25078
rect 59404 25076 60004 25078
rect 95404 25076 96004 25078
rect 131404 25076 132004 25078
rect 167404 25076 168004 25078
rect 203404 25076 204004 25078
rect 239404 25076 240004 25078
rect 275404 25076 276004 25078
rect 311404 25076 312004 25078
rect 347404 25076 348004 25078
rect 383404 25076 384004 25078
rect 419404 25076 420004 25078
rect 455404 25076 456004 25078
rect 491404 25076 492004 25078
rect 527404 25076 528004 25078
rect 563404 25076 564004 25078
rect 588140 25076 588740 25078
rect -4816 25054 588740 25076
rect -4816 24818 -4634 25054
rect -4398 24818 23586 25054
rect 23822 24818 59586 25054
rect 59822 24818 95586 25054
rect 95822 24818 131586 25054
rect 131822 24818 167586 25054
rect 167822 24818 203586 25054
rect 203822 24818 239586 25054
rect 239822 24818 275586 25054
rect 275822 24818 311586 25054
rect 311822 24818 347586 25054
rect 347822 24818 383586 25054
rect 383822 24818 419586 25054
rect 419822 24818 455586 25054
rect 455822 24818 491586 25054
rect 491822 24818 527586 25054
rect 527822 24818 563586 25054
rect 563822 24818 588322 25054
rect 588558 24818 588740 25054
rect -4816 24734 588740 24818
rect -4816 24498 -4634 24734
rect -4398 24498 23586 24734
rect 23822 24498 59586 24734
rect 59822 24498 95586 24734
rect 95822 24498 131586 24734
rect 131822 24498 167586 24734
rect 167822 24498 203586 24734
rect 203822 24498 239586 24734
rect 239822 24498 275586 24734
rect 275822 24498 311586 24734
rect 311822 24498 347586 24734
rect 347822 24498 383586 24734
rect 383822 24498 419586 24734
rect 419822 24498 455586 24734
rect 455822 24498 491586 24734
rect 491822 24498 527586 24734
rect 527822 24498 563586 24734
rect 563822 24498 588322 24734
rect 588558 24498 588740 24734
rect -4816 24476 588740 24498
rect -4816 24474 -4216 24476
rect 23404 24474 24004 24476
rect 59404 24474 60004 24476
rect 95404 24474 96004 24476
rect 131404 24474 132004 24476
rect 167404 24474 168004 24476
rect 203404 24474 204004 24476
rect 239404 24474 240004 24476
rect 275404 24474 276004 24476
rect 311404 24474 312004 24476
rect 347404 24474 348004 24476
rect 383404 24474 384004 24476
rect 419404 24474 420004 24476
rect 455404 24474 456004 24476
rect 491404 24474 492004 24476
rect 527404 24474 528004 24476
rect 563404 24474 564004 24476
rect 588140 24474 588740 24476
rect -2936 21476 -2336 21478
rect 19804 21476 20404 21478
rect 55804 21476 56404 21478
rect 91804 21476 92404 21478
rect 127804 21476 128404 21478
rect 163804 21476 164404 21478
rect 199804 21476 200404 21478
rect 235804 21476 236404 21478
rect 271804 21476 272404 21478
rect 307804 21476 308404 21478
rect 343804 21476 344404 21478
rect 379804 21476 380404 21478
rect 415804 21476 416404 21478
rect 451804 21476 452404 21478
rect 487804 21476 488404 21478
rect 523804 21476 524404 21478
rect 559804 21476 560404 21478
rect 586260 21476 586860 21478
rect -2936 21454 586860 21476
rect -2936 21218 -2754 21454
rect -2518 21218 19986 21454
rect 20222 21218 55986 21454
rect 56222 21218 91986 21454
rect 92222 21218 127986 21454
rect 128222 21218 163986 21454
rect 164222 21218 199986 21454
rect 200222 21218 235986 21454
rect 236222 21218 271986 21454
rect 272222 21218 307986 21454
rect 308222 21218 343986 21454
rect 344222 21218 379986 21454
rect 380222 21218 415986 21454
rect 416222 21218 451986 21454
rect 452222 21218 487986 21454
rect 488222 21218 523986 21454
rect 524222 21218 559986 21454
rect 560222 21218 586442 21454
rect 586678 21218 586860 21454
rect -2936 21134 586860 21218
rect -2936 20898 -2754 21134
rect -2518 20898 19986 21134
rect 20222 20898 55986 21134
rect 56222 20898 91986 21134
rect 92222 20898 127986 21134
rect 128222 20898 163986 21134
rect 164222 20898 199986 21134
rect 200222 20898 235986 21134
rect 236222 20898 271986 21134
rect 272222 20898 307986 21134
rect 308222 20898 343986 21134
rect 344222 20898 379986 21134
rect 380222 20898 415986 21134
rect 416222 20898 451986 21134
rect 452222 20898 487986 21134
rect 488222 20898 523986 21134
rect 524222 20898 559986 21134
rect 560222 20898 586442 21134
rect 586678 20898 586860 21134
rect -2936 20876 586860 20898
rect -2936 20874 -2336 20876
rect 19804 20874 20404 20876
rect 55804 20874 56404 20876
rect 91804 20874 92404 20876
rect 127804 20874 128404 20876
rect 163804 20874 164404 20876
rect 199804 20874 200404 20876
rect 235804 20874 236404 20876
rect 271804 20874 272404 20876
rect 307804 20874 308404 20876
rect 343804 20874 344404 20876
rect 379804 20874 380404 20876
rect 415804 20874 416404 20876
rect 451804 20874 452404 20876
rect 487804 20874 488404 20876
rect 523804 20874 524404 20876
rect 559804 20874 560404 20876
rect 586260 20874 586860 20876
rect -7636 14276 -7036 14278
rect 12604 14276 13204 14278
rect 48604 14276 49204 14278
rect 84604 14276 85204 14278
rect 120604 14276 121204 14278
rect 156604 14276 157204 14278
rect 192604 14276 193204 14278
rect 228604 14276 229204 14278
rect 264604 14276 265204 14278
rect 300604 14276 301204 14278
rect 336604 14276 337204 14278
rect 372604 14276 373204 14278
rect 408604 14276 409204 14278
rect 444604 14276 445204 14278
rect 480604 14276 481204 14278
rect 516604 14276 517204 14278
rect 552604 14276 553204 14278
rect 590960 14276 591560 14278
rect -8576 14254 592500 14276
rect -8576 14018 -7454 14254
rect -7218 14018 12786 14254
rect 13022 14018 48786 14254
rect 49022 14018 84786 14254
rect 85022 14018 120786 14254
rect 121022 14018 156786 14254
rect 157022 14018 192786 14254
rect 193022 14018 228786 14254
rect 229022 14018 264786 14254
rect 265022 14018 300786 14254
rect 301022 14018 336786 14254
rect 337022 14018 372786 14254
rect 373022 14018 408786 14254
rect 409022 14018 444786 14254
rect 445022 14018 480786 14254
rect 481022 14018 516786 14254
rect 517022 14018 552786 14254
rect 553022 14018 591142 14254
rect 591378 14018 592500 14254
rect -8576 13934 592500 14018
rect -8576 13698 -7454 13934
rect -7218 13698 12786 13934
rect 13022 13698 48786 13934
rect 49022 13698 84786 13934
rect 85022 13698 120786 13934
rect 121022 13698 156786 13934
rect 157022 13698 192786 13934
rect 193022 13698 228786 13934
rect 229022 13698 264786 13934
rect 265022 13698 300786 13934
rect 301022 13698 336786 13934
rect 337022 13698 372786 13934
rect 373022 13698 408786 13934
rect 409022 13698 444786 13934
rect 445022 13698 480786 13934
rect 481022 13698 516786 13934
rect 517022 13698 552786 13934
rect 553022 13698 591142 13934
rect 591378 13698 592500 13934
rect -8576 13676 592500 13698
rect -7636 13674 -7036 13676
rect 12604 13674 13204 13676
rect 48604 13674 49204 13676
rect 84604 13674 85204 13676
rect 120604 13674 121204 13676
rect 156604 13674 157204 13676
rect 192604 13674 193204 13676
rect 228604 13674 229204 13676
rect 264604 13674 265204 13676
rect 300604 13674 301204 13676
rect 336604 13674 337204 13676
rect 372604 13674 373204 13676
rect 408604 13674 409204 13676
rect 444604 13674 445204 13676
rect 480604 13674 481204 13676
rect 516604 13674 517204 13676
rect 552604 13674 553204 13676
rect 590960 13674 591560 13676
rect -5756 10676 -5156 10678
rect 9004 10676 9604 10678
rect 45004 10676 45604 10678
rect 81004 10676 81604 10678
rect 117004 10676 117604 10678
rect 153004 10676 153604 10678
rect 189004 10676 189604 10678
rect 225004 10676 225604 10678
rect 261004 10676 261604 10678
rect 297004 10676 297604 10678
rect 333004 10676 333604 10678
rect 369004 10676 369604 10678
rect 405004 10676 405604 10678
rect 441004 10676 441604 10678
rect 477004 10676 477604 10678
rect 513004 10676 513604 10678
rect 549004 10676 549604 10678
rect 589080 10676 589680 10678
rect -6696 10654 590620 10676
rect -6696 10418 -5574 10654
rect -5338 10418 9186 10654
rect 9422 10418 45186 10654
rect 45422 10418 81186 10654
rect 81422 10418 117186 10654
rect 117422 10418 153186 10654
rect 153422 10418 189186 10654
rect 189422 10418 225186 10654
rect 225422 10418 261186 10654
rect 261422 10418 297186 10654
rect 297422 10418 333186 10654
rect 333422 10418 369186 10654
rect 369422 10418 405186 10654
rect 405422 10418 441186 10654
rect 441422 10418 477186 10654
rect 477422 10418 513186 10654
rect 513422 10418 549186 10654
rect 549422 10418 589262 10654
rect 589498 10418 590620 10654
rect -6696 10334 590620 10418
rect -6696 10098 -5574 10334
rect -5338 10098 9186 10334
rect 9422 10098 45186 10334
rect 45422 10098 81186 10334
rect 81422 10098 117186 10334
rect 117422 10098 153186 10334
rect 153422 10098 189186 10334
rect 189422 10098 225186 10334
rect 225422 10098 261186 10334
rect 261422 10098 297186 10334
rect 297422 10098 333186 10334
rect 333422 10098 369186 10334
rect 369422 10098 405186 10334
rect 405422 10098 441186 10334
rect 441422 10098 477186 10334
rect 477422 10098 513186 10334
rect 513422 10098 549186 10334
rect 549422 10098 589262 10334
rect 589498 10098 590620 10334
rect -6696 10076 590620 10098
rect -5756 10074 -5156 10076
rect 9004 10074 9604 10076
rect 45004 10074 45604 10076
rect 81004 10074 81604 10076
rect 117004 10074 117604 10076
rect 153004 10074 153604 10076
rect 189004 10074 189604 10076
rect 225004 10074 225604 10076
rect 261004 10074 261604 10076
rect 297004 10074 297604 10076
rect 333004 10074 333604 10076
rect 369004 10074 369604 10076
rect 405004 10074 405604 10076
rect 441004 10074 441604 10076
rect 477004 10074 477604 10076
rect 513004 10074 513604 10076
rect 549004 10074 549604 10076
rect 589080 10074 589680 10076
rect -3876 7076 -3276 7078
rect 5404 7076 6004 7078
rect 41404 7076 42004 7078
rect 77404 7076 78004 7078
rect 113404 7076 114004 7078
rect 149404 7076 150004 7078
rect 185404 7076 186004 7078
rect 221404 7076 222004 7078
rect 257404 7076 258004 7078
rect 293404 7076 294004 7078
rect 329404 7076 330004 7078
rect 365404 7076 366004 7078
rect 401404 7076 402004 7078
rect 437404 7076 438004 7078
rect 473404 7076 474004 7078
rect 509404 7076 510004 7078
rect 545404 7076 546004 7078
rect 581404 7076 582004 7078
rect 587200 7076 587800 7078
rect -4816 7054 588740 7076
rect -4816 6818 -3694 7054
rect -3458 6818 5586 7054
rect 5822 6818 41586 7054
rect 41822 6818 77586 7054
rect 77822 6818 113586 7054
rect 113822 6818 149586 7054
rect 149822 6818 185586 7054
rect 185822 6818 221586 7054
rect 221822 6818 257586 7054
rect 257822 6818 293586 7054
rect 293822 6818 329586 7054
rect 329822 6818 365586 7054
rect 365822 6818 401586 7054
rect 401822 6818 437586 7054
rect 437822 6818 473586 7054
rect 473822 6818 509586 7054
rect 509822 6818 545586 7054
rect 545822 6818 581586 7054
rect 581822 6818 587382 7054
rect 587618 6818 588740 7054
rect -4816 6734 588740 6818
rect -4816 6498 -3694 6734
rect -3458 6498 5586 6734
rect 5822 6498 41586 6734
rect 41822 6498 77586 6734
rect 77822 6498 113586 6734
rect 113822 6498 149586 6734
rect 149822 6498 185586 6734
rect 185822 6498 221586 6734
rect 221822 6498 257586 6734
rect 257822 6498 293586 6734
rect 293822 6498 329586 6734
rect 329822 6498 365586 6734
rect 365822 6498 401586 6734
rect 401822 6498 437586 6734
rect 437822 6498 473586 6734
rect 473822 6498 509586 6734
rect 509822 6498 545586 6734
rect 545822 6498 581586 6734
rect 581822 6498 587382 6734
rect 587618 6498 588740 6734
rect -4816 6476 588740 6498
rect -3876 6474 -3276 6476
rect 5404 6474 6004 6476
rect 41404 6474 42004 6476
rect 77404 6474 78004 6476
rect 113404 6474 114004 6476
rect 149404 6474 150004 6476
rect 185404 6474 186004 6476
rect 221404 6474 222004 6476
rect 257404 6474 258004 6476
rect 293404 6474 294004 6476
rect 329404 6474 330004 6476
rect 365404 6474 366004 6476
rect 401404 6474 402004 6476
rect 437404 6474 438004 6476
rect 473404 6474 474004 6476
rect 509404 6474 510004 6476
rect 545404 6474 546004 6476
rect 581404 6474 582004 6476
rect 587200 6474 587800 6476
rect -1996 3476 -1396 3478
rect 1804 3476 2404 3478
rect 37804 3476 38404 3478
rect 73804 3476 74404 3478
rect 109804 3476 110404 3478
rect 145804 3476 146404 3478
rect 181804 3476 182404 3478
rect 217804 3476 218404 3478
rect 253804 3476 254404 3478
rect 289804 3476 290404 3478
rect 325804 3476 326404 3478
rect 361804 3476 362404 3478
rect 397804 3476 398404 3478
rect 433804 3476 434404 3478
rect 469804 3476 470404 3478
rect 505804 3476 506404 3478
rect 541804 3476 542404 3478
rect 577804 3476 578404 3478
rect 585320 3476 585920 3478
rect -2936 3454 586860 3476
rect -2936 3218 -1814 3454
rect -1578 3218 1986 3454
rect 2222 3218 37986 3454
rect 38222 3218 73986 3454
rect 74222 3218 109986 3454
rect 110222 3218 145986 3454
rect 146222 3218 181986 3454
rect 182222 3218 217986 3454
rect 218222 3218 253986 3454
rect 254222 3218 289986 3454
rect 290222 3218 325986 3454
rect 326222 3218 361986 3454
rect 362222 3218 397986 3454
rect 398222 3218 433986 3454
rect 434222 3218 469986 3454
rect 470222 3218 505986 3454
rect 506222 3218 541986 3454
rect 542222 3218 577986 3454
rect 578222 3218 585502 3454
rect 585738 3218 586860 3454
rect -2936 3134 586860 3218
rect -2936 2898 -1814 3134
rect -1578 2898 1986 3134
rect 2222 2898 37986 3134
rect 38222 2898 73986 3134
rect 74222 2898 109986 3134
rect 110222 2898 145986 3134
rect 146222 2898 181986 3134
rect 182222 2898 217986 3134
rect 218222 2898 253986 3134
rect 254222 2898 289986 3134
rect 290222 2898 325986 3134
rect 326222 2898 361986 3134
rect 362222 2898 397986 3134
rect 398222 2898 433986 3134
rect 434222 2898 469986 3134
rect 470222 2898 505986 3134
rect 506222 2898 541986 3134
rect 542222 2898 577986 3134
rect 578222 2898 585502 3134
rect 585738 2898 586860 3134
rect -2936 2876 586860 2898
rect -1996 2874 -1396 2876
rect 1804 2874 2404 2876
rect 37804 2874 38404 2876
rect 73804 2874 74404 2876
rect 109804 2874 110404 2876
rect 145804 2874 146404 2876
rect 181804 2874 182404 2876
rect 217804 2874 218404 2876
rect 253804 2874 254404 2876
rect 289804 2874 290404 2876
rect 325804 2874 326404 2876
rect 361804 2874 362404 2876
rect 397804 2874 398404 2876
rect 433804 2874 434404 2876
rect 469804 2874 470404 2876
rect 505804 2874 506404 2876
rect 541804 2874 542404 2876
rect 577804 2874 578404 2876
rect 585320 2874 585920 2876
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 1986 -346
rect 2222 -582 37986 -346
rect 38222 -582 73986 -346
rect 74222 -582 109986 -346
rect 110222 -582 145986 -346
rect 146222 -582 181986 -346
rect 182222 -582 217986 -346
rect 218222 -582 253986 -346
rect 254222 -582 289986 -346
rect 290222 -582 325986 -346
rect 326222 -582 361986 -346
rect 362222 -582 397986 -346
rect 398222 -582 433986 -346
rect 434222 -582 469986 -346
rect 470222 -582 505986 -346
rect 506222 -582 541986 -346
rect 542222 -582 577986 -346
rect 578222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 1986 -666
rect 2222 -902 37986 -666
rect 38222 -902 73986 -666
rect 74222 -902 109986 -666
rect 110222 -902 145986 -666
rect 146222 -902 181986 -666
rect 182222 -902 217986 -666
rect 218222 -902 253986 -666
rect 254222 -902 289986 -666
rect 290222 -902 325986 -666
rect 326222 -902 361986 -666
rect 362222 -902 397986 -666
rect 398222 -902 433986 -666
rect 434222 -902 469986 -666
rect 470222 -902 505986 -666
rect 506222 -902 541986 -666
rect 542222 -902 577986 -666
rect 578222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 19986 -1286
rect 20222 -1522 55986 -1286
rect 56222 -1522 91986 -1286
rect 92222 -1522 127986 -1286
rect 128222 -1522 163986 -1286
rect 164222 -1522 199986 -1286
rect 200222 -1522 235986 -1286
rect 236222 -1522 271986 -1286
rect 272222 -1522 307986 -1286
rect 308222 -1522 343986 -1286
rect 344222 -1522 379986 -1286
rect 380222 -1522 415986 -1286
rect 416222 -1522 451986 -1286
rect 452222 -1522 487986 -1286
rect 488222 -1522 523986 -1286
rect 524222 -1522 559986 -1286
rect 560222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 19986 -1606
rect 20222 -1842 55986 -1606
rect 56222 -1842 91986 -1606
rect 92222 -1842 127986 -1606
rect 128222 -1842 163986 -1606
rect 164222 -1842 199986 -1606
rect 200222 -1842 235986 -1606
rect 236222 -1842 271986 -1606
rect 272222 -1842 307986 -1606
rect 308222 -1842 343986 -1606
rect 344222 -1842 379986 -1606
rect 380222 -1842 415986 -1606
rect 416222 -1842 451986 -1606
rect 452222 -1842 487986 -1606
rect 488222 -1842 523986 -1606
rect 524222 -1842 559986 -1606
rect 560222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 5586 -2226
rect 5822 -2462 41586 -2226
rect 41822 -2462 77586 -2226
rect 77822 -2462 113586 -2226
rect 113822 -2462 149586 -2226
rect 149822 -2462 185586 -2226
rect 185822 -2462 221586 -2226
rect 221822 -2462 257586 -2226
rect 257822 -2462 293586 -2226
rect 293822 -2462 329586 -2226
rect 329822 -2462 365586 -2226
rect 365822 -2462 401586 -2226
rect 401822 -2462 437586 -2226
rect 437822 -2462 473586 -2226
rect 473822 -2462 509586 -2226
rect 509822 -2462 545586 -2226
rect 545822 -2462 581586 -2226
rect 581822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 5586 -2546
rect 5822 -2782 41586 -2546
rect 41822 -2782 77586 -2546
rect 77822 -2782 113586 -2546
rect 113822 -2782 149586 -2546
rect 149822 -2782 185586 -2546
rect 185822 -2782 221586 -2546
rect 221822 -2782 257586 -2546
rect 257822 -2782 293586 -2546
rect 293822 -2782 329586 -2546
rect 329822 -2782 365586 -2546
rect 365822 -2782 401586 -2546
rect 401822 -2782 437586 -2546
rect 437822 -2782 473586 -2546
rect 473822 -2782 509586 -2546
rect 509822 -2782 545586 -2546
rect 545822 -2782 581586 -2546
rect 581822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 23586 -3166
rect 23822 -3402 59586 -3166
rect 59822 -3402 95586 -3166
rect 95822 -3402 131586 -3166
rect 131822 -3402 167586 -3166
rect 167822 -3402 203586 -3166
rect 203822 -3402 239586 -3166
rect 239822 -3402 275586 -3166
rect 275822 -3402 311586 -3166
rect 311822 -3402 347586 -3166
rect 347822 -3402 383586 -3166
rect 383822 -3402 419586 -3166
rect 419822 -3402 455586 -3166
rect 455822 -3402 491586 -3166
rect 491822 -3402 527586 -3166
rect 527822 -3402 563586 -3166
rect 563822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 23586 -3486
rect 23822 -3722 59586 -3486
rect 59822 -3722 95586 -3486
rect 95822 -3722 131586 -3486
rect 131822 -3722 167586 -3486
rect 167822 -3722 203586 -3486
rect 203822 -3722 239586 -3486
rect 239822 -3722 275586 -3486
rect 275822 -3722 311586 -3486
rect 311822 -3722 347586 -3486
rect 347822 -3722 383586 -3486
rect 383822 -3722 419586 -3486
rect 419822 -3722 455586 -3486
rect 455822 -3722 491586 -3486
rect 491822 -3722 527586 -3486
rect 527822 -3722 563586 -3486
rect 563822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 9186 -4106
rect 9422 -4342 45186 -4106
rect 45422 -4342 81186 -4106
rect 81422 -4342 117186 -4106
rect 117422 -4342 153186 -4106
rect 153422 -4342 189186 -4106
rect 189422 -4342 225186 -4106
rect 225422 -4342 261186 -4106
rect 261422 -4342 297186 -4106
rect 297422 -4342 333186 -4106
rect 333422 -4342 369186 -4106
rect 369422 -4342 405186 -4106
rect 405422 -4342 441186 -4106
rect 441422 -4342 477186 -4106
rect 477422 -4342 513186 -4106
rect 513422 -4342 549186 -4106
rect 549422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 9186 -4426
rect 9422 -4662 45186 -4426
rect 45422 -4662 81186 -4426
rect 81422 -4662 117186 -4426
rect 117422 -4662 153186 -4426
rect 153422 -4662 189186 -4426
rect 189422 -4662 225186 -4426
rect 225422 -4662 261186 -4426
rect 261422 -4662 297186 -4426
rect 297422 -4662 333186 -4426
rect 333422 -4662 369186 -4426
rect 369422 -4662 405186 -4426
rect 405422 -4662 441186 -4426
rect 441422 -4662 477186 -4426
rect 477422 -4662 513186 -4426
rect 513422 -4662 549186 -4426
rect 549422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 27186 -5046
rect 27422 -5282 63186 -5046
rect 63422 -5282 99186 -5046
rect 99422 -5282 135186 -5046
rect 135422 -5282 171186 -5046
rect 171422 -5282 207186 -5046
rect 207422 -5282 243186 -5046
rect 243422 -5282 279186 -5046
rect 279422 -5282 315186 -5046
rect 315422 -5282 351186 -5046
rect 351422 -5282 387186 -5046
rect 387422 -5282 423186 -5046
rect 423422 -5282 459186 -5046
rect 459422 -5282 495186 -5046
rect 495422 -5282 531186 -5046
rect 531422 -5282 567186 -5046
rect 567422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 27186 -5366
rect 27422 -5602 63186 -5366
rect 63422 -5602 99186 -5366
rect 99422 -5602 135186 -5366
rect 135422 -5602 171186 -5366
rect 171422 -5602 207186 -5366
rect 207422 -5602 243186 -5366
rect 243422 -5602 279186 -5366
rect 279422 -5602 315186 -5366
rect 315422 -5602 351186 -5366
rect 351422 -5602 387186 -5366
rect 387422 -5602 423186 -5366
rect 423422 -5602 459186 -5366
rect 459422 -5602 495186 -5366
rect 495422 -5602 531186 -5366
rect 531422 -5602 567186 -5366
rect 567422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 12786 -5986
rect 13022 -6222 48786 -5986
rect 49022 -6222 84786 -5986
rect 85022 -6222 120786 -5986
rect 121022 -6222 156786 -5986
rect 157022 -6222 192786 -5986
rect 193022 -6222 228786 -5986
rect 229022 -6222 264786 -5986
rect 265022 -6222 300786 -5986
rect 301022 -6222 336786 -5986
rect 337022 -6222 372786 -5986
rect 373022 -6222 408786 -5986
rect 409022 -6222 444786 -5986
rect 445022 -6222 480786 -5986
rect 481022 -6222 516786 -5986
rect 517022 -6222 552786 -5986
rect 553022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 12786 -6306
rect 13022 -6542 48786 -6306
rect 49022 -6542 84786 -6306
rect 85022 -6542 120786 -6306
rect 121022 -6542 156786 -6306
rect 157022 -6542 192786 -6306
rect 193022 -6542 228786 -6306
rect 229022 -6542 264786 -6306
rect 265022 -6542 300786 -6306
rect 301022 -6542 336786 -6306
rect 337022 -6542 372786 -6306
rect 373022 -6542 408786 -6306
rect 409022 -6542 444786 -6306
rect 445022 -6542 480786 -6306
rect 481022 -6542 516786 -6306
rect 517022 -6542 552786 -6306
rect 553022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 30786 -6926
rect 31022 -7162 66786 -6926
rect 67022 -7162 102786 -6926
rect 103022 -7162 138786 -6926
rect 139022 -7162 174786 -6926
rect 175022 -7162 210786 -6926
rect 211022 -7162 246786 -6926
rect 247022 -7162 282786 -6926
rect 283022 -7162 318786 -6926
rect 319022 -7162 354786 -6926
rect 355022 -7162 390786 -6926
rect 391022 -7162 426786 -6926
rect 427022 -7162 462786 -6926
rect 463022 -7162 498786 -6926
rect 499022 -7162 534786 -6926
rect 535022 -7162 570786 -6926
rect 571022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 30786 -7246
rect 31022 -7482 66786 -7246
rect 67022 -7482 102786 -7246
rect 103022 -7482 138786 -7246
rect 139022 -7482 174786 -7246
rect 175022 -7482 210786 -7246
rect 211022 -7482 246786 -7246
rect 247022 -7482 282786 -7246
rect 283022 -7482 318786 -7246
rect 319022 -7482 354786 -7246
rect 355022 -7482 390786 -7246
rect 391022 -7482 426786 -7246
rect 427022 -7482 462786 -7246
rect 463022 -7482 498786 -7246
rect 499022 -7482 534786 -7246
rect 535022 -7482 570786 -7246
rect 571022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
use adc_wrapper  mprj
timestamp 1626710249
transform 1 0 168000 0 1 338000
box -44936 -1164 268086 140972
<< labels >>
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[10]
port 1 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[11]
port 2 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[12]
port 3 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[8]
port 4 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[9]
port 5 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 6 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 7 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 8 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 9 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 10 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 11 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 12 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 13 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 14 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 15 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 16 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 17 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 18 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[16]
port 19 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[13]
port 20 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[14]
port 21 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[15]
port 22 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 23 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 24 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 25 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 26 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 27 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 28 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 29 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 30 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 31 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 32 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 33 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 34 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 35 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 36 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 37 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 38 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 39 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 40 nsew
rlabel metal2 s 47830 -960 47942 480 4 wbs_adr_i[10]
port 41 nsew
rlabel metal2 s 51326 -960 51438 480 4 wbs_adr_i[11]
port 42 nsew
rlabel metal2 s 54914 -960 55026 480 4 wbs_adr_i[12]
port 43 nsew
rlabel metal2 s 58410 -960 58522 480 4 wbs_adr_i[13]
port 44 nsew
rlabel metal2 s 61998 -960 62110 480 4 wbs_adr_i[14]
port 45 nsew
rlabel metal2 s 65494 -960 65606 480 4 wbs_adr_i[15]
port 46 nsew
rlabel metal2 s 69082 -960 69194 480 4 wbs_adr_i[16]
port 47 nsew
rlabel metal2 s 72578 -960 72690 480 4 wbs_adr_i[17]
port 48 nsew
rlabel metal2 s 12318 -960 12430 480 4 wbs_adr_i[1]
port 49 nsew
rlabel metal2 s 17010 -960 17122 480 4 wbs_adr_i[2]
port 50 nsew
rlabel metal2 s 21794 -960 21906 480 4 wbs_adr_i[3]
port 51 nsew
rlabel metal2 s 26486 -960 26598 480 4 wbs_adr_i[4]
port 52 nsew
rlabel metal2 s 30074 -960 30186 480 4 wbs_adr_i[5]
port 53 nsew
rlabel metal2 s 33570 -960 33682 480 4 wbs_adr_i[6]
port 54 nsew
rlabel metal2 s 37158 -960 37270 480 4 wbs_adr_i[7]
port 55 nsew
rlabel metal2 s 40654 -960 40766 480 4 wbs_adr_i[8]
port 56 nsew
rlabel metal2 s 44242 -960 44354 480 4 wbs_adr_i[9]
port 57 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 58 nsew
rlabel metal2 s 8730 -960 8842 480 4 wbs_dat_i[0]
port 59 nsew
rlabel metal2 s 48934 -960 49046 480 4 wbs_dat_i[10]
port 60 nsew
rlabel metal2 s 52522 -960 52634 480 4 wbs_dat_i[11]
port 61 nsew
rlabel metal2 s 56018 -960 56130 480 4 wbs_dat_i[12]
port 62 nsew
rlabel metal2 s 59606 -960 59718 480 4 wbs_dat_i[13]
port 63 nsew
rlabel metal2 s 63194 -960 63306 480 4 wbs_dat_i[14]
port 64 nsew
rlabel metal2 s 66690 -960 66802 480 4 wbs_dat_i[15]
port 65 nsew
rlabel metal2 s 70278 -960 70390 480 4 wbs_dat_i[16]
port 66 nsew
rlabel metal2 s 13514 -960 13626 480 4 wbs_dat_i[1]
port 67 nsew
rlabel metal2 s 18206 -960 18318 480 4 wbs_dat_i[2]
port 68 nsew
rlabel metal2 s 22990 -960 23102 480 4 wbs_dat_i[3]
port 69 nsew
rlabel metal2 s 27682 -960 27794 480 4 wbs_dat_i[4]
port 70 nsew
rlabel metal2 s 31270 -960 31382 480 4 wbs_dat_i[5]
port 71 nsew
rlabel metal2 s 34766 -960 34878 480 4 wbs_dat_i[6]
port 72 nsew
rlabel metal2 s 38354 -960 38466 480 4 wbs_dat_i[7]
port 73 nsew
rlabel metal2 s 41850 -960 41962 480 4 wbs_dat_i[8]
port 74 nsew
rlabel metal2 s 45438 -960 45550 480 4 wbs_dat_i[9]
port 75 nsew
rlabel metal2 s 9926 -960 10038 480 4 wbs_dat_o[0]
port 76 nsew
rlabel metal2 s 50130 -960 50242 480 4 wbs_dat_o[10]
port 77 nsew
rlabel metal2 s 53718 -960 53830 480 4 wbs_dat_o[11]
port 78 nsew
rlabel metal2 s 57214 -960 57326 480 4 wbs_dat_o[12]
port 79 nsew
rlabel metal2 s 60802 -960 60914 480 4 wbs_dat_o[13]
port 80 nsew
rlabel metal2 s 64298 -960 64410 480 4 wbs_dat_o[14]
port 81 nsew
rlabel metal2 s 67886 -960 67998 480 4 wbs_dat_o[15]
port 82 nsew
rlabel metal2 s 71474 -960 71586 480 4 wbs_dat_o[16]
port 83 nsew
rlabel metal2 s 14710 -960 14822 480 4 wbs_dat_o[1]
port 84 nsew
rlabel metal2 s 19402 -960 19514 480 4 wbs_dat_o[2]
port 85 nsew
rlabel metal2 s 24186 -960 24298 480 4 wbs_dat_o[3]
port 86 nsew
rlabel metal2 s 28878 -960 28990 480 4 wbs_dat_o[4]
port 87 nsew
rlabel metal2 s 32374 -960 32486 480 4 wbs_dat_o[5]
port 88 nsew
rlabel metal2 s 35962 -960 36074 480 4 wbs_dat_o[6]
port 89 nsew
rlabel metal2 s 39550 -960 39662 480 4 wbs_dat_o[7]
port 90 nsew
rlabel metal2 s 43046 -960 43158 480 4 wbs_dat_o[8]
port 91 nsew
rlabel metal2 s 46634 -960 46746 480 4 wbs_dat_o[9]
port 92 nsew
rlabel metal2 s 11122 -960 11234 480 4 wbs_sel_i[0]
port 93 nsew
rlabel metal2 s 15906 -960 16018 480 4 wbs_sel_i[1]
port 94 nsew
rlabel metal2 s 20598 -960 20710 480 4 wbs_sel_i[2]
port 95 nsew
rlabel metal2 s 25290 -960 25402 480 4 wbs_sel_i[3]
port 96 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 97 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 98 nsew
rlabel metal2 s 73774 -960 73886 480 4 wbs_dat_i[17]
port 99 nsew
rlabel metal2 s 77362 -960 77474 480 4 wbs_dat_i[18]
port 100 nsew
rlabel metal2 s 80858 -960 80970 480 4 wbs_dat_i[19]
port 101 nsew
rlabel metal2 s 76166 -960 76278 480 4 wbs_adr_i[18]
port 102 nsew
rlabel metal2 s 84446 -960 84558 480 4 wbs_dat_i[20]
port 103 nsew
rlabel metal2 s 87942 -960 88054 480 4 wbs_dat_i[21]
port 104 nsew
rlabel metal2 s 91530 -960 91642 480 4 wbs_dat_i[22]
port 105 nsew
rlabel metal2 s 95118 -960 95230 480 4 wbs_dat_i[23]
port 106 nsew
rlabel metal2 s 98614 -960 98726 480 4 wbs_dat_i[24]
port 107 nsew
rlabel metal2 s 102202 -960 102314 480 4 wbs_dat_i[25]
port 108 nsew
rlabel metal2 s 105698 -960 105810 480 4 wbs_dat_i[26]
port 109 nsew
rlabel metal2 s 109286 -960 109398 480 4 wbs_dat_i[27]
port 110 nsew
rlabel metal2 s 112782 -960 112894 480 4 wbs_dat_i[28]
port 111 nsew
rlabel metal2 s 116370 -960 116482 480 4 wbs_dat_i[29]
port 112 nsew
rlabel metal2 s 79662 -960 79774 480 4 wbs_adr_i[19]
port 113 nsew
rlabel metal2 s 119866 -960 119978 480 4 wbs_dat_i[30]
port 114 nsew
rlabel metal2 s 123454 -960 123566 480 4 wbs_dat_i[31]
port 115 nsew
rlabel metal2 s 128146 -960 128258 480 4 la_oenb[0]
port 116 nsew
rlabel metal2 s 83250 -960 83362 480 4 wbs_adr_i[20]
port 117 nsew
rlabel metal2 s 86838 -960 86950 480 4 wbs_adr_i[21]
port 118 nsew
rlabel metal2 s 90334 -960 90446 480 4 wbs_adr_i[22]
port 119 nsew
rlabel metal2 s 93922 -960 94034 480 4 wbs_adr_i[23]
port 120 nsew
rlabel metal2 s 97418 -960 97530 480 4 wbs_adr_i[24]
port 121 nsew
rlabel metal2 s 101006 -960 101118 480 4 wbs_adr_i[25]
port 122 nsew
rlabel metal2 s 104502 -960 104614 480 4 wbs_adr_i[26]
port 123 nsew
rlabel metal2 s 108090 -960 108202 480 4 wbs_adr_i[27]
port 124 nsew
rlabel metal2 s 111586 -960 111698 480 4 wbs_adr_i[28]
port 125 nsew
rlabel metal2 s 115174 -960 115286 480 4 wbs_adr_i[29]
port 126 nsew
rlabel metal2 s 131734 -960 131846 480 4 la_oenb[1]
port 127 nsew
rlabel metal2 s 118762 -960 118874 480 4 wbs_adr_i[30]
port 128 nsew
rlabel metal2 s 122258 -960 122370 480 4 wbs_adr_i[31]
port 129 nsew
rlabel metal2 s 135230 -960 135342 480 4 la_oenb[2]
port 130 nsew
rlabel metal2 s 74970 -960 75082 480 4 wbs_dat_o[17]
port 131 nsew
rlabel metal2 s 78558 -960 78670 480 4 wbs_dat_o[18]
port 132 nsew
rlabel metal2 s 82054 -960 82166 480 4 wbs_dat_o[19]
port 133 nsew
rlabel metal2 s 138818 -960 138930 480 4 la_oenb[3]
port 134 nsew
rlabel metal2 s 85642 -960 85754 480 4 wbs_dat_o[20]
port 135 nsew
rlabel metal2 s 89138 -960 89250 480 4 wbs_dat_o[21]
port 136 nsew
rlabel metal2 s 92726 -960 92838 480 4 wbs_dat_o[22]
port 137 nsew
rlabel metal2 s 96222 -960 96334 480 4 wbs_dat_o[23]
port 138 nsew
rlabel metal2 s 99810 -960 99922 480 4 wbs_dat_o[24]
port 139 nsew
rlabel metal2 s 103306 -960 103418 480 4 wbs_dat_o[25]
port 140 nsew
rlabel metal2 s 106894 -960 107006 480 4 wbs_dat_o[26]
port 141 nsew
rlabel metal2 s 110482 -960 110594 480 4 wbs_dat_o[27]
port 142 nsew
rlabel metal2 s 113978 -960 114090 480 4 wbs_dat_o[28]
port 143 nsew
rlabel metal2 s 117566 -960 117678 480 4 wbs_dat_o[29]
port 144 nsew
rlabel metal2 s 142406 -960 142518 480 4 la_oenb[4]
port 145 nsew
rlabel metal2 s 121062 -960 121174 480 4 wbs_dat_o[30]
port 146 nsew
rlabel metal2 s 124650 -960 124762 480 4 wbs_dat_o[31]
port 147 nsew
rlabel metal2 s 145902 -960 146014 480 4 la_oenb[5]
port 148 nsew
rlabel metal2 s 125846 -960 125958 480 4 la_data_in[0]
port 149 nsew
rlabel metal2 s 129342 -960 129454 480 4 la_data_in[1]
port 150 nsew
rlabel metal2 s 132930 -960 133042 480 4 la_data_in[2]
port 151 nsew
rlabel metal2 s 136426 -960 136538 480 4 la_data_in[3]
port 152 nsew
rlabel metal2 s 140014 -960 140126 480 4 la_data_in[4]
port 153 nsew
rlabel metal2 s 143510 -960 143622 480 4 la_data_in[5]
port 154 nsew
rlabel metal2 s 126950 -960 127062 480 4 la_data_out[0]
port 155 nsew
rlabel metal2 s 130538 -960 130650 480 4 la_data_out[1]
port 156 nsew
rlabel metal2 s 134126 -960 134238 480 4 la_data_out[2]
port 157 nsew
rlabel metal2 s 137622 -960 137734 480 4 la_data_out[3]
port 158 nsew
rlabel metal2 s 141210 -960 141322 480 4 la_data_out[4]
port 159 nsew
rlabel metal2 s 144706 -960 144818 480 4 la_data_out[5]
port 160 nsew
rlabel metal2 s 207358 -960 207470 480 4 la_data_in[23]
port 161 nsew
rlabel metal2 s 210946 -960 211058 480 4 la_data_in[24]
port 162 nsew
rlabel metal2 s 214442 -960 214554 480 4 la_data_in[25]
port 163 nsew
rlabel metal2 s 149490 -960 149602 480 4 la_oenb[6]
port 164 nsew
rlabel metal2 s 152986 -960 153098 480 4 la_oenb[7]
port 165 nsew
rlabel metal2 s 156574 -960 156686 480 4 la_oenb[8]
port 166 nsew
rlabel metal2 s 160070 -960 160182 480 4 la_oenb[9]
port 167 nsew
rlabel metal2 s 218030 -960 218142 480 4 la_data_in[26]
port 168 nsew
rlabel metal2 s 164854 -960 164966 480 4 la_data_in[11]
port 169 nsew
rlabel metal2 s 168350 -960 168462 480 4 la_data_in[12]
port 170 nsew
rlabel metal2 s 171938 -960 172050 480 4 la_data_in[13]
port 171 nsew
rlabel metal2 s 175434 -960 175546 480 4 la_data_in[14]
port 172 nsew
rlabel metal2 s 147098 -960 147210 480 4 la_data_in[6]
port 173 nsew
rlabel metal2 s 150594 -960 150706 480 4 la_data_in[7]
port 174 nsew
rlabel metal2 s 154182 -960 154294 480 4 la_data_in[8]
port 175 nsew
rlabel metal2 s 157770 -960 157882 480 4 la_data_in[9]
port 176 nsew
rlabel metal2 s 179022 -960 179134 480 4 la_data_in[15]
port 177 nsew
rlabel metal2 s 162462 -960 162574 480 4 la_data_out[10]
port 178 nsew
rlabel metal2 s 166050 -960 166162 480 4 la_data_out[11]
port 179 nsew
rlabel metal2 s 169546 -960 169658 480 4 la_data_out[12]
port 180 nsew
rlabel metal2 s 173134 -960 173246 480 4 la_data_out[13]
port 181 nsew
rlabel metal2 s 176630 -960 176742 480 4 la_data_out[14]
port 182 nsew
rlabel metal2 s 180218 -960 180330 480 4 la_data_out[15]
port 183 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_out[16]
port 184 nsew
rlabel metal2 s 187302 -960 187414 480 4 la_data_out[17]
port 185 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_out[18]
port 186 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_out[19]
port 187 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_data_in[16]
port 188 nsew
rlabel metal2 s 197882 -960 197994 480 4 la_data_out[20]
port 189 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_out[21]
port 190 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_out[22]
port 191 nsew
rlabel metal2 s 208554 -960 208666 480 4 la_data_out[23]
port 192 nsew
rlabel metal2 s 212142 -960 212254 480 4 la_data_out[24]
port 193 nsew
rlabel metal2 s 215638 -960 215750 480 4 la_data_out[25]
port 194 nsew
rlabel metal2 s 186106 -960 186218 480 4 la_data_in[17]
port 195 nsew
rlabel metal2 s 189694 -960 189806 480 4 la_data_in[18]
port 196 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_data_in[19]
port 197 nsew
rlabel metal2 s 161266 -960 161378 480 4 la_data_in[10]
port 198 nsew
rlabel metal2 s 148294 -960 148406 480 4 la_data_out[6]
port 199 nsew
rlabel metal2 s 151790 -960 151902 480 4 la_data_out[7]
port 200 nsew
rlabel metal2 s 155378 -960 155490 480 4 la_data_out[8]
port 201 nsew
rlabel metal2 s 158874 -960 158986 480 4 la_data_out[9]
port 202 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_data_in[20]
port 203 nsew
rlabel metal2 s 163658 -960 163770 480 4 la_oenb[10]
port 204 nsew
rlabel metal2 s 167154 -960 167266 480 4 la_oenb[11]
port 205 nsew
rlabel metal2 s 170742 -960 170854 480 4 la_oenb[12]
port 206 nsew
rlabel metal2 s 174238 -960 174350 480 4 la_oenb[13]
port 207 nsew
rlabel metal2 s 177826 -960 177938 480 4 la_oenb[14]
port 208 nsew
rlabel metal2 s 181414 -960 181526 480 4 la_oenb[15]
port 209 nsew
rlabel metal2 s 184910 -960 185022 480 4 la_oenb[16]
port 210 nsew
rlabel metal2 s 188498 -960 188610 480 4 la_oenb[17]
port 211 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_oenb[18]
port 212 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_oenb[19]
port 213 nsew
rlabel metal2 s 200274 -960 200386 480 4 la_data_in[21]
port 214 nsew
rlabel metal2 s 199078 -960 199190 480 4 la_oenb[20]
port 215 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_oenb[21]
port 216 nsew
rlabel metal2 s 206162 -960 206274 480 4 la_oenb[22]
port 217 nsew
rlabel metal2 s 209750 -960 209862 480 4 la_oenb[23]
port 218 nsew
rlabel metal2 s 213338 -960 213450 480 4 la_oenb[24]
port 219 nsew
rlabel metal2 s 216834 -960 216946 480 4 la_oenb[25]
port 220 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_data_in[22]
port 221 nsew
rlabel metal2 s 264122 -960 264234 480 4 la_data_in[39]
port 222 nsew
rlabel metal2 s 287766 -960 287878 480 4 la_oenb[45]
port 223 nsew
rlabel metal2 s 267710 -960 267822 480 4 la_data_in[40]
port 224 nsew
rlabel metal2 s 219226 -960 219338 480 4 la_data_out[26]
port 225 nsew
rlabel metal2 s 222722 -960 222834 480 4 la_data_out[27]
port 226 nsew
rlabel metal2 s 226310 -960 226422 480 4 la_data_out[28]
port 227 nsew
rlabel metal2 s 229806 -960 229918 480 4 la_data_out[29]
port 228 nsew
rlabel metal2 s 271206 -960 271318 480 4 la_data_in[41]
port 229 nsew
rlabel metal2 s 233394 -960 233506 480 4 la_data_out[30]
port 230 nsew
rlabel metal2 s 236982 -960 237094 480 4 la_data_out[31]
port 231 nsew
rlabel metal2 s 240478 -960 240590 480 4 la_data_out[32]
port 232 nsew
rlabel metal2 s 244066 -960 244178 480 4 la_data_out[33]
port 233 nsew
rlabel metal2 s 247562 -960 247674 480 4 la_data_out[34]
port 234 nsew
rlabel metal2 s 251150 -960 251262 480 4 la_data_out[35]
port 235 nsew
rlabel metal2 s 254646 -960 254758 480 4 la_data_out[36]
port 236 nsew
rlabel metal2 s 258234 -960 258346 480 4 la_data_out[37]
port 237 nsew
rlabel metal2 s 261730 -960 261842 480 4 la_data_out[38]
port 238 nsew
rlabel metal2 s 265318 -960 265430 480 4 la_data_out[39]
port 239 nsew
rlabel metal2 s 274794 -960 274906 480 4 la_data_in[42]
port 240 nsew
rlabel metal2 s 268814 -960 268926 480 4 la_data_out[40]
port 241 nsew
rlabel metal2 s 272402 -960 272514 480 4 la_data_out[41]
port 242 nsew
rlabel metal2 s 275990 -960 276102 480 4 la_data_out[42]
port 243 nsew
rlabel metal2 s 279486 -960 279598 480 4 la_data_out[43]
port 244 nsew
rlabel metal2 s 283074 -960 283186 480 4 la_data_out[44]
port 245 nsew
rlabel metal2 s 286570 -960 286682 480 4 la_data_out[45]
port 246 nsew
rlabel metal2 s 290158 -960 290270 480 4 la_data_out[46]
port 247 nsew
rlabel metal2 s 278290 -960 278402 480 4 la_data_in[43]
port 248 nsew
rlabel metal2 s 281878 -960 281990 480 4 la_data_in[44]
port 249 nsew
rlabel metal2 s 285374 -960 285486 480 4 la_data_in[45]
port 250 nsew
rlabel metal2 s 288962 -960 289074 480 4 la_data_in[46]
port 251 nsew
rlabel metal2 s 291354 -960 291466 480 4 la_oenb[46]
port 252 nsew
rlabel metal2 s 262926 -960 263038 480 4 la_oenb[38]
port 253 nsew
rlabel metal2 s 266514 -960 266626 480 4 la_oenb[39]
port 254 nsew
rlabel metal2 s 259430 -960 259542 480 4 la_oenb[37]
port 255 nsew
rlabel metal2 s 270010 -960 270122 480 4 la_oenb[40]
port 256 nsew
rlabel metal2 s 273598 -960 273710 480 4 la_oenb[41]
port 257 nsew
rlabel metal2 s 277094 -960 277206 480 4 la_oenb[42]
port 258 nsew
rlabel metal2 s 280682 -960 280794 480 4 la_oenb[43]
port 259 nsew
rlabel metal2 s 221526 -960 221638 480 4 la_data_in[27]
port 260 nsew
rlabel metal2 s 225114 -960 225226 480 4 la_data_in[28]
port 261 nsew
rlabel metal2 s 228702 -960 228814 480 4 la_data_in[29]
port 262 nsew
rlabel metal2 s 284270 -960 284382 480 4 la_oenb[44]
port 263 nsew
rlabel metal2 s 232198 -960 232310 480 4 la_data_in[30]
port 264 nsew
rlabel metal2 s 235786 -960 235898 480 4 la_data_in[31]
port 265 nsew
rlabel metal2 s 239282 -960 239394 480 4 la_data_in[32]
port 266 nsew
rlabel metal2 s 242870 -960 242982 480 4 la_data_in[33]
port 267 nsew
rlabel metal2 s 246366 -960 246478 480 4 la_data_in[34]
port 268 nsew
rlabel metal2 s 249954 -960 250066 480 4 la_data_in[35]
port 269 nsew
rlabel metal2 s 253450 -960 253562 480 4 la_data_in[36]
port 270 nsew
rlabel metal2 s 257038 -960 257150 480 4 la_data_in[37]
port 271 nsew
rlabel metal2 s 220422 -960 220534 480 4 la_oenb[26]
port 272 nsew
rlabel metal2 s 223918 -960 224030 480 4 la_oenb[27]
port 273 nsew
rlabel metal2 s 227506 -960 227618 480 4 la_oenb[28]
port 274 nsew
rlabel metal2 s 231002 -960 231114 480 4 la_oenb[29]
port 275 nsew
rlabel metal2 s 260626 -960 260738 480 4 la_data_in[38]
port 276 nsew
rlabel metal2 s 234590 -960 234702 480 4 la_oenb[30]
port 277 nsew
rlabel metal2 s 238086 -960 238198 480 4 la_oenb[31]
port 278 nsew
rlabel metal2 s 241674 -960 241786 480 4 la_oenb[32]
port 279 nsew
rlabel metal2 s 245170 -960 245282 480 4 la_oenb[33]
port 280 nsew
rlabel metal2 s 248758 -960 248870 480 4 la_oenb[34]
port 281 nsew
rlabel metal2 s 252346 -960 252458 480 4 la_oenb[35]
port 282 nsew
rlabel metal2 s 255842 -960 255954 480 4 la_oenb[36]
port 283 nsew
rlabel metal2 s 294850 -960 294962 480 4 la_oenb[47]
port 284 nsew
rlabel metal2 s 298438 -960 298550 480 4 la_oenb[48]
port 285 nsew
rlabel metal2 s 301934 -960 302046 480 4 la_oenb[49]
port 286 nsew
rlabel metal2 s 305522 -960 305634 480 4 la_oenb[50]
port 287 nsew
rlabel metal2 s 309018 -960 309130 480 4 la_oenb[51]
port 288 nsew
rlabel metal2 s 312606 -960 312718 480 4 la_oenb[52]
port 289 nsew
rlabel metal2 s 316194 -960 316306 480 4 la_oenb[53]
port 290 nsew
rlabel metal2 s 319690 -960 319802 480 4 la_oenb[54]
port 291 nsew
rlabel metal2 s 323278 -960 323390 480 4 la_oenb[55]
port 292 nsew
rlabel metal2 s 326774 -960 326886 480 4 la_oenb[56]
port 293 nsew
rlabel metal2 s 330362 -960 330474 480 4 la_oenb[57]
port 294 nsew
rlabel metal2 s 333858 -960 333970 480 4 la_oenb[58]
port 295 nsew
rlabel metal2 s 337446 -960 337558 480 4 la_oenb[59]
port 296 nsew
rlabel metal2 s 340942 -960 341054 480 4 la_oenb[60]
port 297 nsew
rlabel metal2 s 344530 -960 344642 480 4 la_oenb[61]
port 298 nsew
rlabel metal2 s 348026 -960 348138 480 4 la_oenb[62]
port 299 nsew
rlabel metal2 s 351614 -960 351726 480 4 la_oenb[63]
port 300 nsew
rlabel metal2 s 355202 -960 355314 480 4 la_oenb[64]
port 301 nsew
rlabel metal2 s 358698 -960 358810 480 4 la_oenb[65]
port 302 nsew
rlabel metal2 s 362286 -960 362398 480 4 la_oenb[66]
port 303 nsew
rlabel metal2 s 292550 -960 292662 480 4 la_data_in[47]
port 304 nsew
rlabel metal2 s 296046 -960 296158 480 4 la_data_in[48]
port 305 nsew
rlabel metal2 s 299634 -960 299746 480 4 la_data_in[49]
port 306 nsew
rlabel metal2 s 303130 -960 303242 480 4 la_data_in[50]
port 307 nsew
rlabel metal2 s 306718 -960 306830 480 4 la_data_in[51]
port 308 nsew
rlabel metal2 s 310214 -960 310326 480 4 la_data_in[52]
port 309 nsew
rlabel metal2 s 313802 -960 313914 480 4 la_data_in[53]
port 310 nsew
rlabel metal2 s 317298 -960 317410 480 4 la_data_in[54]
port 311 nsew
rlabel metal2 s 320886 -960 320998 480 4 la_data_in[55]
port 312 nsew
rlabel metal2 s 324382 -960 324494 480 4 la_data_in[56]
port 313 nsew
rlabel metal2 s 327970 -960 328082 480 4 la_data_in[57]
port 314 nsew
rlabel metal2 s 331558 -960 331670 480 4 la_data_in[58]
port 315 nsew
rlabel metal2 s 335054 -960 335166 480 4 la_data_in[59]
port 316 nsew
rlabel metal2 s 338642 -960 338754 480 4 la_data_in[60]
port 317 nsew
rlabel metal2 s 342138 -960 342250 480 4 la_data_in[61]
port 318 nsew
rlabel metal2 s 345726 -960 345838 480 4 la_data_in[62]
port 319 nsew
rlabel metal2 s 349222 -960 349334 480 4 la_data_in[63]
port 320 nsew
rlabel metal2 s 293654 -960 293766 480 4 la_data_out[47]
port 321 nsew
rlabel metal2 s 297242 -960 297354 480 4 la_data_out[48]
port 322 nsew
rlabel metal2 s 300738 -960 300850 480 4 la_data_out[49]
port 323 nsew
rlabel metal2 s 352810 -960 352922 480 4 la_data_in[64]
port 324 nsew
rlabel metal2 s 304326 -960 304438 480 4 la_data_out[50]
port 325 nsew
rlabel metal2 s 307914 -960 308026 480 4 la_data_out[51]
port 326 nsew
rlabel metal2 s 311410 -960 311522 480 4 la_data_out[52]
port 327 nsew
rlabel metal2 s 314998 -960 315110 480 4 la_data_out[53]
port 328 nsew
rlabel metal2 s 318494 -960 318606 480 4 la_data_out[54]
port 329 nsew
rlabel metal2 s 322082 -960 322194 480 4 la_data_out[55]
port 330 nsew
rlabel metal2 s 325578 -960 325690 480 4 la_data_out[56]
port 331 nsew
rlabel metal2 s 329166 -960 329278 480 4 la_data_out[57]
port 332 nsew
rlabel metal2 s 332662 -960 332774 480 4 la_data_out[58]
port 333 nsew
rlabel metal2 s 336250 -960 336362 480 4 la_data_out[59]
port 334 nsew
rlabel metal2 s 356306 -960 356418 480 4 la_data_in[65]
port 335 nsew
rlabel metal2 s 339838 -960 339950 480 4 la_data_out[60]
port 336 nsew
rlabel metal2 s 343334 -960 343446 480 4 la_data_out[61]
port 337 nsew
rlabel metal2 s 346922 -960 347034 480 4 la_data_out[62]
port 338 nsew
rlabel metal2 s 350418 -960 350530 480 4 la_data_out[63]
port 339 nsew
rlabel metal2 s 354006 -960 354118 480 4 la_data_out[64]
port 340 nsew
rlabel metal2 s 357502 -960 357614 480 4 la_data_out[65]
port 341 nsew
rlabel metal2 s 361090 -960 361202 480 4 la_data_out[66]
port 342 nsew
rlabel metal2 s 364586 -960 364698 480 4 la_data_out[67]
port 343 nsew
rlabel metal2 s 359894 -960 360006 480 4 la_data_in[66]
port 344 nsew
rlabel metal2 s 363482 -960 363594 480 4 la_data_in[67]
port 345 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_in[72]
port 346 nsew
rlabel metal2 s 384734 -960 384846 480 4 la_data_in[73]
port 347 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_in[74]
port 348 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_in[75]
port 349 nsew
rlabel metal2 s 395314 -960 395426 480 4 la_data_in[76]
port 350 nsew
rlabel metal2 s 398902 -960 399014 480 4 la_data_in[77]
port 351 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_in[78]
port 352 nsew
rlabel metal2 s 405986 -960 406098 480 4 la_data_in[79]
port 353 nsew
rlabel metal2 s 409574 -960 409686 480 4 la_data_in[80]
port 354 nsew
rlabel metal2 s 413070 -960 413182 480 4 la_data_in[81]
port 355 nsew
rlabel metal2 s 416658 -960 416770 480 4 la_data_in[82]
port 356 nsew
rlabel metal2 s 420154 -960 420266 480 4 la_data_in[83]
port 357 nsew
rlabel metal2 s 423742 -960 423854 480 4 la_data_in[84]
port 358 nsew
rlabel metal2 s 427238 -960 427350 480 4 la_data_in[85]
port 359 nsew
rlabel metal2 s 430826 -960 430938 480 4 la_data_in[86]
port 360 nsew
rlabel metal2 s 434414 -960 434526 480 4 la_data_in[87]
port 361 nsew
rlabel metal2 s 370566 -960 370678 480 4 la_data_in[69]
port 362 nsew
rlabel metal2 s 365782 -960 365894 480 4 la_oenb[67]
port 363 nsew
rlabel metal2 s 369370 -960 369482 480 4 la_oenb[68]
port 364 nsew
rlabel metal2 s 372866 -960 372978 480 4 la_oenb[69]
port 365 nsew
rlabel metal2 s 376454 -960 376566 480 4 la_oenb[70]
port 366 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_oenb[71]
port 367 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_oenb[72]
port 368 nsew
rlabel metal2 s 387126 -960 387238 480 4 la_oenb[73]
port 369 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_oenb[74]
port 370 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_oenb[75]
port 371 nsew
rlabel metal2 s 397706 -960 397818 480 4 la_oenb[76]
port 372 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_oenb[77]
port 373 nsew
rlabel metal2 s 404790 -960 404902 480 4 la_oenb[78]
port 374 nsew
rlabel metal2 s 408378 -960 408490 480 4 la_oenb[79]
port 375 nsew
rlabel metal2 s 411874 -960 411986 480 4 la_oenb[80]
port 376 nsew
rlabel metal2 s 415462 -960 415574 480 4 la_oenb[81]
port 377 nsew
rlabel metal2 s 418958 -960 419070 480 4 la_oenb[82]
port 378 nsew
rlabel metal2 s 422546 -960 422658 480 4 la_oenb[83]
port 379 nsew
rlabel metal2 s 426134 -960 426246 480 4 la_oenb[84]
port 380 nsew
rlabel metal2 s 429630 -960 429742 480 4 la_oenb[85]
port 381 nsew
rlabel metal2 s 433218 -960 433330 480 4 la_oenb[86]
port 382 nsew
rlabel metal2 s 436714 -960 436826 480 4 la_oenb[87]
port 383 nsew
rlabel metal2 s 368174 -960 368286 480 4 la_data_out[68]
port 384 nsew
rlabel metal2 s 371670 -960 371782 480 4 la_data_out[69]
port 385 nsew
rlabel metal2 s 374062 -960 374174 480 4 la_data_in[70]
port 386 nsew
rlabel metal2 s 375258 -960 375370 480 4 la_data_out[70]
port 387 nsew
rlabel metal2 s 378846 -960 378958 480 4 la_data_out[71]
port 388 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_data_out[72]
port 389 nsew
rlabel metal2 s 385930 -960 386042 480 4 la_data_out[73]
port 390 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_data_out[74]
port 391 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_data_out[75]
port 392 nsew
rlabel metal2 s 396510 -960 396622 480 4 la_data_out[76]
port 393 nsew
rlabel metal2 s 400098 -960 400210 480 4 la_data_out[77]
port 394 nsew
rlabel metal2 s 403594 -960 403706 480 4 la_data_out[78]
port 395 nsew
rlabel metal2 s 407182 -960 407294 480 4 la_data_out[79]
port 396 nsew
rlabel metal2 s 377650 -960 377762 480 4 la_data_in[71]
port 397 nsew
rlabel metal2 s 410770 -960 410882 480 4 la_data_out[80]
port 398 nsew
rlabel metal2 s 414266 -960 414378 480 4 la_data_out[81]
port 399 nsew
rlabel metal2 s 417854 -960 417966 480 4 la_data_out[82]
port 400 nsew
rlabel metal2 s 421350 -960 421462 480 4 la_data_out[83]
port 401 nsew
rlabel metal2 s 424938 -960 425050 480 4 la_data_out[84]
port 402 nsew
rlabel metal2 s 428434 -960 428546 480 4 la_data_out[85]
port 403 nsew
rlabel metal2 s 432022 -960 432134 480 4 la_data_out[86]
port 404 nsew
rlabel metal2 s 435518 -960 435630 480 4 la_data_out[87]
port 405 nsew
rlabel metal2 s 366978 -960 367090 480 4 la_data_in[68]
port 406 nsew
rlabel metal2 s 440302 -960 440414 480 4 la_oenb[88]
port 407 nsew
rlabel metal2 s 443798 -960 443910 480 4 la_oenb[89]
port 408 nsew
rlabel metal2 s 447386 -960 447498 480 4 la_oenb[90]
port 409 nsew
rlabel metal2 s 450882 -960 450994 480 4 la_oenb[91]
port 410 nsew
rlabel metal2 s 454470 -960 454582 480 4 la_oenb[92]
port 411 nsew
rlabel metal2 s 458058 -960 458170 480 4 la_oenb[93]
port 412 nsew
rlabel metal2 s 461554 -960 461666 480 4 la_oenb[94]
port 413 nsew
rlabel metal2 s 465142 -960 465254 480 4 la_oenb[95]
port 414 nsew
rlabel metal2 s 468638 -960 468750 480 4 la_oenb[96]
port 415 nsew
rlabel metal2 s 472226 -960 472338 480 4 la_oenb[97]
port 416 nsew
rlabel metal2 s 475722 -960 475834 480 4 la_oenb[98]
port 417 nsew
rlabel metal2 s 479310 -960 479422 480 4 la_oenb[99]
port 418 nsew
rlabel metal2 s 484002 -960 484114 480 4 la_data_in[101]
port 419 nsew
rlabel metal2 s 487590 -960 487702 480 4 la_data_in[102]
port 420 nsew
rlabel metal2 s 491086 -960 491198 480 4 la_data_in[103]
port 421 nsew
rlabel metal2 s 494674 -960 494786 480 4 la_data_in[104]
port 422 nsew
rlabel metal2 s 498170 -960 498282 480 4 la_data_in[105]
port 423 nsew
rlabel metal2 s 501758 -960 501870 480 4 la_data_in[106]
port 424 nsew
rlabel metal2 s 505346 -960 505458 480 4 la_data_in[107]
port 425 nsew
rlabel metal2 s 508842 -960 508954 480 4 la_data_in[108]
port 426 nsew
rlabel metal2 s 480506 -960 480618 480 4 la_data_in[100]
port 427 nsew
rlabel metal2 s 444994 -960 445106 480 4 la_data_in[90]
port 428 nsew
rlabel metal2 s 448582 -960 448694 480 4 la_data_in[91]
port 429 nsew
rlabel metal2 s 452078 -960 452190 480 4 la_data_in[92]
port 430 nsew
rlabel metal2 s 455666 -960 455778 480 4 la_data_in[93]
port 431 nsew
rlabel metal2 s 459162 -960 459274 480 4 la_data_in[94]
port 432 nsew
rlabel metal2 s 462750 -960 462862 480 4 la_data_in[95]
port 433 nsew
rlabel metal2 s 466246 -960 466358 480 4 la_data_in[96]
port 434 nsew
rlabel metal2 s 469834 -960 469946 480 4 la_data_in[97]
port 435 nsew
rlabel metal2 s 473422 -960 473534 480 4 la_data_in[98]
port 436 nsew
rlabel metal2 s 476918 -960 477030 480 4 la_data_in[99]
port 437 nsew
rlabel metal2 s 481702 -960 481814 480 4 la_data_out[100]
port 438 nsew
rlabel metal2 s 485198 -960 485310 480 4 la_data_out[101]
port 439 nsew
rlabel metal2 s 488786 -960 488898 480 4 la_data_out[102]
port 440 nsew
rlabel metal2 s 492282 -960 492394 480 4 la_data_out[103]
port 441 nsew
rlabel metal2 s 495870 -960 495982 480 4 la_data_out[104]
port 442 nsew
rlabel metal2 s 499366 -960 499478 480 4 la_data_out[105]
port 443 nsew
rlabel metal2 s 456862 -960 456974 480 4 la_data_out[93]
port 444 nsew
rlabel metal2 s 502954 -960 503066 480 4 la_data_out[106]
port 445 nsew
rlabel metal2 s 460358 -960 460470 480 4 la_data_out[94]
port 446 nsew
rlabel metal2 s 506450 -960 506562 480 4 la_data_out[107]
port 447 nsew
rlabel metal2 s 463946 -960 464058 480 4 la_data_out[95]
port 448 nsew
rlabel metal2 s 467442 -960 467554 480 4 la_data_out[96]
port 449 nsew
rlabel metal2 s 510038 -960 510150 480 4 la_data_out[108]
port 450 nsew
rlabel metal2 s 471030 -960 471142 480 4 la_data_out[97]
port 451 nsew
rlabel metal2 s 474526 -960 474638 480 4 la_data_out[98]
port 452 nsew
rlabel metal2 s 478114 -960 478226 480 4 la_data_out[99]
port 453 nsew
rlabel metal2 s 453274 -960 453386 480 4 la_data_out[92]
port 454 nsew
rlabel metal2 s 482806 -960 482918 480 4 la_oenb[100]
port 455 nsew
rlabel metal2 s 486394 -960 486506 480 4 la_oenb[101]
port 456 nsew
rlabel metal2 s 489890 -960 490002 480 4 la_oenb[102]
port 457 nsew
rlabel metal2 s 493478 -960 493590 480 4 la_oenb[103]
port 458 nsew
rlabel metal2 s 497066 -960 497178 480 4 la_oenb[104]
port 459 nsew
rlabel metal2 s 500562 -960 500674 480 4 la_oenb[105]
port 460 nsew
rlabel metal2 s 504150 -960 504262 480 4 la_oenb[106]
port 461 nsew
rlabel metal2 s 507646 -960 507758 480 4 la_oenb[107]
port 462 nsew
rlabel metal2 s 437910 -960 438022 480 4 la_data_in[88]
port 463 nsew
rlabel metal2 s 441498 -960 441610 480 4 la_data_in[89]
port 464 nsew
rlabel metal2 s 439106 -960 439218 480 4 la_data_out[88]
port 465 nsew
rlabel metal2 s 442602 -960 442714 480 4 la_data_out[89]
port 466 nsew
rlabel metal2 s 446190 -960 446302 480 4 la_data_out[90]
port 467 nsew
rlabel metal2 s 449778 -960 449890 480 4 la_data_out[91]
port 468 nsew
rlabel metal2 s 547850 -960 547962 480 4 la_data_in[119]
port 469 nsew
rlabel metal2 s 552634 -960 552746 480 4 la_data_out[120]
port 470 nsew
rlabel metal2 s 556130 -960 556242 480 4 la_data_out[121]
port 471 nsew
rlabel metal2 s 559718 -960 559830 480 4 la_data_out[122]
port 472 nsew
rlabel metal2 s 537178 -960 537290 480 4 la_data_in[116]
port 473 nsew
rlabel metal2 s 540766 -960 540878 480 4 la_data_in[117]
port 474 nsew
rlabel metal2 s 563214 -960 563326 480 4 la_data_out[123]
port 475 nsew
rlabel metal2 s 523010 -960 523122 480 4 la_data_in[112]
port 476 nsew
rlabel metal2 s 566802 -960 566914 480 4 la_data_out[124]
port 477 nsew
rlabel metal2 s 570298 -960 570410 480 4 la_data_out[125]
port 478 nsew
rlabel metal2 s 573886 -960 573998 480 4 la_data_out[126]
port 479 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[127]
port 480 nsew
rlabel metal2 s 544354 -960 544466 480 4 la_data_in[118]
port 481 nsew
rlabel metal2 s 514730 -960 514842 480 4 la_oenb[109]
port 482 nsew
rlabel metal2 s 551438 -960 551550 480 4 la_data_in[120]
port 483 nsew
rlabel metal2 s 518318 -960 518430 480 4 la_oenb[110]
port 484 nsew
rlabel metal2 s 554934 -960 555046 480 4 la_data_in[121]
port 485 nsew
rlabel metal2 s 521814 -960 521926 480 4 la_oenb[111]
port 486 nsew
rlabel metal2 s 525402 -960 525514 480 4 la_oenb[112]
port 487 nsew
rlabel metal2 s 528990 -960 529102 480 4 la_oenb[113]
port 488 nsew
rlabel metal2 s 532486 -960 532598 480 4 la_oenb[114]
port 489 nsew
rlabel metal2 s 536074 -960 536186 480 4 la_oenb[115]
port 490 nsew
rlabel metal2 s 539570 -960 539682 480 4 la_oenb[116]
port 491 nsew
rlabel metal2 s 543158 -960 543270 480 4 la_oenb[117]
port 492 nsew
rlabel metal2 s 546654 -960 546766 480 4 la_oenb[118]
port 493 nsew
rlabel metal2 s 550242 -960 550354 480 4 la_oenb[119]
port 494 nsew
rlabel metal2 s 558522 -960 558634 480 4 la_data_in[122]
port 495 nsew
rlabel metal2 s 562018 -960 562130 480 4 la_data_in[123]
port 496 nsew
rlabel metal2 s 553738 -960 553850 480 4 la_oenb[120]
port 497 nsew
rlabel metal2 s 557326 -960 557438 480 4 la_oenb[121]
port 498 nsew
rlabel metal2 s 560822 -960 560934 480 4 la_oenb[122]
port 499 nsew
rlabel metal2 s 564410 -960 564522 480 4 la_oenb[123]
port 500 nsew
rlabel metal2 s 567998 -960 568110 480 4 la_oenb[124]
port 501 nsew
rlabel metal2 s 571494 -960 571606 480 4 la_oenb[125]
port 502 nsew
rlabel metal2 s 575082 -960 575194 480 4 la_oenb[126]
port 503 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oenb[127]
port 504 nsew
rlabel metal2 s 565606 -960 565718 480 4 la_data_in[124]
port 505 nsew
rlabel metal2 s 569102 -960 569214 480 4 la_data_in[125]
port 506 nsew
rlabel metal2 s 572690 -960 572802 480 4 la_data_in[126]
port 507 nsew
rlabel metal2 s 576278 -960 576390 480 4 la_data_in[127]
port 508 nsew
rlabel metal2 s 517122 -960 517234 480 4 la_data_out[110]
port 509 nsew
rlabel metal2 s 579774 -960 579886 480 4 user_clock2
port 510 nsew
rlabel metal2 s 580970 -960 581082 480 4 user_irq[0]
port 511 nsew
rlabel metal2 s 526598 -960 526710 480 4 la_data_in[113]
port 512 nsew
rlabel metal2 s 582166 -960 582278 480 4 user_irq[1]
port 513 nsew
rlabel metal2 s 530094 -960 530206 480 4 la_data_in[114]
port 514 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_irq[2]
port 515 nsew
rlabel metal2 s 520710 -960 520822 480 4 la_data_out[111]
port 516 nsew
rlabel metal2 s 524206 -960 524318 480 4 la_data_out[112]
port 517 nsew
rlabel metal2 s 513534 -960 513646 480 4 la_data_out[109]
port 518 nsew
rlabel metal2 s 512430 -960 512542 480 4 la_data_in[109]
port 519 nsew
rlabel metal2 s 527794 -960 527906 480 4 la_data_out[113]
port 520 nsew
rlabel metal2 s 515926 -960 516038 480 4 la_data_in[110]
port 521 nsew
rlabel metal2 s 531290 -960 531402 480 4 la_data_out[114]
port 522 nsew
rlabel metal2 s 511234 -960 511346 480 4 la_oenb[108]
port 523 nsew
rlabel metal2 s 534878 -960 534990 480 4 la_data_out[115]
port 524 nsew
rlabel metal2 s 538374 -960 538486 480 4 la_data_out[116]
port 525 nsew
rlabel metal2 s 519514 -960 519626 480 4 la_data_in[111]
port 526 nsew
rlabel metal2 s 541962 -960 542074 480 4 la_data_out[117]
port 527 nsew
rlabel metal2 s 533682 -960 533794 480 4 la_data_in[115]
port 528 nsew
rlabel metal2 s 545458 -960 545570 480 4 la_data_out[118]
port 529 nsew
rlabel metal2 s 549046 -960 549158 480 4 la_data_out[119]
port 530 nsew
rlabel metal4 s 433804 598000 434404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 397804 598000 398404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 361804 598000 362404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 325804 598000 326404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 415804 598000 416404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 379804 598000 380404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 343804 598000 344404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 307804 598000 308404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 437404 598000 438004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 401404 598000 402004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 365404 598000 366004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 329404 598000 330004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 293404 598000 294004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 419404 598000 420004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 383404 598000 384004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 347404 598000 348004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 311404 598000 312004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 441004 598000 441604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 405004 598000 405604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 369004 598000 369604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 333004 598000 333604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 297004 598000 297604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 423004 598000 423604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 387004 598000 387604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 351004 598000 351604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 315004 598000 315604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 444604 598000 445204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 408604 598000 409204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 372604 598000 373204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 336604 598000 337204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 300604 598000 301204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 426604 598000 427204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 390604 598000 391204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 354604 598000 355204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 318604 598000 319204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 203404 598000 204004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 167404 598000 168004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 131404 598000 132004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 163804 598000 164404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 127804 598000 128404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 145804 598000 146404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 109804 598000 110404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 289804 598000 290404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 261004 598000 261604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 225004 598000 225604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 189004 598000 189604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 153004 598000 153604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 117004 598000 117604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 253804 598000 254404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 217804 598000 218404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 257404 598000 258004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 221404 598000 222004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 279004 598000 279604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 243004 598000 243604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 207004 598000 207604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 171004 598000 171604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 135004 598000 135604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 185404 598000 186004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 149404 598000 150004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 113404 598000 114004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 181804 598000 182404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 271804 598000 272404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 264604 598000 265204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 228604 598000 229204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 192604 598000 193204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 156604 598000 157204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 120604 598000 121204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 235804 598000 236404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 199804 598000 200404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 275404 598000 276004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 239404 598000 240004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 282604 598000 283204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 246604 598000 247204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 210604 598000 211204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 174604 598000 175204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 138604 598000 139204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 73804 -1864 74404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 37804 -1864 38404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 1804 -1864 2404 705800 4 vccd1
port 531 nsew
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 531 nsew
rlabel metal4 s 289804 -1864 290404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 253804 -1864 254404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 217804 -1864 218404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 181804 -1864 182404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 145804 -1864 146404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 81004 -5624 81604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 45004 -5624 45604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 9004 -5624 9604 709560 4 vdda1
port 535 nsew
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 535 nsew
rlabel metal4 s 261004 -5624 261604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 225004 -5624 225604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 189004 -5624 189604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 153004 -5624 153604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 117004 -5624 117604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 77404 -3744 78004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 41404 -3744 42004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 5404 -3744 6004 707680 4 vccd2
port 533 nsew
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 533 nsew
rlabel metal4 s 257404 -3744 258004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 221404 -3744 222004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 185404 -3744 186004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 149404 -3744 150004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 113404 -3744 114004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 99004 -5624 99604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 63004 -5624 63604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 27004 -5624 27604 709560 4 vssa1
port 536 nsew
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 536 nsew
rlabel metal4 s 279004 -5624 279604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 243004 -5624 243604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 207004 -5624 207604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 171004 -5624 171604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 135004 -5624 135604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 91804 -1864 92404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 55804 -1864 56404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 19804 -1864 20404 705800 4 vssd1
port 532 nsew
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 532 nsew
rlabel metal4 s 271804 -1864 272404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 235804 -1864 236404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 199804 -1864 200404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 163804 -1864 164404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 127804 -1864 128404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 95404 -3744 96004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 84604 -7504 85204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 48604 -7504 49204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 12604 -7504 13204 711440 4 vdda2
port 537 nsew
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 537 nsew
rlabel metal4 s 264604 -7504 265204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 228604 -7504 229204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 192604 -7504 193204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 156604 -7504 157204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 120604 -7504 121204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 59404 -3744 60004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 23404 -3744 24004 707680 4 vssd2
port 534 nsew
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 534 nsew
rlabel metal4 s 275404 -3744 276004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 239404 -3744 240004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 203404 -3744 204004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 167404 -3744 168004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 131404 -3744 132004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 109804 -1864 110404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 102604 -7504 103204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 66604 -7504 67204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 30604 -7504 31204 711440 4 vssa2
port 538 nsew
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 538 nsew
rlabel metal4 s 282604 -7504 283204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 246604 -7504 247204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 210604 -7504 211204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 174604 -7504 175204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 138604 -7504 139204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 586260 -1864 586860 705800 4 vssd1
port 532 nsew
rlabel metal4 s 559804 -1864 560404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 523804 -1864 524404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 487804 -1864 488404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 415804 -1864 416404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 419404 -3744 420004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 383404 -3744 384004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 347404 -3744 348004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 311404 -3744 312004 218000 4 vssd2
port 534 nsew
rlabel metal4 s 423004 -5624 423604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 387004 -5624 387604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 351004 -5624 351604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 315004 -5624 315604 218000 4 vssa1
port 536 nsew
rlabel metal4 s 379804 -1864 380404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 343804 -1864 344404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 307804 -1864 308404 218000 4 vssd1
port 532 nsew
rlabel metal4 s 587200 -2804 587800 706740 4 vccd2
port 533 nsew
rlabel metal4 s 451804 -1864 452404 705800 4 vssd1
port 532 nsew
rlabel metal4 s 552604 -7504 553204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 516604 -7504 517204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 480604 -7504 481204 711440 4 vdda2
port 537 nsew
rlabel metal4 s 549004 -5624 549604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 513004 -5624 513604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 477004 -5624 477604 709560 4 vdda1
port 535 nsew
rlabel metal4 s 437404 -3744 438004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 401404 -3744 402004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 365404 -3744 366004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 329404 -3744 330004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 293404 -3744 294004 218000 4 vccd2
port 533 nsew
rlabel metal4 s 397804 -1864 398404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 361804 -1864 362404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 325804 -1864 326404 218000 4 vccd1
port 531 nsew
rlabel metal4 s 505804 -1864 506404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 581404 -3744 582004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 590960 -6564 591560 710500 4 vdda2
port 537 nsew
rlabel metal4 s 588140 -3744 588740 707680 4 vssd2
port 534 nsew
rlabel metal4 s 444604 -7504 445204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 408604 -7504 409204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 372604 -7504 373204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 336604 -7504 337204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 300604 -7504 301204 218000 4 vdda2
port 537 nsew
rlabel metal4 s 563404 -3744 564004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 527404 -3744 528004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 589080 -4684 589680 708620 4 vdda1
port 535 nsew
rlabel metal4 s 491404 -3744 492004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 441004 -5624 441604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 591900 -7504 592500 711440 4 vssa2
port 538 nsew
rlabel metal4 s 570604 -7504 571204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 534604 -7504 535204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 498604 -7504 499204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 462604 -7504 463204 711440 4 vssa2
port 538 nsew
rlabel metal4 s 405004 -5624 405604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 369004 -5624 369604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 333004 -5624 333604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 297004 -5624 297604 218000 4 vdda1
port 535 nsew
rlabel metal4 s 455404 -3744 456004 707680 4 vssd2
port 534 nsew
rlabel metal4 s 545404 -3744 546004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 509404 -3744 510004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 473404 -3744 474004 707680 4 vccd2
port 533 nsew
rlabel metal4 s 469804 -1864 470404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 590020 -5624 590620 709560 4 vssa1
port 536 nsew
rlabel metal4 s 567004 -5624 567604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 531004 -5624 531604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 495004 -5624 495604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 426604 -7504 427204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 390604 -7504 391204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 354604 -7504 355204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 318604 -7504 319204 218000 4 vssa2
port 538 nsew
rlabel metal4 s 459004 -5624 459604 709560 4 vssa1
port 536 nsew
rlabel metal4 s 577804 -1864 578404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 585320 -924 585920 704860 4 vccd1
port 531 nsew
rlabel metal4 s 541804 -1864 542404 705800 4 vccd1
port 531 nsew
rlabel metal4 s 433804 -1864 434404 218000 4 vccd1
port 531 nsew
rlabel metal3 s 583520 391628 584960 391868 4 analog_io[2]
port 539 nsew
rlabel metal3 s 583520 444668 584960 444908 4 analog_io[3]
port 540 nsew
rlabel metal3 s 583520 497844 584960 498084 4 analog_io[4]
port 541 nsew
rlabel metal3 s 583520 551020 584960 551260 4 analog_io[5]
port 542 nsew
rlabel metal3 s 583520 604060 584960 604300 4 analog_io[6]
port 543 nsew
rlabel metal3 s 583520 657236 584960 657476 4 analog_io[7]
port 544 nsew
rlabel metal3 s 583520 457996 584960 458236 4 io_in[10]
port 545 nsew
rlabel metal3 s 583520 511172 584960 511412 4 io_in[11]
port 546 nsew
rlabel metal3 s 583520 564212 584960 564452 4 io_in[12]
port 547 nsew
rlabel metal3 s 583520 617388 584960 617628 4 io_in[13]
port 548 nsew
rlabel metal3 s 583520 670564 584960 670804 4 io_in[14]
port 549 nsew
rlabel metal3 s 583520 404820 584960 405060 4 io_in[9]
port 550 nsew
rlabel metal3 s 583520 484516 584960 484756 4 io_oeb[10]
port 551 nsew
rlabel metal3 s 583520 537692 584960 537932 4 io_oeb[11]
port 552 nsew
rlabel metal3 s 583520 590868 584960 591108 4 io_oeb[12]
port 553 nsew
rlabel metal3 s 583520 643908 584960 644148 4 io_oeb[13]
port 554 nsew
rlabel metal3 s 583520 697084 584960 697324 4 io_oeb[14]
port 555 nsew
rlabel metal3 s 583520 378300 584960 378540 4 io_oeb[8]
port 556 nsew
rlabel metal3 s 583520 431476 584960 431716 4 io_oeb[9]
port 557 nsew
rlabel metal3 s 583520 471324 584960 471564 4 io_out[10]
port 558 nsew
rlabel metal3 s 583520 524364 584960 524604 4 io_out[11]
port 559 nsew
rlabel metal3 s 583520 577540 584960 577780 4 io_out[12]
port 560 nsew
rlabel metal3 s 583520 630716 584960 630956 4 io_out[13]
port 561 nsew
rlabel metal3 s 583520 683756 584960 683996 4 io_out[14]
port 562 nsew
rlabel metal3 s 583520 364972 584960 365212 4 io_out[8]
port 563 nsew
rlabel metal3 s 583520 418148 584960 418388 4 io_out[9]
port 564 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 565 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 566 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 567 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 568 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 569 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 570 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 571 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 572 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 573 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 574 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 575 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 576 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 577 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 578 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 579 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 580 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 581 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 582 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 583 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 584 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 585 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 586 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 587 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 588 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 589 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 590 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 591 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 592 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 593 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 594 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 595 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 596 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 597 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 598 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 599 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 600 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 601 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 602 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 603 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 604 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 605 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 606 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 607 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 608 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 609 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 610 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 611 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 612 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 613 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 614 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 615 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 616 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 617 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 618 nsew
rlabel metal3 s 583520 351780 584960 352020 4 io_in[8]
port 619 nsew
rlabel metal3 s 583520 338452 584960 338692 4 analog_io[1]
port 620 nsew
rlabel metal3 s 583520 112692 584960 112932 4 io_oeb[2]
port 621 nsew
rlabel metal3 s 583520 32996 584960 33236 4 io_oeb[0]
port 622 nsew
rlabel metal3 s 583520 59516 584960 59756 4 io_out[1]
port 623 nsew
rlabel metal3 s 583520 86036 584960 86276 4 io_in[2]
port 624 nsew
rlabel metal3 s 583520 285276 584960 285516 4 analog_io[0]
port 625 nsew
rlabel metal3 s 583520 46188 584960 46428 4 io_in[1]
port 626 nsew
rlabel metal3 s 583520 6476 584960 6716 4 io_in[0]
port 627 nsew
rlabel metal3 s 583520 125884 584960 126124 4 io_in[3]
port 628 nsew
rlabel metal3 s 583520 72844 584960 73084 4 io_oeb[1]
port 629 nsew
rlabel metal3 s 583520 99364 584960 99604 4 io_out[2]
port 630 nsew
rlabel metal3 s 583520 165732 584960 165972 4 io_in[4]
port 631 nsew
rlabel metal3 s 583520 152540 584960 152780 4 io_oeb[3]
port 632 nsew
rlabel metal3 s 583520 192388 584960 192628 4 io_oeb[4]
port 633 nsew
rlabel metal3 s 583520 232236 584960 232476 4 io_oeb[5]
port 634 nsew
rlabel metal3 s 583520 272084 584960 272324 4 io_oeb[6]
port 635 nsew
rlabel metal3 s 583520 325124 584960 325364 4 io_oeb[7]
port 636 nsew
rlabel metal3 s 583520 205580 584960 205820 4 io_in[5]
port 637 nsew
rlabel metal3 s 583520 245428 584960 245668 4 io_in[6]
port 638 nsew
rlabel metal3 s 583520 139212 584960 139452 4 io_out[3]
port 639 nsew
rlabel metal3 s 583520 179060 584960 179300 4 io_out[4]
port 640 nsew
rlabel metal3 s 583520 218908 584960 219148 4 io_out[5]
port 641 nsew
rlabel metal3 s 583520 258756 584960 258996 4 io_out[6]
port 642 nsew
rlabel metal3 s 583520 311932 584960 312172 4 io_out[7]
port 643 nsew
rlabel metal3 s 583520 19668 584960 19908 4 io_out[0]
port 644 nsew
rlabel metal3 s 583520 298604 584960 298844 4 io_in[7]
port 645 nsew
rlabel metal5 s -1996 704260 585920 704860 4 vccd1
port 531 nsew
rlabel metal5 s -2936 686876 586860 687476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 650876 586860 651476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 614876 586860 615476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 578876 586860 579476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 542876 586860 543476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 506876 586860 507476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 470876 586860 471476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 434876 586860 435476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 398876 586860 399476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 362876 586860 363476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 705200 586860 705800 4 vssd1
port 532 nsew
rlabel metal5 s -2936 668876 586860 669476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 632876 586860 633476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 596876 586860 597476 4 vssd1
port 532 nsew
rlabel metal5 s 425267 560876 586860 561476 4 vssd1
port 532 nsew
rlabel metal5 s 425267 524876 586860 525476 4 vssd1
port 532 nsew
rlabel metal5 s 425267 488876 586860 489476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 452876 586860 453476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 416876 586860 417476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 380876 586860 381476 4 vssd1
port 532 nsew
rlabel metal5 s -3876 706140 587800 706740 4 vccd2
port 533 nsew
rlabel metal5 s -4816 690476 588740 691076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 654476 588740 655076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 618476 588740 619076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 582476 588740 583076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 546476 588740 547076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 510476 588740 511076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 474476 588740 475076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 438476 588740 439076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 402476 588740 403076 4 vccd2
port 533 nsew
rlabel metal5 s 448000 366476 588740 367076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 707080 588740 707680 4 vssd2
port 534 nsew
rlabel metal5 s -4816 672476 588740 673076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 636476 588740 637076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 600476 588740 601076 4 vssd2
port 534 nsew
rlabel metal5 s 407589 564476 588740 565076 4 vssd2
port 534 nsew
rlabel metal5 s 407589 528476 588740 529076 4 vssd2
port 534 nsew
rlabel metal5 s 407589 492476 588740 493076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 456476 588740 457076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 420476 588740 421076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 384476 588740 385076 4 vssd2
port 534 nsew
rlabel metal5 s -5756 708020 589680 708620 4 vdda1
port 535 nsew
rlabel metal5 s -6696 694076 590620 694676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 658076 590620 658676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 622076 590620 622676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 586076 590620 586676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 550076 590620 550676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 514076 590620 514676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 478076 590620 478676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 442076 590620 442676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 406076 590620 406676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 370076 590620 370676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 708960 590620 709560 4 vssa1
port 536 nsew
rlabel metal5 s -6696 676076 590620 676676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 640076 590620 640676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 604076 590620 604676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 568076 590620 568676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 532076 590620 532676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 496076 590620 496676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 460076 590620 460676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 424076 590620 424676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 388076 590620 388676 4 vssa1
port 536 nsew
rlabel metal5 s 448000 352076 590620 352676 4 vssa1
port 536 nsew
rlabel metal5 s -7636 709900 591560 710500 4 vdda2
port 537 nsew
rlabel metal5 s -8576 697676 592500 698276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 661676 592500 662276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 625676 592500 626276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 589676 592500 590276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 553676 592500 554276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 517676 592500 518276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 481676 592500 482276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 445676 592500 446276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 409676 592500 410276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 373676 592500 374276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 710840 592500 711440 4 vssa2
port 538 nsew
rlabel metal5 s -8576 679676 592500 680276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 643676 592500 644276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 607676 592500 608276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 571676 592500 572276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 535676 592500 536276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 499676 592500 500276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 463676 592500 464276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 427676 592500 428276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 391676 592500 392276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 355676 592500 356276 4 vssa2
port 538 nsew
rlabel metal5 s -6696 370076 108000 370676 4 vdda1
port 535 nsew
rlabel metal5 s -2936 416876 108000 417476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 434876 108000 435476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 380876 108000 381476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 506876 151560 507476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 596876 108000 597476 4 vssd1
port 532 nsew
rlabel metal5 s -6696 568076 108000 568676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 564476 108000 565076 4 vssd2
port 534 nsew
rlabel metal5 s -6696 532076 108000 532676 4 vssa1
port 536 nsew
rlabel metal5 s -2936 398876 108000 399476 4 vccd1
port 531 nsew
rlabel metal5 s -6696 496076 108000 496676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 528476 108000 529076 4 vssd2
port 534 nsew
rlabel metal5 s -6696 460076 108000 460676 4 vssa1
port 536 nsew
rlabel metal5 s -2936 560876 108000 561476 4 vssd1
port 532 nsew
rlabel metal5 s -6696 424076 108000 424676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 492476 108000 493076 4 vssd2
port 534 nsew
rlabel metal5 s -6696 388076 108000 388676 4 vssa1
port 536 nsew
rlabel metal5 s -2936 542876 151560 543476 4 vccd1
port 531 nsew
rlabel metal5 s -6696 352076 108000 352676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 456476 108000 457076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 582476 133883 583076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 420476 108000 421076 4 vssd2
port 534 nsew
rlabel metal5 s -2936 524876 108000 525476 4 vssd1
port 532 nsew
rlabel metal5 s -4816 384476 108000 385076 4 vssd2
port 534 nsew
rlabel metal5 s -8576 589676 108000 590276 4 vdda2
port 537 nsew
rlabel metal5 s -4816 546476 133883 547076 4 vccd2
port 533 nsew
rlabel metal5 s -8576 553676 108000 554276 4 vdda2
port 537 nsew
rlabel metal5 s -2936 362876 108000 363476 4 vccd1
port 531 nsew
rlabel metal5 s -8576 517676 108000 518276 4 vdda2
port 537 nsew
rlabel metal5 s -4816 510476 133883 511076 4 vccd2
port 533 nsew
rlabel metal5 s -8576 481676 108000 482276 4 vdda2
port 537 nsew
rlabel metal5 s -2936 488876 108000 489476 4 vssd1
port 532 nsew
rlabel metal5 s -8576 445676 108000 446276 4 vdda2
port 537 nsew
rlabel metal5 s -4816 474476 108000 475076 4 vccd2
port 533 nsew
rlabel metal5 s -8576 409676 108000 410276 4 vdda2
port 537 nsew
rlabel metal5 s -6696 586076 108000 586676 4 vdda1
port 535 nsew
rlabel metal5 s -8576 373676 108000 374276 4 vdda2
port 537 nsew
rlabel metal5 s -2936 470876 108000 471476 4 vccd1
port 531 nsew
rlabel metal5 s -6696 550076 108000 550676 4 vdda1
port 535 nsew
rlabel metal5 s -4816 438476 108000 439076 4 vccd2
port 533 nsew
rlabel metal5 s -6696 514076 108000 514676 4 vdda1
port 535 nsew
rlabel metal5 s -2936 452876 108000 453476 4 vssd1
port 532 nsew
rlabel metal5 s -8576 571676 108000 572276 4 vssa2
port 538 nsew
rlabel metal5 s -6696 478076 108000 478676 4 vdda1
port 535 nsew
rlabel metal5 s -8576 535676 108000 536276 4 vssa2
port 538 nsew
rlabel metal5 s -4816 402476 108000 403076 4 vccd2
port 533 nsew
rlabel metal5 s -8576 499676 108000 500276 4 vssa2
port 538 nsew
rlabel metal5 s -6696 442076 108000 442676 4 vdda1
port 535 nsew
rlabel metal5 s -8576 463676 108000 464276 4 vssa2
port 538 nsew
rlabel metal5 s -2936 578876 151560 579476 4 vccd1
port 531 nsew
rlabel metal5 s -8576 427676 108000 428276 4 vssa2
port 538 nsew
rlabel metal5 s -6696 406076 108000 406676 4 vdda1
port 535 nsew
rlabel metal5 s -8576 391676 108000 392276 4 vssa2
port 538 nsew
rlabel metal5 s -4816 366476 108000 367076 4 vccd2
port 533 nsew
rlabel metal5 s -8576 355676 108000 356276 4 vssa2
port 538 nsew
rlabel metal5 s -4816 312476 108000 313076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 276476 108000 277076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 240476 108000 241076 4 vssd2
port 534 nsew
rlabel metal5 s -2936 272876 108000 273476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 236876 108000 237476 4 vssd1
port 532 nsew
rlabel metal5 s -8576 337676 108000 338276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 301676 108000 302276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 265676 108000 266276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 229676 108000 230276 4 vdda2
port 537 nsew
rlabel metal5 s -6696 334076 108000 334676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 298076 108000 298676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 316076 108000 316676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 280076 108000 280676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 244076 108000 244676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 262076 108000 262676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 226076 108000 226676 4 vdda1
port 535 nsew
rlabel metal5 s -2936 290876 151560 291476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 254876 151560 255476 4 vccd1
port 531 nsew
rlabel metal5 s -4816 330476 133883 331076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 294476 133883 295076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 258476 133883 259076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 222476 108000 223076 4 vccd2
port 533 nsew
rlabel metal5 s -2936 218876 108000 219476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 326876 151560 327476 4 vccd1
port 531 nsew
rlabel metal5 s -2936 344876 108000 345476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 308876 108000 309476 4 vssd1
port 532 nsew
rlabel metal5 s -4816 348476 108000 349076 4 vssd2
port 534 nsew
rlabel metal5 s -8576 319676 108000 320276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 283676 108000 284276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 247676 108000 248276 4 vssa2
port 538 nsew
rlabel metal5 s 407589 312476 588740 313076 4 vssd2
port 534 nsew
rlabel metal5 s -2936 128876 586860 129476 4 vssd1
port 532 nsew
rlabel metal5 s 407589 276476 588740 277076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 330476 588740 331076 4 vccd2
port 533 nsew
rlabel metal5 s 407589 240476 588740 241076 4 vssd2
port 534 nsew
rlabel metal5 s -2936 92876 586860 93476 4 vssd1
port 532 nsew
rlabel metal5 s -4816 204476 588740 205076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 168476 588740 169076 4 vssd2
port 534 nsew
rlabel metal5 s -4816 132476 588740 133076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 316076 590620 316676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 96476 588740 97076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 280076 590620 280676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 60476 588740 61076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 244076 590620 244676 4 vssa1
port 536 nsew
rlabel metal5 s -4816 24476 588740 25076 4 vssd2
port 534 nsew
rlabel metal5 s -6696 208076 590620 208676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 172076 590620 172676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 136076 590620 136676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 100076 590620 100676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 64076 590620 64676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 28076 590620 28676 4 vssa1
port 536 nsew
rlabel metal5 s -6696 -5624 590620 -5024 4 vssa1
port 536 nsew
rlabel metal5 s -4816 -3744 588740 -3144 4 vssd2
port 534 nsew
rlabel metal5 s 448000 294476 588740 295076 4 vccd2
port 533 nsew
rlabel metal5 s -2936 56876 586860 57476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 258476 588740 259076 4 vccd2
port 533 nsew
rlabel metal5 s -2936 20876 586860 21476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 222476 588740 223076 4 vccd2
port 533 nsew
rlabel metal5 s -2936 -1864 586860 -1264 4 vssd1
port 532 nsew
rlabel metal5 s -4816 186476 588740 187076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 150476 588740 151076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 114476 588740 115076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 78476 588740 79076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 42476 588740 43076 4 vccd2
port 533 nsew
rlabel metal5 s -4816 6476 588740 7076 4 vccd2
port 533 nsew
rlabel metal5 s -3876 -2804 587800 -2204 4 vccd2
port 533 nsew
rlabel metal5 s -1996 -924 585920 -324 4 vccd1
port 531 nsew
rlabel metal5 s 448000 254876 586860 255476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 290876 586860 291476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 218876 586860 219476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 337676 592500 338276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 326876 586860 327476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 301676 592500 302276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 334076 590620 334676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 265676 592500 266276 4 vdda2
port 537 nsew
rlabel metal5 s -2936 182876 586860 183476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 229676 592500 230276 4 vdda2
port 537 nsew
rlabel metal5 s 448000 298076 590620 298676 4 vdda1
port 535 nsew
rlabel metal5 s -8576 193676 592500 194276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 157676 592500 158276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 121676 592500 122276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 85676 592500 86276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 49676 592500 50276 4 vdda2
port 537 nsew
rlabel metal5 s -8576 13676 592500 14276 4 vdda2
port 537 nsew
rlabel metal5 s -7636 -6564 591560 -5964 4 vdda2
port 537 nsew
rlabel metal5 s -2936 146876 586860 147476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 262076 590620 262676 4 vdda1
port 535 nsew
rlabel metal5 s 448000 344876 586860 345476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 226076 590620 226676 4 vdda1
port 535 nsew
rlabel metal5 s -2936 110876 586860 111476 4 vccd1
port 531 nsew
rlabel metal5 s -6696 190076 590620 190676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 154076 590620 154676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 118076 590620 118676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 82076 590620 82676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 46076 590620 46676 4 vdda1
port 535 nsew
rlabel metal5 s -6696 10076 590620 10676 4 vdda1
port 535 nsew
rlabel metal5 s -5756 -4684 589680 -4084 4 vdda1
port 535 nsew
rlabel metal5 s 425267 308876 586860 309476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 74876 586860 75476 4 vccd1
port 531 nsew
rlabel metal5 s 425267 272876 586860 273476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 38876 586860 39476 4 vccd1
port 531 nsew
rlabel metal5 s 425267 236876 586860 237476 4 vssd1
port 532 nsew
rlabel metal5 s -2936 2876 586860 3476 4 vccd1
port 531 nsew
rlabel metal5 s 448000 319676 592500 320276 4 vssa2
port 538 nsew
rlabel metal5 s -2936 200876 586860 201476 4 vssd1
port 532 nsew
rlabel metal5 s 448000 283676 592500 284276 4 vssa2
port 538 nsew
rlabel metal5 s 448000 348476 588740 349076 4 vssd2
port 534 nsew
rlabel metal5 s 448000 247676 592500 248276 4 vssa2
port 538 nsew
rlabel metal5 s -2936 164876 586860 165476 4 vssd1
port 532 nsew
rlabel metal5 s -8576 211676 592500 212276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 175676 592500 176276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 139676 592500 140276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 103676 592500 104276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 67676 592500 68276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 31676 592500 32276 4 vssa2
port 538 nsew
rlabel metal5 s -8576 -7504 592500 -6904 4 vssa2
port 538 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string GDS_FILE user_project_wrapper.gds
string GDS_END 15555190
string GDS_START 13561098
<< end >>
