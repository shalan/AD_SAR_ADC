magic
tech sky130A
magscale 1 2
timestamp 1626382392
<< obsli1 >>
rect 1104 2159 259043 157777
<< obsm1 >>
rect 198 1164 259702 158228
<< metal2 >>
rect 3606 159200 3662 160000
rect 10782 159200 10838 160000
rect 18050 159200 18106 160000
rect 25226 159200 25282 160000
rect 32494 159200 32550 160000
rect 39670 159200 39726 160000
rect 46938 159200 46994 160000
rect 54114 159200 54170 160000
rect 61382 159200 61438 160000
rect 68558 159200 68614 160000
rect 75826 159200 75882 160000
rect 83002 159200 83058 160000
rect 90270 159200 90326 160000
rect 97446 159200 97502 160000
rect 104714 159200 104770 160000
rect 111890 159200 111946 160000
rect 119158 159200 119214 160000
rect 126334 159200 126390 160000
rect 133602 159200 133658 160000
rect 140778 159200 140834 160000
rect 148046 159200 148102 160000
rect 155222 159200 155278 160000
rect 162490 159200 162546 160000
rect 169666 159200 169722 160000
rect 176934 159200 176990 160000
rect 184110 159200 184166 160000
rect 191378 159200 191434 160000
rect 198554 159200 198610 160000
rect 205822 159200 205878 160000
rect 212998 159200 213054 160000
rect 220266 159200 220322 160000
rect 227442 159200 227498 160000
rect 234710 159200 234766 160000
rect 241886 159200 241942 160000
rect 249154 159200 249210 160000
rect 256330 159200 256386 160000
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2778 0 2834 800
rect 3330 0 3386 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8022 0 8078 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 10138 0 10194 800
rect 10690 0 10746 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12254 0 12310 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19614 0 19670 800
rect 20166 0 20222 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21730 0 21786 800
rect 22282 0 22338 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25410 0 25466 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30654 0 30710 800
rect 31206 0 31262 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 35990 0 36046 800
rect 36450 0 36506 800
rect 37002 0 37058 800
rect 37554 0 37610 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40682 0 40738 800
rect 41234 0 41290 800
rect 41694 0 41750 800
rect 42246 0 42302 800
rect 42798 0 42854 800
rect 43350 0 43406 800
rect 43810 0 43866 800
rect 44362 0 44418 800
rect 44914 0 44970 800
rect 45374 0 45430 800
rect 45926 0 45982 800
rect 46478 0 46534 800
rect 47030 0 47086 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54390 0 54446 800
rect 54850 0 54906 800
rect 55402 0 55458 800
rect 55954 0 56010 800
rect 56506 0 56562 800
rect 56966 0 57022 800
rect 57518 0 57574 800
rect 58070 0 58126 800
rect 58530 0 58586 800
rect 59082 0 59138 800
rect 59634 0 59690 800
rect 60186 0 60242 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63866 0 63922 800
rect 64326 0 64382 800
rect 64878 0 64934 800
rect 65430 0 65486 800
rect 65982 0 66038 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68006 0 68062 800
rect 68558 0 68614 800
rect 69110 0 69166 800
rect 69662 0 69718 800
rect 70122 0 70178 800
rect 70674 0 70730 800
rect 71226 0 71282 800
rect 71778 0 71834 800
rect 72238 0 72294 800
rect 72790 0 72846 800
rect 73342 0 73398 800
rect 73802 0 73858 800
rect 74354 0 74410 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76470 0 76526 800
rect 77022 0 77078 800
rect 77482 0 77538 800
rect 78034 0 78090 800
rect 78586 0 78642 800
rect 79138 0 79194 800
rect 79598 0 79654 800
rect 80150 0 80206 800
rect 80702 0 80758 800
rect 81162 0 81218 800
rect 81714 0 81770 800
rect 82266 0 82322 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83830 0 83886 800
rect 84382 0 84438 800
rect 84934 0 84990 800
rect 85394 0 85450 800
rect 85946 0 86002 800
rect 86498 0 86554 800
rect 86958 0 87014 800
rect 87510 0 87566 800
rect 88062 0 88118 800
rect 88614 0 88670 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90638 0 90694 800
rect 91190 0 91246 800
rect 91742 0 91798 800
rect 92294 0 92350 800
rect 92754 0 92810 800
rect 93306 0 93362 800
rect 93858 0 93914 800
rect 94318 0 94374 800
rect 94870 0 94926 800
rect 95422 0 95478 800
rect 95974 0 96030 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97538 0 97594 800
rect 98090 0 98146 800
rect 98550 0 98606 800
rect 99102 0 99158 800
rect 99654 0 99710 800
rect 100114 0 100170 800
rect 100666 0 100722 800
rect 101218 0 101274 800
rect 101770 0 101826 800
rect 102230 0 102286 800
rect 102782 0 102838 800
rect 103334 0 103390 800
rect 103794 0 103850 800
rect 104346 0 104402 800
rect 104898 0 104954 800
rect 105450 0 105506 800
rect 105910 0 105966 800
rect 106462 0 106518 800
rect 107014 0 107070 800
rect 107566 0 107622 800
rect 108026 0 108082 800
rect 108578 0 108634 800
rect 109130 0 109186 800
rect 109590 0 109646 800
rect 110142 0 110198 800
rect 110694 0 110750 800
rect 111246 0 111302 800
rect 111706 0 111762 800
rect 112258 0 112314 800
rect 112810 0 112866 800
rect 113270 0 113326 800
rect 113822 0 113878 800
rect 114374 0 114430 800
rect 114926 0 114982 800
rect 115386 0 115442 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 118054 0 118110 800
rect 118606 0 118662 800
rect 119066 0 119122 800
rect 119618 0 119674 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121182 0 121238 800
rect 121734 0 121790 800
rect 122286 0 122342 800
rect 122746 0 122802 800
rect 123298 0 123354 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 125966 0 126022 800
rect 126426 0 126482 800
rect 126978 0 127034 800
rect 127530 0 127586 800
rect 128082 0 128138 800
rect 128542 0 128598 800
rect 129094 0 129150 800
rect 129646 0 129702 800
rect 130198 0 130254 800
rect 130658 0 130714 800
rect 131210 0 131266 800
rect 131762 0 131818 800
rect 132222 0 132278 800
rect 132774 0 132830 800
rect 133326 0 133382 800
rect 133878 0 133934 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135902 0 135958 800
rect 136454 0 136510 800
rect 137006 0 137062 800
rect 137558 0 137614 800
rect 138018 0 138074 800
rect 138570 0 138626 800
rect 139122 0 139178 800
rect 139582 0 139638 800
rect 140134 0 140190 800
rect 140686 0 140742 800
rect 141238 0 141294 800
rect 141698 0 141754 800
rect 142250 0 142306 800
rect 142802 0 142858 800
rect 143354 0 143410 800
rect 143814 0 143870 800
rect 144366 0 144422 800
rect 144918 0 144974 800
rect 145378 0 145434 800
rect 145930 0 145986 800
rect 146482 0 146538 800
rect 147034 0 147090 800
rect 147494 0 147550 800
rect 148046 0 148102 800
rect 148598 0 148654 800
rect 149058 0 149114 800
rect 149610 0 149666 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152278 0 152334 800
rect 152738 0 152794 800
rect 153290 0 153346 800
rect 153842 0 153898 800
rect 154394 0 154450 800
rect 154854 0 154910 800
rect 155406 0 155462 800
rect 155958 0 156014 800
rect 156510 0 156566 800
rect 156970 0 157026 800
rect 157522 0 157578 800
rect 158074 0 158130 800
rect 158534 0 158590 800
rect 159086 0 159142 800
rect 159638 0 159694 800
rect 160190 0 160246 800
rect 160650 0 160706 800
rect 161202 0 161258 800
rect 161754 0 161810 800
rect 162214 0 162270 800
rect 162766 0 162822 800
rect 163318 0 163374 800
rect 163870 0 163926 800
rect 164330 0 164386 800
rect 164882 0 164938 800
rect 165434 0 165490 800
rect 165986 0 166042 800
rect 166446 0 166502 800
rect 166998 0 167054 800
rect 167550 0 167606 800
rect 168010 0 168066 800
rect 168562 0 168618 800
rect 169114 0 169170 800
rect 169666 0 169722 800
rect 170126 0 170182 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171690 0 171746 800
rect 172242 0 172298 800
rect 172794 0 172850 800
rect 173346 0 173402 800
rect 173806 0 173862 800
rect 174358 0 174414 800
rect 174910 0 174966 800
rect 175370 0 175426 800
rect 175922 0 175978 800
rect 176474 0 176530 800
rect 177026 0 177082 800
rect 177486 0 177542 800
rect 178038 0 178094 800
rect 178590 0 178646 800
rect 179142 0 179198 800
rect 179602 0 179658 800
rect 180154 0 180210 800
rect 180706 0 180762 800
rect 181166 0 181222 800
rect 181718 0 181774 800
rect 182270 0 182326 800
rect 182822 0 182878 800
rect 183282 0 183338 800
rect 183834 0 183890 800
rect 184386 0 184442 800
rect 184846 0 184902 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186502 0 186558 800
rect 186962 0 187018 800
rect 187514 0 187570 800
rect 188066 0 188122 800
rect 188526 0 188582 800
rect 189078 0 189134 800
rect 189630 0 189686 800
rect 190182 0 190238 800
rect 190642 0 190698 800
rect 191194 0 191250 800
rect 191746 0 191802 800
rect 192298 0 192354 800
rect 192758 0 192814 800
rect 193310 0 193366 800
rect 193862 0 193918 800
rect 194322 0 194378 800
rect 194874 0 194930 800
rect 195426 0 195482 800
rect 195978 0 196034 800
rect 196438 0 196494 800
rect 196990 0 197046 800
rect 197542 0 197598 800
rect 198002 0 198058 800
rect 198554 0 198610 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200118 0 200174 800
rect 200670 0 200726 800
rect 201222 0 201278 800
rect 201774 0 201830 800
rect 202234 0 202290 800
rect 202786 0 202842 800
rect 203338 0 203394 800
rect 203798 0 203854 800
rect 204350 0 204406 800
rect 204902 0 204958 800
rect 205454 0 205510 800
rect 205914 0 205970 800
rect 206466 0 206522 800
rect 207018 0 207074 800
rect 207478 0 207534 800
rect 208030 0 208086 800
rect 208582 0 208638 800
rect 209134 0 209190 800
rect 209594 0 209650 800
rect 210146 0 210202 800
rect 210698 0 210754 800
rect 211158 0 211214 800
rect 211710 0 211766 800
rect 212262 0 212318 800
rect 212814 0 212870 800
rect 213274 0 213330 800
rect 213826 0 213882 800
rect 214378 0 214434 800
rect 214930 0 214986 800
rect 215390 0 215446 800
rect 215942 0 215998 800
rect 216494 0 216550 800
rect 216954 0 217010 800
rect 217506 0 217562 800
rect 218058 0 218114 800
rect 218610 0 218666 800
rect 219070 0 219126 800
rect 219622 0 219678 800
rect 220174 0 220230 800
rect 220634 0 220690 800
rect 221186 0 221242 800
rect 221738 0 221794 800
rect 222290 0 222346 800
rect 222750 0 222806 800
rect 223302 0 223358 800
rect 223854 0 223910 800
rect 224314 0 224370 800
rect 224866 0 224922 800
rect 225418 0 225474 800
rect 225970 0 226026 800
rect 226430 0 226486 800
rect 226982 0 227038 800
rect 227534 0 227590 800
rect 228086 0 228142 800
rect 228546 0 228602 800
rect 229098 0 229154 800
rect 229650 0 229706 800
rect 230110 0 230166 800
rect 230662 0 230718 800
rect 231214 0 231270 800
rect 231766 0 231822 800
rect 232226 0 232282 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234894 0 234950 800
rect 235446 0 235502 800
rect 235906 0 235962 800
rect 236458 0 236514 800
rect 237010 0 237066 800
rect 237562 0 237618 800
rect 238022 0 238078 800
rect 238574 0 238630 800
rect 239126 0 239182 800
rect 239586 0 239642 800
rect 240138 0 240194 800
rect 240690 0 240746 800
rect 241242 0 241298 800
rect 241702 0 241758 800
rect 242254 0 242310 800
rect 242806 0 242862 800
rect 243266 0 243322 800
rect 243818 0 243874 800
rect 244370 0 244426 800
rect 244922 0 244978 800
rect 245382 0 245438 800
rect 245934 0 245990 800
rect 246486 0 246542 800
rect 246946 0 247002 800
rect 247498 0 247554 800
rect 248050 0 248106 800
rect 248602 0 248658 800
rect 249062 0 249118 800
rect 249614 0 249670 800
rect 250166 0 250222 800
rect 250718 0 250774 800
rect 251178 0 251234 800
rect 251730 0 251786 800
rect 252282 0 252338 800
rect 252742 0 252798 800
rect 253294 0 253350 800
rect 253846 0 253902 800
rect 254398 0 254454 800
rect 254858 0 254914 800
rect 255410 0 255466 800
rect 255962 0 256018 800
rect 256422 0 256478 800
rect 256974 0 257030 800
rect 257526 0 257582 800
rect 258078 0 258134 800
rect 258538 0 258594 800
rect 259090 0 259146 800
rect 259642 0 259698 800
<< obsm2 >>
rect 204 159144 3550 159200
rect 3718 159144 10726 159200
rect 10894 159144 17994 159200
rect 18162 159144 25170 159200
rect 25338 159144 32438 159200
rect 32606 159144 39614 159200
rect 39782 159144 46882 159200
rect 47050 159144 54058 159200
rect 54226 159144 61326 159200
rect 61494 159144 68502 159200
rect 68670 159144 75770 159200
rect 75938 159144 82946 159200
rect 83114 159144 90214 159200
rect 90382 159144 97390 159200
rect 97558 159144 104658 159200
rect 104826 159144 111834 159200
rect 112002 159144 119102 159200
rect 119270 159144 126278 159200
rect 126446 159144 133546 159200
rect 133714 159144 140722 159200
rect 140890 159144 147990 159200
rect 148158 159144 155166 159200
rect 155334 159144 162434 159200
rect 162602 159144 169610 159200
rect 169778 159144 176878 159200
rect 177046 159144 184054 159200
rect 184222 159144 191322 159200
rect 191490 159144 198498 159200
rect 198666 159144 205766 159200
rect 205934 159144 212942 159200
rect 213110 159144 220210 159200
rect 220378 159144 227386 159200
rect 227554 159144 234654 159200
rect 234822 159144 241830 159200
rect 241998 159144 249098 159200
rect 249266 159144 256274 159200
rect 256442 159144 259696 159200
rect 204 856 259696 159144
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1710 856
rect 1878 800 2170 856
rect 2338 800 2722 856
rect 2890 800 3274 856
rect 3442 800 3826 856
rect 3994 800 4286 856
rect 4454 800 4838 856
rect 5006 800 5390 856
rect 5558 800 5850 856
rect 6018 800 6402 856
rect 6570 800 6954 856
rect 7122 800 7506 856
rect 7674 800 7966 856
rect 8134 800 8518 856
rect 8686 800 9070 856
rect 9238 800 9530 856
rect 9698 800 10082 856
rect 10250 800 10634 856
rect 10802 800 11186 856
rect 11354 800 11646 856
rect 11814 800 12198 856
rect 12366 800 12750 856
rect 12918 800 13302 856
rect 13470 800 13762 856
rect 13930 800 14314 856
rect 14482 800 14866 856
rect 15034 800 15326 856
rect 15494 800 15878 856
rect 16046 800 16430 856
rect 16598 800 16982 856
rect 17150 800 17442 856
rect 17610 800 17994 856
rect 18162 800 18546 856
rect 18714 800 19006 856
rect 19174 800 19558 856
rect 19726 800 20110 856
rect 20278 800 20662 856
rect 20830 800 21122 856
rect 21290 800 21674 856
rect 21842 800 22226 856
rect 22394 800 22686 856
rect 22854 800 23238 856
rect 23406 800 23790 856
rect 23958 800 24342 856
rect 24510 800 24802 856
rect 24970 800 25354 856
rect 25522 800 25906 856
rect 26074 800 26458 856
rect 26626 800 26918 856
rect 27086 800 27470 856
rect 27638 800 28022 856
rect 28190 800 28482 856
rect 28650 800 29034 856
rect 29202 800 29586 856
rect 29754 800 30138 856
rect 30306 800 30598 856
rect 30766 800 31150 856
rect 31318 800 31702 856
rect 31870 800 32162 856
rect 32330 800 32714 856
rect 32882 800 33266 856
rect 33434 800 33818 856
rect 33986 800 34278 856
rect 34446 800 34830 856
rect 34998 800 35382 856
rect 35550 800 35934 856
rect 36102 800 36394 856
rect 36562 800 36946 856
rect 37114 800 37498 856
rect 37666 800 37958 856
rect 38126 800 38510 856
rect 38678 800 39062 856
rect 39230 800 39614 856
rect 39782 800 40074 856
rect 40242 800 40626 856
rect 40794 800 41178 856
rect 41346 800 41638 856
rect 41806 800 42190 856
rect 42358 800 42742 856
rect 42910 800 43294 856
rect 43462 800 43754 856
rect 43922 800 44306 856
rect 44474 800 44858 856
rect 45026 800 45318 856
rect 45486 800 45870 856
rect 46038 800 46422 856
rect 46590 800 46974 856
rect 47142 800 47434 856
rect 47602 800 47986 856
rect 48154 800 48538 856
rect 48706 800 49090 856
rect 49258 800 49550 856
rect 49718 800 50102 856
rect 50270 800 50654 856
rect 50822 800 51114 856
rect 51282 800 51666 856
rect 51834 800 52218 856
rect 52386 800 52770 856
rect 52938 800 53230 856
rect 53398 800 53782 856
rect 53950 800 54334 856
rect 54502 800 54794 856
rect 54962 800 55346 856
rect 55514 800 55898 856
rect 56066 800 56450 856
rect 56618 800 56910 856
rect 57078 800 57462 856
rect 57630 800 58014 856
rect 58182 800 58474 856
rect 58642 800 59026 856
rect 59194 800 59578 856
rect 59746 800 60130 856
rect 60298 800 60590 856
rect 60758 800 61142 856
rect 61310 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62706 856
rect 62874 800 63258 856
rect 63426 800 63810 856
rect 63978 800 64270 856
rect 64438 800 64822 856
rect 64990 800 65374 856
rect 65542 800 65926 856
rect 66094 800 66386 856
rect 66554 800 66938 856
rect 67106 800 67490 856
rect 67658 800 67950 856
rect 68118 800 68502 856
rect 68670 800 69054 856
rect 69222 800 69606 856
rect 69774 800 70066 856
rect 70234 800 70618 856
rect 70786 800 71170 856
rect 71338 800 71722 856
rect 71890 800 72182 856
rect 72350 800 72734 856
rect 72902 800 73286 856
rect 73454 800 73746 856
rect 73914 800 74298 856
rect 74466 800 74850 856
rect 75018 800 75402 856
rect 75570 800 75862 856
rect 76030 800 76414 856
rect 76582 800 76966 856
rect 77134 800 77426 856
rect 77594 800 77978 856
rect 78146 800 78530 856
rect 78698 800 79082 856
rect 79250 800 79542 856
rect 79710 800 80094 856
rect 80262 800 80646 856
rect 80814 800 81106 856
rect 81274 800 81658 856
rect 81826 800 82210 856
rect 82378 800 82762 856
rect 82930 800 83222 856
rect 83390 800 83774 856
rect 83942 800 84326 856
rect 84494 800 84878 856
rect 85046 800 85338 856
rect 85506 800 85890 856
rect 86058 800 86442 856
rect 86610 800 86902 856
rect 87070 800 87454 856
rect 87622 800 88006 856
rect 88174 800 88558 856
rect 88726 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90122 856
rect 90290 800 90582 856
rect 90750 800 91134 856
rect 91302 800 91686 856
rect 91854 800 92238 856
rect 92406 800 92698 856
rect 92866 800 93250 856
rect 93418 800 93802 856
rect 93970 800 94262 856
rect 94430 800 94814 856
rect 94982 800 95366 856
rect 95534 800 95918 856
rect 96086 800 96378 856
rect 96546 800 96930 856
rect 97098 800 97482 856
rect 97650 800 98034 856
rect 98202 800 98494 856
rect 98662 800 99046 856
rect 99214 800 99598 856
rect 99766 800 100058 856
rect 100226 800 100610 856
rect 100778 800 101162 856
rect 101330 800 101714 856
rect 101882 800 102174 856
rect 102342 800 102726 856
rect 102894 800 103278 856
rect 103446 800 103738 856
rect 103906 800 104290 856
rect 104458 800 104842 856
rect 105010 800 105394 856
rect 105562 800 105854 856
rect 106022 800 106406 856
rect 106574 800 106958 856
rect 107126 800 107510 856
rect 107678 800 107970 856
rect 108138 800 108522 856
rect 108690 800 109074 856
rect 109242 800 109534 856
rect 109702 800 110086 856
rect 110254 800 110638 856
rect 110806 800 111190 856
rect 111358 800 111650 856
rect 111818 800 112202 856
rect 112370 800 112754 856
rect 112922 800 113214 856
rect 113382 800 113766 856
rect 113934 800 114318 856
rect 114486 800 114870 856
rect 115038 800 115330 856
rect 115498 800 115882 856
rect 116050 800 116434 856
rect 116602 800 116894 856
rect 117062 800 117446 856
rect 117614 800 117998 856
rect 118166 800 118550 856
rect 118718 800 119010 856
rect 119178 800 119562 856
rect 119730 800 120114 856
rect 120282 800 120666 856
rect 120834 800 121126 856
rect 121294 800 121678 856
rect 121846 800 122230 856
rect 122398 800 122690 856
rect 122858 800 123242 856
rect 123410 800 123794 856
rect 123962 800 124346 856
rect 124514 800 124806 856
rect 124974 800 125358 856
rect 125526 800 125910 856
rect 126078 800 126370 856
rect 126538 800 126922 856
rect 127090 800 127474 856
rect 127642 800 128026 856
rect 128194 800 128486 856
rect 128654 800 129038 856
rect 129206 800 129590 856
rect 129758 800 130142 856
rect 130310 800 130602 856
rect 130770 800 131154 856
rect 131322 800 131706 856
rect 131874 800 132166 856
rect 132334 800 132718 856
rect 132886 800 133270 856
rect 133438 800 133822 856
rect 133990 800 134282 856
rect 134450 800 134834 856
rect 135002 800 135386 856
rect 135554 800 135846 856
rect 136014 800 136398 856
rect 136566 800 136950 856
rect 137118 800 137502 856
rect 137670 800 137962 856
rect 138130 800 138514 856
rect 138682 800 139066 856
rect 139234 800 139526 856
rect 139694 800 140078 856
rect 140246 800 140630 856
rect 140798 800 141182 856
rect 141350 800 141642 856
rect 141810 800 142194 856
rect 142362 800 142746 856
rect 142914 800 143298 856
rect 143466 800 143758 856
rect 143926 800 144310 856
rect 144478 800 144862 856
rect 145030 800 145322 856
rect 145490 800 145874 856
rect 146042 800 146426 856
rect 146594 800 146978 856
rect 147146 800 147438 856
rect 147606 800 147990 856
rect 148158 800 148542 856
rect 148710 800 149002 856
rect 149170 800 149554 856
rect 149722 800 150106 856
rect 150274 800 150658 856
rect 150826 800 151118 856
rect 151286 800 151670 856
rect 151838 800 152222 856
rect 152390 800 152682 856
rect 152850 800 153234 856
rect 153402 800 153786 856
rect 153954 800 154338 856
rect 154506 800 154798 856
rect 154966 800 155350 856
rect 155518 800 155902 856
rect 156070 800 156454 856
rect 156622 800 156914 856
rect 157082 800 157466 856
rect 157634 800 158018 856
rect 158186 800 158478 856
rect 158646 800 159030 856
rect 159198 800 159582 856
rect 159750 800 160134 856
rect 160302 800 160594 856
rect 160762 800 161146 856
rect 161314 800 161698 856
rect 161866 800 162158 856
rect 162326 800 162710 856
rect 162878 800 163262 856
rect 163430 800 163814 856
rect 163982 800 164274 856
rect 164442 800 164826 856
rect 164994 800 165378 856
rect 165546 800 165930 856
rect 166098 800 166390 856
rect 166558 800 166942 856
rect 167110 800 167494 856
rect 167662 800 167954 856
rect 168122 800 168506 856
rect 168674 800 169058 856
rect 169226 800 169610 856
rect 169778 800 170070 856
rect 170238 800 170622 856
rect 170790 800 171174 856
rect 171342 800 171634 856
rect 171802 800 172186 856
rect 172354 800 172738 856
rect 172906 800 173290 856
rect 173458 800 173750 856
rect 173918 800 174302 856
rect 174470 800 174854 856
rect 175022 800 175314 856
rect 175482 800 175866 856
rect 176034 800 176418 856
rect 176586 800 176970 856
rect 177138 800 177430 856
rect 177598 800 177982 856
rect 178150 800 178534 856
rect 178702 800 179086 856
rect 179254 800 179546 856
rect 179714 800 180098 856
rect 180266 800 180650 856
rect 180818 800 181110 856
rect 181278 800 181662 856
rect 181830 800 182214 856
rect 182382 800 182766 856
rect 182934 800 183226 856
rect 183394 800 183778 856
rect 183946 800 184330 856
rect 184498 800 184790 856
rect 184958 800 185342 856
rect 185510 800 185894 856
rect 186062 800 186446 856
rect 186614 800 186906 856
rect 187074 800 187458 856
rect 187626 800 188010 856
rect 188178 800 188470 856
rect 188638 800 189022 856
rect 189190 800 189574 856
rect 189742 800 190126 856
rect 190294 800 190586 856
rect 190754 800 191138 856
rect 191306 800 191690 856
rect 191858 800 192242 856
rect 192410 800 192702 856
rect 192870 800 193254 856
rect 193422 800 193806 856
rect 193974 800 194266 856
rect 194434 800 194818 856
rect 194986 800 195370 856
rect 195538 800 195922 856
rect 196090 800 196382 856
rect 196550 800 196934 856
rect 197102 800 197486 856
rect 197654 800 197946 856
rect 198114 800 198498 856
rect 198666 800 199050 856
rect 199218 800 199602 856
rect 199770 800 200062 856
rect 200230 800 200614 856
rect 200782 800 201166 856
rect 201334 800 201718 856
rect 201886 800 202178 856
rect 202346 800 202730 856
rect 202898 800 203282 856
rect 203450 800 203742 856
rect 203910 800 204294 856
rect 204462 800 204846 856
rect 205014 800 205398 856
rect 205566 800 205858 856
rect 206026 800 206410 856
rect 206578 800 206962 856
rect 207130 800 207422 856
rect 207590 800 207974 856
rect 208142 800 208526 856
rect 208694 800 209078 856
rect 209246 800 209538 856
rect 209706 800 210090 856
rect 210258 800 210642 856
rect 210810 800 211102 856
rect 211270 800 211654 856
rect 211822 800 212206 856
rect 212374 800 212758 856
rect 212926 800 213218 856
rect 213386 800 213770 856
rect 213938 800 214322 856
rect 214490 800 214874 856
rect 215042 800 215334 856
rect 215502 800 215886 856
rect 216054 800 216438 856
rect 216606 800 216898 856
rect 217066 800 217450 856
rect 217618 800 218002 856
rect 218170 800 218554 856
rect 218722 800 219014 856
rect 219182 800 219566 856
rect 219734 800 220118 856
rect 220286 800 220578 856
rect 220746 800 221130 856
rect 221298 800 221682 856
rect 221850 800 222234 856
rect 222402 800 222694 856
rect 222862 800 223246 856
rect 223414 800 223798 856
rect 223966 800 224258 856
rect 224426 800 224810 856
rect 224978 800 225362 856
rect 225530 800 225914 856
rect 226082 800 226374 856
rect 226542 800 226926 856
rect 227094 800 227478 856
rect 227646 800 228030 856
rect 228198 800 228490 856
rect 228658 800 229042 856
rect 229210 800 229594 856
rect 229762 800 230054 856
rect 230222 800 230606 856
rect 230774 800 231158 856
rect 231326 800 231710 856
rect 231878 800 232170 856
rect 232338 800 232722 856
rect 232890 800 233274 856
rect 233442 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234838 856
rect 235006 800 235390 856
rect 235558 800 235850 856
rect 236018 800 236402 856
rect 236570 800 236954 856
rect 237122 800 237506 856
rect 237674 800 237966 856
rect 238134 800 238518 856
rect 238686 800 239070 856
rect 239238 800 239530 856
rect 239698 800 240082 856
rect 240250 800 240634 856
rect 240802 800 241186 856
rect 241354 800 241646 856
rect 241814 800 242198 856
rect 242366 800 242750 856
rect 242918 800 243210 856
rect 243378 800 243762 856
rect 243930 800 244314 856
rect 244482 800 244866 856
rect 245034 800 245326 856
rect 245494 800 245878 856
rect 246046 800 246430 856
rect 246598 800 246890 856
rect 247058 800 247442 856
rect 247610 800 247994 856
rect 248162 800 248546 856
rect 248714 800 249006 856
rect 249174 800 249558 856
rect 249726 800 250110 856
rect 250278 800 250662 856
rect 250830 800 251122 856
rect 251290 800 251674 856
rect 251842 800 252226 856
rect 252394 800 252686 856
rect 252854 800 253238 856
rect 253406 800 253790 856
rect 253958 800 254342 856
rect 254510 800 254802 856
rect 254970 800 255354 856
rect 255522 800 255906 856
rect 256074 800 256366 856
rect 256534 800 256918 856
rect 257086 800 257470 856
rect 257638 800 258022 856
rect 258190 800 258482 856
rect 258650 800 259034 856
rect 259202 800 259586 856
<< metal3 >>
rect 0 158312 800 158432
rect 259200 158312 260000 158432
rect 0 155320 800 155440
rect 259200 155320 260000 155440
rect 0 152328 800 152448
rect 259200 152328 260000 152448
rect 0 149336 800 149456
rect 259200 149336 260000 149456
rect 0 146480 800 146600
rect 259200 146344 260000 146464
rect 0 143488 800 143608
rect 259200 143216 260000 143336
rect 0 140496 800 140616
rect 259200 140224 260000 140344
rect 0 137504 800 137624
rect 259200 137232 260000 137352
rect 0 134648 800 134768
rect 259200 134240 260000 134360
rect 0 131656 800 131776
rect 259200 131248 260000 131368
rect 0 128664 800 128784
rect 259200 128120 260000 128240
rect 0 125672 800 125792
rect 259200 125128 260000 125248
rect 0 122680 800 122800
rect 259200 122136 260000 122256
rect 0 119824 800 119944
rect 259200 119144 260000 119264
rect 0 116832 800 116952
rect 259200 116152 260000 116272
rect 0 113840 800 113960
rect 259200 113024 260000 113144
rect 0 110848 800 110968
rect 259200 110032 260000 110152
rect 0 107992 800 108112
rect 259200 107040 260000 107160
rect 0 105000 800 105120
rect 259200 104048 260000 104168
rect 0 102008 800 102128
rect 259200 101056 260000 101176
rect 0 99016 800 99136
rect 259200 98064 260000 98184
rect 0 96024 800 96144
rect 259200 94936 260000 95056
rect 0 93168 800 93288
rect 259200 91944 260000 92064
rect 0 90176 800 90296
rect 259200 88952 260000 89072
rect 0 87184 800 87304
rect 259200 85960 260000 86080
rect 0 84192 800 84312
rect 259200 82968 260000 83088
rect 0 81336 800 81456
rect 259200 79840 260000 79960
rect 0 78344 800 78464
rect 259200 76848 260000 76968
rect 0 75352 800 75472
rect 259200 73856 260000 73976
rect 0 72360 800 72480
rect 259200 70864 260000 70984
rect 0 69368 800 69488
rect 259200 67872 260000 67992
rect 0 66512 800 66632
rect 259200 64744 260000 64864
rect 0 63520 800 63640
rect 259200 61752 260000 61872
rect 0 60528 800 60648
rect 259200 58760 260000 58880
rect 0 57536 800 57656
rect 259200 55768 260000 55888
rect 0 54680 800 54800
rect 259200 52776 260000 52896
rect 0 51688 800 51808
rect 259200 49784 260000 49904
rect 0 48696 800 48816
rect 259200 46656 260000 46776
rect 0 45704 800 45824
rect 259200 43664 260000 43784
rect 0 42712 800 42832
rect 259200 40672 260000 40792
rect 0 39856 800 39976
rect 259200 37680 260000 37800
rect 0 36864 800 36984
rect 259200 34688 260000 34808
rect 0 33872 800 33992
rect 259200 31560 260000 31680
rect 0 30880 800 31000
rect 259200 28568 260000 28688
rect 0 28024 800 28144
rect 259200 25576 260000 25696
rect 0 25032 800 25152
rect 259200 22584 260000 22704
rect 0 22040 800 22160
rect 259200 19592 260000 19712
rect 0 19048 800 19168
rect 259200 16464 260000 16584
rect 0 16056 800 16176
rect 259200 13472 260000 13592
rect 0 13200 800 13320
rect 259200 10480 260000 10600
rect 0 10208 800 10328
rect 259200 7488 260000 7608
rect 0 7216 800 7336
rect 259200 4496 260000 4616
rect 0 4224 800 4344
rect 0 1368 800 1488
rect 259200 1504 260000 1624
<< obsm3 >>
rect 880 158232 259120 158405
rect 800 155520 259200 158232
rect 880 155240 259120 155520
rect 800 152528 259200 155240
rect 880 152248 259120 152528
rect 800 149536 259200 152248
rect 880 149256 259120 149536
rect 800 146680 259200 149256
rect 880 146544 259200 146680
rect 880 146400 259120 146544
rect 800 146264 259120 146400
rect 800 143688 259200 146264
rect 880 143416 259200 143688
rect 880 143408 259120 143416
rect 800 143136 259120 143408
rect 800 140696 259200 143136
rect 880 140424 259200 140696
rect 880 140416 259120 140424
rect 800 140144 259120 140416
rect 800 137704 259200 140144
rect 880 137432 259200 137704
rect 880 137424 259120 137432
rect 800 137152 259120 137424
rect 800 134848 259200 137152
rect 880 134568 259200 134848
rect 800 134440 259200 134568
rect 800 134160 259120 134440
rect 800 131856 259200 134160
rect 880 131576 259200 131856
rect 800 131448 259200 131576
rect 800 131168 259120 131448
rect 800 128864 259200 131168
rect 880 128584 259200 128864
rect 800 128320 259200 128584
rect 800 128040 259120 128320
rect 800 125872 259200 128040
rect 880 125592 259200 125872
rect 800 125328 259200 125592
rect 800 125048 259120 125328
rect 800 122880 259200 125048
rect 880 122600 259200 122880
rect 800 122336 259200 122600
rect 800 122056 259120 122336
rect 800 120024 259200 122056
rect 880 119744 259200 120024
rect 800 119344 259200 119744
rect 800 119064 259120 119344
rect 800 117032 259200 119064
rect 880 116752 259200 117032
rect 800 116352 259200 116752
rect 800 116072 259120 116352
rect 800 114040 259200 116072
rect 880 113760 259200 114040
rect 800 113224 259200 113760
rect 800 112944 259120 113224
rect 800 111048 259200 112944
rect 880 110768 259200 111048
rect 800 110232 259200 110768
rect 800 109952 259120 110232
rect 800 108192 259200 109952
rect 880 107912 259200 108192
rect 800 107240 259200 107912
rect 800 106960 259120 107240
rect 800 105200 259200 106960
rect 880 104920 259200 105200
rect 800 104248 259200 104920
rect 800 103968 259120 104248
rect 800 102208 259200 103968
rect 880 101928 259200 102208
rect 800 101256 259200 101928
rect 800 100976 259120 101256
rect 800 99216 259200 100976
rect 880 98936 259200 99216
rect 800 98264 259200 98936
rect 800 97984 259120 98264
rect 800 96224 259200 97984
rect 880 95944 259200 96224
rect 800 95136 259200 95944
rect 800 94856 259120 95136
rect 800 93368 259200 94856
rect 880 93088 259200 93368
rect 800 92144 259200 93088
rect 800 91864 259120 92144
rect 800 90376 259200 91864
rect 880 90096 259200 90376
rect 800 89152 259200 90096
rect 800 88872 259120 89152
rect 800 87384 259200 88872
rect 880 87104 259200 87384
rect 800 86160 259200 87104
rect 800 85880 259120 86160
rect 800 84392 259200 85880
rect 880 84112 259200 84392
rect 800 83168 259200 84112
rect 800 82888 259120 83168
rect 800 81536 259200 82888
rect 880 81256 259200 81536
rect 800 80040 259200 81256
rect 800 79760 259120 80040
rect 800 78544 259200 79760
rect 880 78264 259200 78544
rect 800 77048 259200 78264
rect 800 76768 259120 77048
rect 800 75552 259200 76768
rect 880 75272 259200 75552
rect 800 74056 259200 75272
rect 800 73776 259120 74056
rect 800 72560 259200 73776
rect 880 72280 259200 72560
rect 800 71064 259200 72280
rect 800 70784 259120 71064
rect 800 69568 259200 70784
rect 880 69288 259200 69568
rect 800 68072 259200 69288
rect 800 67792 259120 68072
rect 800 66712 259200 67792
rect 880 66432 259200 66712
rect 800 64944 259200 66432
rect 800 64664 259120 64944
rect 800 63720 259200 64664
rect 880 63440 259200 63720
rect 800 61952 259200 63440
rect 800 61672 259120 61952
rect 800 60728 259200 61672
rect 880 60448 259200 60728
rect 800 58960 259200 60448
rect 800 58680 259120 58960
rect 800 57736 259200 58680
rect 880 57456 259200 57736
rect 800 55968 259200 57456
rect 800 55688 259120 55968
rect 800 54880 259200 55688
rect 880 54600 259200 54880
rect 800 52976 259200 54600
rect 800 52696 259120 52976
rect 800 51888 259200 52696
rect 880 51608 259200 51888
rect 800 49984 259200 51608
rect 800 49704 259120 49984
rect 800 48896 259200 49704
rect 880 48616 259200 48896
rect 800 46856 259200 48616
rect 800 46576 259120 46856
rect 800 45904 259200 46576
rect 880 45624 259200 45904
rect 800 43864 259200 45624
rect 800 43584 259120 43864
rect 800 42912 259200 43584
rect 880 42632 259200 42912
rect 800 40872 259200 42632
rect 800 40592 259120 40872
rect 800 40056 259200 40592
rect 880 39776 259200 40056
rect 800 37880 259200 39776
rect 800 37600 259120 37880
rect 800 37064 259200 37600
rect 880 36784 259200 37064
rect 800 34888 259200 36784
rect 800 34608 259120 34888
rect 800 34072 259200 34608
rect 880 33792 259200 34072
rect 800 31760 259200 33792
rect 800 31480 259120 31760
rect 800 31080 259200 31480
rect 880 30800 259200 31080
rect 800 28768 259200 30800
rect 800 28488 259120 28768
rect 800 28224 259200 28488
rect 880 27944 259200 28224
rect 800 25776 259200 27944
rect 800 25496 259120 25776
rect 800 25232 259200 25496
rect 880 24952 259200 25232
rect 800 22784 259200 24952
rect 800 22504 259120 22784
rect 800 22240 259200 22504
rect 880 21960 259200 22240
rect 800 19792 259200 21960
rect 800 19512 259120 19792
rect 800 19248 259200 19512
rect 880 18968 259200 19248
rect 800 16664 259200 18968
rect 800 16384 259120 16664
rect 800 16256 259200 16384
rect 880 15976 259200 16256
rect 800 13672 259200 15976
rect 800 13400 259120 13672
rect 880 13392 259120 13400
rect 880 13120 259200 13392
rect 800 10680 259200 13120
rect 800 10408 259120 10680
rect 880 10400 259120 10408
rect 880 10128 259200 10400
rect 800 7688 259200 10128
rect 800 7416 259120 7688
rect 880 7408 259120 7416
rect 880 7136 259200 7408
rect 800 4696 259200 7136
rect 800 4424 259120 4696
rect 880 4416 259120 4424
rect 880 4144 259200 4416
rect 800 1704 259200 4144
rect 800 1568 259120 1704
rect 880 1424 259120 1568
rect 880 1395 259200 1424
<< metal4 >>
rect 4018 2128 4718 157808
rect 5058 2176 5758 157760
rect 8518 2128 9218 157808
rect 9558 2176 10258 157760
rect 13018 2128 13718 157808
rect 14058 2176 14758 157760
rect 17518 2128 18218 157808
rect 18558 16744 19258 157760
rect 22018 16696 22718 157808
rect 23058 16744 23758 157760
rect 26518 16696 27218 157808
rect 27558 16744 28258 157760
rect 31018 16696 31718 157808
rect 32058 16744 32758 157760
rect 35518 16696 36218 157808
rect 36558 16744 37258 157760
rect 40018 2128 40718 157808
rect 41058 2176 41758 157760
rect 44518 2128 45218 157808
rect 45558 2176 46258 157760
rect 49018 2128 49718 157808
rect 50058 2176 50758 157760
rect 53518 2128 54218 157808
rect 54558 2176 55258 157760
rect 58018 2128 58718 157808
rect 59058 2176 59758 157760
rect 62518 2128 63218 157808
rect 63558 2176 64258 157760
rect 67018 2128 67718 157808
rect 68058 2176 68758 157760
rect 71518 2128 72218 157808
rect 72558 2176 73258 157760
rect 76018 2128 76718 157808
rect 77058 2176 77758 157760
rect 80518 2128 81218 157808
rect 81558 2176 82258 157760
rect 85018 2128 85718 157808
rect 86058 2176 86758 157760
rect 89518 2128 90218 157808
rect 90558 2176 91258 157760
rect 94018 2128 94718 157808
rect 95058 2176 95758 157760
rect 98518 2128 99218 157808
rect 99558 2176 100258 157760
rect 103018 2128 103718 157808
rect 104058 2176 104758 157760
rect 107518 2128 108218 157808
rect 108558 2176 109258 157760
rect 112018 2128 112718 157808
rect 113058 2176 113758 157760
rect 116518 91064 117218 157808
rect 117558 91112 118258 157760
rect 121018 91064 121718 157808
rect 122058 91112 122758 157760
rect 125518 91064 126218 157808
rect 126558 91112 127258 157760
rect 130018 91064 130718 157808
rect 131058 91112 131758 157760
rect 134518 91064 135218 157808
rect 135558 91112 136258 157760
rect 139018 91064 139718 157808
rect 140058 91112 140758 157760
rect 143518 91064 144218 157808
rect 144558 91112 145258 157760
rect 148018 91064 148718 157808
rect 149058 91112 149758 157760
rect 152518 91064 153218 157808
rect 153558 91112 154258 157760
rect 157018 91064 157718 157808
rect 158058 91112 158758 157760
rect 161518 91064 162218 157808
rect 162558 91112 163258 157760
rect 166018 91064 166718 157808
rect 167058 91112 167758 157760
rect 170518 91064 171218 157808
rect 171558 91112 172258 157760
rect 175018 91064 175718 157808
rect 176058 91112 176758 157760
rect 179518 91064 180218 157808
rect 180558 91112 181258 157760
rect 184018 91064 184718 157808
rect 185058 91112 185758 157760
rect 188518 91064 189218 157808
rect 189558 91112 190258 157760
rect 193018 91064 193718 157808
rect 194058 91112 194758 157760
rect 197518 91064 198218 157808
rect 198558 91112 199258 157760
rect 202018 91064 202718 157808
rect 203058 91112 203758 157760
rect 206518 91064 207218 157808
rect 207558 91112 208258 157760
rect 211018 91064 211718 157808
rect 212058 91112 212758 157760
rect 215518 91064 216218 157808
rect 216558 91112 217258 157760
rect 220018 91064 220718 157808
rect 221058 91112 221758 157760
rect 116518 2128 117218 21048
rect 117558 2176 118258 21000
rect 121018 2128 121718 21048
rect 122058 2176 122758 21000
rect 125518 2128 126218 21048
rect 126558 2176 127258 21000
rect 130018 2128 130718 21048
rect 131058 2176 131758 21000
rect 134518 2128 135218 21048
rect 135558 2176 136258 21000
rect 139018 2128 139718 21048
rect 140058 2176 140758 21000
rect 143518 2128 144218 21048
rect 144558 2176 145258 21000
rect 148018 2128 148718 21048
rect 149058 2176 149758 21000
rect 152518 2128 153218 21048
rect 153558 2176 154258 21000
rect 157018 2128 157718 21048
rect 158058 2176 158758 21000
rect 161518 2128 162218 21048
rect 162558 2176 163258 21000
rect 166018 2128 166718 21048
rect 167058 2176 167758 21000
rect 170518 2128 171218 21048
rect 171558 2176 172258 21000
rect 175018 2128 175718 21048
rect 176058 2176 176758 21000
rect 179518 2128 180218 21048
rect 180558 2176 181258 21000
rect 184018 2128 184718 21048
rect 185058 2176 185758 21000
rect 188518 2128 189218 21048
rect 189558 2176 190258 21000
rect 193018 2128 193718 21048
rect 194058 2176 194758 21000
rect 197518 2128 198218 21048
rect 198558 2176 199258 21000
rect 202018 2128 202718 21048
rect 203058 2176 203758 21000
rect 206518 2128 207218 21048
rect 207558 2176 208258 21000
rect 211018 2128 211718 21048
rect 212058 2176 212758 21000
rect 215518 2128 216218 21048
rect 216558 2176 217258 21000
rect 220018 2128 220718 21048
rect 221058 2176 221758 21000
rect 224518 2128 225218 157808
rect 225558 2176 226258 157760
rect 229018 2128 229718 157808
rect 230058 2176 230758 157760
rect 233518 2128 234218 157808
rect 234558 2176 235258 157760
rect 238018 2128 238718 157808
rect 239058 2176 239758 157760
rect 242518 2128 243218 157808
rect 243558 2176 244258 157760
rect 247018 2128 247718 157808
rect 248058 2176 248758 157760
rect 251518 2128 252218 157808
rect 252558 2176 253258 157760
rect 256018 2128 256718 157808
rect 257058 2176 257758 157760
<< obsm4 >>
rect 22798 16664 22978 157453
rect 23838 16664 26438 157453
rect 22798 16616 26438 16664
rect 27298 16664 27478 157453
rect 28338 16664 30938 157453
rect 27298 16616 30938 16664
rect 31798 16664 31978 157453
rect 32838 16664 35438 157453
rect 31798 16616 35438 16664
rect 36298 16664 36478 157453
rect 37338 16664 39938 157453
rect 36298 16616 39938 16664
rect 22000 2619 39938 16616
rect 40798 2619 40978 157453
rect 41838 2619 44438 157453
rect 45298 2619 45478 157453
rect 46338 2619 48938 157453
rect 49798 2619 49978 157453
rect 50838 2619 53438 157453
rect 54298 2619 54478 157453
rect 55338 2619 57938 157453
rect 58798 2619 58978 157453
rect 59838 2619 62438 157453
rect 63298 2619 63478 157453
rect 64338 2619 66938 157453
rect 67798 2619 67978 157453
rect 68838 2619 71438 157453
rect 72298 2619 72478 157453
rect 73338 2619 75938 157453
rect 76798 2619 76978 157453
rect 77838 2619 80438 157453
rect 81298 2619 81478 157453
rect 82338 2619 84938 157453
rect 85798 2619 85978 157453
rect 86838 2619 89438 157453
rect 90298 2619 90478 157453
rect 91338 2619 93938 157453
rect 94798 2619 94978 157453
rect 95838 2619 98438 157453
rect 99298 2619 99478 157453
rect 100338 2619 102938 157453
rect 103798 2619 103978 157453
rect 104838 2619 107438 157453
rect 108298 2619 108478 157453
rect 109338 2619 111938 157453
rect 112798 2619 112978 157453
rect 113838 90984 116438 157453
rect 117298 91032 117478 157453
rect 118338 91032 120938 157453
rect 117298 90984 120938 91032
rect 121798 91032 121978 157453
rect 122838 91032 125438 157453
rect 121798 90984 125438 91032
rect 126298 91032 126478 157453
rect 127338 91032 129938 157453
rect 126298 90984 129938 91032
rect 130798 91032 130978 157453
rect 131838 91032 134438 157453
rect 130798 90984 134438 91032
rect 135298 91032 135478 157453
rect 136338 91032 138938 157453
rect 135298 90984 138938 91032
rect 139798 91032 139978 157453
rect 140838 91032 143438 157453
rect 139798 90984 143438 91032
rect 144298 91032 144478 157453
rect 145338 91032 147938 157453
rect 144298 90984 147938 91032
rect 148798 91032 148978 157453
rect 149838 91032 152438 157453
rect 148798 90984 152438 91032
rect 153298 91032 153478 157453
rect 154338 91032 156938 157453
rect 153298 90984 156938 91032
rect 157798 91032 157978 157453
rect 158838 91032 161438 157453
rect 157798 90984 161438 91032
rect 162298 91032 162478 157453
rect 163338 91032 165938 157453
rect 162298 90984 165938 91032
rect 166798 91032 166978 157453
rect 167838 91032 170438 157453
rect 166798 90984 170438 91032
rect 171298 91032 171478 157453
rect 172338 91032 174938 157453
rect 171298 90984 174938 91032
rect 175798 91032 175978 157453
rect 176838 91032 179438 157453
rect 175798 90984 179438 91032
rect 180298 91032 180478 157453
rect 181338 91032 183938 157453
rect 180298 90984 183938 91032
rect 184798 91032 184978 157453
rect 185838 91032 188438 157453
rect 184798 90984 188438 91032
rect 189298 91032 189478 157453
rect 190338 91032 192938 157453
rect 189298 90984 192938 91032
rect 193798 91032 193978 157453
rect 194838 91032 197438 157453
rect 193798 90984 197438 91032
rect 198298 91032 198478 157453
rect 199338 91032 201938 157453
rect 198298 90984 201938 91032
rect 202798 91032 202978 157453
rect 203838 91032 206438 157453
rect 202798 90984 206438 91032
rect 207298 91032 207478 157453
rect 208338 91032 210938 157453
rect 207298 90984 210938 91032
rect 211798 91032 211978 157453
rect 212838 91032 215438 157453
rect 211798 90984 215438 91032
rect 216298 91032 216478 157453
rect 217338 91032 219637 157453
rect 216298 90984 219637 91032
rect 113838 21128 219637 90984
rect 113838 2619 116438 21128
rect 117298 21080 120938 21128
rect 117298 2619 117478 21080
rect 118338 2619 120938 21080
rect 121798 21080 125438 21128
rect 121798 2619 121978 21080
rect 122838 2619 125438 21080
rect 126298 21080 129938 21128
rect 126298 2619 126478 21080
rect 127338 2619 129938 21080
rect 130798 21080 134438 21128
rect 130798 2619 130978 21080
rect 131838 2619 134438 21080
rect 135298 21080 138938 21128
rect 135298 2619 135478 21080
rect 136338 2619 138938 21080
rect 139798 21080 143438 21128
rect 139798 2619 139978 21080
rect 140838 2619 143438 21080
rect 144298 21080 147938 21128
rect 144298 2619 144478 21080
rect 145338 2619 147938 21080
rect 148798 21080 152438 21128
rect 148798 2619 148978 21080
rect 149838 2619 152438 21080
rect 153298 21080 156938 21128
rect 153298 2619 153478 21080
rect 154338 2619 156938 21080
rect 157798 21080 161438 21128
rect 157798 2619 157978 21080
rect 158838 2619 161438 21080
rect 162298 21080 165938 21128
rect 162298 2619 162478 21080
rect 163338 2619 165938 21080
rect 166798 21080 170438 21128
rect 166798 2619 166978 21080
rect 167838 2619 170438 21080
rect 171298 21080 174938 21128
rect 171298 2619 171478 21080
rect 172338 2619 174938 21080
rect 175798 21080 179438 21128
rect 175798 2619 175978 21080
rect 176838 2619 179438 21080
rect 180298 21080 183938 21128
rect 180298 2619 180478 21080
rect 181338 2619 183938 21080
rect 184798 21080 188438 21128
rect 184798 2619 184978 21080
rect 185838 2619 188438 21080
rect 189298 21080 192938 21128
rect 189298 2619 189478 21080
rect 190338 2619 192938 21080
rect 193798 21080 197438 21128
rect 193798 2619 193978 21080
rect 194838 2619 197438 21080
rect 198298 21080 201938 21128
rect 198298 2619 198478 21080
rect 199338 2619 201938 21080
rect 202798 21080 206438 21128
rect 202798 2619 202978 21080
rect 203838 2619 206438 21080
rect 207298 21080 210938 21128
rect 207298 2619 207478 21080
rect 208338 2619 210938 21080
rect 211798 21080 215438 21128
rect 211798 2619 211978 21080
rect 212838 2619 215438 21080
rect 216298 21080 219637 21128
rect 216298 2619 216478 21080
rect 217338 2619 219637 21080
<< metal5 >>
rect 1104 154696 258888 155396
rect 1104 153608 258888 154308
rect 1104 150196 258888 150896
rect 1104 149108 258888 149808
rect 1104 145696 258888 146396
rect 1104 144608 258888 145308
rect 1104 141196 258888 141896
rect 1104 140108 258888 140808
rect 1104 136696 258888 137396
rect 1104 135608 258888 136308
rect 1104 132196 258888 132896
rect 1104 131108 258888 131808
rect 1104 127696 258888 128396
rect 1104 126608 258888 127308
rect 1104 123196 258888 123896
rect 1104 122108 258888 122808
rect 1104 118696 258888 119396
rect 1104 117608 258888 118308
rect 1104 114196 258888 114896
rect 1104 113108 258888 113808
rect 1104 109696 258888 110396
rect 1104 108608 258888 109308
rect 1104 105196 258888 105896
rect 1104 104108 258888 104808
rect 1104 100696 258888 101396
rect 1104 99608 258888 100308
rect 1104 96196 258888 96896
rect 1104 95108 258888 95808
rect 1104 91696 258888 92396
rect 1104 90608 258888 91308
rect 1104 87196 258888 87896
rect 1104 86108 258888 86808
rect 1104 82696 258888 83396
rect 1104 81608 258888 82308
rect 1104 78196 258888 78896
rect 1104 77108 258888 77808
rect 1104 73696 258888 74396
rect 1104 72608 258888 73308
rect 1104 69196 258888 69896
rect 1104 68108 258888 68808
rect 1104 64696 258888 65396
rect 1104 63608 258888 64308
rect 1104 60196 258888 60896
rect 1104 59108 258888 59808
rect 1104 55696 258888 56396
rect 1104 54608 258888 55308
rect 1104 51196 258888 51896
rect 1104 50108 258888 50808
rect 1104 46696 258888 47396
rect 1104 45608 258888 46308
rect 1104 42196 258888 42896
rect 1104 41108 258888 41808
rect 1104 37696 258888 38396
rect 1104 36608 258888 37308
rect 1104 33196 258888 33896
rect 1104 32108 258888 32808
rect 1104 28696 258888 29396
rect 1104 27608 258888 28308
rect 1104 24196 258888 24896
rect 1104 23108 258888 23808
rect 1104 19696 258888 20396
rect 1104 18608 258888 19308
rect 1104 15196 258888 15896
rect 1104 14108 258888 14808
rect 1104 10696 258888 11396
rect 1104 9608 258888 10308
rect 1104 6196 258888 6896
rect 1104 5108 258888 5808
<< labels >>
rlabel metal3 s 259200 64744 260000 64864 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 198554 159200 198610 160000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 169666 159200 169722 160000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 140778 159200 140834 160000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 111890 159200 111946 160000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 83002 159200 83058 160000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 54114 159200 54170 160000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 25226 159200 25282 160000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 158312 800 158432 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 146480 800 146600 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 134648 800 134768 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 259200 76848 260000 76968 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 122680 800 122800 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 110848 800 110968 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 99016 800 99136 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 87184 800 87304 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 75352 800 75472 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 63520 800 63640 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 51688 800 51808 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 39856 800 39976 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 28024 800 28144 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 259200 88952 260000 89072 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 259200 101056 260000 101176 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 259200 113024 260000 113144 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 259200 125128 260000 125248 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 259200 137232 260000 137352 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 259200 149336 260000 149456 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 256330 159200 256386 160000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 227442 159200 227498 160000 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 259200 1504 260000 1624 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 259200 104048 260000 104168 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 259200 116152 260000 116272 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 259200 128120 260000 128240 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 259200 140224 260000 140344 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 259200 152328 260000 152448 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 249154 159200 249210 160000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 220266 159200 220322 160000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 191378 159200 191434 160000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 162490 159200 162546 160000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 133602 159200 133658 160000 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 259200 10480 260000 10600 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 104714 159200 104770 160000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 75826 159200 75882 160000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 46938 159200 46994 160000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 18050 159200 18106 160000 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 155320 800 155440 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 259200 19592 260000 19712 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 259200 28568 260000 28688 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 259200 37680 260000 37800 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 259200 46656 260000 46776 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 259200 55768 260000 55888 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 259200 67872 260000 67992 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 259200 79840 260000 79960 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 259200 91944 260000 92064 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 259200 7488 260000 7608 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 259200 110032 260000 110152 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 259200 122136 260000 122256 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 259200 134240 260000 134360 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 259200 146344 260000 146464 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 259200 158312 260000 158432 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 234710 159200 234766 160000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 205822 159200 205878 160000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 176934 159200 176990 160000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 148046 159200 148102 160000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 119158 159200 119214 160000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 259200 16464 260000 16584 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 90270 159200 90326 160000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 61382 159200 61438 160000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 32494 159200 32550 160000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 3606 159200 3662 160000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 149336 800 149456 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 137504 800 137624 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 113840 800 113960 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 90176 800 90296 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 259200 25576 260000 25696 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 66512 800 66632 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 259200 34688 260000 34808 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 259200 43664 260000 43784 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 259200 52776 260000 52896 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 259200 61752 260000 61872 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 259200 73856 260000 73976 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 259200 85960 260000 86080 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 259200 98064 260000 98184 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 259200 4496 260000 4616 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 259200 107040 260000 107160 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 259200 119144 260000 119264 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 259200 131248 260000 131368 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 259200 143216 260000 143336 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 259200 155320 260000 155440 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 241886 159200 241942 160000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 212998 159200 213054 160000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 184110 159200 184166 160000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 155222 159200 155278 160000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 126334 159200 126390 160000 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 259200 13472 260000 13592 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 97446 159200 97502 160000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 68558 159200 68614 160000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 39670 159200 39726 160000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 10782 159200 10838 160000 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 140496 800 140616 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 128664 800 128784 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 116832 800 116952 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 105000 800 105120 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 259200 22584 260000 22704 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 259200 31560 260000 31680 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 259200 40672 260000 40792 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 259200 49784 260000 49904 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 259200 58760 260000 58880 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 259200 70864 260000 70984 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 259200 82968 260000 83088 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 259200 94936 260000 95056 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 213826 0 213882 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 216954 0 217010 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 220174 0 220230 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 226430 0 226486 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 240690 0 240746 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 246946 0 247002 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 251730 0 251786 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 253294 0 253350 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 254858 0 254914 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 179142 0 179198 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 191746 0 191802 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 193310 0 193366 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 194874 0 194930 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 210698 0 210754 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 214378 0 214434 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 215942 0 215998 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 217506 0 217562 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 219070 0 219126 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 220634 0 220690 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 222290 0 222346 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 223854 0 223910 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 226982 0 227038 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 228546 0 228602 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 230110 0 230166 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 231766 0 231822 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 234894 0 234950 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 238022 0 238078 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 239586 0 239642 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 241242 0 241298 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 244370 0 244426 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 247498 0 247554 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 250718 0 250774 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 252282 0 252338 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 253846 0 253902 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 255410 0 255466 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 256974 0 257030 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 58070 0 58126 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 157522 0 157578 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 168562 0 168618 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 173346 0 173402 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 174910 0 174966 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 179602 0 179658 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 181166 0 181222 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 182822 0 182878 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 196990 0 197046 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 198554 0 198610 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 200118 0 200174 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 204902 0 204958 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 208030 0 208086 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 209594 0 209650 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 212814 0 212870 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 222750 0 222806 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 224314 0 224370 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 229098 0 229154 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 240138 0 240194 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 243266 0 243322 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 246486 0 246542 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 252742 0 252798 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 200670 0 200726 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 210146 0 210202 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 258078 0 258134 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 258538 0 258594 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 259090 0 259146 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 259642 0 259698 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 532 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 256018 2128 256718 157808 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 247018 2128 247718 157808 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 238018 2128 238718 157808 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 229018 2128 229718 157808 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 220018 91064 220718 157808 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 211018 91064 211718 157808 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 202018 91064 202718 157808 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 193018 91064 193718 157808 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 184018 91064 184718 157808 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 175018 91064 175718 157808 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 166018 91064 166718 157808 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 157018 91064 157718 157808 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 148018 91064 148718 157808 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 139018 91064 139718 157808 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 130018 91064 130718 157808 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 121018 91064 121718 157808 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 112018 2128 112718 157808 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 103018 2128 103718 157808 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 94018 2128 94718 157808 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 85018 2128 85718 157808 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 76018 2128 76718 157808 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 67018 2128 67718 157808 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 58018 2128 58718 157808 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 49018 2128 49718 157808 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 40018 2128 40718 157808 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 31018 16696 31718 157808 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 22018 16696 22718 157808 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 13018 2128 13718 157808 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 4018 2128 4718 157808 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 220018 2128 220718 21048 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 211018 2128 211718 21048 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 202018 2128 202718 21048 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 193018 2128 193718 21048 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 184018 2128 184718 21048 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 175018 2128 175718 21048 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 166018 2128 166718 21048 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 157018 2128 157718 21048 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s 148018 2128 148718 21048 6 vccd1
port 675 nsew power bidirectional
rlabel metal4 s 139018 2128 139718 21048 6 vccd1
port 676 nsew power bidirectional
rlabel metal4 s 130018 2128 130718 21048 6 vccd1
port 677 nsew power bidirectional
rlabel metal4 s 121018 2128 121718 21048 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s 1104 149108 258888 149808 6 vccd1
port 679 nsew power bidirectional
rlabel metal5 s 1104 140108 258888 140808 6 vccd1
port 680 nsew power bidirectional
rlabel metal5 s 1104 131108 258888 131808 6 vccd1
port 681 nsew power bidirectional
rlabel metal5 s 1104 122108 258888 122808 6 vccd1
port 682 nsew power bidirectional
rlabel metal5 s 1104 113108 258888 113808 6 vccd1
port 683 nsew power bidirectional
rlabel metal5 s 1104 104108 258888 104808 6 vccd1
port 684 nsew power bidirectional
rlabel metal5 s 1104 95108 258888 95808 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s 1104 86108 258888 86808 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s 1104 77108 258888 77808 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s 1104 68108 258888 68808 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s 1104 59108 258888 59808 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s 1104 50108 258888 50808 6 vccd1
port 690 nsew power bidirectional
rlabel metal5 s 1104 41108 258888 41808 6 vccd1
port 691 nsew power bidirectional
rlabel metal5 s 1104 32108 258888 32808 6 vccd1
port 692 nsew power bidirectional
rlabel metal5 s 1104 23108 258888 23808 6 vccd1
port 693 nsew power bidirectional
rlabel metal5 s 1104 14108 258888 14808 6 vccd1
port 694 nsew power bidirectional
rlabel metal5 s 1104 5108 258888 5808 6 vccd1
port 695 nsew power bidirectional
rlabel metal4 s 251518 2128 252218 157808 6 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s 242518 2128 243218 157808 6 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 233518 2128 234218 157808 6 vssd1
port 698 nsew ground bidirectional
rlabel metal4 s 224518 2128 225218 157808 6 vssd1
port 699 nsew ground bidirectional
rlabel metal4 s 215518 91064 216218 157808 6 vssd1
port 700 nsew ground bidirectional
rlabel metal4 s 206518 91064 207218 157808 6 vssd1
port 701 nsew ground bidirectional
rlabel metal4 s 197518 91064 198218 157808 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 188518 91064 189218 157808 6 vssd1
port 703 nsew ground bidirectional
rlabel metal4 s 179518 91064 180218 157808 6 vssd1
port 704 nsew ground bidirectional
rlabel metal4 s 170518 91064 171218 157808 6 vssd1
port 705 nsew ground bidirectional
rlabel metal4 s 161518 91064 162218 157808 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 152518 91064 153218 157808 6 vssd1
port 707 nsew ground bidirectional
rlabel metal4 s 143518 91064 144218 157808 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s 134518 91064 135218 157808 6 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s 125518 91064 126218 157808 6 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 116518 91064 117218 157808 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 107518 2128 108218 157808 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 98518 2128 99218 157808 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 89518 2128 90218 157808 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 80518 2128 81218 157808 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 71518 2128 72218 157808 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 62518 2128 63218 157808 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 53518 2128 54218 157808 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 44518 2128 45218 157808 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 35518 16696 36218 157808 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 26518 16696 27218 157808 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 17518 2128 18218 157808 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 8518 2128 9218 157808 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 215518 2128 216218 21048 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s 206518 2128 207218 21048 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 197518 2128 198218 21048 6 vssd1
port 726 nsew ground bidirectional
rlabel metal4 s 188518 2128 189218 21048 6 vssd1
port 727 nsew ground bidirectional
rlabel metal4 s 179518 2128 180218 21048 6 vssd1
port 728 nsew ground bidirectional
rlabel metal4 s 170518 2128 171218 21048 6 vssd1
port 729 nsew ground bidirectional
rlabel metal4 s 161518 2128 162218 21048 6 vssd1
port 730 nsew ground bidirectional
rlabel metal4 s 152518 2128 153218 21048 6 vssd1
port 731 nsew ground bidirectional
rlabel metal4 s 143518 2128 144218 21048 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s 134518 2128 135218 21048 6 vssd1
port 733 nsew ground bidirectional
rlabel metal4 s 125518 2128 126218 21048 6 vssd1
port 734 nsew ground bidirectional
rlabel metal4 s 116518 2128 117218 21048 6 vssd1
port 735 nsew ground bidirectional
rlabel metal5 s 1104 153608 258888 154308 6 vssd1
port 736 nsew ground bidirectional
rlabel metal5 s 1104 144608 258888 145308 6 vssd1
port 737 nsew ground bidirectional
rlabel metal5 s 1104 135608 258888 136308 6 vssd1
port 738 nsew ground bidirectional
rlabel metal5 s 1104 126608 258888 127308 6 vssd1
port 739 nsew ground bidirectional
rlabel metal5 s 1104 117608 258888 118308 6 vssd1
port 740 nsew ground bidirectional
rlabel metal5 s 1104 108608 258888 109308 6 vssd1
port 741 nsew ground bidirectional
rlabel metal5 s 1104 99608 258888 100308 6 vssd1
port 742 nsew ground bidirectional
rlabel metal5 s 1104 90608 258888 91308 6 vssd1
port 743 nsew ground bidirectional
rlabel metal5 s 1104 81608 258888 82308 6 vssd1
port 744 nsew ground bidirectional
rlabel metal5 s 1104 72608 258888 73308 6 vssd1
port 745 nsew ground bidirectional
rlabel metal5 s 1104 63608 258888 64308 6 vssd1
port 746 nsew ground bidirectional
rlabel metal5 s 1104 54608 258888 55308 6 vssd1
port 747 nsew ground bidirectional
rlabel metal5 s 1104 45608 258888 46308 6 vssd1
port 748 nsew ground bidirectional
rlabel metal5 s 1104 36608 258888 37308 6 vssd1
port 749 nsew ground bidirectional
rlabel metal5 s 1104 27608 258888 28308 6 vssd1
port 750 nsew ground bidirectional
rlabel metal5 s 1104 18608 258888 19308 6 vssd1
port 751 nsew ground bidirectional
rlabel metal5 s 1104 9608 258888 10308 6 vssd1
port 752 nsew ground bidirectional
rlabel metal4 s 257058 2176 257758 157760 6 vccd2
port 753 nsew power bidirectional
rlabel metal4 s 248058 2176 248758 157760 6 vccd2
port 754 nsew power bidirectional
rlabel metal4 s 239058 2176 239758 157760 6 vccd2
port 755 nsew power bidirectional
rlabel metal4 s 230058 2176 230758 157760 6 vccd2
port 756 nsew power bidirectional
rlabel metal4 s 221058 91112 221758 157760 6 vccd2
port 757 nsew power bidirectional
rlabel metal4 s 212058 91112 212758 157760 6 vccd2
port 758 nsew power bidirectional
rlabel metal4 s 203058 91112 203758 157760 6 vccd2
port 759 nsew power bidirectional
rlabel metal4 s 194058 91112 194758 157760 6 vccd2
port 760 nsew power bidirectional
rlabel metal4 s 185058 91112 185758 157760 6 vccd2
port 761 nsew power bidirectional
rlabel metal4 s 176058 91112 176758 157760 6 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 167058 91112 167758 157760 6 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 158058 91112 158758 157760 6 vccd2
port 764 nsew power bidirectional
rlabel metal4 s 149058 91112 149758 157760 6 vccd2
port 765 nsew power bidirectional
rlabel metal4 s 140058 91112 140758 157760 6 vccd2
port 766 nsew power bidirectional
rlabel metal4 s 131058 91112 131758 157760 6 vccd2
port 767 nsew power bidirectional
rlabel metal4 s 122058 91112 122758 157760 6 vccd2
port 768 nsew power bidirectional
rlabel metal4 s 113058 2176 113758 157760 6 vccd2
port 769 nsew power bidirectional
rlabel metal4 s 104058 2176 104758 157760 6 vccd2
port 770 nsew power bidirectional
rlabel metal4 s 95058 2176 95758 157760 6 vccd2
port 771 nsew power bidirectional
rlabel metal4 s 86058 2176 86758 157760 6 vccd2
port 772 nsew power bidirectional
rlabel metal4 s 77058 2176 77758 157760 6 vccd2
port 773 nsew power bidirectional
rlabel metal4 s 68058 2176 68758 157760 6 vccd2
port 774 nsew power bidirectional
rlabel metal4 s 59058 2176 59758 157760 6 vccd2
port 775 nsew power bidirectional
rlabel metal4 s 50058 2176 50758 157760 6 vccd2
port 776 nsew power bidirectional
rlabel metal4 s 41058 2176 41758 157760 6 vccd2
port 777 nsew power bidirectional
rlabel metal4 s 32058 16744 32758 157760 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 23058 16744 23758 157760 6 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 14058 2176 14758 157760 6 vccd2
port 780 nsew power bidirectional
rlabel metal4 s 5058 2176 5758 157760 6 vccd2
port 781 nsew power bidirectional
rlabel metal4 s 221058 2176 221758 21000 6 vccd2
port 782 nsew power bidirectional
rlabel metal4 s 212058 2176 212758 21000 6 vccd2
port 783 nsew power bidirectional
rlabel metal4 s 203058 2176 203758 21000 6 vccd2
port 784 nsew power bidirectional
rlabel metal4 s 194058 2176 194758 21000 6 vccd2
port 785 nsew power bidirectional
rlabel metal4 s 185058 2176 185758 21000 6 vccd2
port 786 nsew power bidirectional
rlabel metal4 s 176058 2176 176758 21000 6 vccd2
port 787 nsew power bidirectional
rlabel metal4 s 167058 2176 167758 21000 6 vccd2
port 788 nsew power bidirectional
rlabel metal4 s 158058 2176 158758 21000 6 vccd2
port 789 nsew power bidirectional
rlabel metal4 s 149058 2176 149758 21000 6 vccd2
port 790 nsew power bidirectional
rlabel metal4 s 140058 2176 140758 21000 6 vccd2
port 791 nsew power bidirectional
rlabel metal4 s 131058 2176 131758 21000 6 vccd2
port 792 nsew power bidirectional
rlabel metal4 s 122058 2176 122758 21000 6 vccd2
port 793 nsew power bidirectional
rlabel metal5 s 1104 150196 258888 150896 6 vccd2
port 794 nsew power bidirectional
rlabel metal5 s 1104 141196 258888 141896 6 vccd2
port 795 nsew power bidirectional
rlabel metal5 s 1104 132196 258888 132896 6 vccd2
port 796 nsew power bidirectional
rlabel metal5 s 1104 123196 258888 123896 6 vccd2
port 797 nsew power bidirectional
rlabel metal5 s 1104 114196 258888 114896 6 vccd2
port 798 nsew power bidirectional
rlabel metal5 s 1104 105196 258888 105896 6 vccd2
port 799 nsew power bidirectional
rlabel metal5 s 1104 96196 258888 96896 6 vccd2
port 800 nsew power bidirectional
rlabel metal5 s 1104 87196 258888 87896 6 vccd2
port 801 nsew power bidirectional
rlabel metal5 s 1104 78196 258888 78896 6 vccd2
port 802 nsew power bidirectional
rlabel metal5 s 1104 69196 258888 69896 6 vccd2
port 803 nsew power bidirectional
rlabel metal5 s 1104 60196 258888 60896 6 vccd2
port 804 nsew power bidirectional
rlabel metal5 s 1104 51196 258888 51896 6 vccd2
port 805 nsew power bidirectional
rlabel metal5 s 1104 42196 258888 42896 6 vccd2
port 806 nsew power bidirectional
rlabel metal5 s 1104 33196 258888 33896 6 vccd2
port 807 nsew power bidirectional
rlabel metal5 s 1104 24196 258888 24896 6 vccd2
port 808 nsew power bidirectional
rlabel metal5 s 1104 15196 258888 15896 6 vccd2
port 809 nsew power bidirectional
rlabel metal5 s 1104 6196 258888 6896 6 vccd2
port 810 nsew power bidirectional
rlabel metal4 s 252558 2176 253258 157760 6 vssd2
port 811 nsew ground bidirectional
rlabel metal4 s 243558 2176 244258 157760 6 vssd2
port 812 nsew ground bidirectional
rlabel metal4 s 234558 2176 235258 157760 6 vssd2
port 813 nsew ground bidirectional
rlabel metal4 s 225558 2176 226258 157760 6 vssd2
port 814 nsew ground bidirectional
rlabel metal4 s 216558 91112 217258 157760 6 vssd2
port 815 nsew ground bidirectional
rlabel metal4 s 207558 91112 208258 157760 6 vssd2
port 816 nsew ground bidirectional
rlabel metal4 s 198558 91112 199258 157760 6 vssd2
port 817 nsew ground bidirectional
rlabel metal4 s 189558 91112 190258 157760 6 vssd2
port 818 nsew ground bidirectional
rlabel metal4 s 180558 91112 181258 157760 6 vssd2
port 819 nsew ground bidirectional
rlabel metal4 s 171558 91112 172258 157760 6 vssd2
port 820 nsew ground bidirectional
rlabel metal4 s 162558 91112 163258 157760 6 vssd2
port 821 nsew ground bidirectional
rlabel metal4 s 153558 91112 154258 157760 6 vssd2
port 822 nsew ground bidirectional
rlabel metal4 s 144558 91112 145258 157760 6 vssd2
port 823 nsew ground bidirectional
rlabel metal4 s 135558 91112 136258 157760 6 vssd2
port 824 nsew ground bidirectional
rlabel metal4 s 126558 91112 127258 157760 6 vssd2
port 825 nsew ground bidirectional
rlabel metal4 s 117558 91112 118258 157760 6 vssd2
port 826 nsew ground bidirectional
rlabel metal4 s 108558 2176 109258 157760 6 vssd2
port 827 nsew ground bidirectional
rlabel metal4 s 99558 2176 100258 157760 6 vssd2
port 828 nsew ground bidirectional
rlabel metal4 s 90558 2176 91258 157760 6 vssd2
port 829 nsew ground bidirectional
rlabel metal4 s 81558 2176 82258 157760 6 vssd2
port 830 nsew ground bidirectional
rlabel metal4 s 72558 2176 73258 157760 6 vssd2
port 831 nsew ground bidirectional
rlabel metal4 s 63558 2176 64258 157760 6 vssd2
port 832 nsew ground bidirectional
rlabel metal4 s 54558 2176 55258 157760 6 vssd2
port 833 nsew ground bidirectional
rlabel metal4 s 45558 2176 46258 157760 6 vssd2
port 834 nsew ground bidirectional
rlabel metal4 s 36558 16744 37258 157760 6 vssd2
port 835 nsew ground bidirectional
rlabel metal4 s 27558 16744 28258 157760 6 vssd2
port 836 nsew ground bidirectional
rlabel metal4 s 18558 16744 19258 157760 6 vssd2
port 837 nsew ground bidirectional
rlabel metal4 s 9558 2176 10258 157760 6 vssd2
port 838 nsew ground bidirectional
rlabel metal4 s 216558 2176 217258 21000 6 vssd2
port 839 nsew ground bidirectional
rlabel metal4 s 207558 2176 208258 21000 6 vssd2
port 840 nsew ground bidirectional
rlabel metal4 s 198558 2176 199258 21000 6 vssd2
port 841 nsew ground bidirectional
rlabel metal4 s 189558 2176 190258 21000 6 vssd2
port 842 nsew ground bidirectional
rlabel metal4 s 180558 2176 181258 21000 6 vssd2
port 843 nsew ground bidirectional
rlabel metal4 s 171558 2176 172258 21000 6 vssd2
port 844 nsew ground bidirectional
rlabel metal4 s 162558 2176 163258 21000 6 vssd2
port 845 nsew ground bidirectional
rlabel metal4 s 153558 2176 154258 21000 6 vssd2
port 846 nsew ground bidirectional
rlabel metal4 s 144558 2176 145258 21000 6 vssd2
port 847 nsew ground bidirectional
rlabel metal4 s 135558 2176 136258 21000 6 vssd2
port 848 nsew ground bidirectional
rlabel metal4 s 126558 2176 127258 21000 6 vssd2
port 849 nsew ground bidirectional
rlabel metal4 s 117558 2176 118258 21000 6 vssd2
port 850 nsew ground bidirectional
rlabel metal5 s 1104 154696 258888 155396 6 vssd2
port 851 nsew ground bidirectional
rlabel metal5 s 1104 145696 258888 146396 6 vssd2
port 852 nsew ground bidirectional
rlabel metal5 s 1104 136696 258888 137396 6 vssd2
port 853 nsew ground bidirectional
rlabel metal5 s 1104 127696 258888 128396 6 vssd2
port 854 nsew ground bidirectional
rlabel metal5 s 1104 118696 258888 119396 6 vssd2
port 855 nsew ground bidirectional
rlabel metal5 s 1104 109696 258888 110396 6 vssd2
port 856 nsew ground bidirectional
rlabel metal5 s 1104 100696 258888 101396 6 vssd2
port 857 nsew ground bidirectional
rlabel metal5 s 1104 91696 258888 92396 6 vssd2
port 858 nsew ground bidirectional
rlabel metal5 s 1104 82696 258888 83396 6 vssd2
port 859 nsew ground bidirectional
rlabel metal5 s 1104 73696 258888 74396 6 vssd2
port 860 nsew ground bidirectional
rlabel metal5 s 1104 64696 258888 65396 6 vssd2
port 861 nsew ground bidirectional
rlabel metal5 s 1104 55696 258888 56396 6 vssd2
port 862 nsew ground bidirectional
rlabel metal5 s 1104 46696 258888 47396 6 vssd2
port 863 nsew ground bidirectional
rlabel metal5 s 1104 37696 258888 38396 6 vssd2
port 864 nsew ground bidirectional
rlabel metal5 s 1104 28696 258888 29396 6 vssd2
port 865 nsew ground bidirectional
rlabel metal5 s 1104 19696 258888 20396 6 vssd2
port 866 nsew ground bidirectional
rlabel metal5 s 1104 10696 258888 11396 6 vssd2
port 867 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 260000 160000
string LEFview TRUE
string GDS_FILE /project/openlane/adc_wrapper/runs/adc_wrapper/results/magic/adc_wrapper.gds
string GDS_END 19322832
string GDS_START 353128
<< end >>

