magic
tech sky130A
magscale 1 2
timestamp 1626095698
<< viali >>
rect 8335 10859 8369 10893
rect 3735 10723 3769 10757
rect 4379 10723 4413 10757
rect 8151 10723 8185 10757
rect 3919 10587 3953 10621
rect 7231 8751 7265 8785
rect 6035 8615 6069 8649
rect 7139 8615 7173 8649
rect 6127 8547 6161 8581
rect 6219 8547 6253 8581
rect 6495 8547 6529 8581
rect 6587 8547 6621 8581
rect 7047 8547 7081 8581
rect 6311 8479 6345 8513
rect 7323 8479 7357 8513
rect 6587 8207 6621 8241
rect 6863 8139 6897 8173
rect 6587 8071 6621 8105
rect 6679 8071 6713 8105
rect 6955 8071 6989 8105
rect 7047 8071 7081 8105
rect 6311 7663 6345 7697
rect 6587 7527 6621 7561
rect 6311 7459 6345 7493
rect 6403 7459 6437 7493
rect 6725 7119 6759 7153
rect 3735 6983 3769 7017
rect 4379 6983 4413 7017
rect 6622 6983 6656 7017
rect 7783 6983 7817 7017
rect 8427 6983 8461 7017
rect 8243 6847 8277 6881
rect 3919 6779 3953 6813
rect 5161 6575 5195 6609
rect 6035 6575 6069 6609
rect 6725 6575 6759 6609
rect 6127 6439 6161 6473
rect 5090 6371 5124 6405
rect 5667 6371 5701 6405
rect 5851 6371 5885 6405
rect 5943 6371 5977 6405
rect 6219 6371 6253 6405
rect 6796 6371 6830 6405
rect 4563 6235 4597 6269
rect 5575 5691 5609 5725
rect 6035 5487 6069 5521
rect 5115 5419 5149 5453
rect 6127 5351 6161 5385
rect 5667 5283 5701 5317
rect 5851 5283 5885 5317
rect 5943 5283 5977 5317
rect 6219 5283 6253 5317
rect 8151 3855 8185 3889
rect 7691 3719 7725 3753
rect 8335 3719 8369 3753
<< metal1 >>
rect 3430 11072 9134 11094
rect 3430 11020 4209 11072
rect 4261 11020 4273 11072
rect 4325 11020 4337 11072
rect 4389 11020 4401 11072
rect 4453 11020 4465 11072
rect 4517 11020 4529 11072
rect 4581 11020 6140 11072
rect 6192 11020 6204 11072
rect 6256 11020 6268 11072
rect 6320 11020 6332 11072
rect 6384 11020 6396 11072
rect 6448 11020 6460 11072
rect 6512 11020 8070 11072
rect 8122 11020 8134 11072
rect 8186 11020 8198 11072
rect 8250 11020 8262 11072
rect 8314 11020 8326 11072
rect 8378 11020 8390 11072
rect 8442 11020 9134 11072
rect 3430 10998 9134 11020
rect 8323 10893 8381 10899
rect 8323 10859 8335 10893
rect 8369 10890 8381 10893
rect 9332 10890 9338 10902
rect 8369 10862 9338 10890
rect 8369 10859 8381 10862
rect 8323 10853 8381 10859
rect 9332 10850 9338 10862
rect 9390 10850 9396 10902
rect 3352 10714 3358 10766
rect 3410 10754 3416 10766
rect 3723 10757 3781 10763
rect 3723 10754 3735 10757
rect 3410 10726 3735 10754
rect 3410 10714 3416 10726
rect 3723 10723 3735 10726
rect 3769 10754 3781 10757
rect 4367 10757 4425 10763
rect 4367 10754 4379 10757
rect 3769 10726 4379 10754
rect 3769 10723 3781 10726
rect 3723 10717 3781 10723
rect 4367 10723 4379 10726
rect 4413 10723 4425 10757
rect 4367 10717 4425 10723
rect 7584 10714 7590 10766
rect 7642 10754 7648 10766
rect 8139 10757 8197 10763
rect 8139 10754 8151 10757
rect 7642 10726 8151 10754
rect 7642 10714 7648 10726
rect 8139 10723 8151 10726
rect 8185 10723 8197 10757
rect 8139 10717 8197 10723
rect 3907 10621 3965 10627
rect 3907 10587 3919 10621
rect 3953 10618 3965 10621
rect 6572 10618 6578 10630
rect 3953 10590 6578 10618
rect 3953 10587 3965 10590
rect 3907 10581 3965 10587
rect 6572 10578 6578 10590
rect 6630 10578 6636 10630
rect 3430 10528 9134 10550
rect 3430 10476 5174 10528
rect 5226 10476 5238 10528
rect 5290 10476 5302 10528
rect 5354 10476 5366 10528
rect 5418 10476 5430 10528
rect 5482 10476 5494 10528
rect 5546 10476 7105 10528
rect 7157 10476 7169 10528
rect 7221 10476 7233 10528
rect 7285 10476 7297 10528
rect 7349 10476 7361 10528
rect 7413 10476 7425 10528
rect 7477 10476 9134 10528
rect 3430 10454 9134 10476
rect 3430 9984 9134 10006
rect 3430 9932 4209 9984
rect 4261 9932 4273 9984
rect 4325 9932 4337 9984
rect 4389 9932 4401 9984
rect 4453 9932 4465 9984
rect 4517 9932 4529 9984
rect 4581 9932 6140 9984
rect 6192 9932 6204 9984
rect 6256 9932 6268 9984
rect 6320 9932 6332 9984
rect 6384 9932 6396 9984
rect 6448 9932 6460 9984
rect 6512 9932 8070 9984
rect 8122 9932 8134 9984
rect 8186 9932 8198 9984
rect 8250 9932 8262 9984
rect 8314 9932 8326 9984
rect 8378 9932 8390 9984
rect 8442 9932 9134 9984
rect 3430 9910 9134 9932
rect 3430 9440 9134 9462
rect 3430 9388 5174 9440
rect 5226 9388 5238 9440
rect 5290 9388 5302 9440
rect 5354 9388 5366 9440
rect 5418 9388 5430 9440
rect 5482 9388 5494 9440
rect 5546 9388 7105 9440
rect 7157 9388 7169 9440
rect 7221 9388 7233 9440
rect 7285 9388 7297 9440
rect 7349 9388 7361 9440
rect 7413 9388 7425 9440
rect 7477 9388 9134 9440
rect 3430 9366 9134 9388
rect 3430 8896 9134 8918
rect 3430 8844 4209 8896
rect 4261 8844 4273 8896
rect 4325 8844 4337 8896
rect 4389 8844 4401 8896
rect 4453 8844 4465 8896
rect 4517 8844 4529 8896
rect 4581 8844 6140 8896
rect 6192 8844 6204 8896
rect 6256 8844 6268 8896
rect 6320 8844 6332 8896
rect 6384 8844 6396 8896
rect 6448 8844 6460 8896
rect 6512 8844 8070 8896
rect 8122 8844 8134 8896
rect 8186 8844 8198 8896
rect 8250 8844 8262 8896
rect 8314 8844 8326 8896
rect 8378 8844 8390 8896
rect 8442 8844 9134 8896
rect 3430 8822 9134 8844
rect 7219 8785 7277 8791
rect 7219 8751 7231 8785
rect 7265 8782 7277 8785
rect 7584 8782 7590 8794
rect 7265 8754 7590 8782
rect 7265 8751 7277 8754
rect 7219 8745 7277 8751
rect 7584 8742 7590 8754
rect 7642 8742 7648 8794
rect 6572 8714 6578 8726
rect 6498 8686 6578 8714
rect 6020 8646 6026 8658
rect 5981 8618 6026 8646
rect 6020 8606 6026 8618
rect 6078 8606 6084 8658
rect 5928 8538 5934 8590
rect 5986 8578 5992 8590
rect 6498 8587 6526 8686
rect 6572 8674 6578 8686
rect 6630 8674 6636 8726
rect 7127 8649 7185 8655
rect 7127 8646 7139 8649
rect 6590 8618 7139 8646
rect 6590 8590 6618 8618
rect 7127 8615 7139 8618
rect 7173 8615 7185 8649
rect 7127 8609 7185 8615
rect 6115 8581 6173 8587
rect 6115 8578 6127 8581
rect 5986 8550 6127 8578
rect 5986 8538 5992 8550
rect 6115 8547 6127 8550
rect 6161 8578 6173 8581
rect 6207 8581 6265 8587
rect 6207 8578 6219 8581
rect 6161 8550 6219 8578
rect 6161 8547 6173 8550
rect 6115 8541 6173 8547
rect 6207 8547 6219 8550
rect 6253 8547 6265 8581
rect 6207 8541 6265 8547
rect 6483 8581 6541 8587
rect 6483 8547 6495 8581
rect 6529 8547 6541 8581
rect 6483 8541 6541 8547
rect 6572 8538 6578 8590
rect 6630 8578 6636 8590
rect 6630 8550 6723 8578
rect 6630 8538 6636 8550
rect 6848 8538 6854 8590
rect 6906 8578 6912 8590
rect 7035 8581 7093 8587
rect 7035 8578 7047 8581
rect 6906 8550 7047 8578
rect 6906 8538 6912 8550
rect 7035 8547 7047 8550
rect 7081 8547 7093 8581
rect 7035 8541 7093 8547
rect 5836 8470 5842 8522
rect 5894 8510 5900 8522
rect 6299 8513 6357 8519
rect 6299 8510 6311 8513
rect 5894 8482 6311 8510
rect 5894 8470 5900 8482
rect 6299 8479 6311 8482
rect 6345 8479 6357 8513
rect 6299 8473 6357 8479
rect 6756 8470 6762 8522
rect 6814 8510 6820 8522
rect 7311 8513 7369 8519
rect 7311 8510 7323 8513
rect 6814 8482 7323 8510
rect 6814 8470 6820 8482
rect 7311 8479 7323 8482
rect 7357 8479 7369 8513
rect 7311 8473 7369 8479
rect 3430 8352 9134 8374
rect 3430 8300 5174 8352
rect 5226 8300 5238 8352
rect 5290 8300 5302 8352
rect 5354 8300 5366 8352
rect 5418 8300 5430 8352
rect 5482 8300 5494 8352
rect 5546 8300 7105 8352
rect 7157 8300 7169 8352
rect 7221 8300 7233 8352
rect 7285 8300 7297 8352
rect 7349 8300 7361 8352
rect 7413 8300 7425 8352
rect 7477 8300 9134 8352
rect 3430 8278 9134 8300
rect 6572 8238 6578 8250
rect 6533 8210 6578 8238
rect 6572 8198 6578 8210
rect 6630 8198 6636 8250
rect 5836 8130 5842 8182
rect 5894 8170 5900 8182
rect 6851 8173 6909 8179
rect 6851 8170 6863 8173
rect 5894 8142 6863 8170
rect 5894 8130 5900 8142
rect 6851 8139 6863 8142
rect 6897 8139 6909 8173
rect 6851 8133 6909 8139
rect 6020 8062 6026 8114
rect 6078 8102 6084 8114
rect 6575 8105 6633 8111
rect 6575 8102 6587 8105
rect 6078 8074 6587 8102
rect 6078 8062 6084 8074
rect 6575 8071 6587 8074
rect 6621 8071 6633 8105
rect 6575 8065 6633 8071
rect 6664 8062 6670 8114
rect 6722 8102 6728 8114
rect 6940 8102 6946 8114
rect 6722 8074 6767 8102
rect 6901 8074 6946 8102
rect 6722 8062 6728 8074
rect 6940 8062 6946 8074
rect 6998 8102 7004 8114
rect 7035 8105 7093 8111
rect 7035 8102 7047 8105
rect 6998 8074 7047 8102
rect 6998 8062 7004 8074
rect 7035 8071 7047 8074
rect 7081 8071 7093 8105
rect 7035 8065 7093 8071
rect 3430 7808 9134 7830
rect 3430 7756 4209 7808
rect 4261 7756 4273 7808
rect 4325 7756 4337 7808
rect 4389 7756 4401 7808
rect 4453 7756 4465 7808
rect 4517 7756 4529 7808
rect 4581 7756 6140 7808
rect 6192 7756 6204 7808
rect 6256 7756 6268 7808
rect 6320 7756 6332 7808
rect 6384 7756 6396 7808
rect 6448 7756 6460 7808
rect 6512 7756 8070 7808
rect 8122 7756 8134 7808
rect 8186 7756 8198 7808
rect 8250 7756 8262 7808
rect 8314 7756 8326 7808
rect 8378 7756 8390 7808
rect 8442 7756 9134 7808
rect 3430 7734 9134 7756
rect 6299 7697 6357 7703
rect 6299 7663 6311 7697
rect 6345 7694 6357 7697
rect 6848 7694 6854 7706
rect 6345 7666 6854 7694
rect 6345 7663 6357 7666
rect 6299 7657 6357 7663
rect 6848 7654 6854 7666
rect 6906 7654 6912 7706
rect 6575 7561 6633 7567
rect 6575 7527 6587 7561
rect 6621 7558 6633 7561
rect 7584 7558 7590 7570
rect 6621 7530 7590 7558
rect 6621 7527 6633 7530
rect 6575 7521 6633 7527
rect 7584 7518 7590 7530
rect 7642 7518 7648 7570
rect 6020 7450 6026 7502
rect 6078 7490 6084 7502
rect 6299 7493 6357 7499
rect 6299 7490 6311 7493
rect 6078 7462 6311 7490
rect 6078 7450 6084 7462
rect 6299 7459 6311 7462
rect 6345 7459 6357 7493
rect 6299 7453 6357 7459
rect 6391 7493 6449 7499
rect 6391 7459 6403 7493
rect 6437 7490 6449 7493
rect 6664 7490 6670 7502
rect 6437 7462 6670 7490
rect 6437 7459 6449 7462
rect 6391 7453 6449 7459
rect 6664 7450 6670 7462
rect 6722 7450 6728 7502
rect 3430 7264 9134 7286
rect 3430 7212 5174 7264
rect 5226 7212 5238 7264
rect 5290 7212 5302 7264
rect 5354 7212 5366 7264
rect 5418 7212 5430 7264
rect 5482 7212 5494 7264
rect 5546 7212 7105 7264
rect 7157 7212 7169 7264
rect 7221 7212 7233 7264
rect 7285 7212 7297 7264
rect 7349 7212 7361 7264
rect 7413 7212 7425 7264
rect 7477 7212 9134 7264
rect 3430 7190 9134 7212
rect 6756 7159 6762 7162
rect 6713 7153 6762 7159
rect 6713 7119 6725 7153
rect 6759 7119 6762 7153
rect 6713 7113 6762 7119
rect 6756 7110 6762 7113
rect 6814 7110 6820 7162
rect 3352 6974 3358 7026
rect 3410 7014 3416 7026
rect 3723 7017 3781 7023
rect 3723 7014 3735 7017
rect 3410 6986 3735 7014
rect 3410 6974 3416 6986
rect 3723 6983 3735 6986
rect 3769 7014 3781 7017
rect 4367 7017 4425 7023
rect 4367 7014 4379 7017
rect 3769 6986 4379 7014
rect 3769 6983 3781 6986
rect 3723 6977 3781 6983
rect 4367 6983 4379 6986
rect 4413 6983 4425 7017
rect 4367 6977 4425 6983
rect 6572 6974 6578 7026
rect 6630 7023 6636 7026
rect 6630 7017 6668 7023
rect 6656 6983 6668 7017
rect 6630 6977 6668 6983
rect 7771 7017 7829 7023
rect 7771 6983 7783 7017
rect 7817 7014 7829 7017
rect 8415 7017 8473 7023
rect 8415 7014 8427 7017
rect 7817 6986 8427 7014
rect 7817 6983 7829 6986
rect 7771 6977 7829 6983
rect 8415 6983 8427 6986
rect 8461 7014 8473 7017
rect 9332 7014 9338 7026
rect 8461 6986 9338 7014
rect 8461 6983 8473 6986
rect 8415 6977 8473 6983
rect 6630 6974 6636 6977
rect 9332 6974 9338 6986
rect 9390 6974 9396 7026
rect 6020 6838 6026 6890
rect 6078 6878 6084 6890
rect 8231 6881 8289 6887
rect 8231 6878 8243 6881
rect 6078 6850 8243 6878
rect 6078 6838 6084 6850
rect 8231 6847 8243 6850
rect 8277 6847 8289 6881
rect 8231 6841 8289 6847
rect 3907 6813 3965 6819
rect 3907 6779 3919 6813
rect 3953 6810 3965 6813
rect 5928 6810 5934 6822
rect 3953 6782 5934 6810
rect 3953 6779 3965 6782
rect 3907 6773 3965 6779
rect 5928 6770 5934 6782
rect 5986 6770 5992 6822
rect 3430 6720 9134 6742
rect 3430 6668 4209 6720
rect 4261 6668 4273 6720
rect 4325 6668 4337 6720
rect 4389 6668 4401 6720
rect 4453 6668 4465 6720
rect 4517 6668 4529 6720
rect 4581 6668 6140 6720
rect 6192 6668 6204 6720
rect 6256 6668 6268 6720
rect 6320 6668 6332 6720
rect 6384 6668 6396 6720
rect 6448 6668 6460 6720
rect 6512 6668 8070 6720
rect 8122 6668 8134 6720
rect 8186 6668 8198 6720
rect 8250 6668 8262 6720
rect 8314 6668 8326 6720
rect 8378 6668 8390 6720
rect 8442 6668 9134 6720
rect 3430 6646 9134 6668
rect 5149 6609 5207 6615
rect 5149 6575 5161 6609
rect 5195 6606 5207 6609
rect 5836 6606 5842 6618
rect 5195 6578 5842 6606
rect 5195 6575 5207 6578
rect 5149 6569 5207 6575
rect 5836 6566 5842 6578
rect 5894 6566 5900 6618
rect 6023 6609 6081 6615
rect 6023 6575 6035 6609
rect 6069 6606 6081 6609
rect 6572 6606 6578 6618
rect 6069 6578 6578 6606
rect 6069 6575 6081 6578
rect 6023 6569 6081 6575
rect 6572 6566 6578 6578
rect 6630 6566 6636 6618
rect 6664 6566 6670 6618
rect 6722 6615 6728 6618
rect 6722 6609 6771 6615
rect 6722 6575 6725 6609
rect 6759 6575 6771 6609
rect 6722 6569 6771 6575
rect 6722 6566 6728 6569
rect 6020 6430 6026 6482
rect 6078 6470 6084 6482
rect 6115 6473 6173 6479
rect 6115 6470 6127 6473
rect 6078 6442 6127 6470
rect 6078 6430 6084 6442
rect 6115 6439 6127 6442
rect 6161 6470 6173 6473
rect 6161 6442 6250 6470
rect 6161 6439 6173 6442
rect 6115 6433 6173 6439
rect 5078 6405 5136 6411
rect 5078 6371 5090 6405
rect 5124 6402 5136 6405
rect 5655 6405 5713 6411
rect 5124 6371 5146 6402
rect 5078 6365 5146 6371
rect 5655 6371 5667 6405
rect 5701 6402 5713 6405
rect 5744 6402 5750 6414
rect 5701 6374 5750 6402
rect 5701 6371 5713 6374
rect 5655 6365 5713 6371
rect 4551 6269 4609 6275
rect 4551 6235 4563 6269
rect 4597 6266 4609 6269
rect 5118 6266 5146 6365
rect 5744 6362 5750 6374
rect 5802 6362 5808 6414
rect 5839 6405 5897 6411
rect 5839 6371 5851 6405
rect 5885 6371 5897 6405
rect 5839 6365 5897 6371
rect 5854 6334 5882 6365
rect 5928 6362 5934 6414
rect 5986 6402 5992 6414
rect 6222 6411 6250 6442
rect 6207 6405 6265 6411
rect 5986 6374 6031 6402
rect 5986 6362 5992 6374
rect 6207 6371 6219 6405
rect 6253 6371 6265 6405
rect 6784 6405 6842 6411
rect 6784 6402 6796 6405
rect 6207 6365 6265 6371
rect 6314 6374 6796 6402
rect 5670 6306 5882 6334
rect 5670 6278 5698 6306
rect 5652 6266 5658 6278
rect 4597 6238 5658 6266
rect 4597 6235 4609 6238
rect 4551 6229 4609 6235
rect 5652 6226 5658 6238
rect 5710 6226 5716 6278
rect 5744 6226 5750 6278
rect 5802 6266 5808 6278
rect 6314 6266 6342 6374
rect 6784 6371 6796 6374
rect 6830 6371 6842 6405
rect 6784 6365 6842 6371
rect 5802 6238 6342 6266
rect 5802 6226 5808 6238
rect 3430 6176 9134 6198
rect 3430 6124 5174 6176
rect 5226 6124 5238 6176
rect 5290 6124 5302 6176
rect 5354 6124 5366 6176
rect 5418 6124 5430 6176
rect 5482 6124 5494 6176
rect 5546 6124 7105 6176
rect 7157 6124 7169 6176
rect 7221 6124 7233 6176
rect 7285 6124 7297 6176
rect 7349 6124 7361 6176
rect 7413 6124 7425 6176
rect 7477 6124 9134 6176
rect 3430 6102 9134 6124
rect 5563 5725 5621 5731
rect 5563 5691 5575 5725
rect 5609 5722 5621 5725
rect 5652 5722 5658 5734
rect 5609 5694 5658 5722
rect 5609 5691 5621 5694
rect 5563 5685 5621 5691
rect 5652 5682 5658 5694
rect 5710 5682 5716 5734
rect 3430 5632 9134 5654
rect 3430 5580 4209 5632
rect 4261 5580 4273 5632
rect 4325 5580 4337 5632
rect 4389 5580 4401 5632
rect 4453 5580 4465 5632
rect 4517 5580 4529 5632
rect 4581 5580 6140 5632
rect 6192 5580 6204 5632
rect 6256 5580 6268 5632
rect 6320 5580 6332 5632
rect 6384 5580 6396 5632
rect 6448 5580 6460 5632
rect 6512 5580 8070 5632
rect 8122 5580 8134 5632
rect 8186 5580 8198 5632
rect 8250 5580 8262 5632
rect 8314 5580 8326 5632
rect 8378 5580 8390 5632
rect 8442 5580 9134 5632
rect 3430 5558 9134 5580
rect 5744 5478 5750 5530
rect 5802 5518 5808 5530
rect 6023 5521 6081 5527
rect 6023 5518 6035 5521
rect 5802 5490 6035 5518
rect 5802 5478 5808 5490
rect 6023 5487 6035 5490
rect 6069 5487 6081 5521
rect 6023 5481 6081 5487
rect 3352 5410 3358 5462
rect 3410 5450 3416 5462
rect 5103 5453 5161 5459
rect 5103 5450 5115 5453
rect 3410 5422 5115 5450
rect 3410 5410 3416 5422
rect 5103 5419 5115 5422
rect 5149 5450 5161 5453
rect 5652 5450 5658 5462
rect 5149 5422 5658 5450
rect 5149 5419 5161 5422
rect 5103 5413 5161 5419
rect 5652 5410 5658 5422
rect 5710 5410 5716 5462
rect 5670 5382 5698 5410
rect 6115 5385 6173 5391
rect 5670 5354 5882 5382
rect 5854 5323 5882 5354
rect 6115 5351 6127 5385
rect 6161 5351 6173 5385
rect 6115 5345 6173 5351
rect 5655 5317 5713 5323
rect 5655 5283 5667 5317
rect 5701 5283 5713 5317
rect 5655 5277 5713 5283
rect 5839 5317 5897 5323
rect 5839 5283 5851 5317
rect 5885 5283 5897 5317
rect 5839 5277 5897 5283
rect 5670 5246 5698 5277
rect 5928 5274 5934 5326
rect 5986 5314 5992 5326
rect 6130 5314 6158 5345
rect 6207 5317 6265 5323
rect 6207 5314 6219 5317
rect 5986 5286 6031 5314
rect 6130 5286 6219 5314
rect 5986 5274 5992 5286
rect 6207 5283 6219 5286
rect 6253 5314 6265 5317
rect 6940 5314 6946 5326
rect 6253 5286 6946 5314
rect 6253 5283 6265 5286
rect 6207 5277 6265 5283
rect 6940 5274 6946 5286
rect 6998 5314 7004 5326
rect 7860 5314 7866 5326
rect 6998 5286 7866 5314
rect 6998 5274 7004 5286
rect 7860 5274 7866 5286
rect 7918 5274 7924 5326
rect 6572 5246 6578 5258
rect 5670 5218 6578 5246
rect 6572 5206 6578 5218
rect 6630 5206 6636 5258
rect 3430 5088 9134 5110
rect 3430 5036 5174 5088
rect 5226 5036 5238 5088
rect 5290 5036 5302 5088
rect 5354 5036 5366 5088
rect 5418 5036 5430 5088
rect 5482 5036 5494 5088
rect 5546 5036 7105 5088
rect 7157 5036 7169 5088
rect 7221 5036 7233 5088
rect 7285 5036 7297 5088
rect 7349 5036 7361 5088
rect 7413 5036 7425 5088
rect 7477 5036 9134 5088
rect 3430 5014 9134 5036
rect 3430 4544 9134 4566
rect 3430 4492 4209 4544
rect 4261 4492 4273 4544
rect 4325 4492 4337 4544
rect 4389 4492 4401 4544
rect 4453 4492 4465 4544
rect 4517 4492 4529 4544
rect 4581 4492 6140 4544
rect 6192 4492 6204 4544
rect 6256 4492 6268 4544
rect 6320 4492 6332 4544
rect 6384 4492 6396 4544
rect 6448 4492 6460 4544
rect 6512 4492 8070 4544
rect 8122 4492 8134 4544
rect 8186 4492 8198 4544
rect 8250 4492 8262 4544
rect 8314 4492 8326 4544
rect 8378 4492 8390 4544
rect 8442 4492 9134 4544
rect 3430 4470 9134 4492
rect 3430 4000 9134 4022
rect 3430 3948 5174 4000
rect 5226 3948 5238 4000
rect 5290 3948 5302 4000
rect 5354 3948 5366 4000
rect 5418 3948 5430 4000
rect 5482 3948 5494 4000
rect 5546 3948 7105 4000
rect 7157 3948 7169 4000
rect 7221 3948 7233 4000
rect 7285 3948 7297 4000
rect 7349 3948 7361 4000
rect 7413 3948 7425 4000
rect 7477 3948 9134 4000
rect 3430 3926 9134 3948
rect 7860 3846 7866 3898
rect 7918 3886 7924 3898
rect 8139 3889 8197 3895
rect 8139 3886 8151 3889
rect 7918 3858 8151 3886
rect 7918 3846 7924 3858
rect 8139 3855 8151 3858
rect 8185 3855 8197 3889
rect 8139 3849 8197 3855
rect 7679 3753 7737 3759
rect 7679 3719 7691 3753
rect 7725 3750 7737 3753
rect 8323 3753 8381 3759
rect 8323 3750 8335 3753
rect 7725 3722 8335 3750
rect 7725 3719 7737 3722
rect 7679 3713 7737 3719
rect 8323 3719 8335 3722
rect 8369 3750 8381 3753
rect 9332 3750 9338 3762
rect 8369 3722 9338 3750
rect 8369 3719 8381 3722
rect 8323 3713 8381 3719
rect 9332 3710 9338 3722
rect 9390 3710 9396 3762
rect 3430 3456 9134 3478
rect 3430 3404 4209 3456
rect 4261 3404 4273 3456
rect 4325 3404 4337 3456
rect 4389 3404 4401 3456
rect 4453 3404 4465 3456
rect 4517 3404 4529 3456
rect 4581 3404 6140 3456
rect 6192 3404 6204 3456
rect 6256 3404 6268 3456
rect 6320 3404 6332 3456
rect 6384 3404 6396 3456
rect 6448 3404 6460 3456
rect 6512 3404 8070 3456
rect 8122 3404 8134 3456
rect 8186 3404 8198 3456
rect 8250 3404 8262 3456
rect 8314 3404 8326 3456
rect 8378 3404 8390 3456
rect 8442 3404 9134 3456
rect 3430 3382 9134 3404
<< via1 >>
rect 4209 11020 4261 11072
rect 4273 11020 4325 11072
rect 4337 11020 4389 11072
rect 4401 11020 4453 11072
rect 4465 11020 4517 11072
rect 4529 11020 4581 11072
rect 6140 11020 6192 11072
rect 6204 11020 6256 11072
rect 6268 11020 6320 11072
rect 6332 11020 6384 11072
rect 6396 11020 6448 11072
rect 6460 11020 6512 11072
rect 8070 11020 8122 11072
rect 8134 11020 8186 11072
rect 8198 11020 8250 11072
rect 8262 11020 8314 11072
rect 8326 11020 8378 11072
rect 8390 11020 8442 11072
rect 9338 10850 9390 10902
rect 3358 10714 3410 10766
rect 7590 10714 7642 10766
rect 6578 10578 6630 10630
rect 5174 10476 5226 10528
rect 5238 10476 5290 10528
rect 5302 10476 5354 10528
rect 5366 10476 5418 10528
rect 5430 10476 5482 10528
rect 5494 10476 5546 10528
rect 7105 10476 7157 10528
rect 7169 10476 7221 10528
rect 7233 10476 7285 10528
rect 7297 10476 7349 10528
rect 7361 10476 7413 10528
rect 7425 10476 7477 10528
rect 4209 9932 4261 9984
rect 4273 9932 4325 9984
rect 4337 9932 4389 9984
rect 4401 9932 4453 9984
rect 4465 9932 4517 9984
rect 4529 9932 4581 9984
rect 6140 9932 6192 9984
rect 6204 9932 6256 9984
rect 6268 9932 6320 9984
rect 6332 9932 6384 9984
rect 6396 9932 6448 9984
rect 6460 9932 6512 9984
rect 8070 9932 8122 9984
rect 8134 9932 8186 9984
rect 8198 9932 8250 9984
rect 8262 9932 8314 9984
rect 8326 9932 8378 9984
rect 8390 9932 8442 9984
rect 5174 9388 5226 9440
rect 5238 9388 5290 9440
rect 5302 9388 5354 9440
rect 5366 9388 5418 9440
rect 5430 9388 5482 9440
rect 5494 9388 5546 9440
rect 7105 9388 7157 9440
rect 7169 9388 7221 9440
rect 7233 9388 7285 9440
rect 7297 9388 7349 9440
rect 7361 9388 7413 9440
rect 7425 9388 7477 9440
rect 4209 8844 4261 8896
rect 4273 8844 4325 8896
rect 4337 8844 4389 8896
rect 4401 8844 4453 8896
rect 4465 8844 4517 8896
rect 4529 8844 4581 8896
rect 6140 8844 6192 8896
rect 6204 8844 6256 8896
rect 6268 8844 6320 8896
rect 6332 8844 6384 8896
rect 6396 8844 6448 8896
rect 6460 8844 6512 8896
rect 8070 8844 8122 8896
rect 8134 8844 8186 8896
rect 8198 8844 8250 8896
rect 8262 8844 8314 8896
rect 8326 8844 8378 8896
rect 8390 8844 8442 8896
rect 7590 8742 7642 8794
rect 6026 8649 6078 8658
rect 6026 8615 6035 8649
rect 6035 8615 6069 8649
rect 6069 8615 6078 8649
rect 6026 8606 6078 8615
rect 5934 8538 5986 8590
rect 6578 8674 6630 8726
rect 6578 8581 6630 8590
rect 6578 8547 6587 8581
rect 6587 8547 6621 8581
rect 6621 8547 6630 8581
rect 6578 8538 6630 8547
rect 6854 8538 6906 8590
rect 5842 8470 5894 8522
rect 6762 8470 6814 8522
rect 5174 8300 5226 8352
rect 5238 8300 5290 8352
rect 5302 8300 5354 8352
rect 5366 8300 5418 8352
rect 5430 8300 5482 8352
rect 5494 8300 5546 8352
rect 7105 8300 7157 8352
rect 7169 8300 7221 8352
rect 7233 8300 7285 8352
rect 7297 8300 7349 8352
rect 7361 8300 7413 8352
rect 7425 8300 7477 8352
rect 6578 8241 6630 8250
rect 6578 8207 6587 8241
rect 6587 8207 6621 8241
rect 6621 8207 6630 8241
rect 6578 8198 6630 8207
rect 5842 8130 5894 8182
rect 6026 8062 6078 8114
rect 6670 8105 6722 8114
rect 6670 8071 6679 8105
rect 6679 8071 6713 8105
rect 6713 8071 6722 8105
rect 6946 8105 6998 8114
rect 6670 8062 6722 8071
rect 6946 8071 6955 8105
rect 6955 8071 6989 8105
rect 6989 8071 6998 8105
rect 6946 8062 6998 8071
rect 4209 7756 4261 7808
rect 4273 7756 4325 7808
rect 4337 7756 4389 7808
rect 4401 7756 4453 7808
rect 4465 7756 4517 7808
rect 4529 7756 4581 7808
rect 6140 7756 6192 7808
rect 6204 7756 6256 7808
rect 6268 7756 6320 7808
rect 6332 7756 6384 7808
rect 6396 7756 6448 7808
rect 6460 7756 6512 7808
rect 8070 7756 8122 7808
rect 8134 7756 8186 7808
rect 8198 7756 8250 7808
rect 8262 7756 8314 7808
rect 8326 7756 8378 7808
rect 8390 7756 8442 7808
rect 6854 7654 6906 7706
rect 7590 7518 7642 7570
rect 6026 7450 6078 7502
rect 6670 7450 6722 7502
rect 5174 7212 5226 7264
rect 5238 7212 5290 7264
rect 5302 7212 5354 7264
rect 5366 7212 5418 7264
rect 5430 7212 5482 7264
rect 5494 7212 5546 7264
rect 7105 7212 7157 7264
rect 7169 7212 7221 7264
rect 7233 7212 7285 7264
rect 7297 7212 7349 7264
rect 7361 7212 7413 7264
rect 7425 7212 7477 7264
rect 6762 7110 6814 7162
rect 3358 6974 3410 7026
rect 6578 7017 6630 7026
rect 6578 6983 6622 7017
rect 6622 6983 6630 7017
rect 6578 6974 6630 6983
rect 9338 6974 9390 7026
rect 6026 6838 6078 6890
rect 5934 6770 5986 6822
rect 4209 6668 4261 6720
rect 4273 6668 4325 6720
rect 4337 6668 4389 6720
rect 4401 6668 4453 6720
rect 4465 6668 4517 6720
rect 4529 6668 4581 6720
rect 6140 6668 6192 6720
rect 6204 6668 6256 6720
rect 6268 6668 6320 6720
rect 6332 6668 6384 6720
rect 6396 6668 6448 6720
rect 6460 6668 6512 6720
rect 8070 6668 8122 6720
rect 8134 6668 8186 6720
rect 8198 6668 8250 6720
rect 8262 6668 8314 6720
rect 8326 6668 8378 6720
rect 8390 6668 8442 6720
rect 5842 6566 5894 6618
rect 6578 6566 6630 6618
rect 6670 6566 6722 6618
rect 6026 6430 6078 6482
rect 5750 6362 5802 6414
rect 5934 6405 5986 6414
rect 5934 6371 5943 6405
rect 5943 6371 5977 6405
rect 5977 6371 5986 6405
rect 5934 6362 5986 6371
rect 5658 6226 5710 6278
rect 5750 6226 5802 6278
rect 5174 6124 5226 6176
rect 5238 6124 5290 6176
rect 5302 6124 5354 6176
rect 5366 6124 5418 6176
rect 5430 6124 5482 6176
rect 5494 6124 5546 6176
rect 7105 6124 7157 6176
rect 7169 6124 7221 6176
rect 7233 6124 7285 6176
rect 7297 6124 7349 6176
rect 7361 6124 7413 6176
rect 7425 6124 7477 6176
rect 5658 5682 5710 5734
rect 4209 5580 4261 5632
rect 4273 5580 4325 5632
rect 4337 5580 4389 5632
rect 4401 5580 4453 5632
rect 4465 5580 4517 5632
rect 4529 5580 4581 5632
rect 6140 5580 6192 5632
rect 6204 5580 6256 5632
rect 6268 5580 6320 5632
rect 6332 5580 6384 5632
rect 6396 5580 6448 5632
rect 6460 5580 6512 5632
rect 8070 5580 8122 5632
rect 8134 5580 8186 5632
rect 8198 5580 8250 5632
rect 8262 5580 8314 5632
rect 8326 5580 8378 5632
rect 8390 5580 8442 5632
rect 5750 5478 5802 5530
rect 3358 5410 3410 5462
rect 5658 5410 5710 5462
rect 5934 5317 5986 5326
rect 5934 5283 5943 5317
rect 5943 5283 5977 5317
rect 5977 5283 5986 5317
rect 5934 5274 5986 5283
rect 6946 5274 6998 5326
rect 7866 5274 7918 5326
rect 6578 5206 6630 5258
rect 5174 5036 5226 5088
rect 5238 5036 5290 5088
rect 5302 5036 5354 5088
rect 5366 5036 5418 5088
rect 5430 5036 5482 5088
rect 5494 5036 5546 5088
rect 7105 5036 7157 5088
rect 7169 5036 7221 5088
rect 7233 5036 7285 5088
rect 7297 5036 7349 5088
rect 7361 5036 7413 5088
rect 7425 5036 7477 5088
rect 4209 4492 4261 4544
rect 4273 4492 4325 4544
rect 4337 4492 4389 4544
rect 4401 4492 4453 4544
rect 4465 4492 4517 4544
rect 4529 4492 4581 4544
rect 6140 4492 6192 4544
rect 6204 4492 6256 4544
rect 6268 4492 6320 4544
rect 6332 4492 6384 4544
rect 6396 4492 6448 4544
rect 6460 4492 6512 4544
rect 8070 4492 8122 4544
rect 8134 4492 8186 4544
rect 8198 4492 8250 4544
rect 8262 4492 8314 4544
rect 8326 4492 8378 4544
rect 8390 4492 8442 4544
rect 5174 3948 5226 4000
rect 5238 3948 5290 4000
rect 5302 3948 5354 4000
rect 5366 3948 5418 4000
rect 5430 3948 5482 4000
rect 5494 3948 5546 4000
rect 7105 3948 7157 4000
rect 7169 3948 7221 4000
rect 7233 3948 7285 4000
rect 7297 3948 7349 4000
rect 7361 3948 7413 4000
rect 7425 3948 7477 4000
rect 7866 3846 7918 3898
rect 9338 3710 9390 3762
rect 4209 3404 4261 3456
rect 4273 3404 4325 3456
rect 4337 3404 4389 3456
rect 4401 3404 4453 3456
rect 4465 3404 4517 3456
rect 4529 3404 4581 3456
rect 6140 3404 6192 3456
rect 6204 3404 6256 3456
rect 6268 3404 6320 3456
rect 6332 3404 6384 3456
rect 6396 3404 6448 3456
rect 6460 3404 6512 3456
rect 8070 3404 8122 3456
rect 8134 3404 8186 3456
rect 8198 3404 8250 3456
rect 8262 3404 8314 3456
rect 8326 3404 8378 3456
rect 8390 3404 8442 3456
<< metal2 >>
rect 0 14434 460 14476
rect 0 14378 42 14434
rect 98 14378 122 14434
rect 178 14378 202 14434
rect 258 14378 282 14434
rect 338 14378 362 14434
rect 418 14378 460 14434
rect 0 14354 460 14378
rect 0 14298 42 14354
rect 98 14298 122 14354
rect 178 14298 202 14354
rect 258 14298 282 14354
rect 338 14298 362 14354
rect 418 14298 460 14354
rect 0 14274 460 14298
rect 0 14218 42 14274
rect 98 14218 122 14274
rect 178 14218 202 14274
rect 258 14218 282 14274
rect 338 14218 362 14274
rect 418 14218 460 14274
rect 0 14194 460 14218
rect 0 14138 42 14194
rect 98 14138 122 14194
rect 178 14138 202 14194
rect 258 14138 282 14194
rect 338 14138 362 14194
rect 418 14138 460 14194
rect 0 14114 460 14138
rect 0 14058 42 14114
rect 98 14058 122 14114
rect 178 14058 202 14114
rect 258 14058 282 14114
rect 338 14058 362 14114
rect 418 14058 460 14114
rect 0 8628 460 14058
rect 0 8572 42 8628
rect 98 8572 122 8628
rect 178 8572 202 8628
rect 258 8572 282 8628
rect 338 8572 362 8628
rect 418 8572 460 8628
rect 0 8548 460 8572
rect 0 8492 42 8548
rect 98 8492 122 8548
rect 178 8492 202 8548
rect 258 8492 282 8548
rect 338 8492 362 8548
rect 418 8492 460 8548
rect 0 8468 460 8492
rect 0 8412 42 8468
rect 98 8412 122 8468
rect 178 8412 202 8468
rect 258 8412 282 8468
rect 338 8412 362 8468
rect 418 8412 460 8468
rect 0 8388 460 8412
rect 0 8332 42 8388
rect 98 8332 122 8388
rect 178 8332 202 8388
rect 258 8332 282 8388
rect 338 8332 362 8388
rect 418 8332 460 8388
rect 0 6079 460 8332
rect 0 6023 42 6079
rect 98 6023 122 6079
rect 178 6023 202 6079
rect 258 6023 282 6079
rect 338 6023 362 6079
rect 418 6023 460 6079
rect 0 5999 460 6023
rect 0 5943 42 5999
rect 98 5943 122 5999
rect 178 5943 202 5999
rect 258 5943 282 5999
rect 338 5943 362 5999
rect 418 5943 460 5999
rect 0 5919 460 5943
rect 0 5863 42 5919
rect 98 5863 122 5919
rect 178 5863 202 5919
rect 258 5863 282 5919
rect 338 5863 362 5919
rect 418 5863 460 5919
rect 0 5839 460 5863
rect 0 5783 42 5839
rect 98 5783 122 5839
rect 178 5783 202 5839
rect 258 5783 282 5839
rect 338 5783 362 5839
rect 418 5783 460 5839
rect 0 418 460 5783
rect 800 13634 1260 13676
rect 800 13578 842 13634
rect 898 13578 922 13634
rect 978 13578 1002 13634
rect 1058 13578 1082 13634
rect 1138 13578 1162 13634
rect 1218 13578 1260 13634
rect 800 13554 1260 13578
rect 800 13498 842 13554
rect 898 13498 922 13554
rect 978 13498 1002 13554
rect 1058 13498 1082 13554
rect 1138 13498 1162 13554
rect 1218 13498 1260 13554
rect 800 13474 1260 13498
rect 800 13418 842 13474
rect 898 13418 922 13474
rect 978 13418 1002 13474
rect 1058 13418 1082 13474
rect 1138 13418 1162 13474
rect 1218 13418 1260 13474
rect 800 13394 1260 13418
rect 800 13338 842 13394
rect 898 13338 922 13394
rect 978 13338 1002 13394
rect 1058 13338 1082 13394
rect 1138 13338 1162 13394
rect 1218 13338 1260 13394
rect 800 13314 1260 13338
rect 800 13258 842 13314
rect 898 13258 922 13314
rect 978 13258 1002 13314
rect 1058 13258 1082 13314
rect 1138 13258 1162 13314
rect 1218 13258 1260 13314
rect 800 9903 1260 13258
rect 4185 13634 4605 14476
rect 4185 13578 4207 13634
rect 4263 13578 4287 13634
rect 4343 13578 4367 13634
rect 4423 13578 4447 13634
rect 4503 13578 4527 13634
rect 4583 13578 4605 13634
rect 4185 13554 4605 13578
rect 4185 13498 4207 13554
rect 4263 13498 4287 13554
rect 4343 13498 4367 13554
rect 4423 13498 4447 13554
rect 4503 13498 4527 13554
rect 4583 13498 4605 13554
rect 4185 13474 4605 13498
rect 4185 13418 4207 13474
rect 4263 13418 4287 13474
rect 4343 13418 4367 13474
rect 4423 13418 4447 13474
rect 4503 13418 4527 13474
rect 4583 13418 4605 13474
rect 4185 13394 4605 13418
rect 4185 13338 4207 13394
rect 4263 13338 4287 13394
rect 4343 13338 4367 13394
rect 4423 13338 4447 13394
rect 4503 13338 4527 13394
rect 4583 13338 4605 13394
rect 4185 13314 4605 13338
rect 4185 13258 4207 13314
rect 4263 13258 4287 13314
rect 4343 13258 4367 13314
rect 4423 13258 4447 13314
rect 4503 13258 4527 13314
rect 4583 13258 4605 13314
rect 2026 11158 3126 11256
rect 2026 11130 3398 11158
rect 2026 11032 3126 11130
rect 3370 10772 3398 11130
rect 4185 11072 4605 13258
rect 4185 11020 4209 11072
rect 4261 11020 4273 11072
rect 4325 11020 4337 11072
rect 4389 11020 4401 11072
rect 4453 11020 4465 11072
rect 4517 11020 4529 11072
rect 4581 11020 4605 11072
rect 3358 10766 3410 10772
rect 3358 10708 3410 10714
rect 800 9847 842 9903
rect 898 9847 922 9903
rect 978 9847 1002 9903
rect 1058 9847 1082 9903
rect 1138 9847 1162 9903
rect 1218 9847 1260 9903
rect 800 9823 1260 9847
rect 800 9767 842 9823
rect 898 9767 922 9823
rect 978 9767 1002 9823
rect 1058 9767 1082 9823
rect 1138 9767 1162 9823
rect 1218 9767 1260 9823
rect 800 9743 1260 9767
rect 800 9687 842 9743
rect 898 9687 922 9743
rect 978 9687 1002 9743
rect 1058 9687 1082 9743
rect 1138 9687 1162 9743
rect 1218 9687 1260 9743
rect 800 9663 1260 9687
rect 800 9607 842 9663
rect 898 9607 922 9663
rect 978 9607 1002 9663
rect 1058 9607 1082 9663
rect 1138 9607 1162 9663
rect 1218 9607 1260 9663
rect 800 7354 1260 9607
rect 800 7298 842 7354
rect 898 7298 922 7354
rect 978 7298 1002 7354
rect 1058 7298 1082 7354
rect 1138 7298 1162 7354
rect 1218 7298 1260 7354
rect 4185 9984 4605 11020
rect 4185 9932 4209 9984
rect 4261 9932 4273 9984
rect 4325 9932 4337 9984
rect 4389 9932 4401 9984
rect 4453 9932 4465 9984
rect 4517 9932 4529 9984
rect 4581 9932 4605 9984
rect 4185 9903 4605 9932
rect 4185 9847 4207 9903
rect 4263 9847 4287 9903
rect 4343 9847 4367 9903
rect 4423 9847 4447 9903
rect 4503 9847 4527 9903
rect 4583 9847 4605 9903
rect 4185 9823 4605 9847
rect 4185 9767 4207 9823
rect 4263 9767 4287 9823
rect 4343 9767 4367 9823
rect 4423 9767 4447 9823
rect 4503 9767 4527 9823
rect 4583 9767 4605 9823
rect 4185 9743 4605 9767
rect 4185 9687 4207 9743
rect 4263 9687 4287 9743
rect 4343 9687 4367 9743
rect 4423 9687 4447 9743
rect 4503 9687 4527 9743
rect 4583 9687 4605 9743
rect 4185 9663 4605 9687
rect 4185 9607 4207 9663
rect 4263 9607 4287 9663
rect 4343 9607 4367 9663
rect 4423 9607 4447 9663
rect 4503 9607 4527 9663
rect 4583 9607 4605 9663
rect 4185 8896 4605 9607
rect 4185 8844 4209 8896
rect 4261 8844 4273 8896
rect 4325 8844 4337 8896
rect 4389 8844 4401 8896
rect 4453 8844 4465 8896
rect 4517 8844 4529 8896
rect 4581 8844 4605 8896
rect 4185 7808 4605 8844
rect 4185 7756 4209 7808
rect 4261 7756 4273 7808
rect 4325 7756 4337 7808
rect 4389 7756 4401 7808
rect 4453 7756 4465 7808
rect 4517 7756 4529 7808
rect 4581 7756 4605 7808
rect 4185 7354 4605 7756
rect 800 7274 1260 7298
rect 800 7218 842 7274
rect 898 7218 922 7274
rect 978 7218 1002 7274
rect 1058 7218 1082 7274
rect 1138 7218 1162 7274
rect 1218 7218 1260 7274
rect 800 7194 1260 7218
rect 800 7138 842 7194
rect 898 7138 922 7194
rect 978 7138 1002 7194
rect 1058 7138 1082 7194
rect 1138 7138 1162 7194
rect 1218 7138 1260 7194
rect 800 7114 1260 7138
rect 800 7058 842 7114
rect 898 7058 922 7114
rect 978 7058 1002 7114
rect 1058 7058 1082 7114
rect 1138 7058 1162 7114
rect 1218 7058 1260 7114
rect 2026 7202 3126 7300
rect 4185 7298 4207 7354
rect 4263 7298 4287 7354
rect 4343 7298 4367 7354
rect 4423 7298 4447 7354
rect 4503 7298 4527 7354
rect 4583 7298 4605 7354
rect 4185 7274 4605 7298
rect 4185 7218 4207 7274
rect 4263 7218 4287 7274
rect 4343 7218 4367 7274
rect 4423 7218 4447 7274
rect 4503 7218 4527 7274
rect 4583 7218 4605 7274
rect 2026 7174 3398 7202
rect 2026 7076 3126 7174
rect 800 4804 1260 7058
rect 3370 7032 3398 7174
rect 4185 7194 4605 7218
rect 4185 7138 4207 7194
rect 4263 7138 4287 7194
rect 4343 7138 4367 7194
rect 4423 7138 4447 7194
rect 4503 7138 4527 7194
rect 4583 7138 4605 7194
rect 4185 7114 4605 7138
rect 4185 7058 4207 7114
rect 4263 7058 4287 7114
rect 4343 7058 4367 7114
rect 4423 7058 4447 7114
rect 4503 7058 4527 7114
rect 4583 7058 4605 7114
rect 3358 7026 3410 7032
rect 3358 6968 3410 6974
rect 4185 6720 4605 7058
rect 4185 6668 4209 6720
rect 4261 6668 4273 6720
rect 4325 6668 4337 6720
rect 4389 6668 4401 6720
rect 4453 6668 4465 6720
rect 4517 6668 4529 6720
rect 4581 6668 4605 6720
rect 4185 5632 4605 6668
rect 4185 5580 4209 5632
rect 4261 5580 4273 5632
rect 4325 5580 4337 5632
rect 4389 5580 4401 5632
rect 4453 5580 4465 5632
rect 4517 5580 4529 5632
rect 4581 5580 4605 5632
rect 3358 5462 3410 5468
rect 3358 5404 3410 5410
rect 800 4748 842 4804
rect 898 4748 922 4804
rect 978 4748 1002 4804
rect 1058 4748 1082 4804
rect 1138 4748 1162 4804
rect 1218 4748 1260 4804
rect 800 4724 1260 4748
rect 800 4668 842 4724
rect 898 4668 922 4724
rect 978 4668 1002 4724
rect 1058 4668 1082 4724
rect 1138 4668 1162 4724
rect 1218 4668 1260 4724
rect 800 4644 1260 4668
rect 800 4588 842 4644
rect 898 4588 922 4644
rect 978 4588 1002 4644
rect 1058 4588 1082 4644
rect 1138 4588 1162 4644
rect 1218 4588 1260 4644
rect 800 4564 1260 4588
rect 800 4508 842 4564
rect 898 4508 922 4564
rect 978 4508 1002 4564
rect 1058 4508 1082 4564
rect 1138 4508 1162 4564
rect 1218 4508 1260 4564
rect 800 1218 1260 4508
rect 2026 3246 3126 3344
rect 3370 3246 3398 5404
rect 2026 3218 3398 3246
rect 4185 4804 4605 5580
rect 4185 4748 4207 4804
rect 4263 4748 4287 4804
rect 4343 4748 4367 4804
rect 4423 4748 4447 4804
rect 4503 4748 4527 4804
rect 4583 4748 4605 4804
rect 4185 4724 4605 4748
rect 4185 4668 4207 4724
rect 4263 4668 4287 4724
rect 4343 4668 4367 4724
rect 4423 4668 4447 4724
rect 4503 4668 4527 4724
rect 4583 4668 4605 4724
rect 4185 4644 4605 4668
rect 4185 4588 4207 4644
rect 4263 4588 4287 4644
rect 4343 4588 4367 4644
rect 4423 4588 4447 4644
rect 4503 4588 4527 4644
rect 4583 4588 4605 4644
rect 4185 4564 4605 4588
rect 4185 4508 4207 4564
rect 4263 4544 4287 4564
rect 4343 4544 4367 4564
rect 4423 4544 4447 4564
rect 4503 4544 4527 4564
rect 4263 4508 4273 4544
rect 4517 4508 4527 4544
rect 4583 4508 4605 4564
rect 4185 4492 4209 4508
rect 4261 4492 4273 4508
rect 4325 4492 4337 4508
rect 4389 4492 4401 4508
rect 4453 4492 4465 4508
rect 4517 4492 4529 4508
rect 4581 4492 4605 4508
rect 4185 3456 4605 4492
rect 4185 3404 4209 3456
rect 4261 3404 4273 3456
rect 4325 3404 4337 3456
rect 4389 3404 4401 3456
rect 4453 3404 4465 3456
rect 4517 3404 4529 3456
rect 4581 3404 4605 3456
rect 2026 3120 3126 3218
rect 800 1162 842 1218
rect 898 1162 922 1218
rect 978 1162 1002 1218
rect 1058 1162 1082 1218
rect 1138 1162 1162 1218
rect 1218 1162 1260 1218
rect 800 1138 1260 1162
rect 800 1082 842 1138
rect 898 1082 922 1138
rect 978 1082 1002 1138
rect 1058 1082 1082 1138
rect 1138 1082 1162 1138
rect 1218 1082 1260 1138
rect 800 1058 1260 1082
rect 800 1002 842 1058
rect 898 1002 922 1058
rect 978 1002 1002 1058
rect 1058 1002 1082 1058
rect 1138 1002 1162 1058
rect 1218 1002 1260 1058
rect 800 978 1260 1002
rect 800 922 842 978
rect 898 922 922 978
rect 978 922 1002 978
rect 1058 922 1082 978
rect 1138 922 1162 978
rect 1218 922 1260 978
rect 800 898 1260 922
rect 800 842 842 898
rect 898 842 922 898
rect 978 842 1002 898
rect 1058 842 1082 898
rect 1138 842 1162 898
rect 1218 842 1260 898
rect 800 800 1260 842
rect 4185 1218 4605 3404
rect 4185 1162 4207 1218
rect 4263 1162 4287 1218
rect 4343 1162 4367 1218
rect 4423 1162 4447 1218
rect 4503 1162 4527 1218
rect 4583 1162 4605 1218
rect 4185 1138 4605 1162
rect 4185 1082 4207 1138
rect 4263 1082 4287 1138
rect 4343 1082 4367 1138
rect 4423 1082 4447 1138
rect 4503 1082 4527 1138
rect 4583 1082 4605 1138
rect 4185 1058 4605 1082
rect 4185 1002 4207 1058
rect 4263 1002 4287 1058
rect 4343 1002 4367 1058
rect 4423 1002 4447 1058
rect 4503 1002 4527 1058
rect 4583 1002 4605 1058
rect 4185 978 4605 1002
rect 4185 922 4207 978
rect 4263 922 4287 978
rect 4343 922 4367 978
rect 4423 922 4447 978
rect 4503 922 4527 978
rect 4583 922 4605 978
rect 4185 898 4605 922
rect 4185 842 4207 898
rect 4263 842 4287 898
rect 4343 842 4367 898
rect 4423 842 4447 898
rect 4503 842 4527 898
rect 4583 842 4605 898
rect 0 362 42 418
rect 98 362 122 418
rect 178 362 202 418
rect 258 362 282 418
rect 338 362 362 418
rect 418 362 460 418
rect 0 338 460 362
rect 0 282 42 338
rect 98 282 122 338
rect 178 282 202 338
rect 258 282 282 338
rect 338 282 362 338
rect 418 282 460 338
rect 0 258 460 282
rect 0 202 42 258
rect 98 202 122 258
rect 178 202 202 258
rect 258 202 282 258
rect 338 202 362 258
rect 418 202 460 258
rect 0 178 460 202
rect 0 122 42 178
rect 98 122 122 178
rect 178 122 202 178
rect 258 122 282 178
rect 338 122 362 178
rect 418 122 460 178
rect 0 98 460 122
rect 0 42 42 98
rect 98 42 122 98
rect 178 42 202 98
rect 258 42 282 98
rect 338 42 362 98
rect 418 42 460 98
rect 0 0 460 42
rect 4185 0 4605 842
rect 5150 14434 5571 14476
rect 5150 14378 5172 14434
rect 5228 14378 5252 14434
rect 5308 14378 5332 14434
rect 5388 14378 5412 14434
rect 5468 14378 5492 14434
rect 5548 14378 5571 14434
rect 5150 14354 5571 14378
rect 5150 14298 5172 14354
rect 5228 14298 5252 14354
rect 5308 14298 5332 14354
rect 5388 14298 5412 14354
rect 5468 14298 5492 14354
rect 5548 14298 5571 14354
rect 5150 14274 5571 14298
rect 5150 14218 5172 14274
rect 5228 14218 5252 14274
rect 5308 14218 5332 14274
rect 5388 14218 5412 14274
rect 5468 14218 5492 14274
rect 5548 14218 5571 14274
rect 5150 14194 5571 14218
rect 5150 14138 5172 14194
rect 5228 14138 5252 14194
rect 5308 14138 5332 14194
rect 5388 14138 5412 14194
rect 5468 14138 5492 14194
rect 5548 14138 5571 14194
rect 5150 14114 5571 14138
rect 5150 14058 5172 14114
rect 5228 14058 5252 14114
rect 5308 14058 5332 14114
rect 5388 14058 5412 14114
rect 5468 14058 5492 14114
rect 5548 14058 5571 14114
rect 5150 10528 5571 14058
rect 5150 10476 5174 10528
rect 5226 10476 5238 10528
rect 5290 10476 5302 10528
rect 5354 10476 5366 10528
rect 5418 10476 5430 10528
rect 5482 10476 5494 10528
rect 5546 10476 5571 10528
rect 5150 9440 5571 10476
rect 5150 9388 5174 9440
rect 5226 9388 5238 9440
rect 5290 9388 5302 9440
rect 5354 9388 5366 9440
rect 5418 9388 5430 9440
rect 5482 9388 5494 9440
rect 5546 9388 5571 9440
rect 5150 8628 5571 9388
rect 6116 13634 6536 14476
rect 6116 13578 6138 13634
rect 6194 13578 6218 13634
rect 6274 13578 6298 13634
rect 6354 13578 6378 13634
rect 6434 13578 6458 13634
rect 6514 13578 6536 13634
rect 6116 13554 6536 13578
rect 6116 13498 6138 13554
rect 6194 13498 6218 13554
rect 6274 13498 6298 13554
rect 6354 13498 6378 13554
rect 6434 13498 6458 13554
rect 6514 13498 6536 13554
rect 6116 13474 6536 13498
rect 6116 13418 6138 13474
rect 6194 13418 6218 13474
rect 6274 13418 6298 13474
rect 6354 13418 6378 13474
rect 6434 13418 6458 13474
rect 6514 13418 6536 13474
rect 6116 13394 6536 13418
rect 6116 13338 6138 13394
rect 6194 13338 6218 13394
rect 6274 13338 6298 13394
rect 6354 13338 6378 13394
rect 6434 13338 6458 13394
rect 6514 13338 6536 13394
rect 6116 13314 6536 13338
rect 6116 13258 6138 13314
rect 6194 13258 6218 13314
rect 6274 13258 6298 13314
rect 6354 13258 6378 13314
rect 6434 13258 6458 13314
rect 6514 13258 6536 13314
rect 6116 11072 6536 13258
rect 6116 11020 6140 11072
rect 6192 11020 6204 11072
rect 6256 11020 6268 11072
rect 6320 11020 6332 11072
rect 6384 11020 6396 11072
rect 6448 11020 6460 11072
rect 6512 11020 6536 11072
rect 6116 9984 6536 11020
rect 7081 14434 7501 14476
rect 7081 14378 7103 14434
rect 7159 14378 7183 14434
rect 7239 14378 7263 14434
rect 7319 14378 7343 14434
rect 7399 14378 7423 14434
rect 7479 14378 7501 14434
rect 7081 14354 7501 14378
rect 7081 14298 7103 14354
rect 7159 14298 7183 14354
rect 7239 14298 7263 14354
rect 7319 14298 7343 14354
rect 7399 14298 7423 14354
rect 7479 14298 7501 14354
rect 7081 14274 7501 14298
rect 7081 14218 7103 14274
rect 7159 14218 7183 14274
rect 7239 14218 7263 14274
rect 7319 14218 7343 14274
rect 7399 14218 7423 14274
rect 7479 14218 7501 14274
rect 7081 14194 7501 14218
rect 7081 14138 7103 14194
rect 7159 14138 7183 14194
rect 7239 14138 7263 14194
rect 7319 14138 7343 14194
rect 7399 14138 7423 14194
rect 7479 14138 7501 14194
rect 7081 14114 7501 14138
rect 7081 14058 7103 14114
rect 7159 14058 7183 14114
rect 7239 14058 7263 14114
rect 7319 14058 7343 14114
rect 7399 14058 7423 14114
rect 7479 14058 7501 14114
rect 6578 10630 6630 10636
rect 6578 10572 6630 10578
rect 6116 9932 6140 9984
rect 6192 9932 6204 9984
rect 6256 9932 6268 9984
rect 6320 9932 6332 9984
rect 6384 9932 6396 9984
rect 6448 9932 6460 9984
rect 6512 9932 6536 9984
rect 6116 9903 6536 9932
rect 6116 9847 6138 9903
rect 6194 9847 6218 9903
rect 6274 9847 6298 9903
rect 6354 9847 6378 9903
rect 6434 9847 6458 9903
rect 6514 9847 6536 9903
rect 6116 9823 6536 9847
rect 6116 9767 6138 9823
rect 6194 9767 6218 9823
rect 6274 9767 6298 9823
rect 6354 9767 6378 9823
rect 6434 9767 6458 9823
rect 6514 9767 6536 9823
rect 6116 9743 6536 9767
rect 6116 9687 6138 9743
rect 6194 9687 6218 9743
rect 6274 9687 6298 9743
rect 6354 9687 6378 9743
rect 6434 9687 6458 9743
rect 6514 9687 6536 9743
rect 6116 9663 6536 9687
rect 6116 9607 6138 9663
rect 6194 9607 6218 9663
rect 6274 9607 6298 9663
rect 6354 9607 6378 9663
rect 6434 9607 6458 9663
rect 6514 9607 6536 9663
rect 6116 8896 6536 9607
rect 6116 8844 6140 8896
rect 6192 8844 6204 8896
rect 6256 8844 6268 8896
rect 6320 8844 6332 8896
rect 6384 8844 6396 8896
rect 6448 8844 6460 8896
rect 6512 8844 6536 8896
rect 5150 8572 5172 8628
rect 5228 8572 5252 8628
rect 5308 8572 5332 8628
rect 5388 8572 5412 8628
rect 5468 8572 5492 8628
rect 5548 8572 5571 8628
rect 6026 8658 6078 8664
rect 6026 8600 6078 8606
rect 5150 8548 5571 8572
rect 5150 8492 5172 8548
rect 5228 8492 5252 8548
rect 5308 8492 5332 8548
rect 5388 8492 5412 8548
rect 5468 8492 5492 8548
rect 5548 8492 5571 8548
rect 5934 8590 5986 8596
rect 5934 8532 5986 8538
rect 5150 8468 5571 8492
rect 5150 8412 5172 8468
rect 5228 8412 5252 8468
rect 5308 8412 5332 8468
rect 5388 8412 5412 8468
rect 5468 8412 5492 8468
rect 5548 8412 5571 8468
rect 5842 8522 5894 8528
rect 5842 8464 5894 8470
rect 5150 8388 5571 8412
rect 5150 8332 5172 8388
rect 5228 8352 5252 8388
rect 5308 8352 5332 8388
rect 5388 8352 5412 8388
rect 5468 8352 5492 8388
rect 5228 8332 5238 8352
rect 5482 8332 5492 8352
rect 5548 8332 5571 8388
rect 5150 8300 5174 8332
rect 5226 8300 5238 8332
rect 5290 8300 5302 8332
rect 5354 8300 5366 8332
rect 5418 8300 5430 8332
rect 5482 8300 5494 8332
rect 5546 8300 5571 8332
rect 5150 7264 5571 8300
rect 5854 8188 5882 8464
rect 5842 8182 5894 8188
rect 5842 8124 5894 8130
rect 5150 7212 5174 7264
rect 5226 7212 5238 7264
rect 5290 7212 5302 7264
rect 5354 7212 5366 7264
rect 5418 7212 5430 7264
rect 5482 7212 5494 7264
rect 5546 7212 5571 7264
rect 5150 6176 5571 7212
rect 5854 6624 5882 8124
rect 5946 6912 5974 8532
rect 6038 8120 6066 8600
rect 6026 8114 6078 8120
rect 6026 8056 6078 8062
rect 6038 7508 6066 8056
rect 6116 7808 6536 8844
rect 6590 8732 6618 10572
rect 7081 10528 7501 14058
rect 8046 13634 8467 14476
rect 12104 14434 12564 14476
rect 12104 14378 12146 14434
rect 12202 14378 12226 14434
rect 12282 14378 12306 14434
rect 12362 14378 12386 14434
rect 12442 14378 12466 14434
rect 12522 14378 12564 14434
rect 12104 14354 12564 14378
rect 12104 14298 12146 14354
rect 12202 14298 12226 14354
rect 12282 14298 12306 14354
rect 12362 14298 12386 14354
rect 12442 14298 12466 14354
rect 12522 14298 12564 14354
rect 12104 14274 12564 14298
rect 12104 14218 12146 14274
rect 12202 14218 12226 14274
rect 12282 14218 12306 14274
rect 12362 14218 12386 14274
rect 12442 14218 12466 14274
rect 12522 14218 12564 14274
rect 12104 14194 12564 14218
rect 12104 14138 12146 14194
rect 12202 14138 12226 14194
rect 12282 14138 12306 14194
rect 12362 14138 12386 14194
rect 12442 14138 12466 14194
rect 12522 14138 12564 14194
rect 12104 14114 12564 14138
rect 12104 14058 12146 14114
rect 12202 14058 12226 14114
rect 12282 14058 12306 14114
rect 12362 14058 12386 14114
rect 12442 14058 12466 14114
rect 12522 14058 12564 14114
rect 8046 13578 8068 13634
rect 8124 13578 8148 13634
rect 8204 13578 8228 13634
rect 8284 13578 8308 13634
rect 8364 13578 8388 13634
rect 8444 13578 8467 13634
rect 8046 13554 8467 13578
rect 8046 13498 8068 13554
rect 8124 13498 8148 13554
rect 8204 13498 8228 13554
rect 8284 13498 8308 13554
rect 8364 13498 8388 13554
rect 8444 13498 8467 13554
rect 8046 13474 8467 13498
rect 8046 13418 8068 13474
rect 8124 13418 8148 13474
rect 8204 13418 8228 13474
rect 8284 13418 8308 13474
rect 8364 13418 8388 13474
rect 8444 13418 8467 13474
rect 8046 13394 8467 13418
rect 8046 13338 8068 13394
rect 8124 13338 8148 13394
rect 8204 13338 8228 13394
rect 8284 13338 8308 13394
rect 8364 13338 8388 13394
rect 8444 13338 8467 13394
rect 8046 13314 8467 13338
rect 8046 13258 8068 13314
rect 8124 13258 8148 13314
rect 8204 13258 8228 13314
rect 8284 13258 8308 13314
rect 8364 13258 8388 13314
rect 8444 13258 8467 13314
rect 8046 11072 8467 13258
rect 11304 13634 11764 13676
rect 11304 13578 11346 13634
rect 11402 13578 11426 13634
rect 11482 13578 11506 13634
rect 11562 13578 11586 13634
rect 11642 13578 11666 13634
rect 11722 13578 11764 13634
rect 11304 13554 11764 13578
rect 11304 13498 11346 13554
rect 11402 13498 11426 13554
rect 11482 13498 11506 13554
rect 11562 13498 11586 13554
rect 11642 13498 11666 13554
rect 11722 13498 11764 13554
rect 11304 13474 11764 13498
rect 11304 13418 11346 13474
rect 11402 13418 11426 13474
rect 11482 13418 11506 13474
rect 11562 13418 11586 13474
rect 11642 13418 11666 13474
rect 11722 13418 11764 13474
rect 11304 13394 11764 13418
rect 11304 13338 11346 13394
rect 11402 13338 11426 13394
rect 11482 13338 11506 13394
rect 11562 13338 11586 13394
rect 11642 13338 11666 13394
rect 11722 13338 11764 13394
rect 11304 13314 11764 13338
rect 11304 13258 11346 13314
rect 11402 13258 11426 13314
rect 11482 13258 11506 13314
rect 11562 13258 11586 13314
rect 11642 13258 11666 13314
rect 11722 13258 11764 13314
rect 9526 11158 10626 11256
rect 8046 11020 8070 11072
rect 8122 11020 8134 11072
rect 8186 11020 8198 11072
rect 8250 11020 8262 11072
rect 8314 11020 8326 11072
rect 8378 11020 8390 11072
rect 8442 11020 8467 11072
rect 7590 10766 7642 10772
rect 7590 10708 7642 10714
rect 7081 10476 7105 10528
rect 7157 10476 7169 10528
rect 7221 10476 7233 10528
rect 7285 10476 7297 10528
rect 7349 10476 7361 10528
rect 7413 10476 7425 10528
rect 7477 10476 7501 10528
rect 7081 9440 7501 10476
rect 7081 9388 7105 9440
rect 7157 9388 7169 9440
rect 7221 9388 7233 9440
rect 7285 9388 7297 9440
rect 7349 9388 7361 9440
rect 7413 9388 7425 9440
rect 7477 9388 7501 9440
rect 6578 8726 6630 8732
rect 6630 8674 6710 8680
rect 6578 8668 6710 8674
rect 6590 8652 6710 8668
rect 6578 8590 6630 8596
rect 6578 8532 6630 8538
rect 6590 8256 6618 8532
rect 6578 8250 6630 8256
rect 6578 8192 6630 8198
rect 6682 8120 6710 8652
rect 7081 8628 7501 9388
rect 7602 8800 7630 10708
rect 8046 9984 8467 11020
rect 9350 11130 10626 11158
rect 9350 10908 9378 11130
rect 9526 11032 10626 11130
rect 9338 10902 9390 10908
rect 9338 10844 9390 10850
rect 8046 9932 8070 9984
rect 8122 9932 8134 9984
rect 8186 9932 8198 9984
rect 8250 9932 8262 9984
rect 8314 9932 8326 9984
rect 8378 9932 8390 9984
rect 8442 9932 8467 9984
rect 8046 9903 8467 9932
rect 8046 9847 8068 9903
rect 8124 9847 8148 9903
rect 8204 9847 8228 9903
rect 8284 9847 8308 9903
rect 8364 9847 8388 9903
rect 8444 9847 8467 9903
rect 8046 9823 8467 9847
rect 8046 9767 8068 9823
rect 8124 9767 8148 9823
rect 8204 9767 8228 9823
rect 8284 9767 8308 9823
rect 8364 9767 8388 9823
rect 8444 9767 8467 9823
rect 8046 9743 8467 9767
rect 8046 9687 8068 9743
rect 8124 9687 8148 9743
rect 8204 9687 8228 9743
rect 8284 9687 8308 9743
rect 8364 9687 8388 9743
rect 8444 9687 8467 9743
rect 8046 9663 8467 9687
rect 8046 9607 8068 9663
rect 8124 9607 8148 9663
rect 8204 9607 8228 9663
rect 8284 9607 8308 9663
rect 8364 9607 8388 9663
rect 8444 9607 8467 9663
rect 8046 8896 8467 9607
rect 8046 8844 8070 8896
rect 8122 8844 8134 8896
rect 8186 8844 8198 8896
rect 8250 8844 8262 8896
rect 8314 8844 8326 8896
rect 8378 8844 8390 8896
rect 8442 8844 8467 8896
rect 7590 8794 7642 8800
rect 7590 8736 7642 8742
rect 6854 8590 6906 8596
rect 6854 8532 6906 8538
rect 7081 8572 7103 8628
rect 7159 8572 7183 8628
rect 7239 8572 7263 8628
rect 7319 8572 7343 8628
rect 7399 8572 7423 8628
rect 7479 8572 7501 8628
rect 7081 8548 7501 8572
rect 6762 8522 6814 8528
rect 6762 8464 6814 8470
rect 6670 8114 6722 8120
rect 6670 8056 6722 8062
rect 6116 7756 6140 7808
rect 6192 7756 6204 7808
rect 6256 7756 6268 7808
rect 6320 7756 6332 7808
rect 6384 7756 6396 7808
rect 6448 7756 6460 7808
rect 6512 7756 6536 7808
rect 6026 7502 6078 7508
rect 6026 7444 6078 7450
rect 6116 7354 6536 7756
rect 6670 7502 6722 7508
rect 6670 7444 6722 7450
rect 6116 7298 6138 7354
rect 6194 7298 6218 7354
rect 6274 7298 6298 7354
rect 6354 7298 6378 7354
rect 6434 7298 6458 7354
rect 6514 7298 6536 7354
rect 6116 7274 6536 7298
rect 6116 7218 6138 7274
rect 6194 7218 6218 7274
rect 6274 7218 6298 7274
rect 6354 7218 6378 7274
rect 6434 7218 6458 7274
rect 6514 7218 6536 7274
rect 6116 7194 6536 7218
rect 6116 7138 6138 7194
rect 6194 7138 6218 7194
rect 6274 7138 6298 7194
rect 6354 7138 6378 7194
rect 6434 7138 6458 7194
rect 6514 7138 6536 7194
rect 6116 7114 6536 7138
rect 6116 7058 6138 7114
rect 6194 7058 6218 7114
rect 6274 7058 6298 7114
rect 6354 7058 6378 7114
rect 6434 7058 6458 7114
rect 6514 7058 6536 7114
rect 5946 6896 6066 6912
rect 5946 6890 6078 6896
rect 5946 6884 6026 6890
rect 6026 6832 6078 6838
rect 5934 6822 5986 6828
rect 5934 6764 5986 6770
rect 5842 6618 5894 6624
rect 5842 6560 5894 6566
rect 5946 6420 5974 6764
rect 6038 6488 6066 6832
rect 6116 6720 6536 7058
rect 6578 7026 6630 7032
rect 6578 6968 6630 6974
rect 6116 6668 6140 6720
rect 6192 6668 6204 6720
rect 6256 6668 6268 6720
rect 6320 6668 6332 6720
rect 6384 6668 6396 6720
rect 6448 6668 6460 6720
rect 6512 6668 6536 6720
rect 6026 6482 6078 6488
rect 6026 6424 6078 6430
rect 5750 6414 5802 6420
rect 5750 6356 5802 6362
rect 5934 6414 5986 6420
rect 5934 6356 5986 6362
rect 5762 6284 5790 6356
rect 5658 6278 5710 6284
rect 5658 6220 5710 6226
rect 5750 6278 5802 6284
rect 5750 6220 5802 6226
rect 5150 6124 5174 6176
rect 5226 6124 5238 6176
rect 5290 6124 5302 6176
rect 5354 6124 5366 6176
rect 5418 6124 5430 6176
rect 5482 6124 5494 6176
rect 5546 6124 5571 6176
rect 5150 6079 5571 6124
rect 5150 6023 5172 6079
rect 5228 6023 5252 6079
rect 5308 6023 5332 6079
rect 5388 6023 5412 6079
rect 5468 6023 5492 6079
rect 5548 6023 5571 6079
rect 5150 5999 5571 6023
rect 5150 5943 5172 5999
rect 5228 5943 5252 5999
rect 5308 5943 5332 5999
rect 5388 5943 5412 5999
rect 5468 5943 5492 5999
rect 5548 5943 5571 5999
rect 5150 5919 5571 5943
rect 5150 5863 5172 5919
rect 5228 5863 5252 5919
rect 5308 5863 5332 5919
rect 5388 5863 5412 5919
rect 5468 5863 5492 5919
rect 5548 5863 5571 5919
rect 5150 5839 5571 5863
rect 5150 5783 5172 5839
rect 5228 5783 5252 5839
rect 5308 5783 5332 5839
rect 5388 5783 5412 5839
rect 5468 5783 5492 5839
rect 5548 5783 5571 5839
rect 5150 5088 5571 5783
rect 5670 5740 5698 6220
rect 5658 5734 5710 5740
rect 5658 5676 5710 5682
rect 5670 5468 5698 5676
rect 5762 5536 5790 6220
rect 5750 5530 5802 5536
rect 5750 5472 5802 5478
rect 5658 5462 5710 5468
rect 5658 5404 5710 5410
rect 5946 5332 5974 6356
rect 6116 5632 6536 6668
rect 6590 6624 6618 6968
rect 6682 6624 6710 7444
rect 6774 7168 6802 8464
rect 6866 7712 6894 8532
rect 7081 8492 7103 8548
rect 7159 8492 7183 8548
rect 7239 8492 7263 8548
rect 7319 8492 7343 8548
rect 7399 8492 7423 8548
rect 7479 8492 7501 8548
rect 7081 8468 7501 8492
rect 7081 8412 7103 8468
rect 7159 8412 7183 8468
rect 7239 8412 7263 8468
rect 7319 8412 7343 8468
rect 7399 8412 7423 8468
rect 7479 8412 7501 8468
rect 7081 8388 7501 8412
rect 7081 8332 7103 8388
rect 7159 8352 7183 8388
rect 7239 8352 7263 8388
rect 7319 8352 7343 8388
rect 7399 8352 7423 8388
rect 7159 8332 7169 8352
rect 7413 8332 7423 8352
rect 7479 8332 7501 8388
rect 7081 8300 7105 8332
rect 7157 8300 7169 8332
rect 7221 8300 7233 8332
rect 7285 8300 7297 8332
rect 7349 8300 7361 8332
rect 7413 8300 7425 8332
rect 7477 8300 7501 8332
rect 6946 8114 6998 8120
rect 6946 8056 6998 8062
rect 6854 7706 6906 7712
rect 6854 7648 6906 7654
rect 6762 7162 6814 7168
rect 6762 7104 6814 7110
rect 6578 6618 6630 6624
rect 6578 6560 6630 6566
rect 6670 6618 6722 6624
rect 6670 6560 6722 6566
rect 6116 5580 6140 5632
rect 6192 5580 6204 5632
rect 6256 5580 6268 5632
rect 6320 5580 6332 5632
rect 6384 5580 6396 5632
rect 6448 5580 6460 5632
rect 6512 5580 6536 5632
rect 5934 5326 5986 5332
rect 5934 5268 5986 5274
rect 5150 5036 5174 5088
rect 5226 5036 5238 5088
rect 5290 5036 5302 5088
rect 5354 5036 5366 5088
rect 5418 5036 5430 5088
rect 5482 5036 5494 5088
rect 5546 5036 5571 5088
rect 5150 4000 5571 5036
rect 5150 3948 5174 4000
rect 5226 3948 5238 4000
rect 5290 3948 5302 4000
rect 5354 3948 5366 4000
rect 5418 3948 5430 4000
rect 5482 3948 5494 4000
rect 5546 3948 5571 4000
rect 5150 418 5571 3948
rect 5150 362 5172 418
rect 5228 362 5252 418
rect 5308 362 5332 418
rect 5388 362 5412 418
rect 5468 362 5492 418
rect 5548 362 5571 418
rect 5150 338 5571 362
rect 5150 282 5172 338
rect 5228 282 5252 338
rect 5308 282 5332 338
rect 5388 282 5412 338
rect 5468 282 5492 338
rect 5548 282 5571 338
rect 5150 258 5571 282
rect 5150 202 5172 258
rect 5228 202 5252 258
rect 5308 202 5332 258
rect 5388 202 5412 258
rect 5468 202 5492 258
rect 5548 202 5571 258
rect 5150 178 5571 202
rect 5150 122 5172 178
rect 5228 122 5252 178
rect 5308 122 5332 178
rect 5388 122 5412 178
rect 5468 122 5492 178
rect 5548 122 5571 178
rect 5150 98 5571 122
rect 5150 42 5172 98
rect 5228 42 5252 98
rect 5308 42 5332 98
rect 5388 42 5412 98
rect 5468 42 5492 98
rect 5548 42 5571 98
rect 5150 0 5571 42
rect 6116 4804 6536 5580
rect 6590 5264 6618 6560
rect 6958 5332 6986 8056
rect 7081 7264 7501 8300
rect 7602 7576 7630 8736
rect 8046 7808 8467 8844
rect 8046 7756 8070 7808
rect 8122 7756 8134 7808
rect 8186 7756 8198 7808
rect 8250 7756 8262 7808
rect 8314 7756 8326 7808
rect 8378 7756 8390 7808
rect 8442 7756 8467 7808
rect 7590 7570 7642 7576
rect 7590 7512 7642 7518
rect 7081 7212 7105 7264
rect 7157 7212 7169 7264
rect 7221 7212 7233 7264
rect 7285 7212 7297 7264
rect 7349 7212 7361 7264
rect 7413 7212 7425 7264
rect 7477 7212 7501 7264
rect 7081 6176 7501 7212
rect 7081 6124 7105 6176
rect 7157 6124 7169 6176
rect 7221 6124 7233 6176
rect 7285 6124 7297 6176
rect 7349 6124 7361 6176
rect 7413 6124 7425 6176
rect 7477 6124 7501 6176
rect 7081 6079 7501 6124
rect 7081 6023 7103 6079
rect 7159 6023 7183 6079
rect 7239 6023 7263 6079
rect 7319 6023 7343 6079
rect 7399 6023 7423 6079
rect 7479 6023 7501 6079
rect 7081 5999 7501 6023
rect 7081 5943 7103 5999
rect 7159 5943 7183 5999
rect 7239 5943 7263 5999
rect 7319 5943 7343 5999
rect 7399 5943 7423 5999
rect 7479 5943 7501 5999
rect 7081 5919 7501 5943
rect 7081 5863 7103 5919
rect 7159 5863 7183 5919
rect 7239 5863 7263 5919
rect 7319 5863 7343 5919
rect 7399 5863 7423 5919
rect 7479 5863 7501 5919
rect 7081 5839 7501 5863
rect 7081 5783 7103 5839
rect 7159 5783 7183 5839
rect 7239 5783 7263 5839
rect 7319 5783 7343 5839
rect 7399 5783 7423 5839
rect 7479 5783 7501 5839
rect 6946 5326 6998 5332
rect 6946 5268 6998 5274
rect 6578 5258 6630 5264
rect 6578 5200 6630 5206
rect 6116 4748 6138 4804
rect 6194 4748 6218 4804
rect 6274 4748 6298 4804
rect 6354 4748 6378 4804
rect 6434 4748 6458 4804
rect 6514 4748 6536 4804
rect 6116 4724 6536 4748
rect 6116 4668 6138 4724
rect 6194 4668 6218 4724
rect 6274 4668 6298 4724
rect 6354 4668 6378 4724
rect 6434 4668 6458 4724
rect 6514 4668 6536 4724
rect 6116 4644 6536 4668
rect 6116 4588 6138 4644
rect 6194 4588 6218 4644
rect 6274 4588 6298 4644
rect 6354 4588 6378 4644
rect 6434 4588 6458 4644
rect 6514 4588 6536 4644
rect 6116 4564 6536 4588
rect 6116 4508 6138 4564
rect 6194 4544 6218 4564
rect 6274 4544 6298 4564
rect 6354 4544 6378 4564
rect 6434 4544 6458 4564
rect 6194 4508 6204 4544
rect 6448 4508 6458 4544
rect 6514 4508 6536 4564
rect 6116 4492 6140 4508
rect 6192 4492 6204 4508
rect 6256 4492 6268 4508
rect 6320 4492 6332 4508
rect 6384 4492 6396 4508
rect 6448 4492 6460 4508
rect 6512 4492 6536 4508
rect 6116 3456 6536 4492
rect 6116 3404 6140 3456
rect 6192 3404 6204 3456
rect 6256 3404 6268 3456
rect 6320 3404 6332 3456
rect 6384 3404 6396 3456
rect 6448 3404 6460 3456
rect 6512 3404 6536 3456
rect 6116 1218 6536 3404
rect 6116 1162 6138 1218
rect 6194 1162 6218 1218
rect 6274 1162 6298 1218
rect 6354 1162 6378 1218
rect 6434 1162 6458 1218
rect 6514 1162 6536 1218
rect 6116 1138 6536 1162
rect 6116 1082 6138 1138
rect 6194 1082 6218 1138
rect 6274 1082 6298 1138
rect 6354 1082 6378 1138
rect 6434 1082 6458 1138
rect 6514 1082 6536 1138
rect 6116 1058 6536 1082
rect 6116 1002 6138 1058
rect 6194 1002 6218 1058
rect 6274 1002 6298 1058
rect 6354 1002 6378 1058
rect 6434 1002 6458 1058
rect 6514 1002 6536 1058
rect 6116 978 6536 1002
rect 6116 922 6138 978
rect 6194 922 6218 978
rect 6274 922 6298 978
rect 6354 922 6378 978
rect 6434 922 6458 978
rect 6514 922 6536 978
rect 6116 898 6536 922
rect 6116 842 6138 898
rect 6194 842 6218 898
rect 6274 842 6298 898
rect 6354 842 6378 898
rect 6434 842 6458 898
rect 6514 842 6536 898
rect 6116 0 6536 842
rect 7081 5088 7501 5783
rect 8046 7354 8467 7756
rect 8046 7298 8068 7354
rect 8124 7298 8148 7354
rect 8204 7298 8228 7354
rect 8284 7298 8308 7354
rect 8364 7298 8388 7354
rect 8444 7298 8467 7354
rect 11304 9903 11764 13258
rect 11304 9847 11346 9903
rect 11402 9847 11426 9903
rect 11482 9847 11506 9903
rect 11562 9847 11586 9903
rect 11642 9847 11666 9903
rect 11722 9847 11764 9903
rect 11304 9823 11764 9847
rect 11304 9767 11346 9823
rect 11402 9767 11426 9823
rect 11482 9767 11506 9823
rect 11562 9767 11586 9823
rect 11642 9767 11666 9823
rect 11722 9767 11764 9823
rect 11304 9743 11764 9767
rect 11304 9687 11346 9743
rect 11402 9687 11426 9743
rect 11482 9687 11506 9743
rect 11562 9687 11586 9743
rect 11642 9687 11666 9743
rect 11722 9687 11764 9743
rect 11304 9663 11764 9687
rect 11304 9607 11346 9663
rect 11402 9607 11426 9663
rect 11482 9607 11506 9663
rect 11562 9607 11586 9663
rect 11642 9607 11666 9663
rect 11722 9607 11764 9663
rect 11304 7354 11764 9607
rect 8046 7274 8467 7298
rect 8046 7218 8068 7274
rect 8124 7218 8148 7274
rect 8204 7218 8228 7274
rect 8284 7218 8308 7274
rect 8364 7218 8388 7274
rect 8444 7218 8467 7274
rect 8046 7194 8467 7218
rect 9526 7202 10626 7300
rect 8046 7138 8068 7194
rect 8124 7138 8148 7194
rect 8204 7138 8228 7194
rect 8284 7138 8308 7194
rect 8364 7138 8388 7194
rect 8444 7138 8467 7194
rect 8046 7114 8467 7138
rect 8046 7058 8068 7114
rect 8124 7058 8148 7114
rect 8204 7058 8228 7114
rect 8284 7058 8308 7114
rect 8364 7058 8388 7114
rect 8444 7058 8467 7114
rect 8046 6720 8467 7058
rect 9350 7174 10626 7202
rect 9350 7032 9378 7174
rect 9526 7076 10626 7174
rect 11304 7298 11346 7354
rect 11402 7298 11426 7354
rect 11482 7298 11506 7354
rect 11562 7298 11586 7354
rect 11642 7298 11666 7354
rect 11722 7298 11764 7354
rect 11304 7274 11764 7298
rect 11304 7218 11346 7274
rect 11402 7218 11426 7274
rect 11482 7218 11506 7274
rect 11562 7218 11586 7274
rect 11642 7218 11666 7274
rect 11722 7218 11764 7274
rect 11304 7194 11764 7218
rect 11304 7138 11346 7194
rect 11402 7138 11426 7194
rect 11482 7138 11506 7194
rect 11562 7138 11586 7194
rect 11642 7138 11666 7194
rect 11722 7138 11764 7194
rect 11304 7114 11764 7138
rect 11304 7058 11346 7114
rect 11402 7058 11426 7114
rect 11482 7058 11506 7114
rect 11562 7058 11586 7114
rect 11642 7058 11666 7114
rect 11722 7058 11764 7114
rect 9338 7026 9390 7032
rect 9338 6968 9390 6974
rect 8046 6668 8070 6720
rect 8122 6668 8134 6720
rect 8186 6668 8198 6720
rect 8250 6668 8262 6720
rect 8314 6668 8326 6720
rect 8378 6668 8390 6720
rect 8442 6668 8467 6720
rect 8046 5632 8467 6668
rect 8046 5580 8070 5632
rect 8122 5580 8134 5632
rect 8186 5580 8198 5632
rect 8250 5580 8262 5632
rect 8314 5580 8326 5632
rect 8378 5580 8390 5632
rect 8442 5580 8467 5632
rect 7866 5326 7918 5332
rect 7866 5268 7918 5274
rect 7081 5036 7105 5088
rect 7157 5036 7169 5088
rect 7221 5036 7233 5088
rect 7285 5036 7297 5088
rect 7349 5036 7361 5088
rect 7413 5036 7425 5088
rect 7477 5036 7501 5088
rect 7081 4000 7501 5036
rect 7081 3948 7105 4000
rect 7157 3948 7169 4000
rect 7221 3948 7233 4000
rect 7285 3948 7297 4000
rect 7349 3948 7361 4000
rect 7413 3948 7425 4000
rect 7477 3948 7501 4000
rect 7081 418 7501 3948
rect 7878 3904 7906 5268
rect 8046 4804 8467 5580
rect 8046 4748 8068 4804
rect 8124 4748 8148 4804
rect 8204 4748 8228 4804
rect 8284 4748 8308 4804
rect 8364 4748 8388 4804
rect 8444 4748 8467 4804
rect 8046 4724 8467 4748
rect 8046 4668 8068 4724
rect 8124 4668 8148 4724
rect 8204 4668 8228 4724
rect 8284 4668 8308 4724
rect 8364 4668 8388 4724
rect 8444 4668 8467 4724
rect 8046 4644 8467 4668
rect 8046 4588 8068 4644
rect 8124 4588 8148 4644
rect 8204 4588 8228 4644
rect 8284 4588 8308 4644
rect 8364 4588 8388 4644
rect 8444 4588 8467 4644
rect 8046 4564 8467 4588
rect 8046 4508 8068 4564
rect 8124 4544 8148 4564
rect 8204 4544 8228 4564
rect 8284 4544 8308 4564
rect 8364 4544 8388 4564
rect 8124 4508 8134 4544
rect 8378 4508 8388 4544
rect 8444 4508 8467 4564
rect 8046 4492 8070 4508
rect 8122 4492 8134 4508
rect 8186 4492 8198 4508
rect 8250 4492 8262 4508
rect 8314 4492 8326 4508
rect 8378 4492 8390 4508
rect 8442 4492 8467 4508
rect 7866 3898 7918 3904
rect 7866 3840 7918 3846
rect 7081 362 7103 418
rect 7159 362 7183 418
rect 7239 362 7263 418
rect 7319 362 7343 418
rect 7399 362 7423 418
rect 7479 362 7501 418
rect 7081 338 7501 362
rect 7081 282 7103 338
rect 7159 282 7183 338
rect 7239 282 7263 338
rect 7319 282 7343 338
rect 7399 282 7423 338
rect 7479 282 7501 338
rect 7081 258 7501 282
rect 7081 202 7103 258
rect 7159 202 7183 258
rect 7239 202 7263 258
rect 7319 202 7343 258
rect 7399 202 7423 258
rect 7479 202 7501 258
rect 7081 178 7501 202
rect 7081 122 7103 178
rect 7159 122 7183 178
rect 7239 122 7263 178
rect 7319 122 7343 178
rect 7399 122 7423 178
rect 7479 122 7501 178
rect 7081 98 7501 122
rect 7081 42 7103 98
rect 7159 42 7183 98
rect 7239 42 7263 98
rect 7319 42 7343 98
rect 7399 42 7423 98
rect 7479 42 7501 98
rect 7081 0 7501 42
rect 8046 3456 8467 4492
rect 11304 4804 11764 7058
rect 11304 4748 11346 4804
rect 11402 4748 11426 4804
rect 11482 4748 11506 4804
rect 11562 4748 11586 4804
rect 11642 4748 11666 4804
rect 11722 4748 11764 4804
rect 11304 4724 11764 4748
rect 11304 4668 11346 4724
rect 11402 4668 11426 4724
rect 11482 4668 11506 4724
rect 11562 4668 11586 4724
rect 11642 4668 11666 4724
rect 11722 4668 11764 4724
rect 11304 4644 11764 4668
rect 11304 4588 11346 4644
rect 11402 4588 11426 4644
rect 11482 4588 11506 4644
rect 11562 4588 11586 4644
rect 11642 4588 11666 4644
rect 11722 4588 11764 4644
rect 11304 4564 11764 4588
rect 11304 4508 11346 4564
rect 11402 4508 11426 4564
rect 11482 4508 11506 4564
rect 11562 4508 11586 4564
rect 11642 4508 11666 4564
rect 11722 4508 11764 4564
rect 9338 3762 9390 3768
rect 9338 3704 9390 3710
rect 8046 3404 8070 3456
rect 8122 3404 8134 3456
rect 8186 3404 8198 3456
rect 8250 3404 8262 3456
rect 8314 3404 8326 3456
rect 8378 3404 8390 3456
rect 8442 3404 8467 3456
rect 8046 1218 8467 3404
rect 9350 3246 9378 3704
rect 9526 3246 10626 3344
rect 9350 3218 10626 3246
rect 9526 3120 10626 3218
rect 8046 1162 8068 1218
rect 8124 1162 8148 1218
rect 8204 1162 8228 1218
rect 8284 1162 8308 1218
rect 8364 1162 8388 1218
rect 8444 1162 8467 1218
rect 8046 1138 8467 1162
rect 8046 1082 8068 1138
rect 8124 1082 8148 1138
rect 8204 1082 8228 1138
rect 8284 1082 8308 1138
rect 8364 1082 8388 1138
rect 8444 1082 8467 1138
rect 8046 1058 8467 1082
rect 8046 1002 8068 1058
rect 8124 1002 8148 1058
rect 8204 1002 8228 1058
rect 8284 1002 8308 1058
rect 8364 1002 8388 1058
rect 8444 1002 8467 1058
rect 8046 978 8467 1002
rect 8046 922 8068 978
rect 8124 922 8148 978
rect 8204 922 8228 978
rect 8284 922 8308 978
rect 8364 922 8388 978
rect 8444 922 8467 978
rect 8046 898 8467 922
rect 8046 842 8068 898
rect 8124 842 8148 898
rect 8204 842 8228 898
rect 8284 842 8308 898
rect 8364 842 8388 898
rect 8444 842 8467 898
rect 8046 0 8467 842
rect 11304 1218 11764 4508
rect 11304 1162 11346 1218
rect 11402 1162 11426 1218
rect 11482 1162 11506 1218
rect 11562 1162 11586 1218
rect 11642 1162 11666 1218
rect 11722 1162 11764 1218
rect 11304 1138 11764 1162
rect 11304 1082 11346 1138
rect 11402 1082 11426 1138
rect 11482 1082 11506 1138
rect 11562 1082 11586 1138
rect 11642 1082 11666 1138
rect 11722 1082 11764 1138
rect 11304 1058 11764 1082
rect 11304 1002 11346 1058
rect 11402 1002 11426 1058
rect 11482 1002 11506 1058
rect 11562 1002 11586 1058
rect 11642 1002 11666 1058
rect 11722 1002 11764 1058
rect 11304 978 11764 1002
rect 11304 922 11346 978
rect 11402 922 11426 978
rect 11482 922 11506 978
rect 11562 922 11586 978
rect 11642 922 11666 978
rect 11722 922 11764 978
rect 11304 898 11764 922
rect 11304 842 11346 898
rect 11402 842 11426 898
rect 11482 842 11506 898
rect 11562 842 11586 898
rect 11642 842 11666 898
rect 11722 842 11764 898
rect 11304 800 11764 842
rect 12104 8628 12564 14058
rect 12104 8572 12146 8628
rect 12202 8572 12226 8628
rect 12282 8572 12306 8628
rect 12362 8572 12386 8628
rect 12442 8572 12466 8628
rect 12522 8572 12564 8628
rect 12104 8548 12564 8572
rect 12104 8492 12146 8548
rect 12202 8492 12226 8548
rect 12282 8492 12306 8548
rect 12362 8492 12386 8548
rect 12442 8492 12466 8548
rect 12522 8492 12564 8548
rect 12104 8468 12564 8492
rect 12104 8412 12146 8468
rect 12202 8412 12226 8468
rect 12282 8412 12306 8468
rect 12362 8412 12386 8468
rect 12442 8412 12466 8468
rect 12522 8412 12564 8468
rect 12104 8388 12564 8412
rect 12104 8332 12146 8388
rect 12202 8332 12226 8388
rect 12282 8332 12306 8388
rect 12362 8332 12386 8388
rect 12442 8332 12466 8388
rect 12522 8332 12564 8388
rect 12104 6079 12564 8332
rect 12104 6023 12146 6079
rect 12202 6023 12226 6079
rect 12282 6023 12306 6079
rect 12362 6023 12386 6079
rect 12442 6023 12466 6079
rect 12522 6023 12564 6079
rect 12104 5999 12564 6023
rect 12104 5943 12146 5999
rect 12202 5943 12226 5999
rect 12282 5943 12306 5999
rect 12362 5943 12386 5999
rect 12442 5943 12466 5999
rect 12522 5943 12564 5999
rect 12104 5919 12564 5943
rect 12104 5863 12146 5919
rect 12202 5863 12226 5919
rect 12282 5863 12306 5919
rect 12362 5863 12386 5919
rect 12442 5863 12466 5919
rect 12522 5863 12564 5919
rect 12104 5839 12564 5863
rect 12104 5783 12146 5839
rect 12202 5783 12226 5839
rect 12282 5783 12306 5839
rect 12362 5783 12386 5839
rect 12442 5783 12466 5839
rect 12522 5783 12564 5839
rect 12104 418 12564 5783
rect 12104 362 12146 418
rect 12202 362 12226 418
rect 12282 362 12306 418
rect 12362 362 12386 418
rect 12442 362 12466 418
rect 12522 362 12564 418
rect 12104 338 12564 362
rect 12104 282 12146 338
rect 12202 282 12226 338
rect 12282 282 12306 338
rect 12362 282 12386 338
rect 12442 282 12466 338
rect 12522 282 12564 338
rect 12104 258 12564 282
rect 12104 202 12146 258
rect 12202 202 12226 258
rect 12282 202 12306 258
rect 12362 202 12386 258
rect 12442 202 12466 258
rect 12522 202 12564 258
rect 12104 178 12564 202
rect 12104 122 12146 178
rect 12202 122 12226 178
rect 12282 122 12306 178
rect 12362 122 12386 178
rect 12442 122 12466 178
rect 12522 122 12564 178
rect 12104 98 12564 122
rect 12104 42 12146 98
rect 12202 42 12226 98
rect 12282 42 12306 98
rect 12362 42 12386 98
rect 12442 42 12466 98
rect 12522 42 12564 98
rect 12104 0 12564 42
<< via2 >>
rect 42 14378 98 14434
rect 122 14378 178 14434
rect 202 14378 258 14434
rect 282 14378 338 14434
rect 362 14378 418 14434
rect 42 14298 98 14354
rect 122 14298 178 14354
rect 202 14298 258 14354
rect 282 14298 338 14354
rect 362 14298 418 14354
rect 42 14218 98 14274
rect 122 14218 178 14274
rect 202 14218 258 14274
rect 282 14218 338 14274
rect 362 14218 418 14274
rect 42 14138 98 14194
rect 122 14138 178 14194
rect 202 14138 258 14194
rect 282 14138 338 14194
rect 362 14138 418 14194
rect 42 14058 98 14114
rect 122 14058 178 14114
rect 202 14058 258 14114
rect 282 14058 338 14114
rect 362 14058 418 14114
rect 42 8572 98 8628
rect 122 8572 178 8628
rect 202 8572 258 8628
rect 282 8572 338 8628
rect 362 8572 418 8628
rect 42 8492 98 8548
rect 122 8492 178 8548
rect 202 8492 258 8548
rect 282 8492 338 8548
rect 362 8492 418 8548
rect 42 8412 98 8468
rect 122 8412 178 8468
rect 202 8412 258 8468
rect 282 8412 338 8468
rect 362 8412 418 8468
rect 42 8332 98 8388
rect 122 8332 178 8388
rect 202 8332 258 8388
rect 282 8332 338 8388
rect 362 8332 418 8388
rect 42 6023 98 6079
rect 122 6023 178 6079
rect 202 6023 258 6079
rect 282 6023 338 6079
rect 362 6023 418 6079
rect 42 5943 98 5999
rect 122 5943 178 5999
rect 202 5943 258 5999
rect 282 5943 338 5999
rect 362 5943 418 5999
rect 42 5863 98 5919
rect 122 5863 178 5919
rect 202 5863 258 5919
rect 282 5863 338 5919
rect 362 5863 418 5919
rect 42 5783 98 5839
rect 122 5783 178 5839
rect 202 5783 258 5839
rect 282 5783 338 5839
rect 362 5783 418 5839
rect 842 13578 898 13634
rect 922 13578 978 13634
rect 1002 13578 1058 13634
rect 1082 13578 1138 13634
rect 1162 13578 1218 13634
rect 842 13498 898 13554
rect 922 13498 978 13554
rect 1002 13498 1058 13554
rect 1082 13498 1138 13554
rect 1162 13498 1218 13554
rect 842 13418 898 13474
rect 922 13418 978 13474
rect 1002 13418 1058 13474
rect 1082 13418 1138 13474
rect 1162 13418 1218 13474
rect 842 13338 898 13394
rect 922 13338 978 13394
rect 1002 13338 1058 13394
rect 1082 13338 1138 13394
rect 1162 13338 1218 13394
rect 842 13258 898 13314
rect 922 13258 978 13314
rect 1002 13258 1058 13314
rect 1082 13258 1138 13314
rect 1162 13258 1218 13314
rect 4207 13578 4263 13634
rect 4287 13578 4343 13634
rect 4367 13578 4423 13634
rect 4447 13578 4503 13634
rect 4527 13578 4583 13634
rect 4207 13498 4263 13554
rect 4287 13498 4343 13554
rect 4367 13498 4423 13554
rect 4447 13498 4503 13554
rect 4527 13498 4583 13554
rect 4207 13418 4263 13474
rect 4287 13418 4343 13474
rect 4367 13418 4423 13474
rect 4447 13418 4503 13474
rect 4527 13418 4583 13474
rect 4207 13338 4263 13394
rect 4287 13338 4343 13394
rect 4367 13338 4423 13394
rect 4447 13338 4503 13394
rect 4527 13338 4583 13394
rect 4207 13258 4263 13314
rect 4287 13258 4343 13314
rect 4367 13258 4423 13314
rect 4447 13258 4503 13314
rect 4527 13258 4583 13314
rect 842 9847 898 9903
rect 922 9847 978 9903
rect 1002 9847 1058 9903
rect 1082 9847 1138 9903
rect 1162 9847 1218 9903
rect 842 9767 898 9823
rect 922 9767 978 9823
rect 1002 9767 1058 9823
rect 1082 9767 1138 9823
rect 1162 9767 1218 9823
rect 842 9687 898 9743
rect 922 9687 978 9743
rect 1002 9687 1058 9743
rect 1082 9687 1138 9743
rect 1162 9687 1218 9743
rect 842 9607 898 9663
rect 922 9607 978 9663
rect 1002 9607 1058 9663
rect 1082 9607 1138 9663
rect 1162 9607 1218 9663
rect 842 7298 898 7354
rect 922 7298 978 7354
rect 1002 7298 1058 7354
rect 1082 7298 1138 7354
rect 1162 7298 1218 7354
rect 4207 9847 4263 9903
rect 4287 9847 4343 9903
rect 4367 9847 4423 9903
rect 4447 9847 4503 9903
rect 4527 9847 4583 9903
rect 4207 9767 4263 9823
rect 4287 9767 4343 9823
rect 4367 9767 4423 9823
rect 4447 9767 4503 9823
rect 4527 9767 4583 9823
rect 4207 9687 4263 9743
rect 4287 9687 4343 9743
rect 4367 9687 4423 9743
rect 4447 9687 4503 9743
rect 4527 9687 4583 9743
rect 4207 9607 4263 9663
rect 4287 9607 4343 9663
rect 4367 9607 4423 9663
rect 4447 9607 4503 9663
rect 4527 9607 4583 9663
rect 842 7218 898 7274
rect 922 7218 978 7274
rect 1002 7218 1058 7274
rect 1082 7218 1138 7274
rect 1162 7218 1218 7274
rect 842 7138 898 7194
rect 922 7138 978 7194
rect 1002 7138 1058 7194
rect 1082 7138 1138 7194
rect 1162 7138 1218 7194
rect 842 7058 898 7114
rect 922 7058 978 7114
rect 1002 7058 1058 7114
rect 1082 7058 1138 7114
rect 1162 7058 1218 7114
rect 4207 7298 4263 7354
rect 4287 7298 4343 7354
rect 4367 7298 4423 7354
rect 4447 7298 4503 7354
rect 4527 7298 4583 7354
rect 4207 7218 4263 7274
rect 4287 7218 4343 7274
rect 4367 7218 4423 7274
rect 4447 7218 4503 7274
rect 4527 7218 4583 7274
rect 4207 7138 4263 7194
rect 4287 7138 4343 7194
rect 4367 7138 4423 7194
rect 4447 7138 4503 7194
rect 4527 7138 4583 7194
rect 4207 7058 4263 7114
rect 4287 7058 4343 7114
rect 4367 7058 4423 7114
rect 4447 7058 4503 7114
rect 4527 7058 4583 7114
rect 842 4748 898 4804
rect 922 4748 978 4804
rect 1002 4748 1058 4804
rect 1082 4748 1138 4804
rect 1162 4748 1218 4804
rect 842 4668 898 4724
rect 922 4668 978 4724
rect 1002 4668 1058 4724
rect 1082 4668 1138 4724
rect 1162 4668 1218 4724
rect 842 4588 898 4644
rect 922 4588 978 4644
rect 1002 4588 1058 4644
rect 1082 4588 1138 4644
rect 1162 4588 1218 4644
rect 842 4508 898 4564
rect 922 4508 978 4564
rect 1002 4508 1058 4564
rect 1082 4508 1138 4564
rect 1162 4508 1218 4564
rect 4207 4748 4263 4804
rect 4287 4748 4343 4804
rect 4367 4748 4423 4804
rect 4447 4748 4503 4804
rect 4527 4748 4583 4804
rect 4207 4668 4263 4724
rect 4287 4668 4343 4724
rect 4367 4668 4423 4724
rect 4447 4668 4503 4724
rect 4527 4668 4583 4724
rect 4207 4588 4263 4644
rect 4287 4588 4343 4644
rect 4367 4588 4423 4644
rect 4447 4588 4503 4644
rect 4527 4588 4583 4644
rect 4207 4544 4263 4564
rect 4287 4544 4343 4564
rect 4367 4544 4423 4564
rect 4447 4544 4503 4564
rect 4527 4544 4583 4564
rect 4207 4508 4209 4544
rect 4209 4508 4261 4544
rect 4261 4508 4263 4544
rect 4287 4508 4325 4544
rect 4325 4508 4337 4544
rect 4337 4508 4343 4544
rect 4367 4508 4389 4544
rect 4389 4508 4401 4544
rect 4401 4508 4423 4544
rect 4447 4508 4453 4544
rect 4453 4508 4465 4544
rect 4465 4508 4503 4544
rect 4527 4508 4529 4544
rect 4529 4508 4581 4544
rect 4581 4508 4583 4544
rect 842 1162 898 1218
rect 922 1162 978 1218
rect 1002 1162 1058 1218
rect 1082 1162 1138 1218
rect 1162 1162 1218 1218
rect 842 1082 898 1138
rect 922 1082 978 1138
rect 1002 1082 1058 1138
rect 1082 1082 1138 1138
rect 1162 1082 1218 1138
rect 842 1002 898 1058
rect 922 1002 978 1058
rect 1002 1002 1058 1058
rect 1082 1002 1138 1058
rect 1162 1002 1218 1058
rect 842 922 898 978
rect 922 922 978 978
rect 1002 922 1058 978
rect 1082 922 1138 978
rect 1162 922 1218 978
rect 842 842 898 898
rect 922 842 978 898
rect 1002 842 1058 898
rect 1082 842 1138 898
rect 1162 842 1218 898
rect 4207 1162 4263 1218
rect 4287 1162 4343 1218
rect 4367 1162 4423 1218
rect 4447 1162 4503 1218
rect 4527 1162 4583 1218
rect 4207 1082 4263 1138
rect 4287 1082 4343 1138
rect 4367 1082 4423 1138
rect 4447 1082 4503 1138
rect 4527 1082 4583 1138
rect 4207 1002 4263 1058
rect 4287 1002 4343 1058
rect 4367 1002 4423 1058
rect 4447 1002 4503 1058
rect 4527 1002 4583 1058
rect 4207 922 4263 978
rect 4287 922 4343 978
rect 4367 922 4423 978
rect 4447 922 4503 978
rect 4527 922 4583 978
rect 4207 842 4263 898
rect 4287 842 4343 898
rect 4367 842 4423 898
rect 4447 842 4503 898
rect 4527 842 4583 898
rect 42 362 98 418
rect 122 362 178 418
rect 202 362 258 418
rect 282 362 338 418
rect 362 362 418 418
rect 42 282 98 338
rect 122 282 178 338
rect 202 282 258 338
rect 282 282 338 338
rect 362 282 418 338
rect 42 202 98 258
rect 122 202 178 258
rect 202 202 258 258
rect 282 202 338 258
rect 362 202 418 258
rect 42 122 98 178
rect 122 122 178 178
rect 202 122 258 178
rect 282 122 338 178
rect 362 122 418 178
rect 42 42 98 98
rect 122 42 178 98
rect 202 42 258 98
rect 282 42 338 98
rect 362 42 418 98
rect 5172 14378 5228 14434
rect 5252 14378 5308 14434
rect 5332 14378 5388 14434
rect 5412 14378 5468 14434
rect 5492 14378 5548 14434
rect 5172 14298 5228 14354
rect 5252 14298 5308 14354
rect 5332 14298 5388 14354
rect 5412 14298 5468 14354
rect 5492 14298 5548 14354
rect 5172 14218 5228 14274
rect 5252 14218 5308 14274
rect 5332 14218 5388 14274
rect 5412 14218 5468 14274
rect 5492 14218 5548 14274
rect 5172 14138 5228 14194
rect 5252 14138 5308 14194
rect 5332 14138 5388 14194
rect 5412 14138 5468 14194
rect 5492 14138 5548 14194
rect 5172 14058 5228 14114
rect 5252 14058 5308 14114
rect 5332 14058 5388 14114
rect 5412 14058 5468 14114
rect 5492 14058 5548 14114
rect 6138 13578 6194 13634
rect 6218 13578 6274 13634
rect 6298 13578 6354 13634
rect 6378 13578 6434 13634
rect 6458 13578 6514 13634
rect 6138 13498 6194 13554
rect 6218 13498 6274 13554
rect 6298 13498 6354 13554
rect 6378 13498 6434 13554
rect 6458 13498 6514 13554
rect 6138 13418 6194 13474
rect 6218 13418 6274 13474
rect 6298 13418 6354 13474
rect 6378 13418 6434 13474
rect 6458 13418 6514 13474
rect 6138 13338 6194 13394
rect 6218 13338 6274 13394
rect 6298 13338 6354 13394
rect 6378 13338 6434 13394
rect 6458 13338 6514 13394
rect 6138 13258 6194 13314
rect 6218 13258 6274 13314
rect 6298 13258 6354 13314
rect 6378 13258 6434 13314
rect 6458 13258 6514 13314
rect 7103 14378 7159 14434
rect 7183 14378 7239 14434
rect 7263 14378 7319 14434
rect 7343 14378 7399 14434
rect 7423 14378 7479 14434
rect 7103 14298 7159 14354
rect 7183 14298 7239 14354
rect 7263 14298 7319 14354
rect 7343 14298 7399 14354
rect 7423 14298 7479 14354
rect 7103 14218 7159 14274
rect 7183 14218 7239 14274
rect 7263 14218 7319 14274
rect 7343 14218 7399 14274
rect 7423 14218 7479 14274
rect 7103 14138 7159 14194
rect 7183 14138 7239 14194
rect 7263 14138 7319 14194
rect 7343 14138 7399 14194
rect 7423 14138 7479 14194
rect 7103 14058 7159 14114
rect 7183 14058 7239 14114
rect 7263 14058 7319 14114
rect 7343 14058 7399 14114
rect 7423 14058 7479 14114
rect 6138 9847 6194 9903
rect 6218 9847 6274 9903
rect 6298 9847 6354 9903
rect 6378 9847 6434 9903
rect 6458 9847 6514 9903
rect 6138 9767 6194 9823
rect 6218 9767 6274 9823
rect 6298 9767 6354 9823
rect 6378 9767 6434 9823
rect 6458 9767 6514 9823
rect 6138 9687 6194 9743
rect 6218 9687 6274 9743
rect 6298 9687 6354 9743
rect 6378 9687 6434 9743
rect 6458 9687 6514 9743
rect 6138 9607 6194 9663
rect 6218 9607 6274 9663
rect 6298 9607 6354 9663
rect 6378 9607 6434 9663
rect 6458 9607 6514 9663
rect 5172 8572 5228 8628
rect 5252 8572 5308 8628
rect 5332 8572 5388 8628
rect 5412 8572 5468 8628
rect 5492 8572 5548 8628
rect 5172 8492 5228 8548
rect 5252 8492 5308 8548
rect 5332 8492 5388 8548
rect 5412 8492 5468 8548
rect 5492 8492 5548 8548
rect 5172 8412 5228 8468
rect 5252 8412 5308 8468
rect 5332 8412 5388 8468
rect 5412 8412 5468 8468
rect 5492 8412 5548 8468
rect 5172 8352 5228 8388
rect 5252 8352 5308 8388
rect 5332 8352 5388 8388
rect 5412 8352 5468 8388
rect 5492 8352 5548 8388
rect 5172 8332 5174 8352
rect 5174 8332 5226 8352
rect 5226 8332 5228 8352
rect 5252 8332 5290 8352
rect 5290 8332 5302 8352
rect 5302 8332 5308 8352
rect 5332 8332 5354 8352
rect 5354 8332 5366 8352
rect 5366 8332 5388 8352
rect 5412 8332 5418 8352
rect 5418 8332 5430 8352
rect 5430 8332 5468 8352
rect 5492 8332 5494 8352
rect 5494 8332 5546 8352
rect 5546 8332 5548 8352
rect 12146 14378 12202 14434
rect 12226 14378 12282 14434
rect 12306 14378 12362 14434
rect 12386 14378 12442 14434
rect 12466 14378 12522 14434
rect 12146 14298 12202 14354
rect 12226 14298 12282 14354
rect 12306 14298 12362 14354
rect 12386 14298 12442 14354
rect 12466 14298 12522 14354
rect 12146 14218 12202 14274
rect 12226 14218 12282 14274
rect 12306 14218 12362 14274
rect 12386 14218 12442 14274
rect 12466 14218 12522 14274
rect 12146 14138 12202 14194
rect 12226 14138 12282 14194
rect 12306 14138 12362 14194
rect 12386 14138 12442 14194
rect 12466 14138 12522 14194
rect 12146 14058 12202 14114
rect 12226 14058 12282 14114
rect 12306 14058 12362 14114
rect 12386 14058 12442 14114
rect 12466 14058 12522 14114
rect 8068 13578 8124 13634
rect 8148 13578 8204 13634
rect 8228 13578 8284 13634
rect 8308 13578 8364 13634
rect 8388 13578 8444 13634
rect 8068 13498 8124 13554
rect 8148 13498 8204 13554
rect 8228 13498 8284 13554
rect 8308 13498 8364 13554
rect 8388 13498 8444 13554
rect 8068 13418 8124 13474
rect 8148 13418 8204 13474
rect 8228 13418 8284 13474
rect 8308 13418 8364 13474
rect 8388 13418 8444 13474
rect 8068 13338 8124 13394
rect 8148 13338 8204 13394
rect 8228 13338 8284 13394
rect 8308 13338 8364 13394
rect 8388 13338 8444 13394
rect 8068 13258 8124 13314
rect 8148 13258 8204 13314
rect 8228 13258 8284 13314
rect 8308 13258 8364 13314
rect 8388 13258 8444 13314
rect 11346 13578 11402 13634
rect 11426 13578 11482 13634
rect 11506 13578 11562 13634
rect 11586 13578 11642 13634
rect 11666 13578 11722 13634
rect 11346 13498 11402 13554
rect 11426 13498 11482 13554
rect 11506 13498 11562 13554
rect 11586 13498 11642 13554
rect 11666 13498 11722 13554
rect 11346 13418 11402 13474
rect 11426 13418 11482 13474
rect 11506 13418 11562 13474
rect 11586 13418 11642 13474
rect 11666 13418 11722 13474
rect 11346 13338 11402 13394
rect 11426 13338 11482 13394
rect 11506 13338 11562 13394
rect 11586 13338 11642 13394
rect 11666 13338 11722 13394
rect 11346 13258 11402 13314
rect 11426 13258 11482 13314
rect 11506 13258 11562 13314
rect 11586 13258 11642 13314
rect 11666 13258 11722 13314
rect 8068 9847 8124 9903
rect 8148 9847 8204 9903
rect 8228 9847 8284 9903
rect 8308 9847 8364 9903
rect 8388 9847 8444 9903
rect 8068 9767 8124 9823
rect 8148 9767 8204 9823
rect 8228 9767 8284 9823
rect 8308 9767 8364 9823
rect 8388 9767 8444 9823
rect 8068 9687 8124 9743
rect 8148 9687 8204 9743
rect 8228 9687 8284 9743
rect 8308 9687 8364 9743
rect 8388 9687 8444 9743
rect 8068 9607 8124 9663
rect 8148 9607 8204 9663
rect 8228 9607 8284 9663
rect 8308 9607 8364 9663
rect 8388 9607 8444 9663
rect 7103 8572 7159 8628
rect 7183 8572 7239 8628
rect 7263 8572 7319 8628
rect 7343 8572 7399 8628
rect 7423 8572 7479 8628
rect 6138 7298 6194 7354
rect 6218 7298 6274 7354
rect 6298 7298 6354 7354
rect 6378 7298 6434 7354
rect 6458 7298 6514 7354
rect 6138 7218 6194 7274
rect 6218 7218 6274 7274
rect 6298 7218 6354 7274
rect 6378 7218 6434 7274
rect 6458 7218 6514 7274
rect 6138 7138 6194 7194
rect 6218 7138 6274 7194
rect 6298 7138 6354 7194
rect 6378 7138 6434 7194
rect 6458 7138 6514 7194
rect 6138 7058 6194 7114
rect 6218 7058 6274 7114
rect 6298 7058 6354 7114
rect 6378 7058 6434 7114
rect 6458 7058 6514 7114
rect 5172 6023 5228 6079
rect 5252 6023 5308 6079
rect 5332 6023 5388 6079
rect 5412 6023 5468 6079
rect 5492 6023 5548 6079
rect 5172 5943 5228 5999
rect 5252 5943 5308 5999
rect 5332 5943 5388 5999
rect 5412 5943 5468 5999
rect 5492 5943 5548 5999
rect 5172 5863 5228 5919
rect 5252 5863 5308 5919
rect 5332 5863 5388 5919
rect 5412 5863 5468 5919
rect 5492 5863 5548 5919
rect 5172 5783 5228 5839
rect 5252 5783 5308 5839
rect 5332 5783 5388 5839
rect 5412 5783 5468 5839
rect 5492 5783 5548 5839
rect 7103 8492 7159 8548
rect 7183 8492 7239 8548
rect 7263 8492 7319 8548
rect 7343 8492 7399 8548
rect 7423 8492 7479 8548
rect 7103 8412 7159 8468
rect 7183 8412 7239 8468
rect 7263 8412 7319 8468
rect 7343 8412 7399 8468
rect 7423 8412 7479 8468
rect 7103 8352 7159 8388
rect 7183 8352 7239 8388
rect 7263 8352 7319 8388
rect 7343 8352 7399 8388
rect 7423 8352 7479 8388
rect 7103 8332 7105 8352
rect 7105 8332 7157 8352
rect 7157 8332 7159 8352
rect 7183 8332 7221 8352
rect 7221 8332 7233 8352
rect 7233 8332 7239 8352
rect 7263 8332 7285 8352
rect 7285 8332 7297 8352
rect 7297 8332 7319 8352
rect 7343 8332 7349 8352
rect 7349 8332 7361 8352
rect 7361 8332 7399 8352
rect 7423 8332 7425 8352
rect 7425 8332 7477 8352
rect 7477 8332 7479 8352
rect 5172 362 5228 418
rect 5252 362 5308 418
rect 5332 362 5388 418
rect 5412 362 5468 418
rect 5492 362 5548 418
rect 5172 282 5228 338
rect 5252 282 5308 338
rect 5332 282 5388 338
rect 5412 282 5468 338
rect 5492 282 5548 338
rect 5172 202 5228 258
rect 5252 202 5308 258
rect 5332 202 5388 258
rect 5412 202 5468 258
rect 5492 202 5548 258
rect 5172 122 5228 178
rect 5252 122 5308 178
rect 5332 122 5388 178
rect 5412 122 5468 178
rect 5492 122 5548 178
rect 5172 42 5228 98
rect 5252 42 5308 98
rect 5332 42 5388 98
rect 5412 42 5468 98
rect 5492 42 5548 98
rect 7103 6023 7159 6079
rect 7183 6023 7239 6079
rect 7263 6023 7319 6079
rect 7343 6023 7399 6079
rect 7423 6023 7479 6079
rect 7103 5943 7159 5999
rect 7183 5943 7239 5999
rect 7263 5943 7319 5999
rect 7343 5943 7399 5999
rect 7423 5943 7479 5999
rect 7103 5863 7159 5919
rect 7183 5863 7239 5919
rect 7263 5863 7319 5919
rect 7343 5863 7399 5919
rect 7423 5863 7479 5919
rect 7103 5783 7159 5839
rect 7183 5783 7239 5839
rect 7263 5783 7319 5839
rect 7343 5783 7399 5839
rect 7423 5783 7479 5839
rect 6138 4748 6194 4804
rect 6218 4748 6274 4804
rect 6298 4748 6354 4804
rect 6378 4748 6434 4804
rect 6458 4748 6514 4804
rect 6138 4668 6194 4724
rect 6218 4668 6274 4724
rect 6298 4668 6354 4724
rect 6378 4668 6434 4724
rect 6458 4668 6514 4724
rect 6138 4588 6194 4644
rect 6218 4588 6274 4644
rect 6298 4588 6354 4644
rect 6378 4588 6434 4644
rect 6458 4588 6514 4644
rect 6138 4544 6194 4564
rect 6218 4544 6274 4564
rect 6298 4544 6354 4564
rect 6378 4544 6434 4564
rect 6458 4544 6514 4564
rect 6138 4508 6140 4544
rect 6140 4508 6192 4544
rect 6192 4508 6194 4544
rect 6218 4508 6256 4544
rect 6256 4508 6268 4544
rect 6268 4508 6274 4544
rect 6298 4508 6320 4544
rect 6320 4508 6332 4544
rect 6332 4508 6354 4544
rect 6378 4508 6384 4544
rect 6384 4508 6396 4544
rect 6396 4508 6434 4544
rect 6458 4508 6460 4544
rect 6460 4508 6512 4544
rect 6512 4508 6514 4544
rect 6138 1162 6194 1218
rect 6218 1162 6274 1218
rect 6298 1162 6354 1218
rect 6378 1162 6434 1218
rect 6458 1162 6514 1218
rect 6138 1082 6194 1138
rect 6218 1082 6274 1138
rect 6298 1082 6354 1138
rect 6378 1082 6434 1138
rect 6458 1082 6514 1138
rect 6138 1002 6194 1058
rect 6218 1002 6274 1058
rect 6298 1002 6354 1058
rect 6378 1002 6434 1058
rect 6458 1002 6514 1058
rect 6138 922 6194 978
rect 6218 922 6274 978
rect 6298 922 6354 978
rect 6378 922 6434 978
rect 6458 922 6514 978
rect 6138 842 6194 898
rect 6218 842 6274 898
rect 6298 842 6354 898
rect 6378 842 6434 898
rect 6458 842 6514 898
rect 8068 7298 8124 7354
rect 8148 7298 8204 7354
rect 8228 7298 8284 7354
rect 8308 7298 8364 7354
rect 8388 7298 8444 7354
rect 11346 9847 11402 9903
rect 11426 9847 11482 9903
rect 11506 9847 11562 9903
rect 11586 9847 11642 9903
rect 11666 9847 11722 9903
rect 11346 9767 11402 9823
rect 11426 9767 11482 9823
rect 11506 9767 11562 9823
rect 11586 9767 11642 9823
rect 11666 9767 11722 9823
rect 11346 9687 11402 9743
rect 11426 9687 11482 9743
rect 11506 9687 11562 9743
rect 11586 9687 11642 9743
rect 11666 9687 11722 9743
rect 11346 9607 11402 9663
rect 11426 9607 11482 9663
rect 11506 9607 11562 9663
rect 11586 9607 11642 9663
rect 11666 9607 11722 9663
rect 8068 7218 8124 7274
rect 8148 7218 8204 7274
rect 8228 7218 8284 7274
rect 8308 7218 8364 7274
rect 8388 7218 8444 7274
rect 8068 7138 8124 7194
rect 8148 7138 8204 7194
rect 8228 7138 8284 7194
rect 8308 7138 8364 7194
rect 8388 7138 8444 7194
rect 8068 7058 8124 7114
rect 8148 7058 8204 7114
rect 8228 7058 8284 7114
rect 8308 7058 8364 7114
rect 8388 7058 8444 7114
rect 11346 7298 11402 7354
rect 11426 7298 11482 7354
rect 11506 7298 11562 7354
rect 11586 7298 11642 7354
rect 11666 7298 11722 7354
rect 11346 7218 11402 7274
rect 11426 7218 11482 7274
rect 11506 7218 11562 7274
rect 11586 7218 11642 7274
rect 11666 7218 11722 7274
rect 11346 7138 11402 7194
rect 11426 7138 11482 7194
rect 11506 7138 11562 7194
rect 11586 7138 11642 7194
rect 11666 7138 11722 7194
rect 11346 7058 11402 7114
rect 11426 7058 11482 7114
rect 11506 7058 11562 7114
rect 11586 7058 11642 7114
rect 11666 7058 11722 7114
rect 8068 4748 8124 4804
rect 8148 4748 8204 4804
rect 8228 4748 8284 4804
rect 8308 4748 8364 4804
rect 8388 4748 8444 4804
rect 8068 4668 8124 4724
rect 8148 4668 8204 4724
rect 8228 4668 8284 4724
rect 8308 4668 8364 4724
rect 8388 4668 8444 4724
rect 8068 4588 8124 4644
rect 8148 4588 8204 4644
rect 8228 4588 8284 4644
rect 8308 4588 8364 4644
rect 8388 4588 8444 4644
rect 8068 4544 8124 4564
rect 8148 4544 8204 4564
rect 8228 4544 8284 4564
rect 8308 4544 8364 4564
rect 8388 4544 8444 4564
rect 8068 4508 8070 4544
rect 8070 4508 8122 4544
rect 8122 4508 8124 4544
rect 8148 4508 8186 4544
rect 8186 4508 8198 4544
rect 8198 4508 8204 4544
rect 8228 4508 8250 4544
rect 8250 4508 8262 4544
rect 8262 4508 8284 4544
rect 8308 4508 8314 4544
rect 8314 4508 8326 4544
rect 8326 4508 8364 4544
rect 8388 4508 8390 4544
rect 8390 4508 8442 4544
rect 8442 4508 8444 4544
rect 7103 362 7159 418
rect 7183 362 7239 418
rect 7263 362 7319 418
rect 7343 362 7399 418
rect 7423 362 7479 418
rect 7103 282 7159 338
rect 7183 282 7239 338
rect 7263 282 7319 338
rect 7343 282 7399 338
rect 7423 282 7479 338
rect 7103 202 7159 258
rect 7183 202 7239 258
rect 7263 202 7319 258
rect 7343 202 7399 258
rect 7423 202 7479 258
rect 7103 122 7159 178
rect 7183 122 7239 178
rect 7263 122 7319 178
rect 7343 122 7399 178
rect 7423 122 7479 178
rect 7103 42 7159 98
rect 7183 42 7239 98
rect 7263 42 7319 98
rect 7343 42 7399 98
rect 7423 42 7479 98
rect 11346 4748 11402 4804
rect 11426 4748 11482 4804
rect 11506 4748 11562 4804
rect 11586 4748 11642 4804
rect 11666 4748 11722 4804
rect 11346 4668 11402 4724
rect 11426 4668 11482 4724
rect 11506 4668 11562 4724
rect 11586 4668 11642 4724
rect 11666 4668 11722 4724
rect 11346 4588 11402 4644
rect 11426 4588 11482 4644
rect 11506 4588 11562 4644
rect 11586 4588 11642 4644
rect 11666 4588 11722 4644
rect 11346 4508 11402 4564
rect 11426 4508 11482 4564
rect 11506 4508 11562 4564
rect 11586 4508 11642 4564
rect 11666 4508 11722 4564
rect 8068 1162 8124 1218
rect 8148 1162 8204 1218
rect 8228 1162 8284 1218
rect 8308 1162 8364 1218
rect 8388 1162 8444 1218
rect 8068 1082 8124 1138
rect 8148 1082 8204 1138
rect 8228 1082 8284 1138
rect 8308 1082 8364 1138
rect 8388 1082 8444 1138
rect 8068 1002 8124 1058
rect 8148 1002 8204 1058
rect 8228 1002 8284 1058
rect 8308 1002 8364 1058
rect 8388 1002 8444 1058
rect 8068 922 8124 978
rect 8148 922 8204 978
rect 8228 922 8284 978
rect 8308 922 8364 978
rect 8388 922 8444 978
rect 8068 842 8124 898
rect 8148 842 8204 898
rect 8228 842 8284 898
rect 8308 842 8364 898
rect 8388 842 8444 898
rect 11346 1162 11402 1218
rect 11426 1162 11482 1218
rect 11506 1162 11562 1218
rect 11586 1162 11642 1218
rect 11666 1162 11722 1218
rect 11346 1082 11402 1138
rect 11426 1082 11482 1138
rect 11506 1082 11562 1138
rect 11586 1082 11642 1138
rect 11666 1082 11722 1138
rect 11346 1002 11402 1058
rect 11426 1002 11482 1058
rect 11506 1002 11562 1058
rect 11586 1002 11642 1058
rect 11666 1002 11722 1058
rect 11346 922 11402 978
rect 11426 922 11482 978
rect 11506 922 11562 978
rect 11586 922 11642 978
rect 11666 922 11722 978
rect 11346 842 11402 898
rect 11426 842 11482 898
rect 11506 842 11562 898
rect 11586 842 11642 898
rect 11666 842 11722 898
rect 12146 8572 12202 8628
rect 12226 8572 12282 8628
rect 12306 8572 12362 8628
rect 12386 8572 12442 8628
rect 12466 8572 12522 8628
rect 12146 8492 12202 8548
rect 12226 8492 12282 8548
rect 12306 8492 12362 8548
rect 12386 8492 12442 8548
rect 12466 8492 12522 8548
rect 12146 8412 12202 8468
rect 12226 8412 12282 8468
rect 12306 8412 12362 8468
rect 12386 8412 12442 8468
rect 12466 8412 12522 8468
rect 12146 8332 12202 8388
rect 12226 8332 12282 8388
rect 12306 8332 12362 8388
rect 12386 8332 12442 8388
rect 12466 8332 12522 8388
rect 12146 6023 12202 6079
rect 12226 6023 12282 6079
rect 12306 6023 12362 6079
rect 12386 6023 12442 6079
rect 12466 6023 12522 6079
rect 12146 5943 12202 5999
rect 12226 5943 12282 5999
rect 12306 5943 12362 5999
rect 12386 5943 12442 5999
rect 12466 5943 12522 5999
rect 12146 5863 12202 5919
rect 12226 5863 12282 5919
rect 12306 5863 12362 5919
rect 12386 5863 12442 5919
rect 12466 5863 12522 5919
rect 12146 5783 12202 5839
rect 12226 5783 12282 5839
rect 12306 5783 12362 5839
rect 12386 5783 12442 5839
rect 12466 5783 12522 5839
rect 12146 362 12202 418
rect 12226 362 12282 418
rect 12306 362 12362 418
rect 12386 362 12442 418
rect 12466 362 12522 418
rect 12146 282 12202 338
rect 12226 282 12282 338
rect 12306 282 12362 338
rect 12386 282 12442 338
rect 12466 282 12522 338
rect 12146 202 12202 258
rect 12226 202 12282 258
rect 12306 202 12362 258
rect 12386 202 12442 258
rect 12466 202 12522 258
rect 12146 122 12202 178
rect 12226 122 12282 178
rect 12306 122 12362 178
rect 12386 122 12442 178
rect 12466 122 12522 178
rect 12146 42 12202 98
rect 12226 42 12282 98
rect 12306 42 12362 98
rect 12386 42 12442 98
rect 12466 42 12522 98
<< metal3 >>
rect 0 14434 12564 14476
rect 0 14378 42 14434
rect 98 14378 122 14434
rect 178 14378 202 14434
rect 258 14378 282 14434
rect 338 14378 362 14434
rect 418 14378 5172 14434
rect 5228 14378 5252 14434
rect 5308 14378 5332 14434
rect 5388 14378 5412 14434
rect 5468 14378 5492 14434
rect 5548 14378 7103 14434
rect 7159 14378 7183 14434
rect 7239 14378 7263 14434
rect 7319 14378 7343 14434
rect 7399 14378 7423 14434
rect 7479 14378 12146 14434
rect 12202 14378 12226 14434
rect 12282 14378 12306 14434
rect 12362 14378 12386 14434
rect 12442 14378 12466 14434
rect 12522 14378 12564 14434
rect 0 14354 12564 14378
rect 0 14298 42 14354
rect 98 14298 122 14354
rect 178 14298 202 14354
rect 258 14298 282 14354
rect 338 14298 362 14354
rect 418 14298 5172 14354
rect 5228 14298 5252 14354
rect 5308 14298 5332 14354
rect 5388 14298 5412 14354
rect 5468 14298 5492 14354
rect 5548 14298 7103 14354
rect 7159 14298 7183 14354
rect 7239 14298 7263 14354
rect 7319 14298 7343 14354
rect 7399 14298 7423 14354
rect 7479 14298 12146 14354
rect 12202 14298 12226 14354
rect 12282 14298 12306 14354
rect 12362 14298 12386 14354
rect 12442 14298 12466 14354
rect 12522 14298 12564 14354
rect 0 14274 12564 14298
rect 0 14218 42 14274
rect 98 14218 122 14274
rect 178 14218 202 14274
rect 258 14218 282 14274
rect 338 14218 362 14274
rect 418 14218 5172 14274
rect 5228 14218 5252 14274
rect 5308 14218 5332 14274
rect 5388 14218 5412 14274
rect 5468 14218 5492 14274
rect 5548 14218 7103 14274
rect 7159 14218 7183 14274
rect 7239 14218 7263 14274
rect 7319 14218 7343 14274
rect 7399 14218 7423 14274
rect 7479 14218 12146 14274
rect 12202 14218 12226 14274
rect 12282 14218 12306 14274
rect 12362 14218 12386 14274
rect 12442 14218 12466 14274
rect 12522 14218 12564 14274
rect 0 14194 12564 14218
rect 0 14138 42 14194
rect 98 14138 122 14194
rect 178 14138 202 14194
rect 258 14138 282 14194
rect 338 14138 362 14194
rect 418 14138 5172 14194
rect 5228 14138 5252 14194
rect 5308 14138 5332 14194
rect 5388 14138 5412 14194
rect 5468 14138 5492 14194
rect 5548 14138 7103 14194
rect 7159 14138 7183 14194
rect 7239 14138 7263 14194
rect 7319 14138 7343 14194
rect 7399 14138 7423 14194
rect 7479 14138 12146 14194
rect 12202 14138 12226 14194
rect 12282 14138 12306 14194
rect 12362 14138 12386 14194
rect 12442 14138 12466 14194
rect 12522 14138 12564 14194
rect 0 14114 12564 14138
rect 0 14058 42 14114
rect 98 14058 122 14114
rect 178 14058 202 14114
rect 258 14058 282 14114
rect 338 14058 362 14114
rect 418 14058 5172 14114
rect 5228 14058 5252 14114
rect 5308 14058 5332 14114
rect 5388 14058 5412 14114
rect 5468 14058 5492 14114
rect 5548 14058 7103 14114
rect 7159 14058 7183 14114
rect 7239 14058 7263 14114
rect 7319 14058 7343 14114
rect 7399 14058 7423 14114
rect 7479 14058 12146 14114
rect 12202 14058 12226 14114
rect 12282 14058 12306 14114
rect 12362 14058 12386 14114
rect 12442 14058 12466 14114
rect 12522 14058 12564 14114
rect 0 14016 12564 14058
rect 800 13634 11764 13676
rect 800 13578 842 13634
rect 898 13578 922 13634
rect 978 13578 1002 13634
rect 1058 13578 1082 13634
rect 1138 13578 1162 13634
rect 1218 13578 4207 13634
rect 4263 13578 4287 13634
rect 4343 13578 4367 13634
rect 4423 13578 4447 13634
rect 4503 13578 4527 13634
rect 4583 13578 6138 13634
rect 6194 13578 6218 13634
rect 6274 13578 6298 13634
rect 6354 13578 6378 13634
rect 6434 13578 6458 13634
rect 6514 13578 8068 13634
rect 8124 13578 8148 13634
rect 8204 13578 8228 13634
rect 8284 13578 8308 13634
rect 8364 13578 8388 13634
rect 8444 13578 11346 13634
rect 11402 13578 11426 13634
rect 11482 13578 11506 13634
rect 11562 13578 11586 13634
rect 11642 13578 11666 13634
rect 11722 13578 11764 13634
rect 800 13554 11764 13578
rect 800 13498 842 13554
rect 898 13498 922 13554
rect 978 13498 1002 13554
rect 1058 13498 1082 13554
rect 1138 13498 1162 13554
rect 1218 13498 4207 13554
rect 4263 13498 4287 13554
rect 4343 13498 4367 13554
rect 4423 13498 4447 13554
rect 4503 13498 4527 13554
rect 4583 13498 6138 13554
rect 6194 13498 6218 13554
rect 6274 13498 6298 13554
rect 6354 13498 6378 13554
rect 6434 13498 6458 13554
rect 6514 13498 8068 13554
rect 8124 13498 8148 13554
rect 8204 13498 8228 13554
rect 8284 13498 8308 13554
rect 8364 13498 8388 13554
rect 8444 13498 11346 13554
rect 11402 13498 11426 13554
rect 11482 13498 11506 13554
rect 11562 13498 11586 13554
rect 11642 13498 11666 13554
rect 11722 13498 11764 13554
rect 800 13474 11764 13498
rect 800 13418 842 13474
rect 898 13418 922 13474
rect 978 13418 1002 13474
rect 1058 13418 1082 13474
rect 1138 13418 1162 13474
rect 1218 13418 4207 13474
rect 4263 13418 4287 13474
rect 4343 13418 4367 13474
rect 4423 13418 4447 13474
rect 4503 13418 4527 13474
rect 4583 13418 6138 13474
rect 6194 13418 6218 13474
rect 6274 13418 6298 13474
rect 6354 13418 6378 13474
rect 6434 13418 6458 13474
rect 6514 13418 8068 13474
rect 8124 13418 8148 13474
rect 8204 13418 8228 13474
rect 8284 13418 8308 13474
rect 8364 13418 8388 13474
rect 8444 13418 11346 13474
rect 11402 13418 11426 13474
rect 11482 13418 11506 13474
rect 11562 13418 11586 13474
rect 11642 13418 11666 13474
rect 11722 13418 11764 13474
rect 800 13394 11764 13418
rect 800 13338 842 13394
rect 898 13338 922 13394
rect 978 13338 1002 13394
rect 1058 13338 1082 13394
rect 1138 13338 1162 13394
rect 1218 13338 4207 13394
rect 4263 13338 4287 13394
rect 4343 13338 4367 13394
rect 4423 13338 4447 13394
rect 4503 13338 4527 13394
rect 4583 13338 6138 13394
rect 6194 13338 6218 13394
rect 6274 13338 6298 13394
rect 6354 13338 6378 13394
rect 6434 13338 6458 13394
rect 6514 13338 8068 13394
rect 8124 13338 8148 13394
rect 8204 13338 8228 13394
rect 8284 13338 8308 13394
rect 8364 13338 8388 13394
rect 8444 13338 11346 13394
rect 11402 13338 11426 13394
rect 11482 13338 11506 13394
rect 11562 13338 11586 13394
rect 11642 13338 11666 13394
rect 11722 13338 11764 13394
rect 800 13314 11764 13338
rect 800 13258 842 13314
rect 898 13258 922 13314
rect 978 13258 1002 13314
rect 1058 13258 1082 13314
rect 1138 13258 1162 13314
rect 1218 13258 4207 13314
rect 4263 13258 4287 13314
rect 4343 13258 4367 13314
rect 4423 13258 4447 13314
rect 4503 13258 4527 13314
rect 4583 13258 6138 13314
rect 6194 13258 6218 13314
rect 6274 13258 6298 13314
rect 6354 13258 6378 13314
rect 6434 13258 6458 13314
rect 6514 13258 8068 13314
rect 8124 13258 8148 13314
rect 8204 13258 8228 13314
rect 8284 13258 8308 13314
rect 8364 13258 8388 13314
rect 8444 13258 11346 13314
rect 11402 13258 11426 13314
rect 11482 13258 11506 13314
rect 11562 13258 11586 13314
rect 11642 13258 11666 13314
rect 11722 13258 11764 13314
rect 800 13216 11764 13258
rect 0 9903 12564 9935
rect 0 9847 842 9903
rect 898 9847 922 9903
rect 978 9847 1002 9903
rect 1058 9847 1082 9903
rect 1138 9847 1162 9903
rect 1218 9847 4207 9903
rect 4263 9847 4287 9903
rect 4343 9847 4367 9903
rect 4423 9847 4447 9903
rect 4503 9847 4527 9903
rect 4583 9847 6138 9903
rect 6194 9847 6218 9903
rect 6274 9847 6298 9903
rect 6354 9847 6378 9903
rect 6434 9847 6458 9903
rect 6514 9847 8068 9903
rect 8124 9847 8148 9903
rect 8204 9847 8228 9903
rect 8284 9847 8308 9903
rect 8364 9847 8388 9903
rect 8444 9847 11346 9903
rect 11402 9847 11426 9903
rect 11482 9847 11506 9903
rect 11562 9847 11586 9903
rect 11642 9847 11666 9903
rect 11722 9847 12564 9903
rect 0 9823 12564 9847
rect 0 9767 842 9823
rect 898 9767 922 9823
rect 978 9767 1002 9823
rect 1058 9767 1082 9823
rect 1138 9767 1162 9823
rect 1218 9767 4207 9823
rect 4263 9767 4287 9823
rect 4343 9767 4367 9823
rect 4423 9767 4447 9823
rect 4503 9767 4527 9823
rect 4583 9767 6138 9823
rect 6194 9767 6218 9823
rect 6274 9767 6298 9823
rect 6354 9767 6378 9823
rect 6434 9767 6458 9823
rect 6514 9767 8068 9823
rect 8124 9767 8148 9823
rect 8204 9767 8228 9823
rect 8284 9767 8308 9823
rect 8364 9767 8388 9823
rect 8444 9767 11346 9823
rect 11402 9767 11426 9823
rect 11482 9767 11506 9823
rect 11562 9767 11586 9823
rect 11642 9767 11666 9823
rect 11722 9767 12564 9823
rect 0 9743 12564 9767
rect 0 9687 842 9743
rect 898 9687 922 9743
rect 978 9687 1002 9743
rect 1058 9687 1082 9743
rect 1138 9687 1162 9743
rect 1218 9687 4207 9743
rect 4263 9687 4287 9743
rect 4343 9687 4367 9743
rect 4423 9687 4447 9743
rect 4503 9687 4527 9743
rect 4583 9687 6138 9743
rect 6194 9687 6218 9743
rect 6274 9687 6298 9743
rect 6354 9687 6378 9743
rect 6434 9687 6458 9743
rect 6514 9687 8068 9743
rect 8124 9687 8148 9743
rect 8204 9687 8228 9743
rect 8284 9687 8308 9743
rect 8364 9687 8388 9743
rect 8444 9687 11346 9743
rect 11402 9687 11426 9743
rect 11482 9687 11506 9743
rect 11562 9687 11586 9743
rect 11642 9687 11666 9743
rect 11722 9687 12564 9743
rect 0 9663 12564 9687
rect 0 9607 842 9663
rect 898 9607 922 9663
rect 978 9607 1002 9663
rect 1058 9607 1082 9663
rect 1138 9607 1162 9663
rect 1218 9607 4207 9663
rect 4263 9607 4287 9663
rect 4343 9607 4367 9663
rect 4423 9607 4447 9663
rect 4503 9607 4527 9663
rect 4583 9607 6138 9663
rect 6194 9607 6218 9663
rect 6274 9607 6298 9663
rect 6354 9607 6378 9663
rect 6434 9607 6458 9663
rect 6514 9607 8068 9663
rect 8124 9607 8148 9663
rect 8204 9607 8228 9663
rect 8284 9607 8308 9663
rect 8364 9607 8388 9663
rect 8444 9607 11346 9663
rect 11402 9607 11426 9663
rect 11482 9607 11506 9663
rect 11562 9607 11586 9663
rect 11642 9607 11666 9663
rect 11722 9607 12564 9663
rect 0 9575 12564 9607
rect 0 8628 12564 8661
rect 0 8572 42 8628
rect 98 8572 122 8628
rect 178 8572 202 8628
rect 258 8572 282 8628
rect 338 8572 362 8628
rect 418 8572 5172 8628
rect 5228 8572 5252 8628
rect 5308 8572 5332 8628
rect 5388 8572 5412 8628
rect 5468 8572 5492 8628
rect 5548 8572 7103 8628
rect 7159 8572 7183 8628
rect 7239 8572 7263 8628
rect 7319 8572 7343 8628
rect 7399 8572 7423 8628
rect 7479 8572 12146 8628
rect 12202 8572 12226 8628
rect 12282 8572 12306 8628
rect 12362 8572 12386 8628
rect 12442 8572 12466 8628
rect 12522 8572 12564 8628
rect 0 8548 12564 8572
rect 0 8492 42 8548
rect 98 8492 122 8548
rect 178 8492 202 8548
rect 258 8492 282 8548
rect 338 8492 362 8548
rect 418 8492 5172 8548
rect 5228 8492 5252 8548
rect 5308 8492 5332 8548
rect 5388 8492 5412 8548
rect 5468 8492 5492 8548
rect 5548 8492 7103 8548
rect 7159 8492 7183 8548
rect 7239 8492 7263 8548
rect 7319 8492 7343 8548
rect 7399 8492 7423 8548
rect 7479 8492 12146 8548
rect 12202 8492 12226 8548
rect 12282 8492 12306 8548
rect 12362 8492 12386 8548
rect 12442 8492 12466 8548
rect 12522 8492 12564 8548
rect 0 8468 12564 8492
rect 0 8412 42 8468
rect 98 8412 122 8468
rect 178 8412 202 8468
rect 258 8412 282 8468
rect 338 8412 362 8468
rect 418 8412 5172 8468
rect 5228 8412 5252 8468
rect 5308 8412 5332 8468
rect 5388 8412 5412 8468
rect 5468 8412 5492 8468
rect 5548 8412 7103 8468
rect 7159 8412 7183 8468
rect 7239 8412 7263 8468
rect 7319 8412 7343 8468
rect 7399 8412 7423 8468
rect 7479 8412 12146 8468
rect 12202 8412 12226 8468
rect 12282 8412 12306 8468
rect 12362 8412 12386 8468
rect 12442 8412 12466 8468
rect 12522 8412 12564 8468
rect 0 8388 12564 8412
rect 0 8332 42 8388
rect 98 8332 122 8388
rect 178 8332 202 8388
rect 258 8332 282 8388
rect 338 8332 362 8388
rect 418 8332 5172 8388
rect 5228 8332 5252 8388
rect 5308 8332 5332 8388
rect 5388 8332 5412 8388
rect 5468 8332 5492 8388
rect 5548 8332 7103 8388
rect 7159 8332 7183 8388
rect 7239 8332 7263 8388
rect 7319 8332 7343 8388
rect 7399 8332 7423 8388
rect 7479 8332 12146 8388
rect 12202 8332 12226 8388
rect 12282 8332 12306 8388
rect 12362 8332 12386 8388
rect 12442 8332 12466 8388
rect 12522 8332 12564 8388
rect 0 8300 12564 8332
rect 0 7354 12564 7386
rect 0 7298 842 7354
rect 898 7298 922 7354
rect 978 7298 1002 7354
rect 1058 7298 1082 7354
rect 1138 7298 1162 7354
rect 1218 7298 4207 7354
rect 4263 7298 4287 7354
rect 4343 7298 4367 7354
rect 4423 7298 4447 7354
rect 4503 7298 4527 7354
rect 4583 7298 6138 7354
rect 6194 7298 6218 7354
rect 6274 7298 6298 7354
rect 6354 7298 6378 7354
rect 6434 7298 6458 7354
rect 6514 7298 8068 7354
rect 8124 7298 8148 7354
rect 8204 7298 8228 7354
rect 8284 7298 8308 7354
rect 8364 7298 8388 7354
rect 8444 7298 11346 7354
rect 11402 7298 11426 7354
rect 11482 7298 11506 7354
rect 11562 7298 11586 7354
rect 11642 7298 11666 7354
rect 11722 7298 12564 7354
rect 0 7274 12564 7298
rect 0 7218 842 7274
rect 898 7218 922 7274
rect 978 7218 1002 7274
rect 1058 7218 1082 7274
rect 1138 7218 1162 7274
rect 1218 7218 4207 7274
rect 4263 7218 4287 7274
rect 4343 7218 4367 7274
rect 4423 7218 4447 7274
rect 4503 7218 4527 7274
rect 4583 7218 6138 7274
rect 6194 7218 6218 7274
rect 6274 7218 6298 7274
rect 6354 7218 6378 7274
rect 6434 7218 6458 7274
rect 6514 7218 8068 7274
rect 8124 7218 8148 7274
rect 8204 7218 8228 7274
rect 8284 7218 8308 7274
rect 8364 7218 8388 7274
rect 8444 7218 11346 7274
rect 11402 7218 11426 7274
rect 11482 7218 11506 7274
rect 11562 7218 11586 7274
rect 11642 7218 11666 7274
rect 11722 7218 12564 7274
rect 0 7194 12564 7218
rect 0 7138 842 7194
rect 898 7138 922 7194
rect 978 7138 1002 7194
rect 1058 7138 1082 7194
rect 1138 7138 1162 7194
rect 1218 7138 4207 7194
rect 4263 7138 4287 7194
rect 4343 7138 4367 7194
rect 4423 7138 4447 7194
rect 4503 7138 4527 7194
rect 4583 7138 6138 7194
rect 6194 7138 6218 7194
rect 6274 7138 6298 7194
rect 6354 7138 6378 7194
rect 6434 7138 6458 7194
rect 6514 7138 8068 7194
rect 8124 7138 8148 7194
rect 8204 7138 8228 7194
rect 8284 7138 8308 7194
rect 8364 7138 8388 7194
rect 8444 7138 11346 7194
rect 11402 7138 11426 7194
rect 11482 7138 11506 7194
rect 11562 7138 11586 7194
rect 11642 7138 11666 7194
rect 11722 7138 12564 7194
rect 0 7114 12564 7138
rect 0 7058 842 7114
rect 898 7058 922 7114
rect 978 7058 1002 7114
rect 1058 7058 1082 7114
rect 1138 7058 1162 7114
rect 1218 7058 4207 7114
rect 4263 7058 4287 7114
rect 4343 7058 4367 7114
rect 4423 7058 4447 7114
rect 4503 7058 4527 7114
rect 4583 7058 6138 7114
rect 6194 7058 6218 7114
rect 6274 7058 6298 7114
rect 6354 7058 6378 7114
rect 6434 7058 6458 7114
rect 6514 7058 8068 7114
rect 8124 7058 8148 7114
rect 8204 7058 8228 7114
rect 8284 7058 8308 7114
rect 8364 7058 8388 7114
rect 8444 7058 11346 7114
rect 11402 7058 11426 7114
rect 11482 7058 11506 7114
rect 11562 7058 11586 7114
rect 11642 7058 11666 7114
rect 11722 7058 12564 7114
rect 0 7026 12564 7058
rect 0 6079 12564 6111
rect 0 6023 42 6079
rect 98 6023 122 6079
rect 178 6023 202 6079
rect 258 6023 282 6079
rect 338 6023 362 6079
rect 418 6023 5172 6079
rect 5228 6023 5252 6079
rect 5308 6023 5332 6079
rect 5388 6023 5412 6079
rect 5468 6023 5492 6079
rect 5548 6023 7103 6079
rect 7159 6023 7183 6079
rect 7239 6023 7263 6079
rect 7319 6023 7343 6079
rect 7399 6023 7423 6079
rect 7479 6023 12146 6079
rect 12202 6023 12226 6079
rect 12282 6023 12306 6079
rect 12362 6023 12386 6079
rect 12442 6023 12466 6079
rect 12522 6023 12564 6079
rect 0 5999 12564 6023
rect 0 5943 42 5999
rect 98 5943 122 5999
rect 178 5943 202 5999
rect 258 5943 282 5999
rect 338 5943 362 5999
rect 418 5943 5172 5999
rect 5228 5943 5252 5999
rect 5308 5943 5332 5999
rect 5388 5943 5412 5999
rect 5468 5943 5492 5999
rect 5548 5943 7103 5999
rect 7159 5943 7183 5999
rect 7239 5943 7263 5999
rect 7319 5943 7343 5999
rect 7399 5943 7423 5999
rect 7479 5943 12146 5999
rect 12202 5943 12226 5999
rect 12282 5943 12306 5999
rect 12362 5943 12386 5999
rect 12442 5943 12466 5999
rect 12522 5943 12564 5999
rect 0 5919 12564 5943
rect 0 5863 42 5919
rect 98 5863 122 5919
rect 178 5863 202 5919
rect 258 5863 282 5919
rect 338 5863 362 5919
rect 418 5863 5172 5919
rect 5228 5863 5252 5919
rect 5308 5863 5332 5919
rect 5388 5863 5412 5919
rect 5468 5863 5492 5919
rect 5548 5863 7103 5919
rect 7159 5863 7183 5919
rect 7239 5863 7263 5919
rect 7319 5863 7343 5919
rect 7399 5863 7423 5919
rect 7479 5863 12146 5919
rect 12202 5863 12226 5919
rect 12282 5863 12306 5919
rect 12362 5863 12386 5919
rect 12442 5863 12466 5919
rect 12522 5863 12564 5919
rect 0 5839 12564 5863
rect 0 5783 42 5839
rect 98 5783 122 5839
rect 178 5783 202 5839
rect 258 5783 282 5839
rect 338 5783 362 5839
rect 418 5783 5172 5839
rect 5228 5783 5252 5839
rect 5308 5783 5332 5839
rect 5388 5783 5412 5839
rect 5468 5783 5492 5839
rect 5548 5783 7103 5839
rect 7159 5783 7183 5839
rect 7239 5783 7263 5839
rect 7319 5783 7343 5839
rect 7399 5783 7423 5839
rect 7479 5783 12146 5839
rect 12202 5783 12226 5839
rect 12282 5783 12306 5839
rect 12362 5783 12386 5839
rect 12442 5783 12466 5839
rect 12522 5783 12564 5839
rect 0 5751 12564 5783
rect 0 4804 12564 4837
rect 0 4748 842 4804
rect 898 4748 922 4804
rect 978 4748 1002 4804
rect 1058 4748 1082 4804
rect 1138 4748 1162 4804
rect 1218 4748 4207 4804
rect 4263 4748 4287 4804
rect 4343 4748 4367 4804
rect 4423 4748 4447 4804
rect 4503 4748 4527 4804
rect 4583 4748 6138 4804
rect 6194 4748 6218 4804
rect 6274 4748 6298 4804
rect 6354 4748 6378 4804
rect 6434 4748 6458 4804
rect 6514 4748 8068 4804
rect 8124 4748 8148 4804
rect 8204 4748 8228 4804
rect 8284 4748 8308 4804
rect 8364 4748 8388 4804
rect 8444 4748 11346 4804
rect 11402 4748 11426 4804
rect 11482 4748 11506 4804
rect 11562 4748 11586 4804
rect 11642 4748 11666 4804
rect 11722 4748 12564 4804
rect 0 4724 12564 4748
rect 0 4668 842 4724
rect 898 4668 922 4724
rect 978 4668 1002 4724
rect 1058 4668 1082 4724
rect 1138 4668 1162 4724
rect 1218 4668 4207 4724
rect 4263 4668 4287 4724
rect 4343 4668 4367 4724
rect 4423 4668 4447 4724
rect 4503 4668 4527 4724
rect 4583 4668 6138 4724
rect 6194 4668 6218 4724
rect 6274 4668 6298 4724
rect 6354 4668 6378 4724
rect 6434 4668 6458 4724
rect 6514 4668 8068 4724
rect 8124 4668 8148 4724
rect 8204 4668 8228 4724
rect 8284 4668 8308 4724
rect 8364 4668 8388 4724
rect 8444 4668 11346 4724
rect 11402 4668 11426 4724
rect 11482 4668 11506 4724
rect 11562 4668 11586 4724
rect 11642 4668 11666 4724
rect 11722 4668 12564 4724
rect 0 4644 12564 4668
rect 0 4588 842 4644
rect 898 4588 922 4644
rect 978 4588 1002 4644
rect 1058 4588 1082 4644
rect 1138 4588 1162 4644
rect 1218 4588 4207 4644
rect 4263 4588 4287 4644
rect 4343 4588 4367 4644
rect 4423 4588 4447 4644
rect 4503 4588 4527 4644
rect 4583 4588 6138 4644
rect 6194 4588 6218 4644
rect 6274 4588 6298 4644
rect 6354 4588 6378 4644
rect 6434 4588 6458 4644
rect 6514 4588 8068 4644
rect 8124 4588 8148 4644
rect 8204 4588 8228 4644
rect 8284 4588 8308 4644
rect 8364 4588 8388 4644
rect 8444 4588 11346 4644
rect 11402 4588 11426 4644
rect 11482 4588 11506 4644
rect 11562 4588 11586 4644
rect 11642 4588 11666 4644
rect 11722 4588 12564 4644
rect 0 4564 12564 4588
rect 0 4508 842 4564
rect 898 4508 922 4564
rect 978 4508 1002 4564
rect 1058 4508 1082 4564
rect 1138 4508 1162 4564
rect 1218 4508 4207 4564
rect 4263 4508 4287 4564
rect 4343 4508 4367 4564
rect 4423 4508 4447 4564
rect 4503 4508 4527 4564
rect 4583 4508 6138 4564
rect 6194 4508 6218 4564
rect 6274 4508 6298 4564
rect 6354 4508 6378 4564
rect 6434 4508 6458 4564
rect 6514 4508 8068 4564
rect 8124 4508 8148 4564
rect 8204 4508 8228 4564
rect 8284 4508 8308 4564
rect 8364 4508 8388 4564
rect 8444 4508 11346 4564
rect 11402 4508 11426 4564
rect 11482 4508 11506 4564
rect 11562 4508 11586 4564
rect 11642 4508 11666 4564
rect 11722 4508 12564 4564
rect 0 4476 12564 4508
rect 800 1218 11764 1260
rect 800 1162 842 1218
rect 898 1162 922 1218
rect 978 1162 1002 1218
rect 1058 1162 1082 1218
rect 1138 1162 1162 1218
rect 1218 1162 4207 1218
rect 4263 1162 4287 1218
rect 4343 1162 4367 1218
rect 4423 1162 4447 1218
rect 4503 1162 4527 1218
rect 4583 1162 6138 1218
rect 6194 1162 6218 1218
rect 6274 1162 6298 1218
rect 6354 1162 6378 1218
rect 6434 1162 6458 1218
rect 6514 1162 8068 1218
rect 8124 1162 8148 1218
rect 8204 1162 8228 1218
rect 8284 1162 8308 1218
rect 8364 1162 8388 1218
rect 8444 1162 11346 1218
rect 11402 1162 11426 1218
rect 11482 1162 11506 1218
rect 11562 1162 11586 1218
rect 11642 1162 11666 1218
rect 11722 1162 11764 1218
rect 800 1138 11764 1162
rect 800 1082 842 1138
rect 898 1082 922 1138
rect 978 1082 1002 1138
rect 1058 1082 1082 1138
rect 1138 1082 1162 1138
rect 1218 1082 4207 1138
rect 4263 1082 4287 1138
rect 4343 1082 4367 1138
rect 4423 1082 4447 1138
rect 4503 1082 4527 1138
rect 4583 1082 6138 1138
rect 6194 1082 6218 1138
rect 6274 1082 6298 1138
rect 6354 1082 6378 1138
rect 6434 1082 6458 1138
rect 6514 1082 8068 1138
rect 8124 1082 8148 1138
rect 8204 1082 8228 1138
rect 8284 1082 8308 1138
rect 8364 1082 8388 1138
rect 8444 1082 11346 1138
rect 11402 1082 11426 1138
rect 11482 1082 11506 1138
rect 11562 1082 11586 1138
rect 11642 1082 11666 1138
rect 11722 1082 11764 1138
rect 800 1058 11764 1082
rect 800 1002 842 1058
rect 898 1002 922 1058
rect 978 1002 1002 1058
rect 1058 1002 1082 1058
rect 1138 1002 1162 1058
rect 1218 1002 4207 1058
rect 4263 1002 4287 1058
rect 4343 1002 4367 1058
rect 4423 1002 4447 1058
rect 4503 1002 4527 1058
rect 4583 1002 6138 1058
rect 6194 1002 6218 1058
rect 6274 1002 6298 1058
rect 6354 1002 6378 1058
rect 6434 1002 6458 1058
rect 6514 1002 8068 1058
rect 8124 1002 8148 1058
rect 8204 1002 8228 1058
rect 8284 1002 8308 1058
rect 8364 1002 8388 1058
rect 8444 1002 11346 1058
rect 11402 1002 11426 1058
rect 11482 1002 11506 1058
rect 11562 1002 11586 1058
rect 11642 1002 11666 1058
rect 11722 1002 11764 1058
rect 800 978 11764 1002
rect 800 922 842 978
rect 898 922 922 978
rect 978 922 1002 978
rect 1058 922 1082 978
rect 1138 922 1162 978
rect 1218 922 4207 978
rect 4263 922 4287 978
rect 4343 922 4367 978
rect 4423 922 4447 978
rect 4503 922 4527 978
rect 4583 922 6138 978
rect 6194 922 6218 978
rect 6274 922 6298 978
rect 6354 922 6378 978
rect 6434 922 6458 978
rect 6514 922 8068 978
rect 8124 922 8148 978
rect 8204 922 8228 978
rect 8284 922 8308 978
rect 8364 922 8388 978
rect 8444 922 11346 978
rect 11402 922 11426 978
rect 11482 922 11506 978
rect 11562 922 11586 978
rect 11642 922 11666 978
rect 11722 922 11764 978
rect 800 898 11764 922
rect 800 842 842 898
rect 898 842 922 898
rect 978 842 1002 898
rect 1058 842 1082 898
rect 1138 842 1162 898
rect 1218 842 4207 898
rect 4263 842 4287 898
rect 4343 842 4367 898
rect 4423 842 4447 898
rect 4503 842 4527 898
rect 4583 842 6138 898
rect 6194 842 6218 898
rect 6274 842 6298 898
rect 6354 842 6378 898
rect 6434 842 6458 898
rect 6514 842 8068 898
rect 8124 842 8148 898
rect 8204 842 8228 898
rect 8284 842 8308 898
rect 8364 842 8388 898
rect 8444 842 11346 898
rect 11402 842 11426 898
rect 11482 842 11506 898
rect 11562 842 11586 898
rect 11642 842 11666 898
rect 11722 842 11764 898
rect 800 800 11764 842
rect 0 418 12564 460
rect 0 362 42 418
rect 98 362 122 418
rect 178 362 202 418
rect 258 362 282 418
rect 338 362 362 418
rect 418 362 5172 418
rect 5228 362 5252 418
rect 5308 362 5332 418
rect 5388 362 5412 418
rect 5468 362 5492 418
rect 5548 362 7103 418
rect 7159 362 7183 418
rect 7239 362 7263 418
rect 7319 362 7343 418
rect 7399 362 7423 418
rect 7479 362 12146 418
rect 12202 362 12226 418
rect 12282 362 12306 418
rect 12362 362 12386 418
rect 12442 362 12466 418
rect 12522 362 12564 418
rect 0 338 12564 362
rect 0 282 42 338
rect 98 282 122 338
rect 178 282 202 338
rect 258 282 282 338
rect 338 282 362 338
rect 418 282 5172 338
rect 5228 282 5252 338
rect 5308 282 5332 338
rect 5388 282 5412 338
rect 5468 282 5492 338
rect 5548 282 7103 338
rect 7159 282 7183 338
rect 7239 282 7263 338
rect 7319 282 7343 338
rect 7399 282 7423 338
rect 7479 282 12146 338
rect 12202 282 12226 338
rect 12282 282 12306 338
rect 12362 282 12386 338
rect 12442 282 12466 338
rect 12522 282 12564 338
rect 0 258 12564 282
rect 0 202 42 258
rect 98 202 122 258
rect 178 202 202 258
rect 258 202 282 258
rect 338 202 362 258
rect 418 202 5172 258
rect 5228 202 5252 258
rect 5308 202 5332 258
rect 5388 202 5412 258
rect 5468 202 5492 258
rect 5548 202 7103 258
rect 7159 202 7183 258
rect 7239 202 7263 258
rect 7319 202 7343 258
rect 7399 202 7423 258
rect 7479 202 12146 258
rect 12202 202 12226 258
rect 12282 202 12306 258
rect 12362 202 12386 258
rect 12442 202 12466 258
rect 12522 202 12564 258
rect 0 178 12564 202
rect 0 122 42 178
rect 98 122 122 178
rect 178 122 202 178
rect 258 122 282 178
rect 338 122 362 178
rect 418 122 5172 178
rect 5228 122 5252 178
rect 5308 122 5332 178
rect 5388 122 5412 178
rect 5468 122 5492 178
rect 5548 122 7103 178
rect 7159 122 7183 178
rect 7239 122 7263 178
rect 7319 122 7343 178
rect 7399 122 7423 178
rect 7479 122 12146 178
rect 12202 122 12226 178
rect 12282 122 12306 178
rect 12362 122 12386 178
rect 12442 122 12466 178
rect 12522 122 12564 178
rect 0 98 12564 122
rect 0 42 42 98
rect 98 42 122 98
rect 178 42 202 98
rect 258 42 282 98
rect 338 42 362 98
rect 418 42 5172 98
rect 5228 42 5252 98
rect 5308 42 5332 98
rect 5388 42 5412 98
rect 5468 42 5492 98
rect 5548 42 7103 98
rect 7159 42 7183 98
rect 7239 42 7263 98
rect 7319 42 7343 98
rect 7399 42 7423 98
rect 7479 42 12146 98
rect 12202 42 12226 98
rect 12282 42 12306 98
rect 12362 42 12386 98
rect 12442 42 12466 98
rect 12522 42 12564 98
rect 0 0 12564 42
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3706 0 1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1624635492
transform 1 0 3706 0 -1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3430 0 1 3974
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 3430 0 -1 3974
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1624635492
transform 1 0 4810 0 1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1624635492
transform 1 0 4810 0 -1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1624635492
transform 1 0 5914 0 1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1624635492
transform 1 0 6190 0 -1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5914 0 -1 3974
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6098 0 -1 3974
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8122 0 1 3974
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1624635492
transform 1 0 7018 0 1 3974
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7754 0 -1 3974
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42
timestamp 1624635492
transform 1 0 7294 0 -1 3974
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7754 0 -1 3974
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8398 0 -1 3974
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8766 0 1 3974
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1624635492
transform 1 0 8398 0 -1 3974
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_30
timestamp 1624635492
transform 1 0 8674 0 1 3974
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_29
timestamp 1624635492
transform 1 0 8766 0 -1 3974
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 9134 0 1 3974
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 9134 0 -1 3974
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 3706 0 -1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 3430 0 -1 5062
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1624635492
transform 1 0 4810 0 -1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 6190 0 -1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1624635492
transform 1 0 5914 0 -1 5062
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_31
timestamp 1624635492
transform 1 0 6098 0 -1 5062
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1624635492
transform 1 0 7294 0 -1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp 1624635492
transform 1 0 8766 0 -1 5062
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1624635492
transform 1 0 8398 0 -1 5062
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 9134 0 -1 5062
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 3706 0 1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 3430 0 1 5062
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1624635492
transform 1 0 5270 0 1 5062
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp 1624635492
transform 1 0 4810 0 1 5062
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x6_B1
timestamp 1624635492
transform 1 0 5086 0 1 5062
box -38 -48 222 592
use sky130_fd_sc_hd__o221ai_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5638 0 1 5062
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 1624635492
transform 1 0 6282 0 1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1624635492
transform 1 0 7386 0 1 5062
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1624635492
transform 1 0 8766 0 1 5062
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1624635492
transform 1 0 8490 0 1 5062
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_32
timestamp 1624635492
transform 1 0 8674 0 1 5062
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 9134 0 1 5062
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 3706 0 -1 6150
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 3430 0 -1 6150
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1624635492
transform 1 0 5638 0 -1 6150
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_21
timestamp 1624635492
transform 1 0 5362 0 -1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp 1624635492
transform 1 0 4810 0 -1 6150
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x9_B1
timestamp 1624635492
transform 1 0 5454 0 -1 6150
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 6190 0 -1 6150
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1624635492
transform 1 0 6006 0 -1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_33
timestamp 1624635492
transform 1 0 6098 0 -1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 7294 0 -1 6150
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1624635492
transform 1 0 8766 0 -1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_54
timestamp 1624635492
transform 1 0 8398 0 -1 6150
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 9134 0 -1 6150
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3706 0 1 6150
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_x15_A
timestamp 1624635492
transform -1 0 4626 0 1 6150
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 3430 0 1 6150
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp 1624635492
transform 1 0 5270 0 1 6150
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1624635492
transform 1 0 4626 0 1 6150
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_1  x9
timestamp 1624635492
transform 1 0 5638 0 1 6150
box -38 -48 682 592
use sky130_fd_sc_hd__inv_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4994 0 1 6150
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_38
timestamp 1624635492
transform 1 0 6926 0 1 6150
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1624635492
transform 1 0 6282 0 1 6150
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  x2
timestamp 1624635492
transform -1 0 6926 0 1 6150
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1624635492
transform 1 0 8030 0 1 6150
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1624635492
transform 1 0 8766 0 1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1624635492
transform 1 0 8582 0 1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1624635492
transform 1 0 8674 0 1 6150
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 9134 0 1 6150
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 3706 0 1 7238
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_12
timestamp 1624635492
transform 1 0 4534 0 -1 7238
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1624635492
transform 1 0 3982 0 -1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 4534 0 -1 7238
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3982 0 -1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 3430 0 1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 3430 0 -1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 4810 0 1 7238
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1624635492
transform 1 0 5638 0 -1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_35
timestamp 1624635492
transform 1 0 6650 0 1 7238
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1624635492
transform 1 0 5914 0 1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_37
timestamp 1624635492
transform 1 0 6834 0 -1 7238
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1624635492
transform 1 0 6190 0 -1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1624635492
transform 1 0 6006 0 -1 7238
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1624635492
transform 1 0 6098 0 -1 7238
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  x3
timestamp 1624635492
transform 1 0 6558 0 -1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  x11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6282 0 1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1624635492
transform 1 0 7754 0 1 7238
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1624635492
transform 1 0 7846 0 -1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_45
timestamp 1624635492
transform 1 0 7570 0 -1 7238
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 7846 0 -1 7238
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1624635492
transform 1 0 8766 0 1 7238
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1624635492
transform 1 0 8490 0 1 7238
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1624635492
transform 1 0 8490 0 -1 7238
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform -1 0 8490 0 -1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1624635492
transform 1 0 8674 0 1 7238
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 9134 0 1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 9134 0 -1 7238
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 3706 0 -1 8326
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 3430 0 -1 8326
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 4810 0 -1 8326
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1624635492
transform 1 0 6190 0 -1 8326
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 5914 0 -1 8326
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1624635492
transform 1 0 6098 0 -1 8326
box -38 -48 130 592
use sky130_fd_sc_hd__a221oi_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6558 0 -1 8326
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1624635492
transform 1 0 7202 0 -1 8326
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1624635492
transform 1 0 8306 0 -1 8326
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 9134 0 -1 8326
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 3706 0 1 8326
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 3430 0 1 8326
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 4810 0 1 8326
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1624635492
transform 1 0 6650 0 1 8326
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1624635492
transform 1 0 5914 0 1 8326
box -38 -48 130 592
use sky130_fd_sc_hd__a221oi_1  x8
timestamp 1624635492
transform -1 0 6650 0 1 8326
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1624635492
transform 1 0 7386 0 1 8326
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_1  x10
timestamp 1624635492
transform 1 0 7018 0 1 8326
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_58
timestamp 1624635492
transform 1 0 8766 0 1 8326
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1624635492
transform 1 0 8490 0 1 8326
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1624635492
transform 1 0 8674 0 1 8326
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 9134 0 1 8326
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 3706 0 -1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 3430 0 -1 9414
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 4810 0 -1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624635492
transform 1 0 6190 0 -1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 5914 0 -1 9414
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1624635492
transform 1 0 6098 0 -1 9414
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624635492
transform 1 0 7294 0 -1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_58
timestamp 1624635492
transform 1 0 8766 0 -1 9414
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1624635492
transform 1 0 8398 0 -1 9414
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 9134 0 -1 9414
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624635492
transform 1 0 3706 0 1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 3430 0 1 9414
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624635492
transform 1 0 4810 0 1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1624635492
transform 1 0 5914 0 1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1624635492
transform 1 0 8122 0 1 9414
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1624635492
transform 1 0 7018 0 1 9414
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_58
timestamp 1624635492
transform 1 0 8766 0 1 9414
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1624635492
transform 1 0 8674 0 1 9414
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 9134 0 1 9414
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624635492
transform 1 0 3706 0 -1 10502
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 3430 0 -1 10502
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624635492
transform 1 0 4810 0 -1 10502
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624635492
transform 1 0 6190 0 -1 10502
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 5914 0 -1 10502
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1624635492
transform 1 0 6098 0 -1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624635492
transform 1 0 7294 0 -1 10502
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_58
timestamp 1624635492
transform 1 0 8766 0 -1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_54
timestamp 1624635492
transform 1 0 8398 0 -1 10502
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 9134 0 -1 10502
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_12
timestamp 1624635492
transform 1 0 4534 0 1 10502
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1624635492
transform 1 0 3982 0 1 10502
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 4534 0 1 10502
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 3706 0 1 10502
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 3430 0 1 10502
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1624635492
transform 1 0 5638 0 1 10502
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1624635492
transform 1 0 6190 0 1 10502
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_28
timestamp 1624635492
transform 1 0 6006 0 1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1624635492
transform 1 0 6098 0 1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_50
timestamp 1624635492
transform 1 0 8030 0 1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_42
timestamp 1624635492
transform 1 0 7294 0 1 10502
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1624635492
transform 1 0 8122 0 1 10502
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_54
timestamp 1624635492
transform 1 0 8398 0 1 10502
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1624635492
transform 1 0 8766 0 1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 9134 0 1 10502
box -38 -48 314 592
<< labels >>
rlabel metal2 s 9526 7076 10626 7300 6 INN
port 0 nsew signal input
rlabel metal2 s 9526 3120 10626 3344 6 INP
port 1 nsew signal input
rlabel metal2 s 9526 11032 10626 11256 6 Q
port 2 nsew signal tristate
rlabel metal2 s 2026 11032 3126 11256 6 VDD
port 3 nsew signal input
rlabel metal2 s 2026 7076 3126 7300 6 VSS
port 4 nsew signal input
rlabel metal2 s 2026 3120 3126 3344 6 clk
port 5 nsew signal input
rlabel metal2 s 8047 0 8467 14476 6 VPWR
port 6 nsew power bidirectional
rlabel metal2 s 6116 0 6536 14476 6 VPWR
port 7 nsew power bidirectional
rlabel metal2 s 4185 0 4605 14476 6 VPWR
port 8 nsew power bidirectional
rlabel metal2 s 11304 800 11764 13676 6 VPWR
port 9 nsew power bidirectional
rlabel metal2 s 800 800 1260 13676 4 VPWR
port 10 nsew power bidirectional
rlabel metal3 s 800 13216 11764 13676 6 VPWR
port 11 nsew power bidirectional
rlabel metal3 s 0 9575 12564 9935 6 VPWR
port 12 nsew power bidirectional
rlabel metal3 s 0 7026 12564 7386 6 VPWR
port 13 nsew power bidirectional
rlabel metal3 s 0 4477 12564 4837 6 VPWR
port 14 nsew power bidirectional
rlabel metal3 s 800 800 11764 1260 8 VPWR
port 15 nsew power bidirectional
rlabel metal2 s 12104 0 12564 14476 6 VGND
port 16 nsew ground bidirectional
rlabel metal2 s 7081 0 7501 14476 6 VGND
port 17 nsew ground bidirectional
rlabel metal2 s 5151 0 5571 14476 6 VGND
port 18 nsew ground bidirectional
rlabel metal2 s 0 0 460 14476 4 VGND
port 19 nsew ground bidirectional
rlabel metal3 s 0 14016 12564 14476 6 VGND
port 20 nsew ground bidirectional
rlabel metal3 s 0 8301 12564 8661 6 VGND
port 21 nsew ground bidirectional
rlabel metal3 s 0 5751 12564 6111 6 VGND
port 22 nsew ground bidirectional
rlabel metal3 s 0 0 12564 460 8 VGND
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12564 14476
<< end >>
