* NGSPICE file created from ACMP_SAR.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for ACMP abstract view
.subckt ACMP INN INP Q VDD VSS clk vccd2 vssd2
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

.subckt ACMP_SAR INN INP Q clk cmp cmp_sel data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] done rstn start vccd1 vssd1 vccd2 vssd2 vccd1_uq0 vccd1_uq1
+ vssd1_uq0 vssd1_uq1 vccd2_uq0 vccd2_uq1 vssd2_uq0 vssd2_uq1
XFILLER_79_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1707 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_22_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1718 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_50_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_488 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_104_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_93_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_53_280 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_398 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_105_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_169 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_63_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_927 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_949 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1559 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_46_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_84 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_46_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_53_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_83_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_228 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_64_397 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_43_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_702 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_735 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1356 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1378 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_062_ _050_/Y _099_/A _055_/X _058_/X _061_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _119_/D sky130_fd_sc_hd__o311a_2
XFILLER_3_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_2_176 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_2_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_65_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_61_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_6_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_575 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_55_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_559 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_510 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_24_581 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_532 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_587 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ _118_/CLK _114_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _114_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1197 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_109_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_128 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__080__A1 _094_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_25_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_494 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__071__A1 _069_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_45_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_351 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__062__A1 _050_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_35_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_80_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_291 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xoutput7 COMP/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 Q sky130_fd_sc_hd__clkbuf_2
XFILLER_76_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_8_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_134 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_22_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1708 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1719 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_572 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_113_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_113_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_917 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output9_A _114_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_939 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_58_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_96 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_631 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__050__A _111_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_87_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_170 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_83_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XPHY_725 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_COMP_INN input1/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_51_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_758 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_061_ _093_/A _093_/B _112_/Q _119_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _061_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__110__D _110_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_58_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_37_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_37_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_100_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_610 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_120 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_409 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_69_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_626 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_587 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_55_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_511 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_593 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_577 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ _118_/CLK _113_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _113_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1176 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_427 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XANTENNA__074__C1 _073_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_47_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__065__C1 _064_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_37_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_80_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__080__A2 _102_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_111_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_20_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__071__A2 _054_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_341 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_390 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_396 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_47_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__062__A2 _099_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_50_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_627 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_103_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_80_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xoutput8 _113_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[0] sky130_fd_sc_hd__clkbuf_2
Xoutput10 _115_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_76_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_117_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_107 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_94_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1709 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__053__A _082_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_77_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_641 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_9_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XANTENNA__113__D _113_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_95_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_584 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_490 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_907 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_929 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1539 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_109_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_109_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_67 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_117_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_77_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_160 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_73_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_41 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__108__D _108_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_6_643 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_6_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_530 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_726 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_704 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1303 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_748 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1369 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_060_ _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _093_/B sky130_fd_sc_hd__buf_6
XFILLER_109_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_59 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_185 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_30_712 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_10_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__092__B1 _105_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_37_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_472 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_517 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_33_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_132 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_688 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_118_176 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_109_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_638 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_211 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_70_100 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_55_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_501 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_512 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_545 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_567 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_112_ _118_/CLK _112_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _112_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_3_410 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_94_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__074__B1 _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_47_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__120__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_69_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_450 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__065__B1 _058_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_84_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__080__A3 _099_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_80_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__056__A _103_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_106_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_102_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__071__A3 _055_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_101_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_575 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_397 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__116__D _116_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_113_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_105 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_98_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__062__A3 _055_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_34_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_106_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_26_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xoutput9 _114_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[1] sky130_fd_sc_hd__clkbuf_2
Xoutput11 _116_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_350 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_32_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_117_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_501 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_67_512 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_62_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_653 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_58_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_1_596 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_88_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_91_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_83_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_99_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_191 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_908 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1529 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_79 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_117_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_37_76 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_85_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_26_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_53 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_hold1_A hold1/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_110_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_99_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_99_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_150 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_95_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__059__A _059_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_55_345 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_24_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_70_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_727 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_COMP_INP input2/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_738 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_749 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1359 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_48_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_64_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__119__D _119_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_73_197 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__092__A1 _106_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_49_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__092__B2 _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_37_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_37_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_484 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_80_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_529 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_118_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_199 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_106_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_223 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_102_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_18_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_502 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1101 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_557 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_111_ COMP/clk _111_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _111_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_579 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_422 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_407 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__074__A1 _072_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_75_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_34_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_95 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_62_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1690 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_84_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__065__A1 _063_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_92_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_431 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XANTENNA__072__A _107_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_88_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_28 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_88_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_48_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_354 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_587 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_398 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_106_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_111_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xoutput12 _117_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_103_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__110__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_117_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_262 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_53_284 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_41_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_107_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_91_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_17_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_909 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1519 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_117_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_114_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_95_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_162 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_717 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output7_A COMP/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_1305 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__075__A _106_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_1316 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1349 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_722 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_6_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_89_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__092__A2 _083_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_37_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_198 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_21_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_668 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__068__C1 _067_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_56_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_514 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_552 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_503 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1113 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_558 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_110_ _118_/CLK _110_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _110_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1124 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_434 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_419 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__074__A2 _054_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_74_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_74 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_34_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_62_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1691 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__065__A2 _099_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_84_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_1_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_316 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_92_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_300 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_322 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_344 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_366 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_399 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_4_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_113_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_112_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_34_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_0_clk_A clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_89_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__083__A _083_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_21_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_262 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xoutput13 _118_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_103_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_130 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_116 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_4_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_311 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_97_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_7_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__078__A _105_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_38_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_17_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1509 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_81_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_707 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1306 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__086__B1 _111_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_74_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_80_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_111_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__077__B1 _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_49_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_166 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_80_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_179 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_109_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_114_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__068__B1 _058_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_56_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_515 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_564 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_504 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1147 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_446 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_78_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__074__A3 _055_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_74_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_597 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1670 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1681 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__065__A3 _055_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_92_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_65_497 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_21_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_301 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_323 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_361 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_356 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_389 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_74_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_890 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_274 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xoutput14 _119_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_56_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_71_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_131 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_72_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_175 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_72_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_164 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_99_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_67_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ sky130_fd_sc_hd__diode_2
XFILLER_35_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_31_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_623 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_97_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_81_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_81_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__094__A _106_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_22_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_99_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_95_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_35_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_31_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_45_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__086__B2 _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__086__A1 _112_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_74_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_108_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__077__A1 _075_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_64_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_64_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_178 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_21_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_60_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_103 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_118_114 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_88_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_609 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__068__A1 _066_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_18_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_576 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_549 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1159 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__113__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_15_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_42_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1660 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1682 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1693 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_502 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_099_ _099_/A _099_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _104_/D sky130_fd_sc_hd__nor2_8
XFILLER_111_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_489 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_107_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_115_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__097__A _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_56_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_313 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_373 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_52_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_379 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output15_A _120_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_30_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_42_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_880 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1490 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
Xoutput15 _120_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 data[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_107_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_1_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_605 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_112_84 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_71_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_143 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_121 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_72_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_165 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_72_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_154 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_99_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_35_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__094__B _094_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_22_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_107_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_89_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_346 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_195 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_57_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_114_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_input6_A start vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_100_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_101_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_709 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1308 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__086__A2 _098_/A1 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_104_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__077__A2 _054_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_1_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_605 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_87_227 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XANTENNA__068__A2 _099_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_68_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_28_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_517 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_105_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_5 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_93_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_77 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_74_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1661 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_098_ _098_/A1 _099_/B input6/X _101_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _103_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_97_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_41 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_319 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_402 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_107_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_603 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_75_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_614 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_314 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_347 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_870 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
Xoutput16 _093_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 done sky130_fd_sc_hd__clkbuf_2
XANTENNA__103__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_115_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_731 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_17_617 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_112_52 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_21_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_35_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xclkbuf_0_clk clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_31_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_104_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_22_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_22_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_358 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_9_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_185 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_82_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__098__B1 input6/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_380 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_42_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_53_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_649 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_5_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__089__B1 _108_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_78_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_271 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_9_410 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_90_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1309 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_86_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_54_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_80_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_6_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__077__A3 _102_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_1_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_72_191 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_639 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__068__A3 _055_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_68_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_64_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_507 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_24_523 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XPHY_518 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_24_71 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1651 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1695 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_097_ _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _101_/A sky130_fd_sc_hd__inv_2
XFILLER_97_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_53 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_38_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_29_626 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_56_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_68_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_320 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_304 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_871 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_93_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_65_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_65_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_29 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_33_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_233 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_356 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_404 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_64 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_21_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_75_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_35_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_690 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_112_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_22_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_108_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_1_569 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_89_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_610 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_8_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_381 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XANTENNA__098__A1 _098_/A1 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__098__B2 _101_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_145 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_26_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__089__A1 _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__089__B2 _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_78_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__116__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_72_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_422 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_68_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_36_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__103__RESET_B hold1/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_54_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_42_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_6_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_92 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_508 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_535 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_519 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1118 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_109_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_24_83 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_1652 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1696 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_096_ _108_/Q _107_/Q _096_/C _096_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _099_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_97_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_402 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_61_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_102_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_316 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_332 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_349 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_338 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_87_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_872 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_079_ _059_/A _060_/A _106_/Q _113_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _079_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_112_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_210 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_245 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_368 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_102_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_711 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_416 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_76 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_21_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_79_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_50_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output13_A _118_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_15_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_43_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_680 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1290 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_541 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_54_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_268 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_22_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_67_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_32_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_12_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_113_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_393 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_90_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_23_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_98_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__098__A2 _099_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__089__A2 _083_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_76_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_434 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_input4_A cmp_sel vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_98_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_58_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_86_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_6_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_593 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_77_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_33_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_509 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_547 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_51_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1108 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__106__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_117_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1642 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1697 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_095_ _112_/Q _111_/Q _110_/Q _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _096_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_69_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_414 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_344 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_317 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_47_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__070__B1 _116_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_35_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_862 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_078_ _105_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _094_/B sky130_fd_sc_hd__clkinv_4
XFILLER_112_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_222 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_65_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__061__B1 _119_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_33_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_61_450 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_33_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_257 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_115_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_102_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_102_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_69_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_723 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_72_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_25_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_136 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_106_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_670 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_103_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_199 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_69_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_718 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_60_729 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_13_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_12_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_85_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_86_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_383 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_6_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_91_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_84_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_446 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_43_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_4_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_104_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_66_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_729 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_81_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_75 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_1_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_65_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_95_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1109 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_117_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_117_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1643 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1676 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1698 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_094_ _106_/Q _094_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _096_/C sky130_fd_sc_hd__or2_4
XFILLER_109_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_49_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_426 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_426 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_37_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_307 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_378 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_540 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_106_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_27_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__070__A1 _093_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_55_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_304 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_43_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_852 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_077_ _075_/Y _054_/A _102_/X _097_/A _076_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _114_/D sky130_fd_sc_hd__o311a_4
XFILLER_112_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_147 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_643 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__061__A1 _093_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_103_626 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_88_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_104 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_72_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_40_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_106_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__119__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_62_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_16_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_660 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_682 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1292 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_629 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_707 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_103_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xrepeater17 _083_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _098_/A1 sky130_fd_sc_hd__buf_8
XFILLER_52_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_490 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_148 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_395 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_29 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_590 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_118_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_104_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_103_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_103_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_13_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_518 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_8_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_719 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_66_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_10_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_682 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_73_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_114_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1600 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1666 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_093_ _093_/A _093_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _093_/Y sky130_fd_sc_hd__nor2_4
XFILLER_77_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_438 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_407 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xinput1 INN vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_37_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_319 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_563 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_55 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_641 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__070__A2 _093_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_55_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_842 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_1496 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_7_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_076_ _059_/A _060_/A _107_/Q _114_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _076_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_111_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_111_159 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__061__A2 _093_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_34_655 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_119_204 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_46 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_37_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_105 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_138 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_62_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_650 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_683 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1293 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_059_ _059_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _093_/A sky130_fd_sc_hd__buf_4
XFILLER_98_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_319 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_88_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_12_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_32_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_730 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XANTENNA__103__D _103_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_95_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_551 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_0_584 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_341 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_48_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output11_A _116_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_480 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1090 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__109__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_118_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_103_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_77_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_26 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_94_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_45_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_13_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_610 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_60 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_95_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_541 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_89_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_77_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_50 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_114_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__091__B1 _106_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_24_506 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__051__A _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_99_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_input2_A INP vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_59_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_1634 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_1689 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_092_ _106_/Q _083_/A _105_/Q _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _105_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_410 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_712 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_49_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__111__D _111_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_77_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_37_108 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_92_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__073__B1 _115_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_45_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_65_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_419 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_114_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
Xinput2 INP vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__064__B1 _118_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_37_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_303 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_575 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_67 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_653 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_74_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__070__A3 _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_70_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_810 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_832 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_854 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_887 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1486 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__106__D _106_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
X_075_ _106_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _075_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_93_501 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_34_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__061__A3 _112_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_119_216 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_455 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_103_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_36 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_24_100 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_177 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_166 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_46_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_662 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_640 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1250 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1261 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1283 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1294 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_058_ _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _058_/X sky130_fd_sc_hd__buf_6
XFILLER_98_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_107_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_467 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_563 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_88_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_48_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_31_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_470 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_492 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_93_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_10_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__054__A _054_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_89_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__114__D _114_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_4_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_67_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_72 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_95_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_31_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_673 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_85_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_60_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__109__D _109_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_41_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_95 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_114_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__091__B2 _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__091__A1 _107_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_24_518 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_17_581 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1624 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_88 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1657 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1679 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_091_ _107_/Q _083_/A _106_/Q _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _106_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_108_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__073__A1 _059_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_65_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_60_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_418 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xinput3 cmp vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 input3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__064__A1 _093_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_36_142 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_37_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_24_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_52_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_587 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_118_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_79 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_114_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_800 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_833 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1421 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_877 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_855 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_899 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
X_074_ _072_/Y _054_/A _055_/X _097_/A _073_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _115_/D sky130_fd_sc_hd__o311a_1
XFILLER_111_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_228 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_115_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_103_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_329 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_111_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_112 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XANTENNA__057__A _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_52_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_395 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_46_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_62_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_652 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__117__D _117_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_685 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1284 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_057_ _104_/Q _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _097_/A sky130_fd_sc_hd__or2_4
XFILLER_97_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_21_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_115_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_479 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_32_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_570 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_581 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_597 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_31_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_460 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_482 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1070 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_174 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_109_ _118_/CLK _109_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_490 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__100__B1 _120_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_18_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_84 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_75_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_290 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_39_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_460 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_82_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_67_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_57_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_176 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__091__A2 _083_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_17_593 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1625 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1669 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
X_090_ _108_/Q _083_/A _107_/Q _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _107_/D
+ sky130_fd_sc_hd__a22o_4
XFILLER_108_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__073__A2 _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_60_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_14_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
Xinput4 cmp_sel vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _102_/S sky130_fd_sc_hd__buf_4
XFILLER_49_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__064__A2 _093_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_64_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_349 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_74_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_801 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_845 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1422 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_889 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_073_ _059_/A _060_/A _108_/Q _115_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _073_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_104_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_34_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__102__S _102_/S vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_111_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_112_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_71_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_146 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XANTENNA__057__B _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_52_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_108 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_20_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_713 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_101_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_620 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_680 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_642 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1241 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_675 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1274 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_697 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_056_ _103_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _060_/A sky130_fd_sc_hd__buf_6
XFILLER_97_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_672 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_722 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_593 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_35_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_450 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_483 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1093 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_186 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
X_108_ COMP/clk _108_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _108_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_112_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_18 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__100__A1 _081_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_57_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_390 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_68_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_12_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_291 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_69_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_472 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__081__A _112_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_104_511 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_53_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_199 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_70_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_64 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_5_410 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_0_170 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XANTENNA__076__B1 _114_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_49_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__067__B1 _117_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_23_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_11_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1615 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1648 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1659 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_704 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_104_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__073__A3 _108_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_115_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xinput5 rstn vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 hold1/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__064__A3 _111_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_64_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_802 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1478 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_11_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_072_ _107_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _072_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_64_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_109 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_32_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_21_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_725 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_610 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1231 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_692 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_687 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1242 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_698 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1286 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1297 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_055_ _102_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _055_/X sky130_fd_sc_hd__buf_6
XFILLER_97_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_66_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_93_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_61_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_22_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_30_684 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_79_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_345 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_194 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_113_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_28_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_462 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1050 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_473 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1083 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_107_ _118_/CLK _107_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _107_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_165 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_1094 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_112_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_584 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_22_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_103_247 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_89_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__100__A2 _054_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_69_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_72_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_25_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_0_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_90_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_292 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_484 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_82_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_523 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_38_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_26_540 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_72_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_422 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_41 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__076__A1 _059_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_49_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_484 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_36_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_392 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_32_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__067__A1 _093_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1616 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_1649 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_29 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xinput6 start vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_83_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_421 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_36_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__112__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_64_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_105_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_49 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_113_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_825 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1468 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
X_071_ _069_/Y _054_/A _055_/X _058_/X _070_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _116_/D sky130_fd_sc_hd__o311a_1
XFILLER_105_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_65_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_402 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_33_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_284 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_600 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_633 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1243 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1265 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1276 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1298 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_054_ _054_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _099_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_109_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_112_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_30_696 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_0_578 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_87_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_335 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_75_357 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_452 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1040 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_485 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_496 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ COMP/clk _106_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _106_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_1095 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_243 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_50_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__100__A3 _102_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_69_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__095__A _112_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_25_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_8_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XPHY_293 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_98_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_82_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_535 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_1_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_54_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_71 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_434 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_53 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_68_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__076__A2 _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_0_183 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_91_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__067__A2 _093_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_293 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_54_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1606 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_59 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1639 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_330 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_6_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_115_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_102 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_36_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_815 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1469 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_070_ _093_/A _093_/B _109_/Q _116_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _070_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_105_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_80 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_14_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _118_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_21_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_366 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_87_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_601 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_634 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1211 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1266 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_053_ _082_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _054_/A sky130_fd_sc_hd__buf_4
XFILLER_109_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_517 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_19_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_414 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_36_90 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_25_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_552 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_107_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_106_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_568 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_75_369 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_90_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_475 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_497 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_145 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
X_105_ COMP/clk _105_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _105_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1096 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_116_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__095__B _111_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_80_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__088__B1 _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_76_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_261 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_113_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__079__B1 _113_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_94_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_446 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_119_83 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_442 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__076__A3 _107_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_48_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_113_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__067__A3 _110_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XPHY_1607 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1629 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_41 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_512 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_26_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_361 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_91_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_114 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_113_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_827 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1459 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_58_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_61_426 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_389 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_56_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_55_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_55_242 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_602 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_24_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_635 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_668 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1256 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_052_ _059_/A _103_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _082_/A sky130_fd_sc_hd__nand2_8
XFILLER_109_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_529 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_69_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_37_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_37_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_119_564 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_106_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_102_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_186 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_498 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_104_ _118_/CLK _104_/D hold1/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _104_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1086 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 COMP/clk
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1097 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_598 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_116_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_7_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_153 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__095__C _110_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_80_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_473 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_21_462 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_119_361 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__088__A1 _110_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__088__B2 _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_76_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_101 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_102_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_44_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_251 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_33_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_273 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_295 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_113_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__079__A1 _059_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__115__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_94_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_62_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_38_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_58_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_1_620 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_95_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_48_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_454 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_17_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_117_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1619 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_53 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_58_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_524 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_54_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_126 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_605 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_817 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output8_A _113_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_51_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_839 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_73_221 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_73_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_438 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_60 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_418 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_24_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_724 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_118_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_254 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_625 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_658 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_120_ COMP/clk _120_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _120_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1268 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1279 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_051_ _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _059_/A sky130_fd_sc_hd__inv_4
XFILLER_11_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_11_73 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_116_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_165 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_102_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_460 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_477 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_11_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
X_103_ COMP/clk _103_/D hold1/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _103_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1098 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_94_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_360 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_165 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_84_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__095__D _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_80_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_485 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_373 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_5_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_108_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__088__A2 _098_/A1 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_76_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_91_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_230 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_33_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__079__A2 _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
Xhold1 hold1/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_466 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_66_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_58_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_73_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_170 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_119_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_95_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_175 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_466 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_680 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_91_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1609 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_569 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_41_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__105__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_107_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__101__A _101_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_39_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_138 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_17_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_617 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_807 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1406 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_829 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1439 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_117_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_50 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_37_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_102_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_55_266 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_615 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_604 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1203 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_174 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_24_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_648 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_050_ _111_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _050_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_85 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_30_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_188 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_106_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_114_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_199 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_401 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_423 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_494 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_467 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ COMP/Q input3/X _102_/S vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _102_/X sky130_fd_sc_hd__mux2_8
XFILLER_7_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_148 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_7_159 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_113_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_398 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_62_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_990 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_65_383 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_92_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_394 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_21_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_497 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_56_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_44_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_231 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XPHY_242 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_291 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__079__A3 _106_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_3_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_94_445 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_81_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_26_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_12 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_103_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_56 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_88_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_478 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_63_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_86_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_65_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_515 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_53_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_107_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_67_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_629 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_808 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_819 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1429 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_40 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_10_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_118_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_153 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_110_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_610 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_278 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_102_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_605 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_70_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1204 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_186 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_1259 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_97 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_6_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XANTENNA__118__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_92_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_523 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_578 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_9_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_88_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_539 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_318 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_57_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_435 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_101_ _101_/A _101_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _120_/D sky130_fd_sc_hd__or2_2
XPHY_479 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output16_A _093_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_63_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_42_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_980 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_991 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1590 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_160 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_112_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_111_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_38_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_320 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_102_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_88_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_44_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_221 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_31_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_8_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_119_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_107_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_100 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_251 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_95_24 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_340 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_56_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_398 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_71_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_287 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_55_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_104_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_427 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_91_257 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_809 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1419 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_104_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_27_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_41 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_63 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_10_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_96_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_45_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_165 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_114_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_617 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_606 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1205 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_30_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_500 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_92_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_21_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_535 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_425 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_447 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_100_ _081_/Y _054_/A _102_/X _120_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _101_/B
+ sky130_fd_sc_hd__o31a_1
XPHY_1035 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_7_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_1057 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_981 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1580 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1591 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_111_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_271 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_119_332 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_31_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_233 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_52_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_288 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__108__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_99_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_88 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_112 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_1_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_36 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_28_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_266 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_67_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_299 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__090__B1 _107_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_63_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_31_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_65_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_314 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_81_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_336 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_14_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_1_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_49_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_269 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_247 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_45_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1409 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_31_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_614 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_104_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_100_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_31 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_26_152 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_27_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_64 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_26_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_108_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_55_236 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_24_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_607 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_65_512 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_60_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_547 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_107_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_88_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_431 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_415 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_22_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_15_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_960 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1592 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_97_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_93_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_283 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_119_344 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_75_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_71_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_71_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_223 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_256 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_289 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XANTENNA__104__D _104_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_79_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_67_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_75_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_790 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_90 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_98_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_97_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_97_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_470 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_26_515 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_26_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_65_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_119_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_119_185 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_1_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_48 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_146 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__090__B2 _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__090__A1 _108_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_35_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_104_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_89_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_45_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_626 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XANTENNA__052__A _059_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_86_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_21 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_27_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_43 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_76 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_108_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__112__D _112_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_64_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_608 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_668 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_619 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1229 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_7 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__107__D _107_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_108_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_416 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_427 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1048 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1059 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_105_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_321 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_86_181 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_15_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_950 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_089_ _109_/Q _083_/A _108_/Q _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _108_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_97_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_38_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_398 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_61_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_479 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_119_378 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__060__A _060_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_75_107 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_68_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_262 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_235 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_79_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__120__D _120_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_47_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output14_A _119_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_43_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_780 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_30_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_791 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1390 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__055__A _102_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_119_197 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_119_175 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_79_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_0_158 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__115__D _115_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_5_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__090__A2 _083_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_35_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_50_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_140 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_39_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_22_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_108_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_9_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_9_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_50_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__052__B _103_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_input5_A rstn vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_58_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_86_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_227 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_54_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_44 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_6_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_111_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_104_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_113 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_68_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_36_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_609 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1219 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__063__A _110_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_105_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_82_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1720 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_113_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_417 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__058__A _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_1005 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_439 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1016 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1049 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_105_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_193 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_103_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__118__D _118_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_15_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_962 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_175 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_088_ _110_/Q _098_/A1 _109_/Q _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _109_/D
+ sky130_fd_sc_hd__a22o_4
XFILLER_112_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_61_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_83_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_274 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_269 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_770 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_450 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_26_506 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_65_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_61_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_29 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XANTENNA__084__B1 _058_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_28_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_60_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_94_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_85_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_16_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_86_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_86_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_112_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_325 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_494 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_26_369 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_41_317 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XANTENNA__066__A _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_6_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_76_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_409 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_32_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_36_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_12 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_26_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_45 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_67 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_89 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_50_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_66_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_398 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1209 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_1710 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_65_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_33_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_506 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_87_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_407 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_12_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_429 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1006 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_489 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_51_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1039 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_930 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_952 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1584 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1595 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_087_ _111_/Q _098_/A1 _110_/Q _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _110_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_6_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_112_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_69_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_97_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_34_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_61_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_303 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_108_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_102_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__069__A _108_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_25_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_215 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_12_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_43_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_760 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_7_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_93 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_112_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_495 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_0_71 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_186 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_100 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_59 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_18 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_76_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_69_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__084__A1 _081_/Y vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_28_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_57_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_650 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_94_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_62_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_590 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_98_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_26_337 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_392 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XANTENNA__082__A _082_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_108_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_116_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_40_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_598 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_113_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_98_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_26_178 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_54_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_68 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XANTENNA__111__CLK COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_57 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_50_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_91_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_605 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_36_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_117_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_113_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_36_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1700 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_73_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_518 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_61_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_402 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_408 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_419 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1007 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__102__A0 COMP/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_59_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_324 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_368 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_55_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_920 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XPHY_964 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1585 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_6_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_086_ _112_/Q _098_/A1 _111_/Q _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _111_/D
+ sky130_fd_sc_hd__a22o_4
XFILLER_109_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_80_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_102_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_69_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__085__A _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_109_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_772 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_7_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_069_ _108_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _069_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_112_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_198 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_80_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_112 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_103_502 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__084__A2 _098_/A1 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_69_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_541 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_684 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output12_A _117_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XPHY_580 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1190 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_29 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_349 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_91_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_106_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_94_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_26_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_36 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_69 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__093__A _093_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_22_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_105 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_110_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_48_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_639 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_input3_A cmp vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_113_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1701 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_117_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_506 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_37_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_73_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_409 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_1019 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_20_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__102__A1 input3/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_59_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_87_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_74_336 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_27_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_910 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_998 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1586 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
X_085_ _104_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _085_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_88_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_77_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_80_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_349 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_717 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_102_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_84_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_380 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_206 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_233 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_217 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_40_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_33_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__087__B1 _110_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XCOMP input1/X input2/X COMP/Q COMP/VDD COMP/VSS COMP/clk vccd2_uq1 vssd2_uq1 ACMP
XFILLER_58_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_740 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_795 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1394 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_7_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_068_ _066_/Y _099_/A _055_/X _058_/X _067_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _117_/D sky130_fd_sc_hd__o311a_2
XFILLER_98_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_66_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_509 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_9_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_146 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_608 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_203 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_44_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__096__A _108_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_37_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_553 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_40_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_680 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_79_203 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_696 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_570 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_54_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_34_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_62_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_52_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_141 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_113_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_209 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_66_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_37 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_81_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__093__B _093_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_41_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_653 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_103_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_77_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_19 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_66_11 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_103_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_91_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_91_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_51_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_701 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_99_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1702 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_COMP_clk COMP/clk vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_18_423 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_73_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_110_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_109 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_1009 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_20_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_99_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XANTENNA__099__A _099_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_59_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_348 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_27_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_27_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_900 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_944 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1598 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1587 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_084_ _081_/Y _098_/A1 _058_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _112_/D sky130_fd_sc_hd__o21ai_4
XFILLER_88_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_90 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_14_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_103_729 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_88_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_52_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_207 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_24_245 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_37_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_4_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_106_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__087__A1 _111_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__087__B2 _085_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_58_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_74_101 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_730 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_752 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_785 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1395 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_7_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_067_ _093_/A _093_/B _110_/Q _117_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _067_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_38_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_66_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_34_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_158 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_215 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_304 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__114__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA__096__B _107_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_25_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_52_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_80_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_52_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_692 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_403 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_118_191 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_109_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_4_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_215 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XPHY_560 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_8_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_582 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1181 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_119_ COMP/clk _119_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _119_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_34_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_62_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_107_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_103_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_107_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_20 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_95_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_51_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_390 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_8_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_8_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_454 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_81_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_81_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_34_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_10_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_17_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_26_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_95_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_59_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1703 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_435 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_630 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_41_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_99_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__099__B _099_/B vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_59_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_912 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1500 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_945 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_967 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_083_ _083_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _083_/X sky130_fd_sc_hd__buf_1
XFILLER_10_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_12_50 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_88_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_21_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_471 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_88_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_84_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_219 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_12_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_257 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_52_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_3_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_3_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__087__A2 _098_/A1 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_114_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_113 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_360 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_720 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_742 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_753 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_30_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_786 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_11_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_797 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_066_ _109_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _066_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_115_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_227 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_316 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__096__C _096_/C vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_52_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_415 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_107_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_4_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_621 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_79_227 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_95_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_561 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_583 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_118_ _118_/CLK _118_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _118_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_503 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_30_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_115_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_103_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_75_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_16_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_output10_A _115_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ sky130_fd_sc_hd__diode_2
XFILLER_31_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_380 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_573 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__104__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_59_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_81_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_633 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_606 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_41_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_598 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_99_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_113 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_67_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_609 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_70_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_52_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1704 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_92_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_447 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_675 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_642 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_13_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_114_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_118_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_47_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA_input1_A INN vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_86_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_86_199 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_67_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_902 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_42_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_935 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1501 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_601 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_957 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_634 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1578 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_082_ _082_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _083_/A sky130_fd_sc_hd__clkinv_8
XFILLER_12_73 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_111_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_398 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_37_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_33_247 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_525 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_52_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_569 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_103_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_84_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_56_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_52_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_33_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_20_464 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_125 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_710 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_11_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_787 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_475 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_798 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_065_ _063_/Y _099_/A _055_/X _058_/X _064_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _118_/D sky130_fd_sc_hd__o311a_2
XFILLER_78_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_105_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_78_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_486 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_520 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_542 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_66_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_34_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_73_191 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_115_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_88_239 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_17 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_328 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XANTENNA__096__D _096_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_71_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_100_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_0_655 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_48_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_63_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_372 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_562 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_117_ _118_/CLK _117_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _117_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1194 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_515 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_94_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_93_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_93_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_81_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_1_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_526 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_331 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_53_640 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_508 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_96_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_452 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_75_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_29_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_43_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_370 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_585 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_6_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_100_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_607 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_29 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_41_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_645 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_106_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_85_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_18_618 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_106 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_17_139 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_41_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_31_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_544 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_110_648 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_49_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_99_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_98_142 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_100_125 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_82_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_67_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_448 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_70_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_35_481 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1705 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_108_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_104_453 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_681 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_459 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_14_687 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_76_370 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_36_201 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_49_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_407 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_567 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_118_534 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_9_691 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_412 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__117__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_82_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1513 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_613 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_23_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_958 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_646 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1579 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_081_ _112_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _081_/Y sky130_fd_sc_hd__inv_4
XFILLER_12_85 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_88_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_78_624 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_294 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_705 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_33_259 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_721 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_92_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_204 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_52_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_476 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_58_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_102_732 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_101_220 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_101_253 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_286 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_510 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_137 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_114_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_543 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_700 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_733 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_432 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_777 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_799 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1398 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_487 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_064_ _093_/A _093_/B _111_/Q _118_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _064_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_97_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_498 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_532 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_65_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_81_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_565 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_554 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_88 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_34_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_117 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_334 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_6_480 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_367 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_111_562 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_111_595 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_60_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_119_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_667 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_351 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_384 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_56_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_71_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_552 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_116_ _118_/CLK _116_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _116_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_315 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_527 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_104 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_22_516 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__104__RESET_B hold1/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_89_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_89_538 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_115 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_45_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_25_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_652 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__080__C1 _079_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_71_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_715 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_107_676 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_420 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_96_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_0_464 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_192 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_45_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__071__C1 _070_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_43_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_360 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_371 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_54 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_87 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_123 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_112_156 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_446 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_27_619 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_50_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_429 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_657 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_89_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_700 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_15_41 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_5_556 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_589 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_64_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_110 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_86_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_137 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_39_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_54_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_35_493 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_23_622 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1706 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1717 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_237 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_504 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_270 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_537 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_465 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_77_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_100_693 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_14_699 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_13_187 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_96_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_36_213 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_419 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_9_670 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_8_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_118_579 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_105_229 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_424 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_457 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_714 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_157 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_82_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_63_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_249 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_915 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_463 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_948 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_658 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1569 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_10_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
X_080_ _094_/B _102_/X _099_/A _097_/A _079_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1
+ _113_/D sky130_fd_sc_hd__o311a_2
XFILLER_12_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_5_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_636 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_93_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_703 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_505 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_6_651 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_549 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_5_172 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_68_135 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_96_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_68_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_83_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_24_216 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_64_385 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_32_282 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_60_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_87_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_2
XFILLER_101_265 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_298 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_522 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_74_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_114_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_555 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_31_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_701 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_723 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_444 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XPHY_789 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_310 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1388 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1399 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_499 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_109_343 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
X_063_ _110_/Q vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _063_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_571 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_208 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_93_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_65_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_19_577 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_46_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_46_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_42_591 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_119_129 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__107__CLK _118_/CLK vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_89_709 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_492 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_115_379 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_514 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_25_569 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_119_663 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_118_140 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_69_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_0_679 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_87_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_47_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_85_58 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_75_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_18_30 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_28_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_322 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_12_720 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_520 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_1141 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_115_ _118_/CLK _115_/D vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 _115_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1196 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_151 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_109_184 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_539 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_3_451 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_327 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_59_70 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_38_116 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_93_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_19_396 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_22_528 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_61_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_61_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_600 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_69_241 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_97_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_127 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_57_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_55_39 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_355 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_53_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__080__B1 _097_/A vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_53_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_71_27 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_119_460 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_5_727 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_105_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_20_42 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_29_51 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_0_476 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_75_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_90_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_90_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__071__B1 _058_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_45_94 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_43_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XPHY_361 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_394 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_561 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_372 vssd1_uq1 vccd1_uq1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_594 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_61_82 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_66 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_6_99 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_112_168 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_550 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_79_583 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_39_436 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_39_469 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_35_664 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XANTENNA__062__B1 _058_/X vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__diode_2
XFILLER_35_697 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_50_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_108_408 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_116_441 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_2_708 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_104_669 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_106_78 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_58_712 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__fill_1
XFILLER_97_391 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_57_277 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_72_225 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_82_15 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_72_258 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_25_163 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
XFILLER_15_53 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_4
XFILLER_25_196 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_111 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_40_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_64_726 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_6
XFILLER_32_612 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_3
XFILLER_68_3 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_113_400 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_122 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_98_144 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_101_628 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_339 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_12
XFILLER_86_306 vssd1_uq1 vssd1_uq1 vccd1_uq1 vccd1_uq1 sky130_fd_sc_hd__decap_8
.ends

