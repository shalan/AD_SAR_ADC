module ACMP (INN,
    INP,
    Q,
    VDD,
    VSS,
    clk,
    vccd2,
    vssd2);
 input INN;
 input INP;
 output Q;
 input VDD;
 input VSS;
 input clk;
 input vccd2;
 input vssd2;

 sky130_fd_sc_hd__nor3_1 x10 (.A(net5),
    .B(net1),
    .C(net7),
    .Y(net12),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__nor3_1 x11 (.A(net12),
    .B(net6),
    .C(net2),
    .Y(net7),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__inv_1 x15 (.A(clk),
    .Y(clkb),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__inv_1 x2 (.A(net3),
    .Y(net6),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__inv_1 x3 (.A(net4),
    .Y(net5),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__o221ai_1 x6 (.A1(net9),
    .A2(net9),
    .B1(clk),
    .B2(net11),
    .C1(net4),
    .Y(net3),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__a221oi_1 x7 (.A1(net9),
    .A2(net9),
    .B1(clkb),
    .B2(net10),
    .C1(net2),
    .Y(net1),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__a221oi_1 x8 (.A1(net8),
    .A2(net8),
    .B1(clkb),
    .B2(net10),
    .C1(net1),
    .Y(net2),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__o221ai_1 x9 (.A1(net8),
    .A2(net8),
    .B1(clk),
    .B2(net11),
    .C1(net3),
    .Y(net4),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_50 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_51 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_52 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_53 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_54 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_55 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_62 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_63 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_64 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_65 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_66 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_67 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_73 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__buf_1 input1 (.A(INN),
    .X(net8),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__buf_1 input2 (.A(INP),
    .X(net9),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__buf_1 input3 (.A(VDD),
    .X(net10),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(VSS),
    .X(net11),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__buf_1 output5 (.A(net12),
    .X(Q),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(INN),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(INP),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(VDD),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(VSS),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_x9_B1 (.DIODE(clk),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_x6_B1 (.DIODE(clk),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__diode_2 ANTENNA_x15_A (.DIODE(clk),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_0_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_1_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_1_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_2_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_2_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_2_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_2_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_2_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_2_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_2_55 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_3_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_3_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_3_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_3_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_3_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_3_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_4_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_4_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_4_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_4_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_4_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_4_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_4_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_5_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_5_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_5_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_5_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_5_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_5_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_6_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_6_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_6_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_6_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_6_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_6_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_6_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_7_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_7_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_7_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_7_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_7_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_7_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_8_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_8_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_8_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_8_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_8_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_8_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_8_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_9_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_9_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_9_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_9_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_9_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_9_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_10_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_10_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_10_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 FILLER_10_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_10_35 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_10_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_10_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_10_55 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_11_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_11_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_11_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_11_35 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_11_46 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_11_53 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_11_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_12_6 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_12_12 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_12_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_12_28 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_12_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_12_34 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_12_38 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_8 FILLER_12_49 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_12_57 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_13_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_13_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_13_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 FILLER_13_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_8 FILLER_13_49 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_13_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_14_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_14_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_14_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 FILLER_14_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_14_35 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_14_46 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_14_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_14_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_15_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_15_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_15_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_15_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_8 FILLER_15_49 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_15_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_16_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_16_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_16_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_16_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_16_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_16_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_16_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_17_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_17_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_17_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_17_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_17_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_17_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_18_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_18_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_18_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_18_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_18_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_18_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_18_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_19_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_19_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_19_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_19_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_19_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_19_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_20_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_20_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_20_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_20_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_20_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_20_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_20_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_21_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_21_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_21_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_21_39 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_21_51 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_21_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_22_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_22_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_22_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_22_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_22_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_22_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_22_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_23_6 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_23_12 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_23_24 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_23_36 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_23_48 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_23_53 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_23_58 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_24_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_24_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_24_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_24_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_24_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_24_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
endmodule
