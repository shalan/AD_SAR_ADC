VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO adc
  CLASS BLOCK ;
  FOREIGN adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN INN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 124.480 250.000 125.080 ;
    END
  END INN
  PIN INP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 41.520 250.000 42.120 ;
    END
  END INP
  PIN Q
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 208.120 250.000 208.720 ;
    END
  END Q
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END clk
  PIN data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END data[0]
  PIN data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END data[1]
  PIN data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END data[2]
  PIN data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END data[3]
  PIN data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END data[4]
  PIN data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END data[5]
  PIN data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data[6]
  PIN data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END data[7]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END done
  PIN rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END rstn
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END start
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 236.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.880 172.640 236.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.880 122.640 236.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 236.880 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 236.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.880 147.640 236.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.880 97.640 236.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 236.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 244.260 236.880 ;
      LAYER met2 ;
        RECT 6.990 4.280 240.950 237.845 ;
        RECT 6.990 4.000 61.910 4.280 ;
        RECT 62.750 4.000 186.570 4.280 ;
        RECT 187.410 4.000 240.950 4.280 ;
      LAYER met3 ;
        RECT 4.400 236.960 246.000 237.825 ;
        RECT 4.000 213.200 246.000 236.960 ;
        RECT 4.400 211.800 246.000 213.200 ;
        RECT 4.000 209.120 246.000 211.800 ;
        RECT 4.000 207.720 245.600 209.120 ;
        RECT 4.000 188.040 246.000 207.720 ;
        RECT 4.400 186.640 246.000 188.040 ;
        RECT 4.000 162.880 246.000 186.640 ;
        RECT 4.400 161.480 246.000 162.880 ;
        RECT 4.000 138.400 246.000 161.480 ;
        RECT 4.400 137.000 246.000 138.400 ;
        RECT 4.000 125.480 246.000 137.000 ;
        RECT 4.000 124.080 245.600 125.480 ;
        RECT 4.000 113.240 246.000 124.080 ;
        RECT 4.400 111.840 246.000 113.240 ;
        RECT 4.000 88.080 246.000 111.840 ;
        RECT 4.400 86.680 246.000 88.080 ;
        RECT 4.000 62.920 246.000 86.680 ;
        RECT 4.400 61.520 246.000 62.920 ;
        RECT 4.000 42.520 246.000 61.520 ;
        RECT 4.000 41.120 245.600 42.520 ;
        RECT 4.000 37.760 246.000 41.120 ;
        RECT 4.400 36.360 246.000 37.760 ;
        RECT 4.000 13.280 246.000 36.360 ;
        RECT 4.400 11.880 246.000 13.280 ;
        RECT 4.000 10.000 246.000 11.880 ;
  END
END adc
END LIBRARY

