module dac_8bit(
    input wire d0,
    input wire d1,
    input wire d2,
    input wire d3,
    input wire d4,
    input wire d5,
    input wire d6,
    input wire d7,
    
    input wire inp1,
    
    output wire out_v
);



endmodule