magic
tech sky130A
magscale 1 2
timestamp 1626450099
<< checkpaint >>
rect -1260 -1260 101104 65372
<< locali >>
rect 45770 56616 90780 56624
rect 95360 56616 96184 56620
rect 45770 56582 96184 56616
rect 45770 56432 45824 56582
rect 95364 56578 96184 56582
rect 45770 56398 45777 56432
rect 45811 56398 45824 56432
rect 45770 56388 45824 56398
rect 96148 56528 96184 56578
rect 21190 56340 21746 56342
rect 21190 56336 37460 56340
rect 20370 56334 37460 56336
rect 20370 56317 48154 56334
rect 20370 56292 20399 56317
rect 20372 56283 20399 56292
rect 20433 56296 48154 56317
rect 20433 56292 21390 56296
rect 20433 56283 20452 56292
rect 20372 56272 20452 56283
rect 45768 56252 45818 56258
rect 45768 56218 45777 56252
rect 45811 56218 45818 56252
rect 796 55687 854 55734
rect 796 55653 811 55687
rect 845 55653 854 55687
rect 796 55648 854 55653
rect 808 55513 844 55514
rect 808 55479 809 55513
rect 843 55479 844 55513
rect 808 55478 844 55479
rect 20382 55473 20456 55494
rect 20382 55439 20399 55473
rect 20433 55439 20456 55473
rect 20382 54622 20456 55439
rect 45768 54878 45818 56218
rect 48098 55724 48154 56296
rect 48092 55705 48158 55724
rect 48092 55671 48111 55705
rect 48145 55671 48158 55705
rect 48092 55656 48158 55671
rect 48098 55652 48154 55656
rect 48114 55503 48158 55508
rect 48114 55469 48119 55503
rect 48153 55469 48158 55503
rect 48114 55464 48158 55469
rect 20380 31254 20460 54622
rect 45768 32536 45816 54878
rect 96148 54264 96190 56528
rect 96146 32684 96190 54264
rect 96146 32642 96196 32684
rect 43122 31793 43162 32466
rect 43122 31759 43124 31793
rect 43158 31759 43162 31793
rect 43122 31744 43162 31759
rect 90376 31817 90468 32454
rect 90376 31783 90401 31817
rect 90435 31783 90468 31817
rect 90376 31720 90468 31783
rect 43110 31579 43164 31588
rect 43110 31545 43120 31579
rect 43154 31545 43164 31579
rect 43110 31534 43164 31545
rect 20380 31224 20466 31254
rect 20386 7872 20466 31224
rect 43116 30468 43164 31534
rect 43110 29448 43164 30468
rect 43102 28990 43164 29448
rect 90376 31463 90434 31522
rect 90376 31429 90389 31463
rect 90423 31429 90434 31463
rect 20386 7374 20472 7872
rect 20382 7350 20472 7374
rect 20382 6942 20468 7350
rect 20600 7246 20702 7420
rect 20776 6942 20878 7036
rect 20382 6852 20884 6942
rect 20386 6850 20884 6852
rect 21292 3892 21352 5110
rect 24370 4036 24430 5254
rect 27710 4244 27770 5502
rect 31104 4426 31164 5796
rect 34346 4620 34406 6082
rect 37808 4762 37868 6518
rect 43102 6354 43154 28990
rect 67809 7395 68298 7416
rect 67809 7394 67910 7395
rect 67809 7360 67832 7394
rect 67866 7361 67910 7394
rect 67944 7361 67986 7395
rect 68020 7394 68143 7395
rect 68020 7361 68065 7394
rect 67866 7360 68065 7361
rect 68099 7361 68143 7394
rect 68177 7361 68219 7395
rect 68253 7361 68298 7395
rect 68099 7360 68298 7361
rect 67809 7321 68298 7360
rect 67809 7320 67911 7321
rect 67809 7286 67833 7320
rect 67867 7287 67911 7320
rect 67945 7287 67987 7321
rect 68021 7320 68144 7321
rect 68021 7287 68066 7320
rect 67867 7286 68066 7287
rect 68100 7287 68144 7320
rect 68178 7287 68220 7321
rect 68254 7287 68298 7321
rect 68100 7286 68298 7287
rect 67809 7240 68298 7286
rect 67809 7239 67913 7240
rect 67809 7205 67835 7239
rect 67869 7206 67913 7239
rect 67947 7206 67989 7240
rect 68023 7239 68146 7240
rect 68023 7206 68068 7239
rect 67869 7205 68068 7206
rect 68102 7206 68146 7239
rect 68180 7206 68222 7240
rect 68256 7206 68298 7240
rect 68102 7205 68298 7206
rect 67809 7166 68298 7205
rect 67809 7165 67914 7166
rect 67809 7131 67836 7165
rect 67870 7132 67914 7165
rect 67948 7132 67990 7166
rect 68024 7165 68147 7166
rect 68024 7132 68069 7165
rect 67870 7131 68069 7132
rect 68103 7132 68147 7165
rect 68181 7132 68223 7166
rect 68257 7132 68298 7166
rect 68103 7131 68298 7132
rect 67809 7083 68298 7131
rect 43092 4954 43158 6354
rect 48502 5101 48572 5116
rect 78542 5112 78638 5724
rect 81690 5114 81788 6064
rect 85120 5494 85182 6460
rect 85120 5160 85190 5494
rect 85120 5134 85202 5160
rect 85126 5132 85202 5134
rect 48502 5067 48523 5101
rect 48557 5067 48572 5101
rect 48502 5052 48572 5067
rect 78540 5085 78640 5112
rect 78540 5051 78570 5085
rect 78604 5051 78640 5085
rect 81688 5078 81790 5114
rect 81688 5070 81722 5078
rect 78540 5024 78640 5051
rect 81690 5044 81722 5070
rect 81756 5070 81790 5078
rect 85126 5098 85142 5132
rect 85176 5098 85202 5132
rect 85126 5070 85202 5098
rect 81756 5044 81788 5070
rect 85126 5058 85190 5070
rect 78542 5018 78638 5024
rect 81690 5014 81788 5044
rect 88292 4960 89642 4964
rect 90376 4960 90434 31429
rect 93032 31158 93112 32596
rect 96150 32384 96196 32642
rect 96320 32098 96520 32114
rect 96320 32064 96331 32098
rect 96365 32064 96520 32098
rect 96320 32050 96520 32064
rect 93930 31956 93980 31984
rect 93930 31922 93967 31956
rect 93930 31892 93980 31922
rect 96172 31426 96214 31632
rect 96172 31182 96218 31426
rect 96172 31162 96212 31182
rect 93540 31158 96212 31162
rect 93032 31092 96212 31158
rect 93032 31088 93562 31092
rect 88292 4954 90434 4960
rect 43090 4942 90434 4954
rect 43090 4941 44244 4942
rect 43090 4907 44166 4941
rect 44200 4908 44244 4941
rect 44278 4908 44320 4942
rect 44354 4908 90434 4942
rect 44200 4907 90434 4908
rect 43090 4894 90434 4907
rect 43090 4890 85110 4894
rect 85226 4890 90434 4894
rect 43090 4876 43236 4890
rect 88292 4878 90434 4890
rect 85120 4798 85182 4824
rect 85120 4764 85134 4798
rect 85168 4790 85182 4798
rect 85168 4764 85194 4790
rect 37800 4758 63320 4762
rect 85120 4758 85194 4764
rect 37800 4747 85194 4758
rect 37800 4746 38760 4747
rect 37800 4712 38682 4746
rect 38716 4713 38760 4746
rect 38794 4713 38836 4747
rect 38870 4713 85194 4747
rect 38716 4712 85194 4713
rect 37800 4700 85194 4712
rect 37800 4696 85178 4700
rect 37800 4690 63320 4696
rect 37808 4682 37868 4690
rect 34350 4594 34406 4620
rect 81688 4602 81790 4642
rect 44280 4600 81790 4602
rect 44280 4598 81724 4600
rect 39300 4594 81724 4598
rect 34350 4581 81724 4594
rect 34350 4580 35215 4581
rect 34350 4546 35137 4580
rect 35171 4547 35215 4580
rect 35249 4547 35291 4581
rect 35325 4566 81724 4581
rect 81758 4598 81790 4600
rect 81758 4566 81788 4598
rect 35325 4547 81788 4566
rect 35171 4546 81788 4547
rect 34350 4542 81788 4546
rect 34350 4538 81758 4542
rect 34350 4534 70790 4538
rect 34350 4530 44304 4534
rect 34350 4528 39342 4530
rect 34448 4526 39342 4528
rect 31098 4418 36684 4426
rect 42164 4418 57422 4422
rect 31098 4414 65052 4418
rect 31098 4412 72694 4414
rect 31098 4411 31597 4412
rect 31098 4377 31519 4411
rect 31553 4378 31597 4411
rect 31631 4378 31673 4412
rect 31707 4402 72694 4412
rect 78542 4402 78638 4410
rect 31707 4387 78638 4402
rect 31707 4378 78574 4387
rect 31553 4377 78574 4378
rect 31098 4366 78574 4377
rect 31104 4358 31164 4366
rect 36646 4358 78574 4366
rect 42164 4353 78574 4358
rect 78608 4353 78638 4387
rect 42164 4350 78638 4353
rect 57366 4346 78638 4350
rect 65008 4342 78638 4346
rect 78534 4332 78638 4342
rect 27698 4240 33728 4244
rect 27698 4233 75364 4240
rect 27698 4232 27924 4233
rect 27698 4198 27846 4232
rect 27880 4199 27924 4232
rect 27958 4199 28000 4233
rect 28034 4227 75364 4233
rect 28034 4199 75311 4227
rect 27880 4198 75311 4199
rect 27698 4193 75311 4198
rect 75345 4196 75364 4227
rect 75345 4193 75362 4196
rect 27698 4186 75362 4193
rect 27710 4176 27770 4186
rect 75290 4178 75362 4186
rect 71794 4036 71862 4040
rect 24370 4034 71862 4036
rect 24370 4031 71812 4034
rect 24370 4030 24856 4031
rect 24370 3996 24778 4030
rect 24812 3997 24856 4030
rect 24890 3997 24932 4031
rect 24966 4000 71812 4031
rect 71846 4000 71862 4034
rect 24966 3997 58626 4000
rect 24812 3996 58626 3997
rect 24370 3994 58626 3996
rect 24370 3992 39590 3994
rect 71794 3990 71862 4000
rect 46996 3892 48574 3902
rect 21286 3890 27752 3892
rect 40626 3890 48574 3892
rect 21286 3885 48574 3890
rect 21286 3880 48521 3885
rect 21286 3879 21382 3880
rect 21286 3845 21304 3879
rect 21338 3846 21382 3879
rect 21416 3846 21458 3880
rect 21492 3851 48521 3880
rect 48555 3851 48574 3885
rect 21492 3846 48574 3851
rect 21338 3845 48574 3846
rect 21286 3838 48574 3845
rect 21286 3832 47092 3838
rect 21424 3830 26450 3832
rect 27734 3830 40650 3832
<< viali >>
rect 45777 56398 45811 56432
rect 20399 56283 20433 56317
rect 45777 56218 45811 56252
rect 811 55653 845 55687
rect 809 55479 843 55513
rect 20399 55439 20433 55473
rect 48111 55671 48145 55705
rect 48119 55469 48153 55503
rect 43124 31759 43158 31793
rect 90401 31783 90435 31817
rect 43120 31545 43154 31579
rect 90389 31429 90423 31463
rect 67832 7360 67866 7394
rect 67910 7361 67944 7395
rect 67986 7361 68020 7395
rect 68065 7360 68099 7394
rect 68143 7361 68177 7395
rect 68219 7361 68253 7395
rect 67833 7286 67867 7320
rect 67911 7287 67945 7321
rect 67987 7287 68021 7321
rect 68066 7286 68100 7320
rect 68144 7287 68178 7321
rect 68220 7287 68254 7321
rect 67835 7205 67869 7239
rect 67913 7206 67947 7240
rect 67989 7206 68023 7240
rect 68068 7205 68102 7239
rect 68146 7206 68180 7240
rect 68222 7206 68256 7240
rect 67836 7131 67870 7165
rect 67914 7132 67948 7166
rect 67990 7132 68024 7166
rect 68069 7131 68103 7165
rect 68147 7132 68181 7166
rect 68223 7132 68257 7166
rect 48523 5067 48557 5101
rect 78570 5051 78604 5085
rect 81722 5044 81756 5078
rect 85142 5098 85176 5132
rect 96331 32064 96365 32098
rect 93967 31922 94001 31956
rect 44166 4907 44200 4941
rect 44244 4908 44278 4942
rect 44320 4908 44354 4942
rect 85134 4764 85168 4798
rect 38682 4712 38716 4746
rect 38760 4713 38794 4747
rect 38836 4713 38870 4747
rect 35137 4546 35171 4580
rect 35215 4547 35249 4581
rect 35291 4547 35325 4581
rect 81724 4566 81758 4600
rect 31519 4377 31553 4411
rect 31597 4378 31631 4412
rect 31673 4378 31707 4412
rect 78574 4353 78608 4387
rect 27846 4198 27880 4232
rect 27924 4199 27958 4233
rect 28000 4199 28034 4233
rect 75311 4193 75345 4227
rect 24778 3996 24812 4030
rect 24856 3997 24890 4031
rect 24932 3997 24966 4031
rect 71812 4000 71846 4034
rect 21304 3845 21338 3879
rect 21382 3846 21416 3880
rect 21458 3846 21492 3880
rect 48521 3851 48555 3885
<< metal1 >>
rect 45766 56434 45824 56446
rect 45764 56432 45824 56434
rect 45764 56398 45777 56432
rect 45811 56398 45824 56432
rect 45764 56388 45824 56398
rect 20376 56317 20450 56338
rect 20376 56283 20399 56317
rect 20433 56283 20450 56317
rect 625 56021 1160 56042
rect 625 55854 634 56021
rect 803 56020 1160 56021
rect 625 55853 806 55854
rect 1149 55853 1160 56020
rect 625 55847 1160 55853
rect 796 55687 854 55847
rect 796 55653 811 55687
rect 845 55653 854 55687
rect 796 55513 854 55653
rect 796 55479 809 55513
rect 843 55479 854 55513
rect 796 55466 854 55479
rect 20376 55473 20450 56283
rect 45768 56254 45822 56388
rect 45766 56252 45822 56254
rect 45766 56218 45777 56252
rect 45811 56218 45822 56252
rect 45766 56202 45822 56218
rect 48092 55720 48158 55724
rect 48092 55705 48168 55720
rect 48092 55671 48111 55705
rect 48145 55671 48168 55705
rect 48092 55656 48168 55671
rect 48100 55518 48168 55656
rect 20376 55439 20399 55473
rect 20433 55439 20450 55473
rect 48098 55503 48168 55518
rect 48098 55469 48119 55503
rect 48153 55474 48168 55503
rect 48153 55469 48164 55474
rect 48098 55450 48164 55469
rect 20376 55420 20450 55439
rect 94792 32416 94880 32428
rect 94792 32364 94825 32416
rect 94877 32364 94880 32416
rect 94792 32352 94880 32364
rect 96320 32109 96658 32115
rect 96320 32098 96390 32109
rect 96320 32064 96331 32098
rect 96365 32064 96390 32098
rect 96320 32057 96390 32064
rect 96572 32057 96658 32109
rect 96320 32049 96658 32057
rect 96320 32048 96386 32049
rect 93703 31964 94020 31984
rect 93703 31912 93710 31964
rect 93813 31956 94020 31964
rect 93813 31922 93967 31956
rect 94001 31922 94020 31956
rect 93813 31912 94020 31922
rect 93703 31889 94020 31912
rect 43116 31804 43162 31820
rect 90362 31817 90468 31854
rect 43116 31793 43164 31804
rect 43116 31759 43124 31793
rect 43158 31759 43164 31793
rect 43116 31748 43164 31759
rect 90362 31783 90401 31817
rect 90435 31783 90468 31817
rect 43116 31588 43162 31748
rect 43110 31579 43162 31588
rect 43110 31545 43120 31579
rect 43154 31545 43162 31579
rect 43110 31534 43162 31545
rect 43116 31532 43162 31534
rect 90362 31463 90468 31783
rect 94048 31640 94160 31692
rect 94048 31588 94073 31640
rect 94125 31588 94160 31640
rect 94048 31554 94160 31588
rect 90362 31429 90389 31463
rect 90423 31429 90468 31463
rect 90362 31402 90468 31429
rect 67808 7395 68300 7473
rect 67808 7394 67910 7395
rect 67808 7360 67832 7394
rect 67866 7361 67910 7394
rect 67944 7361 67986 7395
rect 68020 7394 68143 7395
rect 68020 7361 68065 7394
rect 67866 7360 68065 7361
rect 68099 7361 68143 7394
rect 68177 7361 68219 7395
rect 68253 7361 68300 7395
rect 68099 7360 68300 7361
rect 67808 7321 68300 7360
rect 67808 7320 67911 7321
rect 67808 7286 67833 7320
rect 67867 7287 67911 7320
rect 67945 7287 67987 7321
rect 68021 7320 68144 7321
rect 68021 7287 68066 7320
rect 67867 7286 68066 7287
rect 68100 7287 68144 7320
rect 68178 7287 68220 7321
rect 68254 7287 68300 7321
rect 68100 7286 68300 7287
rect 67808 7240 68300 7286
rect 67808 7239 67913 7240
rect 67808 7205 67835 7239
rect 67869 7206 67913 7239
rect 67947 7206 67989 7240
rect 68023 7239 68146 7240
rect 68023 7206 68068 7239
rect 67869 7205 68068 7206
rect 68102 7206 68146 7239
rect 68180 7206 68222 7240
rect 68256 7206 68300 7240
rect 68102 7205 68300 7206
rect 67808 7166 68300 7205
rect 67808 7165 67914 7166
rect 67808 7131 67836 7165
rect 67870 7132 67914 7165
rect 67948 7132 67990 7166
rect 68024 7165 68147 7166
rect 68024 7132 68069 7165
rect 67870 7131 68069 7132
rect 68103 7132 68147 7165
rect 68181 7132 68223 7166
rect 68257 7132 68300 7166
rect 68103 7131 68300 7132
rect 48502 5108 48572 5116
rect 48502 5101 48574 5108
rect 48502 5067 48523 5101
rect 48557 5067 48574 5101
rect 48502 5052 48574 5067
rect 44152 4942 44376 4963
rect 44152 4941 44244 4942
rect 44152 4907 44166 4941
rect 44200 4908 44244 4941
rect 44278 4908 44320 4942
rect 44354 4908 44376 4942
rect 44200 4907 44376 4908
rect 38663 4747 38887 4762
rect 38663 4746 38760 4747
rect 38663 4712 38682 4746
rect 38716 4713 38760 4746
rect 38794 4713 38836 4747
rect 38870 4713 38887 4747
rect 38716 4712 38887 4713
rect 35118 4581 35342 4594
rect 35118 4580 35215 4581
rect 35118 4546 35137 4580
rect 35171 4547 35215 4580
rect 35249 4547 35291 4581
rect 35325 4547 35342 4581
rect 35171 4546 35342 4547
rect 31501 4412 31725 4426
rect 31501 4411 31597 4412
rect 31501 4377 31519 4411
rect 31553 4378 31597 4411
rect 31631 4378 31673 4412
rect 31707 4378 31725 4412
rect 31553 4377 31725 4378
rect 27829 4233 28053 4244
rect 27829 4232 27924 4233
rect 27829 4198 27846 4232
rect 27880 4199 27924 4232
rect 27958 4199 28000 4233
rect 28034 4199 28053 4233
rect 27880 4198 28053 4199
rect 24766 4031 24990 4042
rect 24766 4030 24856 4031
rect 24766 3996 24778 4030
rect 24812 3997 24856 4030
rect 24890 3997 24932 4031
rect 24966 3997 24990 4031
rect 24812 3996 24990 3997
rect 21287 3880 21511 3892
rect 21287 3879 21382 3880
rect 21287 3845 21304 3879
rect 21338 3846 21382 3879
rect 21416 3846 21458 3880
rect 21492 3846 21511 3880
rect 21338 3845 21511 3846
rect 21287 2237 21511 3845
rect 21287 2070 21314 2237
rect 21483 2070 21511 2237
rect 21287 2056 21511 2070
rect 24766 2237 24990 3996
rect 24766 2070 24793 2237
rect 24962 2070 24990 2237
rect 24766 2056 24990 2070
rect 27829 2236 28053 4198
rect 27829 2069 27856 2236
rect 28025 2069 28053 2236
rect 27829 2055 28053 2069
rect 31501 2236 31725 4377
rect 31501 2069 31528 2236
rect 31697 2069 31725 2236
rect 31501 2055 31725 2069
rect 35118 2235 35342 4546
rect 35118 2068 35145 2235
rect 35314 2068 35342 2235
rect 35118 2054 35342 2068
rect 38663 2235 38887 4712
rect 38663 2068 38690 2235
rect 38859 2068 38887 2235
rect 38663 2054 38887 2068
rect 44152 2236 44376 4907
rect 48512 3900 48574 5052
rect 48506 3885 48574 3900
rect 48506 3851 48521 3885
rect 48555 3851 48574 3885
rect 48506 3838 48574 3851
rect 44152 2069 44179 2236
rect 44348 2069 44376 2236
rect 44152 2055 44376 2069
rect 67808 2214 68300 7131
rect 71798 4040 71858 5234
rect 75288 4282 75364 5498
rect 85122 5160 85186 5188
rect 85122 5132 85202 5160
rect 78540 5085 78640 5112
rect 78540 5051 78570 5085
rect 78604 5051 78640 5085
rect 81688 5104 81790 5114
rect 81688 5078 81792 5104
rect 81688 5070 81722 5078
rect 78540 5024 78640 5051
rect 81694 5044 81722 5070
rect 81756 5044 81792 5078
rect 78542 4387 78638 5024
rect 81694 4600 81792 5044
rect 85122 5098 85142 5132
rect 85176 5098 85202 5132
rect 85122 5070 85202 5098
rect 85122 4856 85186 5070
rect 85114 4798 85186 4856
rect 85114 4764 85134 4798
rect 85168 4790 85186 4798
rect 85168 4764 85194 4790
rect 85114 4700 85194 4764
rect 85114 4684 85178 4700
rect 81694 4566 81724 4600
rect 81758 4566 81792 4600
rect 81694 4528 81792 4566
rect 78542 4370 78574 4387
rect 78540 4353 78574 4370
rect 78608 4353 78638 4387
rect 78540 4332 78638 4353
rect 75288 4240 75360 4282
rect 75288 4227 75364 4240
rect 75288 4193 75311 4227
rect 75345 4196 75364 4227
rect 75345 4193 75362 4196
rect 75288 4190 75362 4193
rect 75290 4178 75362 4190
rect 71794 4034 71862 4040
rect 71794 4000 71812 4034
rect 71846 4000 71862 4034
rect 71794 3990 71862 4000
rect 67808 2056 67823 2214
rect 67875 2213 68300 2214
rect 67932 2212 68053 2213
rect 68105 2212 68300 2213
rect 67808 2055 67880 2056
rect 68039 2055 68053 2212
rect 68269 2055 68300 2212
rect 67808 2053 68300 2055
<< via1 >>
rect 634 56020 803 56021
rect 634 55854 1149 56020
rect 806 55853 1149 55854
rect 94825 32364 94877 32416
rect 96390 32057 96572 32109
rect 93710 31912 93813 31964
rect 94073 31588 94125 31640
rect 21314 2070 21483 2237
rect 24793 2070 24962 2237
rect 27856 2069 28025 2236
rect 31528 2069 31697 2236
rect 35145 2068 35314 2235
rect 38690 2068 38859 2235
rect 44179 2069 44348 2236
rect 67823 2213 67875 2214
rect 67823 2212 67932 2213
rect 68053 2212 68105 2213
rect 67823 2056 68039 2212
rect 67880 2055 68039 2056
rect 68053 2055 68269 2212
<< metal2 >>
rect 799 63712 977 64112
rect 625 56021 1160 63712
rect 625 55854 634 56021
rect 803 56020 1160 56021
rect 625 55853 806 55854
rect 1149 55853 1160 56020
rect 24290 55972 25152 55982
rect 24290 55968 58282 55972
rect 24290 55916 58400 55968
rect 24290 55912 58282 55916
rect 25120 55910 58282 55912
rect 625 55847 1160 55853
rect 94810 32498 94880 32508
rect 94810 32442 94816 32498
rect 94872 32442 94880 32498
rect 94810 32416 94880 32442
rect 94810 32364 94825 32416
rect 94877 32364 94880 32416
rect 94810 32354 94880 32364
rect 96320 32152 97000 32200
rect 96320 32109 96668 32152
rect 96320 32057 96390 32109
rect 96572 32096 96668 32109
rect 96724 32096 96748 32152
rect 96804 32096 96828 32152
rect 96884 32096 96908 32152
rect 96964 32096 97000 32152
rect 96572 32057 97000 32096
rect 96320 32049 97000 32057
rect 93584 31964 93820 31984
rect 93584 31963 93710 31964
rect 93584 31907 93629 31963
rect 93685 31907 93709 31963
rect 93813 31912 93820 31964
rect 93765 31907 93820 31912
rect 93584 31889 93820 31907
rect 93934 31648 94146 31654
rect 93914 31640 94146 31648
rect 93914 31588 94073 31640
rect 94125 31588 94146 31640
rect 93914 31562 94146 31588
rect 93914 31302 93954 31562
rect 91012 31300 93958 31302
rect 90500 31264 93958 31300
rect 90500 31262 92030 31264
rect 90500 31260 91014 31262
rect 21288 2237 21509 2265
rect 21288 2070 21314 2237
rect 21483 2070 21509 2237
rect 21288 1169 21509 2070
rect 24767 2237 24988 2265
rect 24767 2070 24793 2237
rect 24962 2070 24988 2237
rect 24767 1169 24988 2070
rect 27830 2236 28051 2264
rect 27830 2069 27856 2236
rect 28025 2069 28051 2236
rect 27830 1169 28051 2069
rect 31502 2236 31723 2264
rect 31502 2069 31528 2236
rect 31697 2069 31723 2236
rect 31502 1169 31723 2069
rect 35119 2235 35340 2263
rect 35119 2068 35145 2235
rect 35314 2068 35340 2235
rect 35119 1169 35340 2068
rect 38664 2235 38885 2263
rect 38664 2068 38690 2235
rect 38859 2068 38885 2235
rect 38664 1169 38885 2068
rect 44153 2236 44374 2264
rect 44153 2069 44179 2236
rect 44348 2069 44374 2236
rect 44153 1169 44374 2069
rect 67808 2214 68300 2218
rect 67808 2056 67823 2214
rect 67875 2213 68300 2214
rect 67932 2212 68053 2213
rect 68105 2212 68300 2213
rect 67808 2055 67880 2056
rect 68039 2055 68053 2212
rect 68269 2055 68300 2212
rect 67808 1172 68300 2055
rect 21343 800 21458 1169
rect 24820 800 24935 1169
rect 21342 0 21458 800
rect 24819 0 24935 800
rect 27876 0 27992 1169
rect 31555 0 31671 1169
rect 35169 0 35285 1169
rect 38704 0 38820 1169
rect 44192 0 44308 1169
rect 67957 0 68073 1172
<< via2 >>
rect 11049 55906 11105 55963
rect 11136 55906 11192 55962
rect 11223 55906 11426 55963
rect 11453 55906 11509 55964
rect 11622 55963 11908 55964
rect 11540 55906 11596 55963
rect 11622 55906 11984 55963
rect 94816 32442 94872 32498
rect 96668 32096 96724 32152
rect 96748 32096 96804 32152
rect 96828 32096 96884 32152
rect 96908 32096 96964 32152
rect 93629 31907 93685 31963
rect 93709 31912 93710 31963
rect 93710 31912 93765 31963
rect 93709 31907 93765 31912
<< metal3 >>
rect 11020 56446 12070 56463
rect 11020 56445 11883 56446
rect 11020 56444 11818 56445
rect 11020 56443 11740 56444
rect 11020 56442 11609 56443
rect 11020 56441 11473 56442
rect 11020 56440 11408 56441
rect 11020 56439 11330 56440
rect 11020 56438 11194 56439
rect 11020 56369 11050 56438
rect 12018 56382 12070 56446
rect 11020 56302 11049 56369
rect 12017 56313 12070 56382
rect 11020 56238 11048 56302
rect 12016 56246 12070 56313
rect 11880 56245 12070 56246
rect 11802 56244 12070 56245
rect 11737 56243 12070 56244
rect 11606 56242 12070 56243
rect 11470 56241 12070 56242
rect 11392 56240 12070 56241
rect 11327 56239 12070 56240
rect 11191 56238 12070 56239
rect 2837 56146 3901 56164
rect 2837 56145 3724 56146
rect 2837 56144 3659 56145
rect 2837 56143 3581 56144
rect 2837 56142 3450 56143
rect 2837 56141 3314 56142
rect 2837 56140 3249 56141
rect 2837 56139 3171 56140
rect 2837 56138 3035 56139
rect 2837 56069 2891 56138
rect 3859 56082 3901 56146
rect 2837 56005 2890 56069
rect 3858 56013 3901 56082
rect 3722 56012 3901 56013
rect 3644 56011 3901 56012
rect 3579 56010 3901 56011
rect 3448 56009 3901 56010
rect 3312 56008 3901 56009
rect 3234 56007 3901 56008
rect 3169 56006 3901 56007
rect 3033 56005 3901 56006
rect 2837 55995 3901 56005
rect 2837 55994 3724 55995
rect 2837 55993 3659 55994
rect 2837 55992 3581 55993
rect 2837 55991 3450 55992
rect 2837 55990 3314 55991
rect 2837 55989 3249 55990
rect 2837 55988 3171 55989
rect 2837 55987 3035 55988
rect 2837 55918 2891 55987
rect 3859 55931 3901 55995
rect 2837 55854 2890 55918
rect 3858 55862 3901 55931
rect 11020 55964 12070 56238
rect 11020 55963 11453 55964
rect 11020 55906 11049 55963
rect 11105 55962 11223 55963
rect 11105 55906 11136 55962
rect 11192 55906 11223 55962
rect 11426 55906 11453 55963
rect 11509 55963 11622 55964
rect 11908 55963 12070 55964
rect 11509 55906 11540 55963
rect 11596 55906 11622 55963
rect 11984 55906 12070 55963
rect 11020 55862 12070 55906
rect 3722 55861 3901 55862
rect 3644 55860 3901 55861
rect 3579 55859 3901 55860
rect 3448 55858 3901 55859
rect 3312 55857 3901 55858
rect 3234 55856 3901 55857
rect 3169 55855 3901 55856
rect 3033 55854 3901 55855
rect 2837 55464 3901 55854
rect 2837 55400 2866 55464
rect 2930 55400 2946 55464
rect 3010 55400 3026 55464
rect 3090 55400 3106 55464
rect 3170 55400 3199 55464
rect 3263 55400 3279 55464
rect 3343 55400 3359 55464
rect 3423 55400 3439 55464
rect 3503 55400 3534 55464
rect 3598 55400 3614 55464
rect 3678 55400 3694 55464
rect 3758 55400 3774 55464
rect 3838 55400 3901 55464
rect 2837 55381 3901 55400
rect 94810 32592 94890 32600
rect 94810 32528 94820 32592
rect 94884 32528 94890 32592
rect 94810 32518 94890 32528
rect 94810 32498 94880 32518
rect 94810 32442 94816 32498
rect 94872 32442 94880 32498
rect 94810 32434 94880 32442
rect 96515 32152 99401 33311
rect 96515 32096 96668 32152
rect 96724 32096 96748 32152
rect 96804 32096 96828 32152
rect 96884 32096 96908 32152
rect 96964 32141 99401 32152
rect 96964 32096 99844 32141
rect 96515 32021 99844 32096
rect 93584 31963 93817 31984
rect 93584 31907 93629 31963
rect 93685 31907 93709 31963
rect 93765 31907 93817 31963
rect 93584 30257 93817 31907
rect 96515 31051 99401 32021
rect 93584 30014 99416 30257
rect 93584 29854 99844 30014
rect 93584 29683 99416 29854
rect 93584 29682 93817 29683
<< via3 >>
rect 11883 56445 12018 56446
rect 11818 56444 12018 56445
rect 11740 56443 12018 56444
rect 11609 56442 12018 56443
rect 11473 56441 12018 56442
rect 11408 56440 12018 56441
rect 11330 56439 12018 56440
rect 11194 56438 12018 56439
rect 11050 56382 12018 56438
rect 11050 56369 12017 56382
rect 11049 56313 12017 56369
rect 11049 56302 12016 56313
rect 11048 56246 12016 56302
rect 11048 56245 11880 56246
rect 11048 56244 11802 56245
rect 11048 56243 11737 56244
rect 11048 56242 11606 56243
rect 11048 56241 11470 56242
rect 11048 56240 11392 56241
rect 11048 56239 11327 56240
rect 11048 56238 11191 56239
rect 3724 56145 3859 56146
rect 3659 56144 3859 56145
rect 3581 56143 3859 56144
rect 3450 56142 3859 56143
rect 3314 56141 3859 56142
rect 3249 56140 3859 56141
rect 3171 56139 3859 56140
rect 3035 56138 3859 56139
rect 2891 56082 3859 56138
rect 2891 56069 3858 56082
rect 2890 56013 3858 56069
rect 2890 56012 3722 56013
rect 2890 56011 3644 56012
rect 2890 56010 3579 56011
rect 2890 56009 3448 56010
rect 2890 56008 3312 56009
rect 2890 56007 3234 56008
rect 2890 56006 3169 56007
rect 2890 56005 3033 56006
rect 3724 55994 3859 55995
rect 3659 55993 3859 55994
rect 3581 55992 3859 55993
rect 3450 55991 3859 55992
rect 3314 55990 3859 55991
rect 3249 55989 3859 55990
rect 3171 55988 3859 55989
rect 3035 55987 3859 55988
rect 2891 55931 3859 55987
rect 2891 55918 3858 55931
rect 2890 55862 3858 55918
rect 2890 55861 3722 55862
rect 2890 55860 3644 55861
rect 2890 55859 3579 55860
rect 2890 55858 3448 55859
rect 2890 55857 3312 55858
rect 2890 55856 3234 55857
rect 2890 55855 3169 55856
rect 2890 55854 3033 55855
rect 2866 55400 2930 55464
rect 2946 55400 3010 55464
rect 3026 55400 3090 55464
rect 3106 55400 3170 55464
rect 3199 55400 3263 55464
rect 3279 55400 3343 55464
rect 3359 55400 3423 55464
rect 3439 55400 3503 55464
rect 3534 55400 3598 55464
rect 3614 55400 3678 55464
rect 3694 55400 3758 55464
rect 3774 55400 3838 55464
rect 94820 32528 94884 32592
<< metal4 >>
rect 2837 56146 3901 64112
rect 11006 56446 12070 64112
rect 23762 56558 49764 56562
rect 22752 56496 49764 56558
rect 22752 56494 23808 56496
rect 11006 56445 11883 56446
rect 11006 56444 11818 56445
rect 11006 56443 11740 56444
rect 11006 56442 11609 56443
rect 11006 56441 11473 56442
rect 11006 56440 11408 56441
rect 11006 56439 11330 56440
rect 11006 56438 11194 56439
rect 11006 56369 11050 56438
rect 12018 56382 12070 56446
rect 11006 56302 11049 56369
rect 12017 56313 12070 56382
rect 11006 56238 11048 56302
rect 12016 56246 12070 56313
rect 11880 56245 12070 56246
rect 11802 56244 12070 56245
rect 11737 56243 12070 56244
rect 11606 56242 12070 56243
rect 11470 56241 12070 56242
rect 11392 56240 12070 56241
rect 11327 56239 12070 56240
rect 11191 56238 12070 56239
rect 11006 56201 12070 56238
rect 2837 56145 3724 56146
rect 2837 56144 3659 56145
rect 2837 56143 3581 56144
rect 2837 56142 3450 56143
rect 2837 56141 3314 56142
rect 2837 56140 3249 56141
rect 2837 56139 3171 56140
rect 2837 56138 3035 56139
rect 2837 56069 2891 56138
rect 3859 56082 3901 56146
rect 2837 56005 2890 56069
rect 3858 56013 3901 56082
rect 3722 56012 3901 56013
rect 3644 56011 3901 56012
rect 3579 56010 3901 56011
rect 3448 56009 3901 56010
rect 3312 56008 3901 56009
rect 3234 56007 3901 56008
rect 3169 56006 3901 56007
rect 3033 56005 3901 56006
rect 2837 55995 3901 56005
rect 2837 55994 3724 55995
rect 2837 55993 3659 55994
rect 2837 55992 3581 55993
rect 2837 55991 3450 55992
rect 2837 55990 3314 55991
rect 2837 55989 3249 55990
rect 2837 55988 3171 55989
rect 2837 55987 3035 55988
rect 2837 55918 2891 55987
rect 3859 55931 3901 55995
rect 2837 55854 2890 55918
rect 3858 55862 3901 55931
rect 3722 55861 3901 55862
rect 3644 55860 3901 55861
rect 3579 55859 3901 55860
rect 3448 55858 3901 55859
rect 3312 55857 3901 55858
rect 3234 55856 3901 55857
rect 3169 55855 3901 55856
rect 3033 55854 3901 55855
rect 2837 55826 3901 55854
rect 22764 55684 22848 56494
rect 49692 55376 49762 56496
rect 91334 33132 94890 33202
rect 94816 32652 94890 33132
rect 94810 32646 94890 32652
rect 94810 32592 94888 32646
rect 94810 32528 94820 32592
rect 94884 32528 94888 32592
rect 94810 32522 94888 32528
use switch_layout  switch_layout_0
timestamp 1626450099
transform 1 0 93914 0 1 31372
box 40 154 2460 1180
use 7bitdac_layout  7bitdac_layout_0
timestamp 1626450099
transform 1 0 47558 0 1 7506
box -252 -2456 45562 48686
use 7bitdac_layout  7bitdac_layout_1
timestamp 1626450099
transform 1 0 252 0 1 7518
box -252 -2456 45562 48686
use res250_layout  res250_layout_0
timestamp 1626450099
transform 1 0 20392 0 1 7364
box 202 -342 510 -90
<< labels >>
rlabel locali s 21316 4998 21316 4998 4 d0
port 1 nsew
rlabel locali s 24396 5102 24396 5102 4 d1
port 2 nsew
rlabel locali s 27736 5214 27736 5214 4 d2
port 3 nsew
rlabel locali s 31132 5548 31132 5548 4 d3
port 4 nsew
rlabel locali s 34364 5674 34364 5674 4 d4
port 5 nsew
rlabel locali s 37842 4844 37842 4844 4 d5
port 6 nsew
rlabel locali s 43126 5106 43126 5106 4 d6
port 7 nsew
rlabel locali s 96200 31450 96200 31450 4 x2_out_v
port 8 nsew
rlabel locali s 96176 32606 96176 32606 4 x1_out_v
port 9 nsew
rlabel locali s 96452 32076 96452 32076 4 out_v
port 10 nsew
rlabel locali s 93952 31924 93952 31924 4 d7
port 11 nsew
rlabel locali s 804 55726 804 55726 4 inp1
port 12 nsew
rlabel locali s 20812 6930 20812 6930 4 x2_vref1
port 13 nsew
rlabel locali s 20652 7326 20652 7326 4 x1_vref5
port 14 nsew
rlabel metal2 s 799 62919 977 64112 4 inp1
port 12 nsew
rlabel metal2 s 93978 31602 93978 31602 4 gnd!
port 15 nsew
rlabel metal2 s 38704 0 38820 800 4 d5
port 6 nsew
rlabel metal2 s 35169 0 35285 800 4 d4
port 5 nsew
rlabel metal2 s 31555 0 31671 800 4 d3
port 4 nsew
rlabel metal2 s 27876 0 27992 800 4 d2
port 3 nsew
rlabel metal2 s 24819 0 24935 800 4 d1
port 2 nsew
rlabel metal2 s 21342 0 21458 800 4 d0
port 1 nsew
rlabel metal2 s 67957 0 68073 800 4 inp2
port 16 nsew
rlabel metal2 s 44192 0 44308 800 4 d6
port 7 nsew
rlabel metal3 s 99044 29854 99844 30014 4 d7
port 11 nsew
rlabel metal3 s 99044 32021 99844 32141 4 out_v
port 10 nsew
rlabel metal4 s 94864 32616 94864 32616 4 vdd!
port 17 nsew
rlabel metal4 s 11006 56201 12070 64112 4 gnd
port 18 nsew
rlabel metal4 s 2837 55826 3901 64112 4 vdd
port 19 nsew
<< properties >>
string FIXED_BBOX 0 0 99844 64112
string GDS_FILE gds/adc_wrapper.gds
string GDS_END 196322
string GDS_START 157834
<< end >>
